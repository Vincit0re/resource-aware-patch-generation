module top ( g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 );
input g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 ;
output g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 ;

wire n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , 
     n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , 
     n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , 
     n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , 
     n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , 
     n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , 
     n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , 
     n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , 
     n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , 
     n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , 
     n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , 
     n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , 
     n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , 
     n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , 
     n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , 
     n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , 
     n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , 
     n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , 
     n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , 
     n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , 
     n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , 
     n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , 
     n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , 
     n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , 
     n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , 
     n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , 
     n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , 
     n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , 
     n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , 
     n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , 
     n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , 
     n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , 
     n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , 
     n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , 
     n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , 
     n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , 
     n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , 
     n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , 
     n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , 
     n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , 
     n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , 
     n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , 
     n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , 
     n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , 
     n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , 
     n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , 
     n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , 
     n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , 
     n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , 
     n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , 
     n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , 
     n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , 
     n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , 
     n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , 
     n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , 
     n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , 
     n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , 
     n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , 
     n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , 
     n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , 
     n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , 
     n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , 
     n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , 
     n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , 
     n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , 
     n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , 
     n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , 
     n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , 
     n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , 
     n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , 
     n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , 
     n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , 
     n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , 
     n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , 
     n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , 
     n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , 
     n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , 
     n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , 
     n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , 
     n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , 
     n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , 
     n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , 
     n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , 
     n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , 
     n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , 
     n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , 
     n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , 
     n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , 
     n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , 
     n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , 
     n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , 
     n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , 
     n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , 
     n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , 
     n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , 
     n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , 
     n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , 
     n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , 
     n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , 
     n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , 
     n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , 
     n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , 
     n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , 
     n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , 
     n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , 
     n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , 
     n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , 
     n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , 
     n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , 
     n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , 
     n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , 
     n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , 
     n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , 
     n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , 
     n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , 
     n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , 
     n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , 
     n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , 
     n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , 
     n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , 
     n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , 
     n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , 
     n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , 
     n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , 
     n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , 
     n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , 
     n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , 
     n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , 
     n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , 
     n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , 
     n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , 
     n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , 
     n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , 
     n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , 
     n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , 
     n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , 
     n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , 
     n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , 
     n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , 
     n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , 
     n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , 
     n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , 
     n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , 
     n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , 
     n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , 
     n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , 
     n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , 
     n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , 
     n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , 
     n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , 
     n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , 
     n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , 
     n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , 
     n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , 
     n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , 
     n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , 
     n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , 
     n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , 
     n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , 
     n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , 
     n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , 
     n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , 
     n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , 
     n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , 
     n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , 
     n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , 
     n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , 
     n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , 
     n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , 
     n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , 
     n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , 
     n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , 
     n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , 
     n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , 
     n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , 
     n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , 
     n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , 
     n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , 
     n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , 
     n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , 
     n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , 
     n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , 
     n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , 
     n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , 
     n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , 
     n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , 
     n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , 
     n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , 
     n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , 
     n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , 
     n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , 
     n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , 
     n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , 
     n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , 
     n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , 
     n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , 
     n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , 
     n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , 
     n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , 
     n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , 
     n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , 
     n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , 
     n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , 
     n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , 
     n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , 
     n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , 
     n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , 
     n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , 
     n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , 
     n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , 
     n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , 
     n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , 
     n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 ;
buf ( n1  , g0 );
buf ( n2  , g1 );
buf ( n3  , g2 );
buf ( n4  , g3 );
buf ( n5  , g4 );
buf ( n6  , g5 );
buf ( n7  , g6 );
buf ( n8  , g7 );
buf ( n9  , g8 );
buf ( n10  , g9 );
buf ( n11  , g10 );
buf ( n12  , g11 );
buf ( n13  , g12 );
buf ( n14  , g13 );
buf ( n15  , g14 );
buf ( n16  , g15 );
buf ( n17  , g16 );
buf ( n18  , g17 );
buf ( n19  , g18 );
buf ( n20  , g19 );
buf ( n21  , g20 );
buf ( n22  , g21 );
buf ( n23  , g22 );
buf ( n24  , g23 );
buf ( n25  , g24 );
buf ( n26  , g25 );
buf ( n27  , g26 );
buf ( n28  , g27 );
buf ( n29  , g28 );
buf ( n30  , g29 );
buf ( n31  , g30 );
buf ( n32  , g31 );
buf ( n33  , g32 );
buf ( n34  , g33 );
buf ( n35  , g34 );
buf ( n36  , g35 );
buf ( n37  , g36 );
buf ( n38  , g37 );
buf ( n39  , g38 );
buf ( n40  , g39 );
buf ( n41  , g40 );
buf ( n42  , g41 );
buf ( n43  , g42 );
buf ( n44  , g43 );
buf ( n45  , g44 );
buf ( n46  , g45 );
buf ( n47  , g46 );
buf ( n48  , g47 );
buf ( g48 , n49  );
buf ( g49 , n50  );
buf ( g50 , n51  );
buf ( g51 , n52  );
buf ( g52 , n53  );
buf ( g53 , n54  );
buf ( g54 , n55  );
buf ( g55 , n56  );
buf ( g56 , n57  );
buf ( g57 , n58  );
buf ( g58 , n59  );
buf ( g59 , n60  );
buf ( g60 , n61  );
buf ( g61 , n62  );
buf ( g62 , n63  );
buf ( g63 , n64  );
buf ( g64 , n65  );
buf ( g65 , n66  );
buf ( g66 , n67  );
buf ( g67 , n68  );
buf ( g68 , n69  );
buf ( g69 , n70  );
buf ( g70 , n71  );
buf ( g71 , n72  );
buf ( g72 , n73  );
buf ( g73 , n74  );
buf ( g74 , n75  );
buf ( g75 , n76  );
buf ( g76 , n77  );
buf ( g77 , n78  );
buf ( g78 , n79  );
buf ( g79 , n80  );
buf ( g80 , n81  );
buf ( g81 , n82  );
buf ( g82 , n83  );
buf ( g83 , n84  );
buf ( g84 , n85  );
buf ( g85 , n86  );
buf ( g86 , n87  );
buf ( g87 , n88  );
buf ( g88 , n89  );
buf ( g89 , n90  );
buf ( g90 , n91  );
buf ( g91 , n92  );
buf ( g92 , n93  );
buf ( g93 , n94  );
buf ( g94 , n95  );
buf ( g95 , n96  );
buf ( g96 , n97  );
buf ( g97 , n98  );
buf ( n49 , 1'b0 );
buf ( n50 , 1'b0 );
buf ( n51 , 1'b0 );
buf ( n52 , 1'b0 );
buf ( n53 , 1'b0 );
buf ( n54 , 1'b0 );
buf ( n55 , 1'b0 );
buf ( n56 , 1'b0 );
buf ( n57 , 1'b0 );
buf ( n58 , 1'b0 );
buf ( n59 , 1'b0 );
buf ( n60 , 1'b0 );
buf ( n61 , 1'b0 );
buf ( n62 , 1'b0 );
buf ( n63 , 1'b0 );
buf ( n64 , 1'b0 );
buf ( n65 , 1'b0 );
buf ( n66 , 1'b0 );
buf ( n67 , n1722 );
buf ( n68 , n2127 );
buf ( n69 , n1959 );
buf ( n70 , n1928 );
buf ( n71 , n1981 );
buf ( n72 , n1942 );
buf ( n73 , n2014 );
buf ( n74 , n2005 );
buf ( n75 , n2024 );
buf ( n76 , n2043 );
buf ( n77 , n2062 );
buf ( n78 , n2079 );
buf ( n79 , n2094 );
buf ( n80 , n2122 );
buf ( n81 , n2112 );
buf ( n82 , n2118 );
buf ( n83 , n1947 );
buf ( n84 , n1913 );
buf ( n85 , n1950 );
buf ( n86 , n1965 );
buf ( n87 , n1970 );
buf ( n88 , n1984 );
buf ( n89 , n1990 );
buf ( n90 , n1998 );
buf ( n91 , n2029 );
buf ( n92 , n2051 );
buf ( n93 , n2068 );
buf ( n94 , n2073 );
buf ( n95 , n2084 );
buf ( n96 , n2100 );
buf ( n97 , n2121 );
buf ( n98 , n2129 );
nand ( n119 , n7 , n17 );
nand ( n120 , n1 , n23 );
xor ( n121 , n119 , n120 );
and ( n122 , n5 , n20 );
and ( n123 , n6 , n19 );
nor ( n124 , n122 , n123 );
not ( n125 , n124 );
nand ( n126 , n7 , n18 );
not ( n127 , n126 );
and ( n128 , n125 , n127 );
nand ( n129 , n5 , n19 );
nand ( n130 , n6 , n20 );
nor ( n131 , n129 , n130 );
nor ( n132 , n128 , n131 );
and ( n133 , n121 , n132 );
and ( n134 , n119 , n120 );
or ( n135 , n133 , n134 );
nand ( n136 , n6 , n18 );
nor ( n137 , n136 , n129 );
not ( n138 , n137 );
nand ( n139 , n136 , n129 );
nand ( n140 , n138 , n139 );
nand ( n141 , n3 , n22 );
nand ( n142 , n2 , n23 );
xor ( n143 , n141 , n142 );
nand ( n144 , n4 , n21 );
and ( n145 , n143 , n144 );
and ( n146 , n141 , n142 );
or ( n147 , n145 , n146 );
xor ( n148 , n140 , n147 );
nand ( n149 , n3 , n20 );
not ( n150 , n149 );
not ( n151 , n150 );
not ( n152 , n144 );
not ( n153 , n152 );
or ( n154 , n151 , n153 );
not ( n155 , n20 );
not ( n156 , n4 );
or ( n157 , n155 , n156 );
nand ( n158 , n3 , n21 );
nand ( n159 , n157 , n158 );
nand ( n160 , n154 , n159 );
nand ( n161 , n2 , n22 );
and ( n162 , n160 , n161 );
not ( n163 , n160 );
not ( n164 , n161 );
and ( n165 , n163 , n164 );
nor ( n166 , n162 , n165 );
not ( n167 , n166 );
and ( n168 , n148 , n167 );
and ( n169 , n140 , n147 );
nor ( n170 , n168 , n169 );
not ( n171 , n170 );
and ( n172 , n1 , n22 );
and ( n173 , n5 , n18 );
nor ( n174 , n172 , n173 );
not ( n175 , n174 );
nand ( n176 , n5 , n22 );
nand ( n177 , n1 , n18 );
or ( n178 , n176 , n177 );
nand ( n179 , n175 , n178 );
not ( n180 , n179 );
and ( n181 , n6 , n17 );
not ( n182 , n181 );
and ( n183 , n180 , n182 );
and ( n184 , n179 , n181 );
nor ( n185 , n183 , n184 );
not ( n186 , n185 );
and ( n187 , n171 , n186 );
and ( n188 , n170 , n185 );
nor ( n189 , n187 , n188 );
not ( n190 , n189 );
buf ( n191 , n137 );
not ( n192 , n191 );
and ( n193 , n4 , n19 );
not ( n194 , n193 );
not ( n195 , n21 );
not ( n196 , n2 );
or ( n197 , n195 , n196 );
nand ( n198 , n197 , n149 );
not ( n199 , n198 );
nand ( n200 , n2 , n20 );
nor ( n201 , n200 , n158 );
nor ( n202 , n199 , n201 );
not ( n203 , n202 );
or ( n204 , n194 , n203 );
or ( n205 , n202 , n193 );
nand ( n206 , n204 , n205 );
not ( n207 , n206 );
or ( n208 , n192 , n207 );
or ( n209 , n206 , n191 );
nand ( n210 , n208 , n209 );
not ( n211 , n210 );
not ( n212 , n159 );
not ( n213 , n212 );
not ( n214 , n161 );
and ( n215 , n213 , n214 );
not ( n216 , n150 );
nor ( n217 , n216 , n144 );
nor ( n218 , n215 , n217 );
not ( n219 , n218 );
and ( n220 , n211 , n219 );
and ( n221 , n210 , n218 );
nor ( n222 , n220 , n221 );
not ( n223 , n222 );
and ( n224 , n190 , n223 );
and ( n225 , n189 , n222 );
nor ( n226 , n224 , n225 );
not ( n227 , n226 );
xor ( n228 , n135 , n227 );
nor ( n229 , n131 , n124 );
and ( n230 , n229 , n127 );
not ( n231 , n229 );
and ( n232 , n231 , n126 );
or ( n233 , n230 , n232 );
not ( n234 , n233 );
not ( n235 , n234 );
nand ( n236 , n4 , n22 );
not ( n237 , n236 );
not ( n238 , n237 );
not ( n239 , n3 );
not ( n240 , n23 );
or ( n241 , n239 , n240 );
nand ( n242 , n2 , n24 );
nand ( n243 , n241 , n242 );
not ( n244 , n243 );
or ( n245 , n238 , n244 );
nand ( n246 , n3 , n24 );
not ( n247 , n246 );
not ( n248 , n142 );
nand ( n249 , n247 , n248 );
nand ( n250 , n245 , n249 );
not ( n251 , n250 );
xor ( n252 , n141 , n142 );
xor ( n253 , n252 , n144 );
not ( n254 , n253 );
or ( n255 , n251 , n254 );
or ( n256 , n253 , n250 );
nand ( n257 , n255 , n256 );
not ( n258 , n257 );
not ( n259 , n258 );
not ( n260 , n259 );
or ( n261 , n235 , n260 );
not ( n262 , n253 );
nand ( n263 , n262 , n250 );
nand ( n264 , n261 , n263 );
not ( n265 , n264 );
xor ( n266 , n119 , n120 );
xor ( n267 , n266 , n132 );
not ( n268 , n148 );
not ( n269 , n166 );
and ( n270 , n268 , n269 );
and ( n271 , n148 , n166 );
nor ( n272 , n270 , n271 );
xnor ( n273 , n267 , n272 );
not ( n274 , n273 );
or ( n275 , n265 , n274 );
not ( n276 , n267 );
nand ( n277 , n276 , n272 );
nand ( n278 , n275 , n277 );
not ( n279 , n278 );
xnor ( n280 , n228 , n279 );
not ( n281 , n280 );
nand ( n282 , n8 , n24 );
nand ( n283 , n1 , n17 );
nor ( n284 , n282 , n283 );
not ( n285 , n284 );
not ( n286 , n285 );
nand ( n287 , n4 , n23 );
not ( n288 , n287 );
not ( n289 , n288 );
nor ( n290 , n289 , n246 );
not ( n291 , n290 );
nand ( n292 , n5 , n21 );
xor ( n293 , n292 , n236 );
nand ( n294 , n249 , n243 );
xnor ( n295 , n293 , n294 );
not ( n296 , n295 );
or ( n297 , n291 , n296 );
not ( n298 , n292 );
and ( n299 , n294 , n236 );
not ( n300 , n294 );
and ( n301 , n300 , n237 );
nor ( n302 , n299 , n301 );
nand ( n303 , n298 , n302 );
nand ( n304 , n297 , n303 );
not ( n305 , n304 );
and ( n306 , n1 , n24 );
and ( n307 , n8 , n17 );
nor ( n308 , n306 , n307 );
nor ( n309 , n284 , n308 );
xor ( n310 , n309 , n233 );
xnor ( n311 , n310 , n257 );
not ( n312 , n311 );
or ( n313 , n305 , n312 );
nand ( n314 , n258 , n234 );
not ( n315 , n314 );
nand ( n316 , n259 , n233 );
not ( n317 , n316 );
or ( n318 , n315 , n317 );
nand ( n319 , n318 , n309 );
nand ( n320 , n313 , n319 );
not ( n321 , n320 );
not ( n322 , n321 );
not ( n323 , n264 );
xor ( n324 , n267 , n272 );
not ( n325 , n324 );
or ( n326 , n323 , n325 );
not ( n327 , n264 );
nand ( n328 , n273 , n327 );
nand ( n329 , n326 , n328 );
not ( n330 , n329 );
or ( n331 , n322 , n330 );
or ( n332 , n321 , n329 );
nand ( n333 , n331 , n332 );
not ( n334 , n333 );
or ( n335 , n286 , n334 );
not ( n336 , n329 );
nand ( n337 , n336 , n321 );
nand ( n338 , n335 , n337 );
buf ( n339 , n338 );
xor ( n340 , n281 , n339 );
not ( n341 , n340 );
xor ( n342 , n285 , n320 );
xnor ( n343 , n342 , n329 );
nand ( n344 , n7 , n19 );
nand ( n345 , n6 , n20 );
nor ( n346 , n344 , n345 );
not ( n347 , n346 );
nand ( n348 , n8 , n18 );
and ( n349 , n347 , n348 );
nand ( n350 , n344 , n345 );
not ( n351 , n350 );
nor ( n352 , n349 , n351 );
and ( n353 , n311 , n304 );
not ( n354 , n311 );
not ( n355 , n304 );
and ( n356 , n354 , n355 );
nor ( n357 , n353 , n356 );
xor ( n358 , n352 , n357 );
not ( n359 , n176 );
xor ( n360 , n288 , n246 );
not ( n361 , n360 );
or ( n362 , n359 , n361 );
nand ( n363 , n6 , n22 );
not ( n364 , n363 );
not ( n365 , n364 );
not ( n366 , n5 );
not ( n367 , n23 );
or ( n368 , n366 , n367 );
nand ( n369 , n4 , n24 );
nand ( n370 , n368 , n369 );
not ( n371 , n370 );
or ( n372 , n365 , n371 );
nand ( n373 , n5 , n24 );
not ( n374 , n373 );
nand ( n375 , n374 , n288 );
nand ( n376 , n372 , n375 );
nand ( n377 , n362 , n376 );
not ( n378 , n176 );
not ( n379 , n360 );
nand ( n380 , n378 , n379 );
nand ( n381 , n377 , n380 );
not ( n382 , n381 );
not ( n383 , n346 );
nand ( n384 , n383 , n350 );
xnor ( n385 , n384 , n348 );
xor ( n386 , n290 , n385 );
xnor ( n387 , n386 , n295 );
not ( n388 , n387 );
or ( n389 , n382 , n388 );
xor ( n390 , n292 , n290 );
xor ( n391 , n390 , n302 );
or ( n392 , n385 , n391 );
nand ( n393 , n389 , n392 );
and ( n394 , n358 , n393 );
and ( n395 , n352 , n357 );
or ( n396 , n394 , n395 );
and ( n397 , n343 , n396 );
not ( n398 , n343 );
not ( n399 , n396 );
and ( n400 , n398 , n399 );
nor ( n401 , n397 , n400 );
not ( n402 , n401 );
xor ( n403 , n352 , n357 );
xor ( n404 , n403 , n393 );
xor ( n405 , n385 , n381 );
xnor ( n406 , n405 , n391 );
not ( n407 , n406 );
not ( n408 , n407 );
nand ( n409 , n7 , n21 );
nor ( n410 , n409 , n130 );
buf ( n411 , n410 );
not ( n412 , n411 );
and ( n413 , n6 , n21 );
and ( n414 , n7 , n20 );
nor ( n415 , n413 , n414 );
nor ( n416 , n410 , n415 );
xor ( n417 , n176 , n416 );
not ( n418 , n379 );
not ( n419 , n376 );
not ( n420 , n419 );
or ( n421 , n418 , n420 );
nand ( n422 , n376 , n360 );
nand ( n423 , n421 , n422 );
xnor ( n424 , n417 , n423 );
nand ( n425 , n5 , n24 );
nand ( n426 , n6 , n23 );
nor ( n427 , n425 , n426 );
not ( n428 , n427 );
nand ( n429 , n425 , n426 );
nand ( n430 , n7 , n22 );
not ( n431 , n430 );
nand ( n432 , n429 , n431 );
nand ( n433 , n428 , n432 );
not ( n434 , n433 );
xor ( n435 , n409 , n363 );
nand ( n436 , n375 , n370 );
xnor ( n437 , n435 , n436 );
not ( n438 , n437 );
or ( n439 , n434 , n438 );
not ( n440 , n409 );
and ( n441 , n436 , n363 );
not ( n442 , n436 );
and ( n443 , n442 , n364 );
nor ( n444 , n441 , n443 );
nand ( n445 , n440 , n444 );
nand ( n446 , n439 , n445 );
nand ( n447 , n424 , n446 );
not ( n448 , n447 );
not ( n449 , n448 );
or ( n450 , n412 , n449 );
or ( n451 , n411 , n448 );
nand ( n452 , n450 , n451 );
not ( n453 , n176 );
buf ( n454 , n423 );
not ( n455 , n454 );
or ( n456 , n453 , n455 );
or ( n457 , n454 , n176 );
nand ( n458 , n456 , n457 );
nand ( n459 , n458 , n416 );
nand ( n460 , n452 , n459 );
not ( n461 , n460 );
or ( n462 , n408 , n461 );
nand ( n463 , n448 , n411 );
nand ( n464 , n462 , n463 );
nand ( n465 , n404 , n464 );
not ( n466 , n465 );
nor ( n467 , n424 , n446 );
not ( n468 , n467 );
nand ( n469 , n468 , n447 );
nand ( n470 , n8 , n20 );
not ( n471 , n470 );
not ( n472 , n471 );
nand ( n473 , n7 , n23 );
nand ( n474 , n6 , n24 );
nor ( n475 , n473 , n474 );
not ( n476 , n475 );
nand ( n477 , n8 , n22 );
not ( n478 , n477 );
nand ( n479 , n473 , n474 );
nand ( n480 , n478 , n479 );
nand ( n481 , n476 , n480 );
not ( n482 , n481 );
nand ( n483 , n8 , n21 );
xor ( n484 , n430 , n483 );
not ( n485 , n427 );
nand ( n486 , n485 , n429 );
xnor ( n487 , n484 , n486 );
not ( n488 , n487 );
or ( n489 , n482 , n488 );
not ( n490 , n483 );
not ( n491 , n486 );
nand ( n492 , n491 , n431 );
not ( n493 , n431 );
nand ( n494 , n493 , n486 );
nand ( n495 , n490 , n492 , n494 );
nand ( n496 , n489 , n495 );
not ( n497 , n496 );
or ( n498 , n472 , n497 );
not ( n499 , n437 );
not ( n500 , n433 );
xnor ( n501 , n499 , n500 );
nand ( n502 , n498 , n501 );
not ( n503 , n496 );
nand ( n504 , n503 , n470 );
nand ( n505 , n502 , n504 );
nor ( n506 , n469 , n505 );
buf ( n507 , n506 );
not ( n508 , n407 );
not ( n509 , n460 );
not ( n510 , n509 );
or ( n511 , n508 , n510 );
nand ( n512 , n460 , n406 );
nand ( n513 , n511 , n512 );
xor ( n514 , n507 , n513 );
not ( n515 , n503 );
not ( n516 , n515 );
xor ( n517 , n471 , n500 );
xnor ( n518 , n517 , n499 );
not ( n519 , n518 );
or ( n520 , n516 , n519 );
or ( n521 , n518 , n515 );
nand ( n522 , n520 , n521 );
buf ( n523 , n487 );
not ( n524 , n481 );
and ( n525 , n523 , n524 );
not ( n526 , n523 );
and ( n527 , n526 , n481 );
nor ( n528 , n525 , n527 );
not ( n529 , n479 );
nor ( n530 , n529 , n475 );
xor ( n531 , n530 , n477 );
not ( n532 , n531 );
not ( n533 , n473 );
not ( n534 , n282 );
nand ( n535 , n533 , n534 );
not ( n536 , n535 );
nand ( n537 , n532 , n536 );
nor ( n538 , n528 , n537 );
nand ( n539 , n522 , n538 );
not ( n540 , n539 );
not ( n541 , n540 );
nand ( n542 , n469 , n505 );
not ( n543 , n542 );
nor ( n544 , n543 , n506 );
not ( n545 , n544 );
or ( n546 , n541 , n545 );
nand ( n547 , n8 , n19 );
not ( n548 , n547 );
nand ( n549 , n542 , n548 );
not ( n550 , n549 );
not ( n551 , n506 );
and ( n552 , n550 , n551 );
nor ( n553 , n539 , n547 );
nor ( n554 , n552 , n553 );
nand ( n555 , n546 , n554 );
and ( n556 , n514 , n555 );
and ( n557 , n507 , n513 );
nor ( n558 , n556 , n557 );
not ( n559 , n558 );
or ( n560 , n466 , n559 );
not ( n561 , n404 );
not ( n562 , n464 );
nand ( n563 , n561 , n562 );
nand ( n564 , n560 , n563 );
not ( n565 , n564 );
not ( n566 , n565 );
or ( n567 , n402 , n566 );
nand ( n568 , n343 , n396 );
nand ( n569 , n567 , n568 );
not ( n570 , n569 );
or ( n571 , n341 , n570 );
not ( n572 , n338 );
nand ( n573 , n572 , n280 );
buf ( n574 , n573 );
nand ( n575 , n571 , n574 );
not ( n576 , n179 );
and ( n577 , n576 , n181 );
not ( n578 , n178 );
nor ( n579 , n577 , n578 );
not ( n580 , n218 );
not ( n581 , n580 );
not ( n582 , n210 );
or ( n583 , n581 , n582 );
not ( n584 , n206 );
nand ( n585 , n584 , n191 );
nand ( n586 , n583 , n585 );
not ( n587 , n586 );
and ( n588 , n5 , n17 );
and ( n589 , n1 , n21 );
nor ( n590 , n588 , n589 );
not ( n591 , n590 );
or ( n592 , n292 , n283 );
nand ( n593 , n591 , n592 );
nand ( n594 , n4 , n18 );
and ( n595 , n593 , n594 );
not ( n596 , n593 );
not ( n597 , n594 );
and ( n598 , n596 , n597 );
or ( n599 , n595 , n598 );
not ( n600 , n599 );
nand ( n601 , n3 , n19 );
not ( n602 , n200 );
xor ( n603 , n601 , n602 );
not ( n604 , n193 );
not ( n605 , n198 );
or ( n606 , n604 , n605 );
not ( n607 , n201 );
nand ( n608 , n606 , n607 );
xnor ( n609 , n603 , n608 );
not ( n610 , n609 );
or ( n611 , n600 , n610 );
or ( n612 , n609 , n599 );
nand ( n613 , n611 , n612 );
not ( n614 , n613 );
not ( n615 , n614 );
or ( n616 , n587 , n615 );
not ( n617 , n586 );
nand ( n618 , n613 , n617 );
nand ( n619 , n616 , n618 );
xor ( n620 , n579 , n619 );
not ( n621 , n189 );
and ( n622 , n621 , n222 );
not ( n623 , n185 );
nor ( n624 , n623 , n170 );
nor ( n625 , n622 , n624 );
xnor ( n626 , n620 , n625 );
not ( n627 , n135 );
nand ( n628 , n278 , n226 );
not ( n629 , n628 );
or ( n630 , n627 , n629 );
nand ( n631 , n279 , n227 );
nand ( n632 , n630 , n631 );
xnor ( n633 , n626 , n632 );
buf ( n634 , n633 );
not ( n635 , n634 );
and ( n636 , n575 , n635 );
not ( n637 , n575 );
and ( n638 , n637 , n634 );
nor ( n639 , n636 , n638 );
not ( n640 , n340 );
and ( n641 , n569 , n640 );
not ( n642 , n569 );
and ( n643 , n642 , n340 );
nor ( n644 , n641 , n643 );
nor ( n645 , n639 , n644 );
xor ( n646 , n555 , n514 );
nand ( n647 , n16 , n32 );
nand ( n648 , n8 , n24 );
nor ( n649 , n647 , n648 );
not ( n650 , n649 );
nand ( n651 , n282 , n647 );
nand ( n652 , n650 , n651 );
not ( n653 , n652 );
not ( n654 , n653 );
buf ( n655 , n654 );
not ( n656 , n655 );
xor ( n657 , n2 , n10 );
not ( n658 , n11 );
not ( n659 , n12 );
nor ( n660 , n7 , n15 );
not ( n661 , n6 );
nor ( n662 , n660 , n661 );
not ( n663 , n662 );
nand ( n664 , n7 , n15 );
nand ( n665 , n8 , n16 );
nand ( n666 , n664 , n665 );
not ( n667 , n666 );
or ( n668 , n663 , n667 );
not ( n669 , n14 );
nand ( n670 , n668 , n669 );
not ( n671 , n660 );
not ( n672 , n671 );
not ( n673 , n666 );
or ( n674 , n672 , n673 );
nand ( n675 , n674 , n661 );
nand ( n676 , n670 , n675 );
nand ( n677 , n5 , n13 );
and ( n678 , n676 , n677 );
nor ( n679 , n5 , n13 );
nor ( n680 , n678 , n679 );
not ( n681 , n680 );
or ( n682 , n659 , n681 );
xor ( n683 , n680 , n12 );
nand ( n684 , n683 , n4 );
nand ( n685 , n682 , n684 );
not ( n686 , n685 );
or ( n687 , n658 , n686 );
not ( n688 , n11 );
not ( n689 , n688 );
not ( n690 , n685 );
or ( n691 , n689 , n690 );
or ( n692 , n685 , n688 );
nand ( n693 , n691 , n692 );
nand ( n694 , n693 , n3 );
nand ( n695 , n687 , n694 );
xnor ( n696 , n657 , n695 );
and ( n697 , n656 , n696 );
not ( n698 , n656 );
xor ( n699 , n18 , n26 );
not ( n700 , n27 );
not ( n701 , n28 );
not ( n702 , n29 );
not ( n703 , n21 );
or ( n704 , n702 , n703 );
nand ( n705 , n24 , n32 );
nor ( n706 , n23 , n31 );
or ( n707 , n705 , n706 );
nand ( n708 , n23 , n31 );
nand ( n709 , n707 , n708 );
not ( n710 , n22 );
not ( n711 , n30 );
nor ( n712 , n710 , n711 );
or ( n713 , n709 , n712 );
or ( n714 , n22 , n30 );
nand ( n715 , n713 , n714 );
nand ( n716 , n704 , n715 );
or ( n717 , n21 , n29 );
nand ( n718 , n716 , n717 );
not ( n719 , n718 );
not ( n720 , n719 );
or ( n721 , n701 , n720 );
xnor ( n722 , n718 , n28 );
nand ( n723 , n722 , n20 );
nand ( n724 , n721 , n723 );
not ( n725 , n724 );
or ( n726 , n700 , n725 );
or ( n727 , n724 , n27 );
nand ( n728 , n727 , n19 );
nand ( n729 , n726 , n728 );
xnor ( n730 , n699 , n729 );
and ( n731 , n698 , n730 );
nor ( n732 , n697 , n731 );
nand ( n733 , n646 , n732 );
not ( n734 , n733 );
xor ( n735 , n19 , n27 );
xnor ( n736 , n735 , n724 );
and ( n737 , n655 , n736 );
not ( n738 , n655 );
xor ( n739 , n3 , n11 );
xnor ( n740 , n739 , n685 );
and ( n741 , n738 , n740 );
nor ( n742 , n737 , n741 );
xor ( n743 , n547 , n540 );
xnor ( n744 , n743 , n544 );
xor ( n745 , n742 , n744 );
or ( n746 , n722 , n20 );
nand ( n747 , n746 , n723 );
and ( n748 , n654 , n747 );
not ( n749 , n654 );
or ( n750 , n4 , n683 );
nand ( n751 , n750 , n684 );
and ( n752 , n749 , n751 );
nor ( n753 , n748 , n752 );
not ( n754 , n753 );
xor ( n755 , n5 , n13 );
xnor ( n756 , n755 , n676 );
and ( n757 , n653 , n756 );
not ( n758 , n653 );
xor ( n759 , n21 , n29 );
and ( n760 , n709 , n711 );
not ( n761 , n709 );
and ( n762 , n761 , n30 );
nor ( n763 , n760 , n762 );
nor ( n764 , n763 , n710 );
and ( n765 , n709 , n30 );
nor ( n766 , n764 , n765 );
xnor ( n767 , n759 , n766 );
and ( n768 , n758 , n767 );
nor ( n769 , n757 , n768 );
not ( n770 , n769 );
not ( n771 , n531 );
not ( n772 , n536 );
and ( n773 , n771 , n772 );
and ( n774 , n531 , n536 );
nor ( n775 , n773 , n774 );
not ( n776 , n775 );
not ( n777 , n652 );
xnor ( n778 , n23 , n31 );
and ( n779 , n778 , n705 );
not ( n780 , n778 );
not ( n781 , n705 );
and ( n782 , n780 , n781 );
nor ( n783 , n779 , n782 );
not ( n784 , n783 );
or ( n785 , n777 , n784 );
xor ( n786 , n15 , n7 );
and ( n787 , n786 , n665 );
not ( n788 , n786 );
not ( n789 , n665 );
and ( n790 , n788 , n789 );
nor ( n791 , n787 , n790 );
or ( n792 , n652 , n791 );
nand ( n793 , n785 , n792 );
nor ( n794 , n282 , n16 );
nand ( n795 , n793 , n794 );
nand ( n796 , n8 , n23 );
nand ( n797 , n7 , n24 );
nand ( n798 , n796 , n797 );
nand ( n799 , n535 , n798 );
and ( n800 , n795 , n799 );
nor ( n801 , n793 , n794 );
nor ( n802 , n800 , n801 );
xor ( n803 , n776 , n802 );
not ( n804 , n652 );
not ( n805 , n6 );
not ( n806 , n789 );
not ( n807 , n671 );
or ( n808 , n806 , n807 );
nand ( n809 , n808 , n664 );
and ( n810 , n809 , n14 );
not ( n811 , n809 );
and ( n812 , n811 , n669 );
nor ( n813 , n810 , n812 );
not ( n814 , n813 );
or ( n815 , n805 , n814 );
or ( n816 , n813 , n6 );
nand ( n817 , n815 , n816 );
and ( n818 , n804 , n817 );
not ( n819 , n804 );
not ( n820 , n763 );
or ( n821 , n820 , n22 );
not ( n822 , n764 );
nand ( n823 , n821 , n822 );
and ( n824 , n819 , n823 );
nor ( n825 , n818 , n824 );
and ( n826 , n803 , n825 );
and ( n827 , n776 , n802 );
nor ( n828 , n826 , n827 );
not ( n829 , n828 );
or ( n830 , n770 , n829 );
or ( n831 , n828 , n769 );
not ( n832 , n538 );
nand ( n833 , n528 , n537 );
nand ( n834 , n832 , n833 );
nand ( n835 , n831 , n834 );
nand ( n836 , n830 , n835 );
not ( n837 , n836 );
not ( n838 , n538 );
not ( n839 , n838 );
not ( n840 , n522 );
not ( n841 , n840 );
or ( n842 , n839 , n841 );
nand ( n843 , n842 , n539 );
not ( n844 , n843 );
not ( n845 , n844 );
or ( n846 , n837 , n845 );
or ( n847 , n844 , n836 );
nand ( n848 , n846 , n847 );
not ( n849 , n848 );
or ( n850 , n754 , n849 );
not ( n851 , n836 );
nand ( n852 , n851 , n844 );
nand ( n853 , n850 , n852 );
and ( n854 , n745 , n853 );
and ( n855 , n742 , n744 );
nor ( n856 , n854 , n855 );
not ( n857 , n856 );
or ( n858 , n734 , n857 );
not ( n859 , n732 );
not ( n860 , n646 );
nand ( n861 , n859 , n860 );
nand ( n862 , n858 , n861 );
not ( n863 , n862 );
not ( n864 , n863 );
nor ( n865 , n564 , n401 );
not ( n866 , n865 );
nand ( n867 , n564 , n401 );
nand ( n868 , n866 , n867 );
xor ( n869 , n9 , n1 );
not ( n870 , n10 );
not ( n871 , n695 );
or ( n872 , n870 , n871 );
not ( n873 , n10 );
not ( n874 , n873 );
not ( n875 , n695 );
or ( n876 , n874 , n875 );
or ( n877 , n695 , n873 );
nand ( n878 , n876 , n877 );
nand ( n879 , n878 , n2 );
nand ( n880 , n872 , n879 );
and ( n881 , n869 , n880 );
and ( n882 , n9 , n1 );
or ( n883 , n881 , n882 );
not ( n884 , n883 );
not ( n885 , n655 );
and ( n886 , n884 , n885 );
not ( n887 , n26 );
not ( n888 , n729 );
or ( n889 , n887 , n888 );
or ( n890 , n729 , n26 );
nand ( n891 , n890 , n18 );
nand ( n892 , n889 , n891 );
or ( n893 , n892 , n25 );
nand ( n894 , n893 , n17 );
and ( n895 , n892 , n25 );
nor ( n896 , n895 , n656 );
and ( n897 , n894 , n896 );
nor ( n898 , n886 , n897 );
nand ( n899 , n868 , n898 );
not ( n900 , n558 );
not ( n901 , n464 );
not ( n902 , n404 );
not ( n903 , n902 );
or ( n904 , n901 , n903 );
nand ( n905 , n404 , n562 );
nand ( n906 , n904 , n905 );
not ( n907 , n906 );
and ( n908 , n900 , n907 );
not ( n909 , n900 );
and ( n910 , n909 , n906 );
nor ( n911 , n908 , n910 );
nand ( n912 , n864 , n899 , n911 );
not ( n913 , n868 );
not ( n914 , n898 );
nand ( n915 , n913 , n914 );
nand ( n916 , n912 , n915 );
not ( n917 , n916 );
not ( n918 , n862 );
not ( n919 , n911 );
nand ( n920 , n918 , n919 );
xor ( n921 , n9 , n1 );
xor ( n922 , n921 , n880 );
or ( n923 , n922 , n655 );
xor ( n924 , n17 , n25 );
xnor ( n925 , n924 , n892 );
nand ( n926 , n925 , n655 );
nand ( n927 , n923 , n926 );
nand ( n928 , n920 , n899 , n927 );
and ( n929 , n645 , n917 , n928 );
not ( n930 , n929 );
and ( n931 , n2 , n19 );
and ( n932 , n3 , n18 );
nor ( n933 , n931 , n932 );
not ( n934 , n933 );
nand ( n935 , n4 , n17 );
not ( n936 , n935 );
and ( n937 , n934 , n936 );
nand ( n938 , n2 , n18 );
nor ( n939 , n601 , n938 );
nor ( n940 , n937 , n939 );
nand ( n941 , n3 , n17 );
xor ( n942 , n940 , n941 );
and ( n943 , n942 , n938 );
and ( n944 , n940 , n941 );
nor ( n945 , n943 , n944 );
nand ( n946 , n2 , n17 );
not ( n947 , n946 );
and ( n948 , n945 , n947 );
not ( n949 , n945 );
and ( n950 , n949 , n946 );
nor ( n951 , n948 , n950 );
not ( n952 , n177 );
and ( n953 , n951 , n952 );
and ( n954 , n945 , n947 );
nor ( n955 , n953 , n954 );
xor ( n956 , n955 , n283 );
not ( n957 , n956 );
nor ( n958 , n939 , n933 );
xor ( n959 , n958 , n935 );
not ( n960 , n959 );
not ( n961 , n602 );
not ( n962 , n601 );
not ( n963 , n608 );
or ( n964 , n962 , n963 );
or ( n965 , n608 , n601 );
nand ( n966 , n964 , n965 );
not ( n967 , n966 );
or ( n968 , n961 , n967 );
not ( n969 , n601 );
nand ( n970 , n969 , n608 );
nand ( n971 , n968 , n970 );
not ( n972 , n971 );
not ( n973 , n972 );
or ( n974 , n960 , n973 );
and ( n975 , n592 , n594 );
nor ( n976 , n975 , n590 );
not ( n977 , n976 );
not ( n978 , n959 );
not ( n979 , n971 );
or ( n980 , n978 , n979 );
or ( n981 , n971 , n959 );
nand ( n982 , n980 , n981 );
nand ( n983 , n977 , n982 );
nand ( n984 , n974 , n983 );
nand ( n985 , n1 , n19 );
xnor ( n986 , n984 , n985 );
xor ( n987 , n940 , n941 );
xor ( n988 , n987 , n938 );
xor ( n989 , n986 , n988 );
nand ( n990 , n1 , n20 );
not ( n991 , n990 );
not ( n992 , n991 );
xor ( n993 , n976 , n959 );
xnor ( n994 , n993 , n971 );
not ( n995 , n994 );
or ( n996 , n992 , n995 );
not ( n997 , n994 );
not ( n998 , n990 );
and ( n999 , n997 , n998 );
and ( n1000 , n994 , n990 );
nor ( n1001 , n999 , n1000 );
not ( n1002 , n1001 );
or ( n1003 , n614 , n617 );
not ( n1004 , n609 );
or ( n1005 , n1004 , n599 );
nand ( n1006 , n1003 , n1005 );
nand ( n1007 , n1002 , n1006 );
nand ( n1008 , n996 , n1007 );
xor ( n1009 , n989 , n1008 );
nand ( n1010 , n573 , n568 );
not ( n1011 , n343 );
nand ( n1012 , n1011 , n399 );
nor ( n1013 , n1010 , n1012 );
not ( n1014 , n281 );
not ( n1015 , n339 );
or ( n1016 , n1014 , n1015 );
nand ( n1017 , n1016 , n633 );
or ( n1018 , n1013 , n1017 );
not ( n1019 , n626 );
nor ( n1020 , n632 , n1019 );
not ( n1021 , n1020 );
nand ( n1022 , n1018 , n1021 );
not ( n1023 , n1010 );
nand ( n1024 , n900 , n906 );
not ( n1025 , n465 );
nor ( n1026 , n1025 , n1020 );
nand ( n1027 , n1023 , n1024 , n1026 );
nand ( n1028 , n1022 , n1027 );
xor ( n1029 , n625 , n619 );
not ( n1030 , n579 );
and ( n1031 , n1029 , n1030 );
and ( n1032 , n625 , n619 );
or ( n1033 , n1031 , n1032 );
not ( n1034 , n1001 );
not ( n1035 , n1006 );
and ( n1036 , n1034 , n1035 );
and ( n1037 , n1001 , n1006 );
nor ( n1038 , n1036 , n1037 );
xor ( n1039 , n1033 , n1038 );
or ( n1040 , n1028 , n1039 );
not ( n1041 , n1038 );
nand ( n1042 , n1041 , n1033 );
nand ( n1043 , n1040 , n1042 );
and ( n1044 , n1009 , n1043 );
and ( n1045 , n989 , n1008 );
or ( n1046 , n1044 , n1045 );
xor ( n1047 , n951 , n952 );
or ( n1048 , n986 , n988 );
or ( n1049 , n984 , n985 );
nand ( n1050 , n1048 , n1049 );
xor ( n1051 , n1047 , n1050 );
and ( n1052 , n1046 , n1051 );
and ( n1053 , n1047 , n1050 );
nor ( n1054 , n1052 , n1053 );
and ( n1055 , n957 , n1054 );
xor ( n1056 , n989 , n1008 );
xor ( n1057 , n1056 , n1043 );
buf ( n1058 , n1028 );
and ( n1059 , n1058 , n1039 );
not ( n1060 , n1058 );
not ( n1061 , n1039 );
and ( n1062 , n1060 , n1061 );
nor ( n1063 , n1059 , n1062 );
nand ( n1064 , n1057 , n1063 );
not ( n1065 , n1064 );
xor ( n1066 , n1046 , n1051 );
nand ( n1067 , n1065 , n1066 );
nor ( n1068 , n1055 , n1067 );
not ( n1069 , n1068 );
or ( n1070 , n930 , n1069 );
not ( n1071 , n955 );
not ( n1072 , n283 );
and ( n1073 , n1071 , n1072 );
not ( n1074 , n1054 );
and ( n1075 , n1074 , n956 );
nor ( n1076 , n1073 , n1075 );
nand ( n1077 , n1070 , n1076 );
nand ( n1078 , n9 , n25 );
and ( n1079 , n11 , n26 );
and ( n1080 , n10 , n27 );
nor ( n1081 , n1079 , n1080 );
not ( n1082 , n1081 );
nand ( n1083 , n12 , n25 );
not ( n1084 , n1083 );
and ( n1085 , n1082 , n1084 );
nand ( n1086 , n11 , n27 );
nand ( n1087 , n10 , n26 );
nor ( n1088 , n1086 , n1087 );
nor ( n1089 , n1085 , n1088 );
nand ( n1090 , n11 , n25 );
xor ( n1091 , n1089 , n1090 );
and ( n1092 , n1091 , n1087 );
and ( n1093 , n1089 , n1090 );
nor ( n1094 , n1092 , n1093 );
not ( n1095 , n1094 );
nand ( n1096 , n10 , n25 );
not ( n1097 , n1096 );
and ( n1098 , n1095 , n1097 );
and ( n1099 , n1094 , n1096 );
nor ( n1100 , n1098 , n1099 );
nand ( n1101 , n9 , n26 );
or ( n1102 , n1100 , n1101 );
not ( n1103 , n1094 );
or ( n1104 , n1103 , n1096 );
nand ( n1105 , n1102 , n1104 );
xnor ( n1106 , n1078 , n1105 );
not ( n1107 , n1106 );
and ( n1108 , n12 , n32 , n11 , n31 );
not ( n1109 , n1108 );
not ( n1110 , n1109 );
not ( n1111 , n1110 );
nand ( n1112 , n10 , n32 );
not ( n1113 , n1112 );
and ( n1114 , n11 , n31 );
not ( n1115 , n1114 );
or ( n1116 , n1113 , n1115 );
and ( n1117 , n11 , n31 );
nand ( n1118 , n10 , n32 );
or ( n1119 , n1117 , n1118 );
nand ( n1120 , n1116 , n1119 );
nand ( n1121 , n12 , n30 );
nand ( n1122 , n1120 , n1121 );
or ( n1123 , n1121 , n1120 );
nand ( n1124 , n13 , n29 );
nand ( n1125 , n1122 , n1123 , n1124 );
not ( n1126 , n1125 );
or ( n1127 , n1111 , n1126 );
not ( n1128 , n1124 );
not ( n1129 , n1121 );
not ( n1130 , n1120 );
or ( n1131 , n1129 , n1130 );
nand ( n1132 , n1131 , n1123 );
nand ( n1133 , n1128 , n1132 );
nand ( n1134 , n1127 , n1133 );
not ( n1135 , n1134 );
nand ( n1136 , n16 , n32 );
nor ( n1137 , n1078 , n1136 );
and ( n1138 , n9 , n32 );
and ( n1139 , n16 , n25 );
nor ( n1140 , n1138 , n1139 );
nor ( n1141 , n1137 , n1140 );
not ( n1142 , n14 );
not ( n1143 , n27 );
or ( n1144 , n1142 , n1143 );
nand ( n1145 , n13 , n28 );
nand ( n1146 , n1144 , n1145 );
not ( n1147 , n1146 );
nand ( n1148 , n13 , n27 );
nand ( n1149 , n14 , n28 );
nor ( n1150 , n1148 , n1149 );
nor ( n1151 , n1147 , n1150 );
nand ( n1152 , n15 , n26 );
not ( n1153 , n1152 );
and ( n1154 , n1151 , n1153 );
not ( n1155 , n1151 );
and ( n1156 , n1155 , n1152 );
or ( n1157 , n1154 , n1156 );
xor ( n1158 , n1141 , n1157 );
and ( n1159 , n11 , n31 );
not ( n1160 , n1159 );
not ( n1161 , n1118 );
not ( n1162 , n1161 );
or ( n1163 , n1160 , n1162 );
not ( n1164 , n1117 );
not ( n1165 , n1164 );
not ( n1166 , n1118 );
or ( n1167 , n1165 , n1166 );
not ( n1168 , n1121 );
nand ( n1169 , n1167 , n1168 );
nand ( n1170 , n1163 , n1169 );
nand ( n1171 , n10 , n30 );
not ( n1172 , n1171 );
not ( n1173 , n1172 );
not ( n1174 , n1117 );
or ( n1175 , n1173 , n1174 );
not ( n1176 , n11 );
not ( n1177 , n30 );
or ( n1178 , n1176 , n1177 );
nand ( n1179 , n10 , n31 );
nand ( n1180 , n1178 , n1179 );
nand ( n1181 , n1175 , n1180 );
nand ( n1182 , n12 , n29 );
and ( n1183 , n1181 , n1182 );
not ( n1184 , n1181 );
not ( n1185 , n1182 );
and ( n1186 , n1184 , n1185 );
nor ( n1187 , n1183 , n1186 );
xor ( n1188 , n1170 , n1187 );
xnor ( n1189 , n1158 , n1188 );
not ( n1190 , n1189 );
or ( n1191 , n1135 , n1190 );
not ( n1192 , n1188 );
not ( n1193 , n1157 );
and ( n1194 , n1192 , n1193 );
and ( n1195 , n1188 , n1157 );
nor ( n1196 , n1194 , n1195 );
not ( n1197 , n1196 );
nand ( n1198 , n1197 , n1141 );
nand ( n1199 , n1191 , n1198 );
not ( n1200 , n1199 );
nand ( n1201 , n1172 , n1159 );
nand ( n1202 , n1185 , n1180 );
and ( n1203 , n1201 , n1202 );
nand ( n1204 , n15 , n25 );
nand ( n1205 , n9 , n31 );
xor ( n1206 , n1204 , n1205 );
and ( n1207 , n1153 , n1146 );
nor ( n1208 , n1207 , n1150 );
xor ( n1209 , n1206 , n1208 );
xor ( n1210 , n1203 , n1209 );
nand ( n1211 , n11 , n29 );
xor ( n1212 , n1211 , n1171 );
nand ( n1213 , n12 , n28 );
xor ( n1214 , n1212 , n1213 );
not ( n1215 , n1214 );
nand ( n1216 , n14 , n26 );
and ( n1217 , n1216 , n1148 );
nor ( n1218 , n1216 , n1148 );
nor ( n1219 , n1217 , n1218 );
not ( n1220 , n1219 );
and ( n1221 , n1215 , n1220 );
and ( n1222 , n1214 , n1219 );
nor ( n1223 , n1221 , n1222 );
xnor ( n1224 , n1210 , n1223 );
not ( n1225 , n1224 );
not ( n1226 , n1157 );
not ( n1227 , n1226 );
not ( n1228 , n1188 );
or ( n1229 , n1227 , n1228 );
nand ( n1230 , n1187 , n1170 );
nand ( n1231 , n1229 , n1230 );
not ( n1232 , n1231 );
not ( n1233 , n1232 );
or ( n1234 , n1225 , n1233 );
or ( n1235 , n1224 , n1232 );
nand ( n1236 , n1234 , n1235 );
not ( n1237 , n1236 );
not ( n1238 , n1237 );
or ( n1239 , n1200 , n1238 );
not ( n1240 , n1199 );
nand ( n1241 , n1240 , n1236 );
nand ( n1242 , n1239 , n1241 );
not ( n1243 , n1242 );
not ( n1244 , n1137 );
nand ( n1245 , n1243 , n1244 );
nand ( n1246 , n1242 , n1137 );
xor ( n1247 , n1141 , n1134 );
xnor ( n1248 , n1247 , n1196 );
not ( n1249 , n1248 );
xor ( n1250 , n1121 , n1108 );
xnor ( n1251 , n1250 , n1120 );
not ( n1252 , n1251 );
not ( n1253 , n1124 );
and ( n1254 , n1252 , n1253 );
and ( n1255 , n1251 , n1124 );
nor ( n1256 , n1254 , n1255 );
not ( n1257 , n1256 );
not ( n1258 , n1257 );
nand ( n1259 , n15 , n27 );
nand ( n1260 , n14 , n28 );
xor ( n1261 , n1259 , n1260 );
nand ( n1262 , n16 , n26 );
xor ( n1263 , n1261 , n1262 );
not ( n1264 , n1263 );
not ( n1265 , n1264 );
or ( n1266 , n1258 , n1265 );
not ( n1267 , n1263 );
not ( n1268 , n1256 );
or ( n1269 , n1267 , n1268 );
not ( n1270 , n11 );
not ( n1271 , n32 );
or ( n1272 , n1270 , n1271 );
nand ( n1273 , n12 , n31 );
nand ( n1274 , n1272 , n1273 );
and ( n1275 , n1274 , n1109 );
not ( n1276 , n1275 );
nand ( n1277 , n13 , n30 );
not ( n1278 , n1277 );
not ( n1279 , n1278 );
not ( n1280 , n31 );
not ( n1281 , n13 );
or ( n1282 , n1280 , n1281 );
nand ( n1283 , n12 , n32 );
nand ( n1284 , n1282 , n1283 );
nand ( n1285 , n14 , n30 );
not ( n1286 , n1285 );
and ( n1287 , n1284 , n1286 );
nand ( n1288 , n13 , n32 );
nor ( n1289 , n1273 , n1288 );
nor ( n1290 , n1287 , n1289 );
not ( n1291 , n1290 );
or ( n1292 , n1279 , n1291 );
and ( n1293 , n1284 , n1286 );
nor ( n1294 , n1293 , n1289 );
or ( n1295 , n1294 , n1278 );
nand ( n1296 , n1292 , n1295 );
not ( n1297 , n1296 );
or ( n1298 , n1276 , n1297 );
not ( n1299 , n1294 );
nand ( n1300 , n1299 , n1278 );
nand ( n1301 , n1298 , n1300 );
buf ( n1302 , n1301 );
nand ( n1303 , n1269 , n1302 );
nand ( n1304 , n1266 , n1303 );
not ( n1305 , n1304 );
xor ( n1306 , n1259 , n1260 );
and ( n1307 , n1306 , n1262 );
and ( n1308 , n1259 , n1260 );
or ( n1309 , n1307 , n1308 );
nand ( n1310 , n1305 , n1309 );
not ( n1311 , n1310 );
or ( n1312 , n1249 , n1311 );
not ( n1313 , n1309 );
nand ( n1314 , n1313 , n1304 );
nand ( n1315 , n1312 , n1314 );
buf ( n1316 , n1315 );
nand ( n1317 , n1245 , n1246 , n1316 );
not ( n1318 , n1317 );
xor ( n1319 , n1137 , n1315 );
xnor ( n1320 , n1319 , n1242 );
not ( n1321 , n1320 );
or ( n1322 , n1318 , n1321 );
not ( n1323 , n1244 );
not ( n1324 , n1242 );
or ( n1325 , n1323 , n1324 );
not ( n1326 , n1199 );
nand ( n1327 , n1326 , n1237 );
nand ( n1328 , n1325 , n1327 );
not ( n1329 , n1328 );
xor ( n1330 , n1204 , n1205 );
and ( n1331 , n1330 , n1208 );
and ( n1332 , n1204 , n1205 );
or ( n1333 , n1331 , n1332 );
not ( n1334 , n1231 );
not ( n1335 , n1224 );
or ( n1336 , n1334 , n1335 );
not ( n1337 , n1209 );
xnor ( n1338 , n1214 , n1219 );
not ( n1339 , n1338 );
nand ( n1340 , n1339 , n1203 );
not ( n1341 , n1203 );
nand ( n1342 , n1341 , n1338 );
nand ( n1343 , n1337 , n1340 , n1342 );
nand ( n1344 , n1336 , n1343 );
not ( n1345 , n1344 );
xor ( n1346 , n1333 , n1345 );
nor ( n1347 , n1277 , n1101 );
and ( n1348 , n9 , n30 );
and ( n1349 , n13 , n26 );
nor ( n1350 , n1348 , n1349 );
nor ( n1351 , n1347 , n1350 );
and ( n1352 , n14 , n25 );
xnor ( n1353 , n1351 , n1352 );
not ( n1354 , n1353 );
not ( n1355 , n1203 );
not ( n1356 , n1223 );
not ( n1357 , n1356 );
or ( n1358 , n1355 , n1357 );
not ( n1359 , n1219 );
nand ( n1360 , n1359 , n1214 );
nand ( n1361 , n1358 , n1360 );
not ( n1362 , n1361 );
not ( n1363 , n1362 );
or ( n1364 , n1354 , n1363 );
not ( n1365 , n1353 );
nand ( n1366 , n1365 , n1361 );
nand ( n1367 , n1364 , n1366 );
xor ( n1368 , n1211 , n1171 );
and ( n1369 , n1368 , n1213 );
and ( n1370 , n1211 , n1171 );
or ( n1371 , n1369 , n1370 );
nand ( n1372 , n12 , n27 );
xor ( n1373 , n1372 , n1218 );
not ( n1374 , n1211 );
nand ( n1375 , n10 , n28 );
not ( n1376 , n1375 );
nand ( n1377 , n1374 , n1376 );
not ( n1378 , n11 );
not ( n1379 , n28 );
or ( n1380 , n1378 , n1379 );
nand ( n1381 , n10 , n29 );
nand ( n1382 , n1380 , n1381 );
nand ( n1383 , n1377 , n1382 );
xor ( n1384 , n1373 , n1383 );
and ( n1385 , n1371 , n1384 );
not ( n1386 , n1371 );
not ( n1387 , n1384 );
and ( n1388 , n1386 , n1387 );
or ( n1389 , n1385 , n1388 );
xor ( n1390 , n1367 , n1389 );
xnor ( n1391 , n1346 , n1390 );
not ( n1392 , n1391 );
not ( n1393 , n1392 );
or ( n1394 , n1329 , n1393 );
not ( n1395 , n1391 );
or ( n1396 , n1395 , n1328 );
nand ( n1397 , n1394 , n1396 );
nand ( n1398 , n1322 , n1397 );
not ( n1399 , n1328 );
nand ( n1400 , n1399 , n1395 );
nand ( n1401 , n1398 , n1400 );
nand ( n1402 , n11 , n32 );
not ( n1403 , n1402 );
not ( n1404 , n1273 );
or ( n1405 , n1403 , n1404 );
nand ( n1406 , n1405 , n1109 );
not ( n1407 , n1260 );
nand ( n1408 , n15 , n29 );
not ( n1409 , n1408 );
and ( n1410 , n1407 , n1409 );
and ( n1411 , n14 , n29 );
and ( n1412 , n15 , n28 );
nor ( n1413 , n1411 , n1412 );
nor ( n1414 , n1410 , n1413 );
xor ( n1415 , n1406 , n1414 );
xnor ( n1416 , n1415 , n1296 );
nand ( n1417 , n15 , n30 );
not ( n1418 , n1417 );
not ( n1419 , n1418 );
nand ( n1420 , n14 , n31 );
nand ( n1421 , n13 , n32 );
nand ( n1422 , n1420 , n1421 );
not ( n1423 , n1422 );
or ( n1424 , n1419 , n1423 );
nor ( n1425 , n1421 , n1420 );
not ( n1426 , n1425 );
nand ( n1427 , n1424 , n1426 );
not ( n1428 , n1427 );
buf ( n1429 , n1285 );
xor ( n1430 , n1408 , n1429 );
not ( n1431 , n1289 );
nand ( n1432 , n1431 , n1284 );
xnor ( n1433 , n1430 , n1432 );
not ( n1434 , n1433 );
or ( n1435 , n1428 , n1434 );
not ( n1436 , n1408 );
xnor ( n1437 , n1286 , n1432 );
nand ( n1438 , n1436 , n1437 );
nand ( n1439 , n1435 , n1438 );
xnor ( n1440 , n1416 , n1439 );
not ( n1441 , n1440 );
and ( n1442 , n16 , n28 );
not ( n1443 , n1442 );
nand ( n1444 , n15 , n31 );
nand ( n1445 , n14 , n32 );
nand ( n1446 , n1444 , n1445 );
nand ( n1447 , n16 , n30 );
not ( n1448 , n1447 );
nand ( n1449 , n1446 , n1448 );
nor ( n1450 , n1444 , n1445 );
not ( n1451 , n1450 );
nand ( n1452 , n1449 , n1451 );
not ( n1453 , n1452 );
and ( n1454 , n16 , n29 );
xor ( n1455 , n1417 , n1454 );
not ( n1456 , n1425 );
nand ( n1457 , n1456 , n1422 );
xor ( n1458 , n1455 , n1457 );
not ( n1459 , n1458 );
or ( n1460 , n1453 , n1459 );
not ( n1461 , n1457 );
nand ( n1462 , n1461 , n1418 );
nand ( n1463 , n1457 , n1417 );
nand ( n1464 , n1462 , n1463 , n1454 );
nand ( n1465 , n1460 , n1464 );
not ( n1466 , n1465 );
or ( n1467 , n1443 , n1466 );
or ( n1468 , n1442 , n1465 );
not ( n1469 , n1433 );
not ( n1470 , n1427 );
and ( n1471 , n1469 , n1470 );
not ( n1472 , n1469 );
and ( n1473 , n1472 , n1427 );
nor ( n1474 , n1471 , n1473 );
nand ( n1475 , n1468 , n1474 );
nand ( n1476 , n1467 , n1475 );
buf ( n1477 , n1476 );
nand ( n1478 , n1441 , n1477 );
not ( n1479 , n1478 );
nor ( n1480 , n1260 , n1408 );
xor ( n1481 , n1263 , n1301 );
xnor ( n1482 , n1481 , n1256 );
xor ( n1483 , n1480 , n1482 );
not ( n1484 , n1439 );
not ( n1485 , n1416 );
or ( n1486 , n1484 , n1485 );
buf ( n1487 , n1296 );
not ( n1488 , n1487 );
nand ( n1489 , n1488 , n1275 );
not ( n1490 , n1489 );
nand ( n1491 , n1487 , n1406 );
not ( n1492 , n1491 );
or ( n1493 , n1490 , n1492 );
nand ( n1494 , n1493 , n1414 );
nand ( n1495 , n1486 , n1494 );
xnor ( n1496 , n1483 , n1495 );
xor ( n1497 , n1479 , n1496 );
not ( n1498 , n1478 );
not ( n1499 , n1477 );
and ( n1500 , n1440 , n1499 );
nand ( n1501 , n16 , n27 );
nor ( n1502 , n1500 , n1501 );
not ( n1503 , n1502 );
or ( n1504 , n1498 , n1503 );
xor ( n1505 , n1501 , n1476 );
xnor ( n1506 , n1505 , n1440 );
buf ( n1507 , n1465 );
not ( n1508 , n1507 );
xor ( n1509 , n1442 , n1470 );
xnor ( n1510 , n1509 , n1469 );
not ( n1511 , n1510 );
or ( n1512 , n1508 , n1511 );
or ( n1513 , n1510 , n1507 );
nand ( n1514 , n1512 , n1513 );
buf ( n1515 , n1458 );
not ( n1516 , n1446 );
not ( n1517 , n1448 );
or ( n1518 , n1516 , n1517 );
nand ( n1519 , n1518 , n1451 );
and ( n1520 , n1515 , n1519 );
not ( n1521 , n1515 );
not ( n1522 , n1452 );
and ( n1523 , n1521 , n1522 );
nor ( n1524 , n1520 , n1523 );
not ( n1525 , n1444 );
not ( n1526 , n1136 );
nand ( n1527 , n1525 , n1526 );
not ( n1528 , n1527 );
not ( n1529 , n1450 );
nand ( n1530 , n1529 , n1446 );
not ( n1531 , n1530 );
not ( n1532 , n1447 );
and ( n1533 , n1531 , n1532 );
and ( n1534 , n1530 , n1447 );
nor ( n1535 , n1533 , n1534 );
and ( n1536 , n1528 , n1535 );
nand ( n1537 , n1524 , n1536 );
not ( n1538 , n1537 );
nand ( n1539 , n1514 , n1538 );
or ( n1540 , n1506 , n1539 );
nand ( n1541 , n1504 , n1540 );
and ( n1542 , n1497 , n1541 );
and ( n1543 , n1479 , n1496 );
or ( n1544 , n1542 , n1543 );
not ( n1545 , n1304 );
xor ( n1546 , n1309 , n1545 );
xnor ( n1547 , n1546 , n1248 );
not ( n1548 , n1547 );
not ( n1549 , n1480 );
not ( n1550 , n1482 );
not ( n1551 , n1495 );
or ( n1552 , n1550 , n1551 );
buf ( n1553 , n1482 );
or ( n1554 , n1553 , n1495 );
nand ( n1555 , n1552 , n1554 );
not ( n1556 , n1555 );
or ( n1557 , n1549 , n1556 );
not ( n1558 , n1553 );
nand ( n1559 , n1558 , n1495 );
nand ( n1560 , n1557 , n1559 );
not ( n1561 , n1560 );
or ( n1562 , n1548 , n1561 );
or ( n1563 , n1560 , n1547 );
nand ( n1564 , n1562 , n1563 );
nand ( n1565 , n1544 , n1564 );
not ( n1566 , n1547 );
nand ( n1567 , n1566 , n1560 );
nand ( n1568 , n1565 , n1317 , n1400 , n1567 );
nand ( n1569 , n1401 , n1568 );
and ( n1570 , n1351 , n1352 );
nor ( n1571 , n1570 , n1347 );
xor ( n1572 , n1086 , n1376 );
not ( n1573 , n1372 );
nand ( n1574 , n1573 , n1382 );
nand ( n1575 , n1377 , n1574 );
xnor ( n1576 , n1572 , n1575 );
and ( n1577 , n9 , n29 );
and ( n1578 , n13 , n25 );
nor ( n1579 , n1577 , n1578 );
not ( n1580 , n1579 );
or ( n1581 , n1124 , n1078 );
nand ( n1582 , n1580 , n1581 );
nand ( n1583 , n12 , n26 );
xor ( n1584 , n1582 , n1583 );
and ( n1585 , n1576 , n1584 );
not ( n1586 , n1576 );
not ( n1587 , n1584 );
and ( n1588 , n1586 , n1587 );
nor ( n1589 , n1585 , n1588 );
not ( n1590 , n1589 );
not ( n1591 , n1371 );
nand ( n1592 , n1591 , n1384 );
or ( n1593 , n1383 , n1372 );
nand ( n1594 , n1383 , n1372 );
nand ( n1595 , n1593 , n1594 , n1218 );
and ( n1596 , n1592 , n1595 );
not ( n1597 , n1596 );
and ( n1598 , n1590 , n1597 );
and ( n1599 , n1589 , n1596 );
nor ( n1600 , n1598 , n1599 );
xor ( n1601 , n1571 , n1600 );
not ( n1602 , n1389 );
not ( n1603 , n1602 );
not ( n1604 , n1367 );
or ( n1605 , n1603 , n1604 );
nand ( n1606 , n1361 , n1353 );
nand ( n1607 , n1605 , n1606 );
xnor ( n1608 , n1601 , n1607 );
not ( n1609 , n1608 );
not ( n1610 , n1333 );
nand ( n1611 , n1390 , n1344 );
not ( n1612 , n1611 );
or ( n1613 , n1610 , n1612 );
not ( n1614 , n1390 );
nand ( n1615 , n1614 , n1345 );
nand ( n1616 , n1613 , n1615 );
not ( n1617 , n1616 );
or ( n1618 , n1609 , n1617 );
or ( n1619 , n1616 , n1608 );
nand ( n1620 , n1618 , n1619 );
not ( n1621 , n1620 );
or ( n1622 , n1569 , n1621 );
nand ( n1623 , n9 , n28 );
not ( n1624 , n1623 );
not ( n1625 , n1624 );
and ( n1626 , n1581 , n1583 );
nor ( n1627 , n1626 , n1579 );
nor ( n1628 , n1088 , n1081 );
xor ( n1629 , n1083 , n1628 );
xor ( n1630 , n1627 , n1629 );
not ( n1631 , n1376 );
not ( n1632 , n1086 );
not ( n1633 , n1575 );
or ( n1634 , n1632 , n1633 );
or ( n1635 , n1575 , n1086 );
nand ( n1636 , n1634 , n1635 );
not ( n1637 , n1636 );
or ( n1638 , n1631 , n1637 );
not ( n1639 , n1086 );
nand ( n1640 , n1639 , n1575 );
nand ( n1641 , n1638 , n1640 );
xnor ( n1642 , n1630 , n1641 );
not ( n1643 , n1642 );
not ( n1644 , n1643 );
or ( n1645 , n1625 , n1644 );
nand ( n1646 , n1642 , n1623 );
nand ( n1647 , n1645 , n1646 );
not ( n1648 , n1589 );
not ( n1649 , n1648 );
not ( n1650 , n1596 );
and ( n1651 , n1649 , n1650 );
and ( n1652 , n1576 , n1584 );
nor ( n1653 , n1651 , n1652 );
xor ( n1654 , n1647 , n1653 );
not ( n1655 , n1654 );
xor ( n1656 , n1600 , n1607 );
and ( n1657 , n1656 , n1571 );
and ( n1658 , n1600 , n1607 );
nor ( n1659 , n1657 , n1658 );
nand ( n1660 , n1655 , n1659 );
not ( n1661 , n1616 );
nand ( n1662 , n1661 , n1608 );
and ( n1663 , n1660 , n1662 );
nand ( n1664 , n1622 , n1663 );
not ( n1665 , n1647 );
or ( n1666 , n1665 , n1653 );
or ( n1667 , n1643 , n1623 );
nand ( n1668 , n1666 , n1667 );
nand ( n1669 , n9 , n27 );
not ( n1670 , n1627 );
not ( n1671 , n1670 );
not ( n1672 , n1629 );
not ( n1673 , n1641 );
or ( n1674 , n1672 , n1673 );
or ( n1675 , n1641 , n1629 );
nand ( n1676 , n1674 , n1675 );
not ( n1677 , n1676 );
or ( n1678 , n1671 , n1677 );
not ( n1679 , n1641 );
nand ( n1680 , n1679 , n1629 );
nand ( n1681 , n1678 , n1680 );
xor ( n1682 , n1669 , n1681 );
xor ( n1683 , n1089 , n1090 );
xor ( n1684 , n1683 , n1087 );
xor ( n1685 , n1682 , n1684 );
xor ( n1686 , n1668 , n1685 );
not ( n1687 , n1654 );
not ( n1688 , n1659 );
or ( n1689 , n1687 , n1688 );
or ( n1690 , n1659 , n1654 );
nand ( n1691 , n1689 , n1690 );
not ( n1692 , n1660 );
nor ( n1693 , n1691 , n1692 );
nor ( n1694 , n1686 , n1693 );
and ( n1695 , n1664 , n1694 );
not ( n1696 , n1668 );
nor ( n1697 , n1696 , n1685 );
nor ( n1698 , n1695 , n1697 );
not ( n1699 , n1698 );
not ( n1700 , n1684 );
not ( n1701 , n1700 );
not ( n1702 , n1682 );
or ( n1703 , n1701 , n1702 );
or ( n1704 , n1681 , n1669 );
nand ( n1705 , n1703 , n1704 );
xor ( n1706 , n1101 , n1100 );
xnor ( n1707 , n1705 , n1706 );
not ( n1708 , n1707 );
and ( n1709 , n1699 , n1708 );
and ( n1710 , n1705 , n1706 );
nor ( n1711 , n1709 , n1710 );
not ( n1712 , n1711 );
not ( n1713 , n1712 );
or ( n1714 , n1107 , n1713 );
not ( n1715 , n1078 );
nand ( n1716 , n1715 , n1105 );
nand ( n1717 , n1714 , n1716 );
and ( n1718 , n1077 , n1717 );
not ( n1719 , n1077 );
not ( n1720 , n1717 );
and ( n1721 , n1719 , n1720 );
nor ( n1722 , n1718 , n1721 );
xnor ( n1723 , n1698 , n1707 );
not ( n1724 , n1723 );
not ( n1725 , n1724 );
not ( n1726 , n868 );
not ( n1727 , n799 );
and ( n1728 , n15 , n32 );
and ( n1729 , n16 , n31 );
nor ( n1730 , n1728 , n1729 );
not ( n1731 , n1730 );
and ( n1732 , n1527 , n1731 );
not ( n1733 , n1732 );
or ( n1734 , n1727 , n1733 );
or ( n1735 , n1732 , n799 );
nand ( n1736 , n1734 , n1735 );
not ( n1737 , n1736 );
buf ( n1738 , n649 );
not ( n1739 , n1738 );
and ( n1740 , n1737 , n1739 );
and ( n1741 , n1736 , n1738 );
nor ( n1742 , n1740 , n1741 );
not ( n1743 , n1742 );
not ( n1744 , n1743 );
buf ( n1745 , n1744 );
nand ( n1746 , n1726 , n1745 );
not ( n1747 , n1746 );
not ( n1748 , n1567 );
not ( n1749 , n1544 );
not ( n1750 , n1749 );
or ( n1751 , n1748 , n1750 );
not ( n1752 , n1560 );
nand ( n1753 , n1752 , n1547 );
nand ( n1754 , n1751 , n1753 );
buf ( n1755 , n1320 );
and ( n1756 , n1754 , n1755 );
not ( n1757 , n1754 );
not ( n1758 , n1755 );
and ( n1759 , n1757 , n1758 );
nor ( n1760 , n1756 , n1759 );
not ( n1761 , n1760 );
or ( n1762 , n1747 , n1761 );
not ( n1763 , n1744 );
not ( n1764 , n744 );
or ( n1765 , n1763 , n1764 );
not ( n1766 , n1506 );
nand ( n1767 , n1766 , n1539 );
not ( n1768 , n1767 );
not ( n1769 , n1539 );
and ( n1770 , n1506 , n1769 );
nor ( n1771 , n1768 , n1770 );
nand ( n1772 , n1765 , n1771 );
or ( n1773 , n1514 , n1538 );
nand ( n1774 , n1773 , n1539 );
not ( n1775 , n1774 );
nor ( n1776 , n1524 , n1536 );
not ( n1777 , n1776 );
nand ( n1778 , n1777 , n1537 );
not ( n1779 , n1778 );
not ( n1780 , n1779 );
xor ( n1781 , n1528 , n1535 );
not ( n1782 , n1781 );
not ( n1783 , n799 );
nand ( n1784 , n1783 , n1738 , n1732 );
nand ( n1785 , n1782 , n1784 );
not ( n1786 , n1785 );
not ( n1787 , n1784 );
not ( n1788 , n1787 );
not ( n1789 , n1781 );
or ( n1790 , n1788 , n1789 );
nand ( n1791 , n1790 , n775 );
not ( n1792 , n1791 );
or ( n1793 , n1786 , n1792 );
nand ( n1794 , n1793 , n1742 );
not ( n1795 , n1794 );
or ( n1796 , n1780 , n1795 );
nand ( n1797 , n1796 , n834 );
not ( n1798 , n1742 );
not ( n1799 , n1791 );
not ( n1800 , n1799 );
or ( n1801 , n1798 , n1800 );
nand ( n1802 , n1801 , n1785 );
nand ( n1803 , n1802 , n1778 );
nand ( n1804 , n1797 , n1742 , n844 , n1803 );
not ( n1805 , n1804 );
or ( n1806 , n1775 , n1805 );
nand ( n1807 , n1778 , n1743 );
nand ( n1808 , n1797 , n1803 , n1807 );
nand ( n1809 , n843 , n1808 , n1742 );
nand ( n1810 , n1806 , n1809 );
not ( n1811 , n744 );
nand ( n1812 , n1810 , n1811 , n1744 );
nand ( n1813 , n1810 , n1771 );
nand ( n1814 , n1772 , n1812 , n1813 );
or ( n1815 , n646 , n1743 );
xor ( n1816 , n1479 , n1496 );
xor ( n1817 , n1816 , n1541 );
nand ( n1818 , n1815 , n1817 );
and ( n1819 , n1814 , n1818 );
and ( n1820 , n646 , n1744 );
nor ( n1821 , n1820 , n1817 );
nor ( n1822 , n1819 , n1821 );
and ( n1823 , n911 , n1745 );
not ( n1824 , n1749 );
not ( n1825 , n1564 );
and ( n1826 , n1824 , n1825 );
buf ( n1827 , n1749 );
and ( n1828 , n1564 , n1827 );
nor ( n1829 , n1826 , n1828 );
nor ( n1830 , n1823 , n1829 );
or ( n1831 , n1822 , n1830 );
nand ( n1832 , n919 , n1745 );
nand ( n1833 , n1832 , n1829 );
nand ( n1834 , n1831 , n1833 );
nand ( n1835 , n1762 , n1834 );
not ( n1836 , n1835 );
not ( n1837 , n1836 );
not ( n1838 , n1837 );
not ( n1839 , n1621 );
nand ( n1840 , n1569 , n1839 );
not ( n1841 , n1840 );
nand ( n1842 , n1401 , n1568 , n1620 );
nand ( n1843 , n1842 , n1662 );
buf ( n1844 , n1691 );
and ( n1845 , n1843 , n1844 );
not ( n1846 , n1843 );
not ( n1847 , n1844 );
and ( n1848 , n1846 , n1847 );
nor ( n1849 , n1845 , n1848 );
nand ( n1850 , n1841 , n1849 );
not ( n1851 , n1663 );
not ( n1852 , n1842 );
or ( n1853 , n1851 , n1852 );
not ( n1854 , n1693 );
nand ( n1855 , n1853 , n1854 );
not ( n1856 , n1686 );
and ( n1857 , n1855 , n1856 );
not ( n1858 , n1855 );
and ( n1859 , n1858 , n1686 );
nor ( n1860 , n1857 , n1859 );
not ( n1861 , n1745 );
not ( n1862 , n868 );
or ( n1863 , n1861 , n1862 );
not ( n1864 , n1760 );
nand ( n1865 , n1863 , n1864 );
not ( n1866 , n1397 );
not ( n1867 , n1866 );
or ( n1868 , n1754 , n1755 );
buf ( n1869 , n1317 );
nand ( n1870 , n1868 , n1869 );
not ( n1871 , n1870 );
or ( n1872 , n1867 , n1871 );
or ( n1873 , n1866 , n1870 );
nand ( n1874 , n1872 , n1873 );
nand ( n1875 , n1865 , n1874 );
nor ( n1876 , n1850 , n1860 , n1875 );
not ( n1877 , n1876 );
or ( n1878 , n1838 , n1877 );
nor ( n1879 , n1836 , n1875 );
not ( n1880 , n1849 );
nor ( n1881 , n1880 , n1860 );
nand ( n1882 , n1398 , n1400 );
nand ( n1883 , n1882 , n1568 );
nor ( n1884 , n1883 , n1839 );
nand ( n1885 , n1879 , n1881 , n1884 );
nand ( n1886 , n1878 , n1885 );
not ( n1887 , n1886 );
or ( n1888 , n1725 , n1887 );
not ( n1889 , n957 );
not ( n1890 , n1074 );
or ( n1891 , n1889 , n1890 );
nand ( n1892 , n1054 , n956 );
nand ( n1893 , n1891 , n1892 );
and ( n1894 , n1711 , n1106 );
not ( n1895 , n1711 );
not ( n1896 , n1106 );
and ( n1897 , n1895 , n1896 );
nor ( n1898 , n1894 , n1897 );
nor ( n1899 , n1893 , n1898 );
nand ( n1900 , n1888 , n1899 );
not ( n1901 , n1893 );
not ( n1902 , n1881 );
nor ( n1903 , n1902 , n1723 );
nand ( n1904 , n1835 , n1865 );
not ( n1905 , n1904 );
not ( n1906 , n1840 );
nor ( n1907 , n1906 , n1884 );
not ( n1908 , n1874 );
nor ( n1909 , n1907 , n1908 );
nand ( n1910 , n1905 , n1909 );
not ( n1911 , n1910 );
nand ( n1912 , n1901 , n1903 , n1911 , n1898 );
nand ( n1913 , n1900 , n1912 );
not ( n1914 , n1064 );
nand ( n1915 , n1914 , n929 );
not ( n1916 , n1915 );
and ( n1917 , n928 , n912 );
not ( n1918 , n915 );
not ( n1919 , n1063 );
nor ( n1920 , n1918 , n1919 );
and ( n1921 , n1917 , n645 , n1920 );
nor ( n1922 , n1921 , n1057 );
nor ( n1923 , n1916 , n1922 );
not ( n1924 , n1860 );
and ( n1925 , n1923 , n1924 );
not ( n1926 , n1923 );
and ( n1927 , n1926 , n1860 );
nor ( n1928 , n1925 , n1927 );
not ( n1929 , n644 );
not ( n1930 , n928 );
nor ( n1931 , n1930 , n916 );
nand ( n1932 , n1929 , n1931 );
not ( n1933 , n1932 );
not ( n1934 , n639 );
or ( n1935 , n1933 , n1934 );
not ( n1936 , n929 );
nand ( n1937 , n1935 , n1936 );
and ( n1938 , n1937 , n1907 );
not ( n1939 , n1937 );
not ( n1940 , n1907 );
and ( n1941 , n1939 , n1940 );
nor ( n1942 , n1938 , n1941 );
not ( n1943 , n1898 );
nand ( n1944 , n1886 , n1943 , n1724 );
and ( n1945 , n1944 , n1720 );
not ( n1946 , n1076 );
nor ( n1947 , n1945 , n1946 );
xor ( n1948 , n1886 , n1723 );
buf ( n1949 , n1066 );
nor ( n1950 , n1948 , n1949 );
and ( n1951 , n1066 , n1724 );
not ( n1952 , n1066 );
and ( n1953 , n1952 , n1723 );
nor ( n1954 , n1951 , n1953 );
not ( n1955 , n1954 );
not ( n1956 , n1915 );
or ( n1957 , n1955 , n1956 );
or ( n1958 , n1915 , n1954 );
nand ( n1959 , n1957 , n1958 );
buf ( n1960 , n1849 );
not ( n1961 , n1960 );
not ( n1962 , n1961 );
and ( n1963 , n1911 , n1962 );
nor ( n1964 , n1963 , n1924 );
nor ( n1965 , n1964 , n1886 , n1057 );
and ( n1966 , n1961 , n1911 );
not ( n1967 , n1961 );
and ( n1968 , n1967 , n1910 );
nor ( n1969 , n1966 , n1968 );
nor ( n1970 , n1969 , n1063 );
nand ( n1971 , n1916 , n1949 );
not ( n1972 , n1971 );
and ( n1973 , n1960 , n1919 );
not ( n1974 , n1960 );
and ( n1975 , n1974 , n1063 );
nor ( n1976 , n1973 , n1975 );
and ( n1977 , n1936 , n1976 );
not ( n1978 , n1936 );
not ( n1979 , n1976 );
and ( n1980 , n1978 , n1979 );
nor ( n1981 , n1977 , n1980 );
or ( n1982 , n1940 , n1879 );
nand ( n1983 , n1982 , n639 );
nor ( n1984 , n1983 , n1911 );
and ( n1985 , n1904 , n1874 );
not ( n1986 , n1904 );
and ( n1987 , n1986 , n1908 );
nor ( n1988 , n1985 , n1987 );
not ( n1989 , n644 );
nor ( n1990 , n1988 , n1989 );
not ( n1991 , n1745 );
not ( n1992 , n1829 );
nand ( n1993 , n1991 , n1992 );
and ( n1994 , n1905 , n1993 );
not ( n1995 , n1834 );
or ( n1996 , n1995 , n1760 );
nand ( n1997 , n1996 , n913 );
nor ( n1998 , n1994 , n1997 );
xnor ( n1999 , n1760 , n914 );
xor ( n2000 , n913 , n1999 );
not ( n2001 , n927 );
xor ( n2002 , n919 , n863 );
nand ( n2003 , n2001 , n2002 );
nand ( n2004 , n2003 , n920 );
xnor ( n2005 , n2000 , n2004 );
and ( n2006 , n644 , n1874 );
not ( n2007 , n644 );
and ( n2008 , n2007 , n1908 );
nor ( n2009 , n2006 , n2008 );
not ( n2010 , n2009 );
and ( n2011 , n1931 , n2010 );
not ( n2012 , n1931 );
and ( n2013 , n2012 , n2009 );
nor ( n2014 , n2011 , n2013 );
not ( n2015 , n2002 );
and ( n2016 , n927 , n1829 );
not ( n2017 , n927 );
and ( n2018 , n2017 , n1992 );
nor ( n2019 , n2016 , n2018 );
not ( n2020 , n2019 );
and ( n2021 , n2015 , n2020 );
not ( n2022 , n2015 );
and ( n2023 , n2022 , n2019 );
nor ( n2024 , n2021 , n2023 );
nand ( n2025 , n1817 , n1991 );
and ( n2026 , n1995 , n2025 );
or ( n2027 , n1992 , n1822 );
nand ( n2028 , n2027 , n911 );
nor ( n2029 , n2026 , n2028 );
and ( n2030 , n856 , n646 );
not ( n2031 , n856 );
and ( n2032 , n2031 , n860 );
nor ( n2033 , n2030 , n2032 );
not ( n2034 , n1817 );
and ( n2035 , n732 , n2034 );
not ( n2036 , n732 );
and ( n2037 , n2036 , n1817 );
nor ( n2038 , n2035 , n2037 );
and ( n2039 , n2033 , n2038 );
not ( n2040 , n2033 );
not ( n2041 , n2038 );
and ( n2042 , n2040 , n2041 );
nor ( n2043 , n2039 , n2042 );
not ( n2044 , n1771 );
nand ( n2045 , n2044 , n1991 );
and ( n2046 , n2045 , n1822 );
not ( n2047 , n2034 );
not ( n2048 , n1814 );
or ( n2049 , n2047 , n2048 );
nand ( n2050 , n2049 , n860 );
nor ( n2051 , n2046 , n2050 );
not ( n2052 , n1771 );
not ( n2053 , n853 );
or ( n2054 , n2052 , n2053 );
or ( n2055 , n1771 , n853 );
nand ( n2056 , n2054 , n2055 );
not ( n2057 , n2056 );
not ( n2058 , n745 );
not ( n2059 , n2058 );
or ( n2060 , n2057 , n2059 );
or ( n2061 , n2058 , n2056 );
nand ( n2062 , n2060 , n2061 );
not ( n2063 , n1774 );
not ( n2064 , n1745 );
and ( n2065 , n2063 , n2064 );
nor ( n2066 , n2065 , n1814 );
not ( n2067 , n1813 );
nor ( n2068 , n2066 , n2067 , n744 );
not ( n2069 , n1810 );
nand ( n2070 , n1779 , n1743 );
and ( n2071 , n2069 , n2070 );
and ( n2072 , n1808 , n1774 );
nor ( n2073 , n2071 , n2072 , n844 );
xor ( n2074 , n1774 , n753 );
not ( n2075 , n2074 );
not ( n2076 , n848 );
or ( n2077 , n2075 , n2076 );
or ( n2078 , n848 , n2074 );
nand ( n2079 , n2077 , n2078 );
and ( n2080 , n1808 , n1803 );
nor ( n2081 , n2070 , n1802 );
nor ( n2082 , n2080 , n2081 );
not ( n2083 , n834 );
nor ( n2084 , n2082 , n2083 );
and ( n2085 , n828 , n834 );
not ( n2086 , n828 );
and ( n2087 , n2086 , n2083 );
nor ( n2088 , n2085 , n2087 );
not ( n2089 , n2088 );
xor ( n2090 , n1779 , n769 );
not ( n2091 , n2090 );
or ( n2092 , n2089 , n2091 );
or ( n2093 , n2090 , n2088 );
nand ( n2094 , n2092 , n2093 );
and ( n2095 , n1742 , n1781 );
not ( n2096 , n1738 );
nand ( n2097 , n2096 , n1736 );
and ( n2098 , n2097 , n1732 );
nor ( n2099 , n2095 , n2098 );
nor ( n2100 , n2099 , n1791 );
not ( n2101 , n1782 );
not ( n2102 , n825 );
or ( n2103 , n2101 , n2102 );
or ( n2104 , n1782 , n825 );
nand ( n2105 , n2103 , n2104 );
not ( n2106 , n801 );
nand ( n2107 , n2106 , n795 );
not ( n2108 , n2107 );
not ( n2109 , n1736 );
or ( n2110 , n2108 , n2109 );
or ( n2111 , n1736 , n2107 );
nand ( n2112 , n2110 , n2111 );
or ( n2113 , n24 , n32 );
nand ( n2114 , n2113 , n665 );
or ( n2115 , n653 , n2114 , n781 );
not ( n2116 , n2114 );
or ( n2117 , n654 , n2116 );
nand ( n2118 , n2115 , n2117 );
buf ( n2119 , n1136 );
and ( n2120 , n1730 , n2119 );
nor ( n2121 , n2120 , n1783 );
xor ( n2122 , n2105 , n803 );
xor ( n2123 , n1893 , n1898 );
and ( n2124 , n2123 , n1971 );
not ( n2125 , n2123 );
and ( n2126 , n2125 , n1972 );
nor ( n2127 , n2124 , n2126 );
not ( n2128 , n1736 );
nor ( n2129 , n2128 , n534 , n2119 );
endmodule
