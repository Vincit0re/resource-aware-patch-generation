module top (out_0, out_1, out_2, out_3, out_4, out_5, out_6, out_7, out_8, out_9, out_10, out_11, out_12, out_13, out_14, in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14);
	input in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14;
	output out_0, out_1, out_2, out_3, out_4, out_5, out_6, out_7, out_8, out_9, out_10, out_11, out_12, out_13, out_14;
	wire gm_n100, gm_n1000, gm_n1001, gm_n1002, gm_n1003, gm_n1004, gm_n1005, gm_n1006, gm_n1007, gm_n1008, gm_n1009, gm_n101, gm_n1010, gm_n1011, gm_n1012, gm_n1013, gm_n1014, gm_n1015, gm_n1016, gm_n1017, gm_n1018, gm_n1019, gm_n102, gm_n1020, gm_n1021, gm_n1022, gm_n1023, gm_n1024, gm_n1025, gm_n1026, gm_n1027, gm_n1028, gm_n1029, gm_n103, gm_n1031, gm_n1032, gm_n1033, gm_n1034, gm_n1035, gm_n1036, gm_n1037, gm_n1038, gm_n1039, gm_n104, gm_n1040, gm_n1041, gm_n1042, gm_n1043, gm_n1044, gm_n1045, gm_n1046, gm_n1047, gm_n1048, gm_n1049, gm_n105, gm_n1050, gm_n1051, gm_n1052, gm_n1053, gm_n1054, gm_n1055, gm_n1056, gm_n1057, gm_n1058, gm_n1059, gm_n106, gm_n1060, gm_n1061, gm_n1062, gm_n1063, gm_n1064, gm_n1065, gm_n1066, gm_n1067, gm_n1068, gm_n1069, gm_n107, gm_n1070, gm_n1071, gm_n1072, gm_n1073, gm_n1074, gm_n1075, gm_n1076, gm_n1077, gm_n1078, gm_n1079, gm_n108, gm_n1080, gm_n1081, gm_n1082, gm_n1083, gm_n1084, gm_n1085, gm_n1086, gm_n1087, gm_n1088, gm_n1089, gm_n109, gm_n1090, gm_n1091, gm_n1092, gm_n1093, gm_n1094, gm_n1095, gm_n1096, gm_n1097, gm_n1098, gm_n1099, gm_n110, gm_n1100, gm_n1101, gm_n1102, gm_n1103, gm_n1104, gm_n1105, gm_n1106, gm_n1107, gm_n1108, gm_n1109, gm_n111, gm_n1110, gm_n1111, gm_n1112, gm_n1113, gm_n1114, gm_n1115, gm_n1116, gm_n1117, gm_n1118, gm_n1119, gm_n112, gm_n1120, gm_n1121, gm_n1122, gm_n1123, gm_n1124, gm_n1125, gm_n1126, gm_n1127, gm_n1128, gm_n1129, gm_n113, gm_n1130, gm_n1131, gm_n1132, gm_n1133, gm_n1134, gm_n1135, gm_n1136, gm_n1137, gm_n1138, gm_n1139, gm_n114, gm_n1140, gm_n1141, gm_n1142, gm_n1143, gm_n1144, gm_n1145, gm_n1146, gm_n1147, gm_n1148, gm_n1149, gm_n115, gm_n1150, gm_n1151, gm_n1152, gm_n1153, gm_n1154, gm_n1155, gm_n1156, gm_n1157, gm_n1158, gm_n1159, gm_n116, gm_n1160, gm_n1161, gm_n1162, gm_n1163, gm_n1164, gm_n1165, gm_n1166, gm_n1167, gm_n1168, gm_n1169, gm_n117, gm_n1171, gm_n1172, gm_n1173, gm_n1174, gm_n1175, gm_n1176, gm_n1177, gm_n1178, gm_n1179, gm_n118, gm_n1180, gm_n1181, gm_n1182, gm_n1183, gm_n1184, gm_n1185, gm_n1186, gm_n1187, gm_n1188, gm_n1189, gm_n119, gm_n1190, gm_n1191, gm_n1192, gm_n1193, gm_n1194, gm_n1195, gm_n1196, gm_n1197, gm_n1198, gm_n1199, gm_n120, gm_n1200, gm_n1201, gm_n1202, gm_n1203, gm_n1204, gm_n1205, gm_n1206, gm_n1207, gm_n1208, gm_n1209, gm_n121, gm_n1210, gm_n1211, gm_n1212, gm_n1213, gm_n1214, gm_n1215, gm_n1216, gm_n1217, gm_n1218, gm_n1219, gm_n122, gm_n1220, gm_n1221, gm_n1222, gm_n1223, gm_n1224, gm_n1225, gm_n1226, gm_n1227, gm_n1228, gm_n1229, gm_n123, gm_n1230, gm_n1231, gm_n1232, gm_n1233, gm_n1234, gm_n1235, gm_n1236, gm_n1237, gm_n1238, gm_n1239, gm_n124, gm_n1240, gm_n1241, gm_n1242, gm_n1243, gm_n1244, gm_n1245, gm_n1246, gm_n1247, gm_n1248, gm_n1249, gm_n125, gm_n1250, gm_n1251, gm_n1252, gm_n1253, gm_n1254, gm_n1255, gm_n1256, gm_n1257, gm_n1258, gm_n1259, gm_n126, gm_n1260, gm_n1261, gm_n1262, gm_n1263, gm_n1264, gm_n1265, gm_n1266, gm_n1267, gm_n1268, gm_n1269, gm_n127, gm_n1270, gm_n1271, gm_n1272, gm_n1273, gm_n1274, gm_n1275, gm_n1276, gm_n1277, gm_n1278, gm_n1279, gm_n128, gm_n1280, gm_n1281, gm_n1282, gm_n1283, gm_n1284, gm_n1285, gm_n1286, gm_n1287, gm_n1288, gm_n1289, gm_n129, gm_n1290, gm_n1291, gm_n1292, gm_n1293, gm_n1294, gm_n1295, gm_n1296, gm_n1297, gm_n1298, gm_n1299, gm_n130, gm_n1300, gm_n1301, gm_n1302, gm_n1303, gm_n1304, gm_n1305, gm_n1306, gm_n1307, gm_n1308, gm_n1309, gm_n131, gm_n1310, gm_n1311, gm_n1312, gm_n1313, gm_n1314, gm_n1315, gm_n1316, gm_n1317, gm_n1318, gm_n1319, gm_n132, gm_n1320, gm_n1321, gm_n1322, gm_n1323, gm_n1324, gm_n1325, gm_n1326, gm_n1327, gm_n1328, gm_n133, gm_n1330, gm_n1331, gm_n1332, gm_n1333, gm_n1334, gm_n1335, gm_n1336, gm_n1337, gm_n1338, gm_n1339, gm_n134, gm_n1340, gm_n1341, gm_n1342, gm_n1343, gm_n1344, gm_n1345, gm_n1346, gm_n1347, gm_n1348, gm_n1349, gm_n135, gm_n1350, gm_n1351, gm_n1352, gm_n1353, gm_n1354, gm_n1355, gm_n1356, gm_n1357, gm_n1358, gm_n1359, gm_n136, gm_n1360, gm_n1361, gm_n1362, gm_n1363, gm_n1364, gm_n1365, gm_n1366, gm_n1367, gm_n1368, gm_n1369, gm_n137, gm_n1370, gm_n1371, gm_n1372, gm_n1373, gm_n1374, gm_n1375, gm_n1376, gm_n1377, gm_n1378, gm_n1379, gm_n138, gm_n1380, gm_n1381, gm_n1382, gm_n1383, gm_n1384, gm_n1385, gm_n1386, gm_n1387, gm_n1388, gm_n1389, gm_n139, gm_n1390, gm_n1391, gm_n1392, gm_n1393, gm_n1394, gm_n1395, gm_n1396, gm_n1397, gm_n1398, gm_n1399, gm_n140, gm_n1400, gm_n1401, gm_n1402, gm_n1403, gm_n1404, gm_n1405, gm_n1406, gm_n1407, gm_n1408, gm_n1409, gm_n141, gm_n1410, gm_n1411, gm_n1412, gm_n1413, gm_n1414, gm_n1415, gm_n1416, gm_n1417, gm_n1418, gm_n1419, gm_n142, gm_n1420, gm_n1421, gm_n1422, gm_n1423, gm_n1424, gm_n1425, gm_n1426, gm_n1427, gm_n1428, gm_n1429, gm_n143, gm_n1431, gm_n1432, gm_n1433, gm_n1434, gm_n1435, gm_n1436, gm_n1437, gm_n1438, gm_n1439, gm_n144, gm_n1440, gm_n1441, gm_n1442, gm_n1443, gm_n1444, gm_n1445, gm_n1446, gm_n1447, gm_n1448, gm_n1449, gm_n145, gm_n1450, gm_n1451, gm_n1452, gm_n1453, gm_n1454, gm_n1455, gm_n1456, gm_n1457, gm_n1458, gm_n1459, gm_n146, gm_n1460, gm_n1461, gm_n1462, gm_n1463, gm_n1464, gm_n1465, gm_n1466, gm_n1467, gm_n1468, gm_n1469, gm_n147, gm_n1470, gm_n1471, gm_n1472, gm_n1473, gm_n1474, gm_n1475, gm_n1476, gm_n1477, gm_n1478, gm_n1479, gm_n148, gm_n1480, gm_n1481, gm_n1482, gm_n1483, gm_n1484, gm_n1485, gm_n1486, gm_n1487, gm_n1488, gm_n1489, gm_n149, gm_n1490, gm_n1491, gm_n1492, gm_n1493, gm_n1494, gm_n1495, gm_n1496, gm_n1497, gm_n1498, gm_n1499, gm_n150, gm_n1500, gm_n1501, gm_n1502, gm_n1503, gm_n1504, gm_n1505, gm_n1506, gm_n1507, gm_n1508, gm_n1509, gm_n151, gm_n1510, gm_n1511, gm_n1512, gm_n1513, gm_n1514, gm_n1515, gm_n1516, gm_n1517, gm_n1518, gm_n1519, gm_n152, gm_n1520, gm_n1521, gm_n1522, gm_n1523, gm_n1524, gm_n1525, gm_n1526, gm_n1527, gm_n1528, gm_n1529, gm_n153, gm_n1530, gm_n1531, gm_n1532, gm_n1533, gm_n1534, gm_n1535, gm_n1536, gm_n1537, gm_n1538, gm_n1539, gm_n154, gm_n1540, gm_n1541, gm_n1542, gm_n1543, gm_n1544, gm_n1545, gm_n1546, gm_n1547, gm_n1548, gm_n1549, gm_n155, gm_n1550, gm_n1551, gm_n1552, gm_n1553, gm_n1554, gm_n1555, gm_n1556, gm_n1557, gm_n1558, gm_n1559, gm_n156, gm_n1560, gm_n1561, gm_n1562, gm_n1563, gm_n1564, gm_n1565, gm_n1566, gm_n1567, gm_n1568, gm_n1569, gm_n157, gm_n1570, gm_n1571, gm_n1572, gm_n1573, gm_n1574, gm_n1575, gm_n1576, gm_n1577, gm_n1578, gm_n1579, gm_n158, gm_n1580, gm_n1581, gm_n1582, gm_n1583, gm_n1584, gm_n1585, gm_n1586, gm_n1587, gm_n1589, gm_n159, gm_n1590, gm_n1591, gm_n1592, gm_n1593, gm_n1594, gm_n1595, gm_n1596, gm_n1597, gm_n1598, gm_n1599, gm_n160, gm_n1600, gm_n1601, gm_n1602, gm_n1603, gm_n1604, gm_n1605, gm_n1606, gm_n1607, gm_n1608, gm_n1609, gm_n161, gm_n1610, gm_n1611, gm_n1612, gm_n1613, gm_n1614, gm_n1615, gm_n1616, gm_n1617, gm_n1618, gm_n1619, gm_n162, gm_n1620, gm_n1621, gm_n1622, gm_n1623, gm_n1624, gm_n1625, gm_n1626, gm_n1627, gm_n1628, gm_n1629, gm_n163, gm_n1630, gm_n1631, gm_n1632, gm_n1633, gm_n1634, gm_n1635, gm_n1636, gm_n1637, gm_n1638, gm_n1639, gm_n164, gm_n1640, gm_n1641, gm_n1642, gm_n1643, gm_n1644, gm_n1645, gm_n1646, gm_n1647, gm_n1648, gm_n1649, gm_n165, gm_n1650, gm_n1651, gm_n1652, gm_n1653, gm_n1654, gm_n1655, gm_n1656, gm_n1657, gm_n1658, gm_n1659, gm_n166, gm_n1660, gm_n1661, gm_n1662, gm_n1663, gm_n1664, gm_n1665, gm_n1666, gm_n1667, gm_n1668, gm_n1669, gm_n167, gm_n1670, gm_n1671, gm_n1672, gm_n1673, gm_n1674, gm_n1675, gm_n1676, gm_n1677, gm_n1678, gm_n1679, gm_n168, gm_n1680, gm_n1681, gm_n1682, gm_n1683, gm_n1684, gm_n1685, gm_n1686, gm_n1687, gm_n1688, gm_n1689, gm_n169, gm_n1690, gm_n1691, gm_n1692, gm_n1693, gm_n1694, gm_n1695, gm_n1696, gm_n1697, gm_n1698, gm_n1699, gm_n170, gm_n1700, gm_n1701, gm_n1702, gm_n1703, gm_n1704, gm_n1705, gm_n1706, gm_n1707, gm_n1708, gm_n1709, gm_n171, gm_n1710, gm_n1711, gm_n1712, gm_n1713, gm_n1714, gm_n1715, gm_n1716, gm_n1717, gm_n1718, gm_n1719, gm_n172, gm_n1720, gm_n1721, gm_n1722, gm_n1723, gm_n1724, gm_n1725, gm_n1726, gm_n1727, gm_n1728, gm_n1729, gm_n173, gm_n1730, gm_n1731, gm_n1732, gm_n1733, gm_n1734, gm_n1735, gm_n1736, gm_n1737, gm_n1739, gm_n174, gm_n1740, gm_n1741, gm_n1742, gm_n1743, gm_n1744, gm_n1745, gm_n1746, gm_n1747, gm_n1748, gm_n1749, gm_n175, gm_n1750, gm_n1751, gm_n1752, gm_n1753, gm_n1754, gm_n1755, gm_n1756, gm_n1757, gm_n1758, gm_n1759, gm_n176, gm_n1760, gm_n1761, gm_n1762, gm_n1763, gm_n1764, gm_n1765, gm_n1766, gm_n1767, gm_n1768, gm_n1769, gm_n177, gm_n1770, gm_n1771, gm_n1772, gm_n1773, gm_n1774, gm_n1775, gm_n1776, gm_n1777, gm_n1778, gm_n1779, gm_n178, gm_n1780, gm_n1781, gm_n1782, gm_n1783, gm_n1784, gm_n1785, gm_n1787, gm_n1788, gm_n1789, gm_n179, gm_n1790, gm_n1791, gm_n1792, gm_n1793, gm_n1794, gm_n1795, gm_n1796, gm_n1797, gm_n1798, gm_n1799, gm_n180, gm_n1800, gm_n1801, gm_n1802, gm_n1803, gm_n1804, gm_n1805, gm_n1806, gm_n1807, gm_n1808, gm_n1809, gm_n181, gm_n1810, gm_n1811, gm_n1812, gm_n1813, gm_n1814, gm_n1815, gm_n1816, gm_n1817, gm_n1818, gm_n1819, gm_n182, gm_n1820, gm_n1821, gm_n1822, gm_n1823, gm_n1824, gm_n1825, gm_n1826, gm_n1827, gm_n1828, gm_n1829, gm_n183, gm_n1830, gm_n1831, gm_n1832, gm_n1833, gm_n1834, gm_n1835, gm_n1836, gm_n1837, gm_n1838, gm_n1839, gm_n184, gm_n1840, gm_n1841, gm_n1842, gm_n1843, gm_n1844, gm_n1845, gm_n1846, gm_n1847, gm_n1848, gm_n1849, gm_n185, gm_n1850, gm_n1851, gm_n1852, gm_n1853, gm_n1854, gm_n1855, gm_n1856, gm_n1857, gm_n1858, gm_n1859, gm_n186, gm_n1860, gm_n1861, gm_n1862, gm_n1863, gm_n1864, gm_n1865, gm_n1866, gm_n1867, gm_n1868, gm_n1869, gm_n187, gm_n1870, gm_n1871, gm_n1872, gm_n1873, gm_n1874, gm_n1875, gm_n1876, gm_n1877, gm_n1878, gm_n1879, gm_n188, gm_n1880, gm_n1881, gm_n1882, gm_n1883, gm_n1884, gm_n1885, gm_n1886, gm_n1887, gm_n1888, gm_n1889, gm_n189, gm_n1890, gm_n1891, gm_n1892, gm_n1893, gm_n1894, gm_n1895, gm_n1896, gm_n1897, gm_n1898, gm_n1899, gm_n190, gm_n1900, gm_n1901, gm_n1902, gm_n1903, gm_n1904, gm_n1905, gm_n1906, gm_n1907, gm_n1908, gm_n1909, gm_n191, gm_n1910, gm_n1911, gm_n1912, gm_n1913, gm_n1914, gm_n1915, gm_n1916, gm_n1917, gm_n1918, gm_n1919, gm_n192, gm_n1920, gm_n1921, gm_n1922, gm_n1923, gm_n1924, gm_n1925, gm_n1926, gm_n1927, gm_n1928, gm_n1929, gm_n193, gm_n1930, gm_n1931, gm_n1932, gm_n1933, gm_n1935, gm_n1936, gm_n1937, gm_n1938, gm_n1939, gm_n194, gm_n1940, gm_n1941, gm_n1942, gm_n1943, gm_n1944, gm_n1945, gm_n1946, gm_n1947, gm_n1948, gm_n1949, gm_n195, gm_n1950, gm_n1951, gm_n1952, gm_n1953, gm_n1954, gm_n1955, gm_n1956, gm_n1957, gm_n1958, gm_n1959, gm_n196, gm_n1960, gm_n1961, gm_n1962, gm_n1963, gm_n1964, gm_n1965, gm_n1966, gm_n1967, gm_n1968, gm_n1969, gm_n197, gm_n1970, gm_n1971, gm_n1972, gm_n1973, gm_n1974, gm_n1975, gm_n1976, gm_n1977, gm_n1978, gm_n1979, gm_n198, gm_n1980, gm_n1981, gm_n1982, gm_n1983, gm_n1984, gm_n1985, gm_n1986, gm_n1987, gm_n1988, gm_n1989, gm_n199, gm_n1990, gm_n1991, gm_n1992, gm_n1993, gm_n1994, gm_n1995, gm_n1996, gm_n1997, gm_n1998, gm_n1999, gm_n200, gm_n2000, gm_n2001, gm_n2002, gm_n2003, gm_n2004, gm_n2005, gm_n2006, gm_n2007, gm_n2008, gm_n2009, gm_n201, gm_n2010, gm_n2011, gm_n2012, gm_n2013, gm_n2014, gm_n2015, gm_n2016, gm_n2017, gm_n2018, gm_n2019, gm_n202, gm_n2020, gm_n2021, gm_n2022, gm_n2023, gm_n2024, gm_n2025, gm_n2026, gm_n2027, gm_n2028, gm_n2029, gm_n203, gm_n2030, gm_n2031, gm_n2032, gm_n2033, gm_n2034, gm_n2035, gm_n2036, gm_n2037, gm_n2038, gm_n2039, gm_n204, gm_n2040, gm_n2041, gm_n2042, gm_n2043, gm_n2044, gm_n2045, gm_n2046, gm_n2047, gm_n2048, gm_n2049, gm_n205, gm_n2050, gm_n2051, gm_n2052, gm_n2053, gm_n2054, gm_n2055, gm_n2056, gm_n2057, gm_n2058, gm_n2059, gm_n206, gm_n2060, gm_n2061, gm_n2062, gm_n2063, gm_n2064, gm_n2065, gm_n2066, gm_n2067, gm_n2068, gm_n2069, gm_n207, gm_n2070, gm_n2071, gm_n2072, gm_n2073, gm_n2074, gm_n2075, gm_n2076, gm_n208, gm_n209, gm_n210, gm_n211, gm_n212, gm_n213, gm_n214, gm_n216, gm_n217, gm_n218, gm_n219, gm_n220, gm_n221, gm_n222, gm_n223, gm_n224, gm_n225, gm_n226, gm_n227, gm_n228, gm_n229, gm_n230, gm_n231, gm_n232, gm_n233, gm_n234, gm_n235, gm_n236, gm_n237, gm_n238, gm_n239, gm_n240, gm_n241, gm_n242, gm_n243, gm_n244, gm_n245, gm_n246, gm_n247, gm_n248, gm_n249, gm_n250, gm_n251, gm_n252, gm_n253, gm_n254, gm_n255, gm_n256, gm_n257, gm_n258, gm_n259, gm_n260, gm_n261, gm_n262, gm_n263, gm_n264, gm_n265, gm_n266, gm_n267, gm_n268, gm_n269, gm_n270, gm_n271, gm_n272, gm_n273, gm_n274, gm_n275, gm_n276, gm_n277, gm_n278, gm_n279, gm_n280, gm_n281, gm_n282, gm_n283, gm_n284, gm_n285, gm_n286, gm_n287, gm_n288, gm_n289, gm_n290, gm_n291, gm_n292, gm_n293, gm_n294, gm_n295, gm_n296, gm_n297, gm_n298, gm_n299, gm_n300, gm_n301, gm_n302, gm_n303, gm_n304, gm_n305, gm_n306, gm_n307, gm_n308, gm_n309, gm_n310, gm_n311, gm_n312, gm_n313, gm_n314, gm_n315, gm_n316, gm_n317, gm_n318, gm_n319, gm_n320, gm_n321, gm_n322, gm_n323, gm_n324, gm_n325, gm_n326, gm_n327, gm_n328, gm_n329, gm_n330, gm_n331, gm_n332, gm_n333, gm_n334, gm_n335, gm_n336, gm_n337, gm_n338, gm_n339, gm_n340, gm_n341, gm_n342, gm_n343, gm_n344, gm_n345, gm_n346, gm_n347, gm_n348, gm_n349, gm_n350, gm_n351, gm_n352, gm_n353, gm_n354, gm_n355, gm_n356, gm_n357, gm_n358, gm_n359, gm_n360, gm_n361, gm_n362, gm_n363, gm_n364, gm_n365, gm_n366, gm_n367, gm_n368, gm_n369, gm_n370, gm_n371, gm_n372, gm_n373, gm_n374, gm_n375, gm_n376, gm_n377, gm_n378, gm_n379, gm_n380, gm_n381, gm_n382, gm_n383, gm_n384, gm_n385, gm_n386, gm_n387, gm_n388, gm_n389, gm_n390, gm_n391, gm_n392, gm_n393, gm_n394, gm_n395, gm_n396, gm_n397, gm_n398, gm_n399, gm_n400, gm_n401, gm_n402, gm_n403, gm_n404, gm_n405, gm_n406, gm_n407, gm_n408, gm_n409, gm_n41, gm_n410, gm_n411, gm_n412, gm_n413, gm_n414, gm_n415, gm_n416, gm_n417, gm_n418, gm_n419, gm_n42, gm_n420, gm_n421, gm_n422, gm_n423, gm_n424, gm_n425, gm_n426, gm_n427, gm_n428, gm_n429, gm_n43, gm_n430, gm_n431, gm_n432, gm_n433, gm_n434, gm_n435, gm_n436, gm_n437, gm_n438, gm_n439, gm_n44, gm_n440, gm_n441, gm_n442, gm_n443, gm_n444, gm_n445, gm_n446, gm_n447, gm_n448, gm_n449, gm_n45, gm_n450, gm_n451, gm_n452, gm_n453, gm_n454, gm_n455, gm_n456, gm_n457, gm_n458, gm_n459, gm_n46, gm_n460, gm_n461, gm_n463, gm_n464, gm_n465, gm_n466, gm_n467, gm_n468, gm_n469, gm_n47, gm_n470, gm_n471, gm_n472, gm_n473, gm_n474, gm_n475, gm_n476, gm_n477, gm_n478, gm_n479, gm_n48, gm_n480, gm_n481, gm_n482, gm_n483, gm_n484, gm_n485, gm_n486, gm_n487, gm_n488, gm_n489, gm_n49, gm_n490, gm_n491, gm_n492, gm_n493, gm_n494, gm_n495, gm_n496, gm_n497, gm_n498, gm_n499, gm_n50, gm_n500, gm_n501, gm_n502, gm_n503, gm_n504, gm_n505, gm_n506, gm_n507, gm_n508, gm_n509, gm_n51, gm_n510, gm_n511, gm_n512, gm_n513, gm_n514, gm_n515, gm_n516, gm_n517, gm_n518, gm_n519, gm_n52, gm_n520, gm_n521, gm_n522, gm_n523, gm_n524, gm_n525, gm_n526, gm_n527, gm_n528, gm_n529, gm_n53, gm_n530, gm_n531, gm_n532, gm_n533, gm_n534, gm_n535, gm_n536, gm_n537, gm_n538, gm_n539, gm_n54, gm_n540, gm_n541, gm_n542, gm_n543, gm_n544, gm_n545, gm_n546, gm_n547, gm_n548, gm_n549, gm_n55, gm_n550, gm_n551, gm_n552, gm_n553, gm_n554, gm_n555, gm_n556, gm_n557, gm_n558, gm_n559, gm_n56, gm_n560, gm_n561, gm_n562, gm_n563, gm_n564, gm_n565, gm_n566, gm_n567, gm_n568, gm_n569, gm_n57, gm_n570, gm_n571, gm_n572, gm_n573, gm_n574, gm_n575, gm_n576, gm_n577, gm_n578, gm_n579, gm_n58, gm_n580, gm_n581, gm_n582, gm_n583, gm_n584, gm_n585, gm_n586, gm_n587, gm_n588, gm_n589, gm_n59, gm_n590, gm_n591, gm_n592, gm_n593, gm_n594, gm_n595, gm_n596, gm_n597, gm_n598, gm_n599, gm_n60, gm_n600, gm_n601, gm_n602, gm_n603, gm_n604, gm_n605, gm_n606, gm_n607, gm_n608, gm_n609, gm_n61, gm_n610, gm_n611, gm_n612, gm_n613, gm_n614, gm_n615, gm_n616, gm_n617, gm_n618, gm_n619, gm_n62, gm_n620, gm_n621, gm_n622, gm_n623, gm_n624, gm_n625, gm_n626, gm_n627, gm_n628, gm_n629, gm_n63, gm_n630, gm_n631, gm_n632, gm_n633, gm_n634, gm_n635, gm_n636, gm_n637, gm_n638, gm_n639, gm_n64, gm_n640, gm_n641, gm_n642, gm_n643, gm_n644, gm_n645, gm_n646, gm_n647, gm_n648, gm_n649, gm_n65, gm_n650, gm_n651, gm_n652, gm_n653, gm_n654, gm_n655, gm_n656, gm_n657, gm_n658, gm_n659, gm_n66, gm_n660, gm_n662, gm_n663, gm_n664, gm_n665, gm_n666, gm_n667, gm_n668, gm_n669, gm_n67, gm_n670, gm_n671, gm_n672, gm_n673, gm_n674, gm_n675, gm_n676, gm_n677, gm_n678, gm_n679, gm_n68, gm_n680, gm_n681, gm_n682, gm_n683, gm_n684, gm_n685, gm_n686, gm_n687, gm_n688, gm_n689, gm_n69, gm_n690, gm_n691, gm_n692, gm_n693, gm_n694, gm_n695, gm_n696, gm_n697, gm_n698, gm_n699, gm_n70, gm_n700, gm_n701, gm_n702, gm_n703, gm_n704, gm_n705, gm_n706, gm_n707, gm_n708, gm_n709, gm_n71, gm_n710, gm_n711, gm_n712, gm_n713, gm_n714, gm_n715, gm_n716, gm_n717, gm_n718, gm_n719, gm_n72, gm_n720, gm_n721, gm_n722, gm_n723, gm_n724, gm_n725, gm_n726, gm_n727, gm_n728, gm_n729, gm_n73, gm_n730, gm_n731, gm_n732, gm_n733, gm_n734, gm_n735, gm_n736, gm_n737, gm_n738, gm_n739, gm_n74, gm_n740, gm_n741, gm_n742, gm_n744, gm_n745, gm_n746, gm_n747, gm_n748, gm_n749, gm_n75, gm_n750, gm_n751, gm_n752, gm_n753, gm_n754, gm_n755, gm_n756, gm_n757, gm_n758, gm_n759, gm_n76, gm_n760, gm_n761, gm_n762, gm_n763, gm_n764, gm_n765, gm_n766, gm_n767, gm_n768, gm_n769, gm_n77, gm_n770, gm_n771, gm_n772, gm_n773, gm_n774, gm_n775, gm_n776, gm_n777, gm_n778, gm_n779, gm_n78, gm_n780, gm_n781, gm_n782, gm_n783, gm_n784, gm_n785, gm_n786, gm_n787, gm_n788, gm_n789, gm_n79, gm_n790, gm_n791, gm_n792, gm_n793, gm_n794, gm_n795, gm_n796, gm_n797, gm_n798, gm_n799, gm_n80, gm_n800, gm_n801, gm_n802, gm_n803, gm_n804, gm_n805, gm_n806, gm_n807, gm_n808, gm_n809, gm_n81, gm_n810, gm_n811, gm_n812, gm_n813, gm_n814, gm_n815, gm_n816, gm_n817, gm_n818, gm_n82, gm_n820, gm_n821, gm_n822, gm_n823, gm_n824, gm_n825, gm_n826, gm_n827, gm_n828, gm_n829, gm_n83, gm_n830, gm_n831, gm_n832, gm_n833, gm_n834, gm_n835, gm_n836, gm_n837, gm_n838, gm_n839, gm_n84, gm_n840, gm_n841, gm_n842, gm_n843, gm_n844, gm_n845, gm_n846, gm_n847, gm_n848, gm_n849, gm_n85, gm_n850, gm_n851, gm_n852, gm_n853, gm_n854, gm_n855, gm_n856, gm_n857, gm_n858, gm_n859, gm_n86, gm_n860, gm_n861, gm_n862, gm_n863, gm_n864, gm_n865, gm_n867, gm_n868, gm_n869, gm_n87, gm_n870, gm_n871, gm_n872, gm_n873, gm_n874, gm_n875, gm_n876, gm_n877, gm_n878, gm_n879, gm_n88, gm_n880, gm_n881, gm_n882, gm_n883, gm_n884, gm_n885, gm_n886, gm_n887, gm_n888, gm_n889, gm_n89, gm_n890, gm_n891, gm_n892, gm_n893, gm_n894, gm_n895, gm_n896, gm_n897, gm_n898, gm_n899, gm_n90, gm_n900, gm_n901, gm_n902, gm_n903, gm_n904, gm_n905, gm_n906, gm_n907, gm_n908, gm_n909, gm_n91, gm_n910, gm_n911, gm_n912, gm_n913, gm_n914, gm_n915, gm_n916, gm_n917, gm_n918, gm_n919, gm_n92, gm_n920, gm_n921, gm_n922, gm_n923, gm_n924, gm_n925, gm_n926, gm_n927, gm_n928, gm_n929, gm_n93, gm_n930, gm_n931, gm_n932, gm_n933, gm_n934, gm_n935, gm_n936, gm_n937, gm_n938, gm_n939, gm_n94, gm_n940, gm_n941, gm_n942, gm_n943, gm_n944, gm_n945, gm_n946, gm_n947, gm_n948, gm_n949, gm_n95, gm_n950, gm_n951, gm_n952, gm_n953, gm_n954, gm_n955, gm_n956, gm_n957, gm_n958, gm_n959, gm_n96, gm_n960, gm_n961, gm_n962, gm_n963, gm_n964, gm_n965, gm_n966, gm_n967, gm_n968, gm_n969, gm_n97, gm_n970, gm_n971, gm_n972, gm_n973, gm_n974, gm_n975, gm_n976, gm_n977, gm_n978, gm_n979, gm_n98, gm_n980, gm_n981, gm_n982, gm_n983, gm_n984, gm_n985, gm_n986, gm_n987, gm_n988, gm_n989, gm_n99, gm_n990, gm_n991, gm_n992, gm_n993, gm_n994, gm_n995, gm_n996, gm_n997, gm_n998, gm_n999;
	wire t_8, t_7, t_1, t_9, t_2, t_0, t_6, t_3, t_5, t_4;
	not (gm_n41, in_12);
	not (gm_n42, in_10);
	not (gm_n43, in_11);
	nor (gm_n44, gm_n43, gm_n42, in_9);
	not (gm_n45, in_8);
	nor (gm_n46, in_7, in_6, in_5);
	not (gm_n47, gm_n46);
	not (gm_n48, in_0);
	not (gm_n49, in_1);
	nand (gm_n50, in_2, gm_n49, gm_n48, in_4, in_3);
	nor (gm_n51, gm_n50, gm_n47, gm_n45);
	and (gm_n52, in_14, in_13, gm_n41, gm_n51, gm_n44);
	and (gm_n53, in_11, in_10, in_9);
	not (gm_n54, in_2);
	not (gm_n55, in_3);
	not (gm_n56, in_4);
	nand (gm_n57, gm_n54, in_1, gm_n48, gm_n56, gm_n55);
	not (gm_n58, in_7);
	nand (gm_n59, gm_n58, in_6, in_5);
	nor (gm_n60, gm_n59, gm_n57, gm_n45);
	nand (gm_n61, in_14, in_13, in_12, gm_n60, gm_n53);
	not (gm_n62, in_13);
	nand (gm_n63, gm_n43, in_10, in_9);
	not (gm_n64, in_5);
	nor (gm_n65, gm_n58, in_6, gm_n64);
	nor (gm_n66, in_2, in_1, gm_n48, in_4, gm_n55);
	nand (gm_n67, gm_n66, gm_n65, gm_n45);
	nor (gm_n68, in_14, gm_n62, gm_n41, gm_n67, gm_n63);
	not (gm_n69, in_14);
	not (gm_n70, in_9);
	nand (gm_n71, in_11, in_10, gm_n70);
	nor (gm_n72, gm_n58, in_6, in_5);
	nor (gm_n73, in_2, in_1, gm_n48, gm_n56, in_3);
	nand (gm_n74, gm_n73, gm_n72, gm_n45);
	nor (gm_n75, gm_n69, gm_n62, in_12, gm_n74, gm_n71);
	nand (gm_n76, in_11, in_10, in_9);
	nand (gm_n77, gm_n69, in_13, in_12);
	or (gm_n78, gm_n76, gm_n47, in_8, gm_n77, gm_n57);
	not (gm_n79, in_6);
	nor (gm_n80, gm_n58, gm_n79, in_5);
	nor (gm_n81, in_2, in_1, gm_n48, in_4, in_3);
	nand (gm_n82, gm_n81, gm_n80, in_8);
	nor (gm_n83, gm_n62, gm_n41, in_11);
	not (gm_n84, gm_n83);
	or (gm_n85, gm_n69, in_10, in_9, gm_n84, gm_n82);
	and (gm_n86, in_13, in_12, in_11);
	not (gm_n87, gm_n86);
	and (gm_n88, in_7, in_6, in_5);
	not (gm_n89, gm_n88);
	nand (gm_n90, gm_n54, in_1, in_0, in_4, gm_n55);
	or (gm_n91, gm_n42, gm_n70, gm_n45, gm_n90, gm_n89);
	nor (gm_n92, gm_n91, gm_n87, in_14);
	nor (gm_n93, gm_n43, in_10, in_9);
	nand (gm_n94, gm_n58, in_6, gm_n64);
	nand (gm_n95, in_2, gm_n49, in_0, gm_n56, in_3);
	nor (gm_n96, gm_n95, gm_n94, in_8);
	and (gm_n97, in_14, in_13, gm_n41, gm_n96, gm_n93);
	nor (gm_n98, in_11, in_10, gm_n70);
	nor (gm_n99, gm_n95, gm_n89, in_8);
	nand (gm_n100, in_14, in_13, in_12, gm_n99, gm_n98);
	nor (gm_n101, in_13, in_12, in_11);
	nor (gm_n102, in_10, in_9, gm_n45, gm_n90, gm_n47);
	nand (gm_n103, gm_n102, gm_n101, gm_n69);
	nor (gm_n104, gm_n69, in_13, in_12);
	nor (gm_n105, in_2, in_1, gm_n48, gm_n56, gm_n55);
	nor (gm_n106, in_10, in_9, in_8);
	nand (gm_n107, gm_n104, gm_n65, gm_n43, gm_n106, gm_n105);
	not (gm_n108, gm_n101);
	nor (gm_n109, in_7, gm_n79, gm_n64);
	nor (gm_n110, gm_n54, gm_n49, in_0, gm_n56, gm_n55);
	nand (gm_n111, gm_n110, gm_n109, gm_n45);
	or (gm_n112, in_14, gm_n42, in_9, gm_n111, gm_n108);
	nand (gm_n113, gm_n103, gm_n100, t_5, gm_n112, gm_n107);
	nor (gm_n114, in_2, in_1, in_0, in_3);
	and (gm_n115, gm_n79, gm_n64, in_4, gm_n114, gm_n58);
	nor (gm_n116, gm_n42, in_9, in_8);
	nor (gm_n117, gm_n69, in_13, gm_n41);
	nand (gm_n118, gm_n116, gm_n115, in_11, gm_n117);
	nand (gm_n119, gm_n62, in_12, in_11);
	or (gm_n120, in_2, in_1, in_0);
	or (gm_n121, gm_n64, in_4, gm_n55, gm_n120, in_6);
	nand (gm_n122, in_9, in_8, gm_n58);
	or (gm_n123, gm_n119, gm_n69, in_10, gm_n122, gm_n121);
	and (gm_n124, in_2, in_1, in_0, in_4, in_3);
	and (gm_n125, in_7, in_6, gm_n64, gm_n124, gm_n45);
	nor (gm_n126, gm_n43, in_10, gm_n70);
	nand (gm_n127, in_14, in_13, gm_n41, gm_n126, gm_n125);
	nand (gm_n128, gm_n127, gm_n123, gm_n118);
	nor (gm_n129, in_2, gm_n49, gm_n48, gm_n56, gm_n55);
	and (gm_n130, gm_n129, gm_n88, in_8);
	nor (gm_n131, in_11, gm_n42, in_9);
	and (gm_n132, gm_n69, gm_n62, in_12, gm_n131, gm_n130);
	nor (gm_n133, gm_n54, in_1, in_0, gm_n56, in_3);
	nand (gm_n134, gm_n133, gm_n88, gm_n45);
	nor (gm_n135, in_14, in_13, gm_n41, gm_n134, gm_n63);
	nor (gm_n136, in_13, gm_n41, in_11);
	nand (gm_n137, in_2, in_1, in_0);
	nor (gm_n138, gm_n64, in_4, in_3, gm_n137, gm_n79);
	nor (gm_n139, gm_n70, in_8, in_7);
	and (gm_n140, gm_n136, in_14, gm_n42, gm_n139, gm_n138);
	or (gm_n141, gm_n140, gm_n135, gm_n132);
	nor (gm_n142, gm_n113, gm_n97, gm_n92, gm_n141, gm_n128);
	or (gm_n143, in_5, gm_n56, gm_n55, gm_n120, in_6);
	and (gm_n144, in_9, in_8, in_7);
	not (gm_n145, gm_n144);
	nor (gm_n146, gm_n119, gm_n69, in_10, gm_n145, gm_n143);
	nand (gm_n147, in_2, in_1, gm_n48, in_4, gm_n55);
	nor (gm_n148, gm_n147, gm_n94, gm_n45);
	and (gm_n149, in_14, gm_n62, gm_n41, gm_n148, gm_n98);
	nand (gm_n150, in_7, in_6, gm_n64);
	or (gm_n151, in_10, gm_n70, in_8, gm_n147, gm_n150);
	nor (gm_n152, gm_n151, gm_n87, gm_n69);
	nor (gm_n153, gm_n152, gm_n149, gm_n146);
	not (gm_n154, gm_n104);
	not (gm_n155, gm_n138);
	nand (gm_n156, in_10, gm_n70, in_8);
	nor (gm_n157, gm_n154, in_11, gm_n58, gm_n156, gm_n155);
	nor (gm_n158, gm_n54, gm_n49, in_0, gm_n56, in_3);
	nand (gm_n159, gm_n44, gm_n41, in_8, gm_n158, gm_n109);
	nor (gm_n160, gm_n159, in_14, gm_n62);
	nor (gm_n161, in_7, gm_n79, in_5);
	nand (gm_n162, in_10, in_9, gm_n45);
	not (gm_n163, gm_n162);
	nor (gm_n164, in_14, in_13, gm_n41);
	and (gm_n165, gm_n133, gm_n161, gm_n43, gm_n164, gm_n163);
	nor (gm_n166, gm_n165, gm_n160, gm_n157);
	nand (gm_n167, gm_n142, gm_n85, gm_n78, gm_n166, gm_n153);
	and (gm_n168, in_14, in_13, in_12);
	nor (gm_n169, in_10, gm_n70, gm_n45);
	nor (gm_n170, gm_n54, in_1, gm_n48, in_4, in_3);
	nand (gm_n171, gm_n168, gm_n88, in_11, gm_n170, gm_n169);
	and (gm_n172, gm_n42, in_9, in_8, gm_n105, gm_n72);
	nand (gm_n173, gm_n172, gm_n86, in_14);
	nor (gm_n174, gm_n69, gm_n62, in_12);
	nand (gm_n175, gm_n161, gm_n44, in_8, gm_n174, gm_n105);
	nand (gm_n176, gm_n175, gm_n173, gm_n171);
	nand (gm_n177, in_13, gm_n41, gm_n43);
	not (gm_n178, gm_n177);
	nor (gm_n179, gm_n89, gm_n57, in_8);
	nand (gm_n180, in_14, gm_n42, gm_n70, gm_n179, gm_n178);
	nor (gm_n181, gm_n90, gm_n47, in_8);
	nand (gm_n182, in_14, in_13, in_12, gm_n181, gm_n93);
	nor (gm_n183, in_7, in_6, gm_n64);
	nor (gm_n184, gm_n54, gm_n49, in_0, in_4, gm_n55);
	and (gm_n185, gm_n184, gm_n183, gm_n45);
	nand (gm_n186, in_14, in_13, gm_n41, gm_n185, gm_n53);
	nand (gm_n187, gm_n186, gm_n182, gm_n180);
	nor (gm_n188, gm_n167, gm_n75, gm_n68, gm_n187, gm_n176);
	or (gm_n189, in_2, in_1, in_0, in_4, in_3);
	nor (gm_n190, gm_n58, gm_n79, gm_n64, gm_n189, gm_n45);
	nor (gm_n191, in_11, in_10, in_9);
	nand (gm_n192, gm_n69, in_13, in_12, gm_n191, gm_n190);
	nand (gm_n193, gm_n54, in_1, in_0, gm_n56, gm_n55);
	nor (gm_n194, gm_n193, gm_n94, in_8);
	nand (gm_n195, in_14, gm_n62, in_12, gm_n194, gm_n93);
	nor (gm_n196, gm_n58, gm_n79, gm_n64, gm_n189, in_8);
	nand (gm_n197, gm_n69, in_10, gm_n70, gm_n196, gm_n136);
	nand (gm_n198, gm_n192, gm_n188, gm_n61, gm_n197, gm_n195);
	nor (gm_n199, in_2, gm_n49, in_0, in_4, gm_n55);
	nand (gm_n200, gm_n169, gm_n136, in_14, gm_n199, gm_n183);
	nand (gm_n201, in_2, gm_n49, gm_n48, gm_n56, gm_n55);
	nor (gm_n202, gm_n201, gm_n150, in_8);
	nand (gm_n203, gm_n69, in_10, in_9, gm_n202, gm_n178);
	and (gm_n204, gm_n199, gm_n80, in_8);
	nand (gm_n205, in_14, gm_n62, gm_n41, gm_n204, gm_n44);
	nand (gm_n206, gm_n205, gm_n203, gm_n200);
	nand (gm_n207, gm_n80, gm_n53, gm_n45, gm_n168, gm_n133);
	nand (gm_n208, gm_n58, gm_n79, in_5);
	nor (gm_n209, gm_n208, gm_n57, gm_n45);
	nand (gm_n210, in_14, in_13, in_12, gm_n209, gm_n93);
	nor (gm_n211, in_5, gm_n56, in_3, gm_n137, gm_n79);
	nor (gm_n212, in_9, in_8, in_7);
	nand (gm_n213, gm_n178, gm_n69, gm_n42, gm_n212, gm_n211);
	nand (gm_n214, gm_n213, gm_n210, gm_n207);
	nor (out_0, gm_n206, gm_n198, gm_n52, gm_n214);
	nand (gm_n216, in_11, gm_n42, gm_n70);
	nand (gm_n217, gm_n133, gm_n109, gm_n45);
	nor (gm_n218, gm_n69, gm_n62, in_12, gm_n217, gm_n216);
	nand (gm_n219, gm_n54, gm_n49, in_0, gm_n56, in_3);
	nor (gm_n220, gm_n150, gm_n219, gm_n45);
	nand (gm_n221, gm_n69, gm_n62, in_12, gm_n220, gm_n44);
	nor (gm_n222, gm_n90, gm_n59, gm_n45);
	nand (gm_n223, gm_n69, in_13, gm_n41, gm_n222, gm_n93);
	nor (gm_n224, in_14, in_13, in_12);
	not (gm_n225, gm_n224);
	nand (gm_n226, gm_n42, gm_n70, in_8);
	nand (gm_n227, in_2, gm_n49, in_0, in_4, in_3);
	nor (gm_n228, gm_n225, gm_n59, in_11, gm_n227, gm_n226);
	nand (gm_n229, gm_n69, gm_n62, in_12);
	not (gm_n230, gm_n191);
	nand (gm_n231, gm_n54, in_1, in_0, gm_n56, in_3);
	nor (gm_n232, gm_n229, gm_n59, in_8, gm_n231, gm_n230);
	and (gm_n233, in_10, in_9, in_8);
	nand (gm_n234, gm_n124, gm_n109, in_11, gm_n233, gm_n164);
	and (gm_n235, gm_n53, gm_n41, in_8, gm_n129, gm_n72);
	nand (gm_n236, gm_n235, in_14, in_13);
	or (gm_n237, in_5, in_4, in_3, gm_n137, gm_n79);
	nor (gm_n238, gm_n87, in_14, in_10, gm_n237, gm_n145);
	nand (gm_n239, gm_n62, gm_n41, in_11);
	and (gm_n240, in_2, in_1, in_0, in_3);
	nand (gm_n241, gm_n79, gm_n64, gm_n56, gm_n240, in_7);
	nor (gm_n242, gm_n239, gm_n162, in_14, gm_n241);
	nor (gm_n243, in_14, gm_n62, gm_n41);
	nand (gm_n244, gm_n243, gm_n65, in_11, gm_n184, gm_n163);
	not (gm_n245, gm_n119);
	nor (gm_n246, in_2, gm_n49, in_0, gm_n56, in_3);
	and (gm_n247, in_10, in_9, in_8, gm_n246, gm_n46);
	nand (gm_n248, gm_n247, gm_n245, in_14);
	not (gm_n249, gm_n106);
	nor (gm_n250, gm_n154, gm_n150, gm_n43, gm_n189, gm_n249);
	nor (gm_n251, gm_n231, gm_n59, gm_n45);
	and (gm_n252, gm_n69, gm_n62, gm_n41, gm_n251, gm_n93);
	and (gm_n253, in_6, gm_n64, gm_n56, gm_n240, in_7);
	nand (gm_n254, gm_n174, gm_n116, in_11, gm_n253);
	nor (gm_n255, gm_n54, gm_n49, in_0, in_4, in_3);
	nand (gm_n256, gm_n255, gm_n161, gm_n45);
	or (gm_n257, in_14, gm_n62, gm_n41, gm_n256, gm_n63);
	nor (gm_n258, gm_n64, gm_n56, gm_n55, gm_n120, in_6);
	not (gm_n259, gm_n258);
	nor (gm_n260, gm_n108, gm_n69, in_10, gm_n259, gm_n122);
	nand (gm_n261, in_11, gm_n42, in_9);
	nand (gm_n262, gm_n158, gm_n88, in_8);
	nor (gm_n263, gm_n69, in_13, in_12, gm_n262, gm_n261);
	and (gm_n264, gm_n105, gm_n80, in_8);
	nand (gm_n265, gm_n69, gm_n62, in_12, gm_n264, gm_n98);
	nor (gm_n266, in_10, gm_n70, in_8);
	nand (gm_n267, gm_n86, gm_n72, gm_n69, gm_n266, gm_n199);
	nor (gm_n268, in_2, gm_n49, in_0, gm_n56, gm_n55);
	nand (gm_n269, gm_n42, in_9, in_8, gm_n268, gm_n80);
	nor (gm_n270, gm_n269, gm_n239, gm_n69);
	nand (gm_n271, in_13, gm_n41, in_11);
	nand (gm_n272, gm_n42, gm_n70, gm_n45, gm_n129, gm_n46);
	nor (gm_n273, gm_n272, gm_n271, in_14);
	nor (gm_n274, gm_n54, in_1, in_0, in_4, gm_n55);
	and (gm_n275, gm_n161, in_12, gm_n45, gm_n274, gm_n126);
	nand (gm_n276, gm_n275, gm_n69, in_13);
	nor (gm_n277, gm_n54, in_1, gm_n48, gm_n56, in_3);
	and (gm_n278, gm_n277, gm_n109, gm_n45);
	nand (gm_n279, gm_n69, gm_n42, in_9, gm_n278, gm_n178);
	nand (gm_n280, in_2, in_1, gm_n48, in_4, in_3);
	nor (gm_n281, gm_n77, gm_n59, gm_n43, gm_n156, gm_n280);
	nand (gm_n282, gm_n161, gm_n73, in_8);
	nor (gm_n283, gm_n69, in_10, in_9, gm_n282, gm_n87);
	nor (gm_n284, in_10, in_9, gm_n45);
	and (gm_n285, gm_n81, gm_n65, gm_n43, gm_n284, gm_n168);
	nand (gm_n286, gm_n70, in_8, in_7);
	or (gm_n287, gm_n64, gm_n56, in_3, gm_n137, gm_n79);
	nor (gm_n288, gm_n108, gm_n69, in_10, gm_n287, gm_n286);
	nor (gm_n289, in_9, gm_n45, gm_n58);
	nand (gm_n290, gm_n110, gm_n79, in_5, gm_n289);
	nor (gm_n291, gm_n108, in_14, in_10, gm_n290);
	nor (gm_n292, gm_n285, gm_n283, gm_n281, gm_n291, gm_n288);
	nand (gm_n293, gm_n277, gm_n183, in_8);
	nor (gm_n294, in_14, in_13, gm_n41, gm_n293, gm_n63);
	nor (gm_n295, in_14, gm_n62, in_12);
	and (gm_n296, gm_n183, gm_n131, in_8, gm_n295, gm_n246);
	or (gm_n297, gm_n76, in_12, in_8, gm_n231, gm_n208);
	nor (gm_n298, gm_n297, gm_n69, gm_n62);
	nor (gm_n299, gm_n298, gm_n296, gm_n294);
	nor (gm_n300, in_13, in_12, gm_n43);
	nand (gm_n301, in_2, gm_n49, gm_n48, gm_n56, in_3);
	nand (gm_n302, gm_n70, in_8, gm_n58);
	nor (gm_n303, gm_n301, in_6, gm_n64, gm_n302);
	and (gm_n304, gm_n300, in_14, gm_n42, gm_n303);
	or (gm_n305, in_5, gm_n56, in_3, gm_n137, in_6);
	nor (gm_n306, gm_n122, gm_n69, gm_n42, gm_n305, gm_n271);
	nand (gm_n307, in_9, gm_n45, in_7);
	nor (gm_n308, gm_n239, in_14, in_10, gm_n307, gm_n287);
	nor (gm_n309, gm_n308, gm_n306, gm_n304);
	nand (gm_n310, gm_n292, gm_n279, gm_n276, gm_n309, gm_n299);
	and (gm_n311, in_6, in_5, gm_n56, gm_n240, gm_n58);
	nand (gm_n312, gm_n163, gm_n243, in_11, gm_n311);
	nor (gm_n313, gm_n201, gm_n150, gm_n45);
	nand (gm_n314, in_14, gm_n62, gm_n41, gm_n313, gm_n98);
	nor (gm_n315, gm_n150, gm_n41, in_8, gm_n280, gm_n216);
	nand (gm_n316, gm_n315, gm_n69, in_13);
	nand (gm_n317, gm_n316, gm_n314, gm_n312);
	and (gm_n318, gm_n81, gm_n65, gm_n45);
	nand (gm_n319, gm_n69, in_13, gm_n41, gm_n318, gm_n93);
	nor (gm_n320, in_2, gm_n49, gm_n48, gm_n56, in_3);
	nand (gm_n321, gm_n161, gm_n320, in_11, gm_n174, gm_n106);
	not (gm_n322, gm_n122);
	nor (gm_n323, gm_n64, gm_n56, gm_n55, gm_n120, gm_n79);
	nand (gm_n324, gm_n86, in_14, gm_n42, gm_n323, gm_n322);
	nand (gm_n325, gm_n324, gm_n321, gm_n319);
	nor (gm_n326, gm_n310, gm_n273, gm_n270, gm_n325, gm_n317);
	nand (gm_n327, gm_n43, in_10, gm_n70);
	nor (gm_n328, gm_n69, in_13, in_12, gm_n134, gm_n327);
	nor (gm_n329, gm_n64, gm_n56, in_3, gm_n137, in_6);
	not (gm_n330, gm_n329);
	nor (gm_n331, gm_n122, in_14, gm_n42, gm_n330, gm_n239);
	and (gm_n332, gm_n163, gm_n72, gm_n43, gm_n268, gm_n168);
	nor (gm_n333, gm_n332, gm_n331, gm_n328);
	and (gm_n334, gm_n98, gm_n109, gm_n45, gm_n133, gm_n117);
	nand (gm_n335, in_7, gm_n79, in_5, gm_n124, gm_n45);
	nor (gm_n336, gm_n69, in_13, in_12, gm_n335, gm_n76);
	and (gm_n337, gm_n83, in_14, in_10, gm_n258, gm_n212);
	nor (gm_n338, gm_n337, gm_n336, gm_n334);
	nand (gm_n339, gm_n326, gm_n267, gm_n265, gm_n338, gm_n333);
	nor (gm_n340, in_7, in_6, gm_n64, gm_n189, gm_n45);
	nand (gm_n341, gm_n340, gm_n295, gm_n93);
	nand (gm_n342, gm_n43, gm_n42, in_9);
	nand (gm_n343, gm_n170, gm_n109, in_8);
	or (gm_n344, in_14, in_13, in_12, gm_n343, gm_n342);
	not (gm_n345, gm_n271);
	nor (gm_n346, in_5, in_4, gm_n55, gm_n120, in_6);
	nand (gm_n347, gm_n345, in_14, gm_n42, gm_n346, gm_n289);
	nand (gm_n348, gm_n347, gm_n344, gm_n341);
	nor (gm_n349, in_11, gm_n42, gm_n70);
	nand (gm_n350, gm_n69, in_13, gm_n41, gm_n313, gm_n349);
	nand (gm_n351, in_7, gm_n79, in_5);
	or (gm_n352, in_10, gm_n70, in_8, gm_n189, gm_n351);
	or (gm_n353, gm_n352, gm_n271, in_14);
	nand (gm_n354, gm_n131, gm_n72, in_8, gm_n295, gm_n246);
	nand (gm_n355, gm_n354, gm_n353, gm_n350);
	nor (gm_n356, gm_n339, gm_n263, gm_n260, gm_n355, gm_n348);
	and (gm_n357, gm_n110, gm_n88, in_14, gm_n300, gm_n169);
	nor (gm_n358, gm_n231, gm_n150, gm_n45);
	and (gm_n359, in_14, in_10, gm_n70, gm_n358, gm_n300);
	nand (gm_n360, gm_n158, gm_n46, in_8);
	nor (gm_n361, in_14, in_13, in_12, gm_n360, gm_n63);
	nor (gm_n362, gm_n361, gm_n359, gm_n357);
	nand (gm_n363, gm_n161, gm_n243, in_8, gm_n191, gm_n184);
	nand (gm_n364, gm_n255, gm_n46, in_8);
	or (gm_n365, in_14, in_13, gm_n41, gm_n364, gm_n76);
	nand (gm_n366, gm_n184, gm_n46, in_8);
	or (gm_n367, gm_n69, gm_n42, in_9, gm_n366, gm_n271);
	and (gm_n368, gm_n367, gm_n365, gm_n363);
	nand (gm_n369, gm_n356, gm_n257, gm_n254, gm_n368, gm_n362);
	nor (gm_n370, gm_n54, in_1, in_0, gm_n56, gm_n55);
	and (gm_n371, gm_n370, gm_n41, gm_n45, gm_n191, gm_n65);
	nand (gm_n372, gm_n371, in_14, in_13);
	and (gm_n373, in_6, in_5, in_4, gm_n114, gm_n58);
	nand (gm_n374, gm_n295, gm_n284, in_11, gm_n373);
	nand (gm_n375, gm_n69, gm_n42, in_9, gm_n278, gm_n345);
	nand (gm_n376, gm_n375, gm_n374, gm_n372);
	nand (gm_n377, gm_n161, gm_n370, gm_n45);
	or (gm_n378, gm_n69, gm_n62, gm_n41, gm_n377, gm_n63);
	nor (gm_n379, gm_n227, gm_n89, gm_n45);
	nand (gm_n380, gm_n69, in_13, in_12, gm_n379, gm_n131);
	nor (gm_n381, in_2, gm_n49, gm_n48, in_4, gm_n55);
	nand (gm_n382, gm_n136, gm_n65, in_14, gm_n266, gm_n381);
	nand (gm_n383, gm_n382, gm_n380, gm_n378);
	nor (gm_n384, gm_n369, gm_n252, gm_n250, gm_n383, gm_n376);
	nand (gm_n385, in_7, gm_n79, gm_n64);
	nor (gm_n386, gm_n227, gm_n385, gm_n45);
	and (gm_n387, in_14, in_13, gm_n41, gm_n386, gm_n98);
	nand (gm_n388, gm_n73, gm_n46, in_8);
	nor (gm_n389, gm_n69, gm_n42, in_9, gm_n388, gm_n119);
	and (gm_n390, gm_n371, gm_n69, gm_n62);
	nor (gm_n391, gm_n390, gm_n389, gm_n387);
	and (gm_n392, gm_n79, in_5, gm_n56, gm_n240, gm_n58);
	and (gm_n393, gm_n116, gm_n104, in_11, gm_n392);
	and (gm_n394, gm_n246, gm_n88, in_8);
	and (gm_n395, in_14, in_10, gm_n70, gm_n394, gm_n345);
	nand (gm_n396, in_2, gm_n49, in_0, gm_n56, gm_n55);
	nor (gm_n397, gm_n396, gm_n351, in_8);
	and (gm_n398, in_14, in_13, in_12, gm_n397, gm_n93);
	nor (gm_n399, gm_n398, gm_n395, gm_n393);
	nand (gm_n400, gm_n384, gm_n248, gm_n244, gm_n399, gm_n391);
	or (gm_n401, gm_n69, gm_n62, in_12, gm_n335, gm_n230);
	nand (gm_n402, gm_n243, gm_n44, in_8, gm_n81, gm_n80);
	and (gm_n403, gm_n129, gm_n80, in_8);
	nand (gm_n404, in_14, in_13, gm_n41, gm_n403, gm_n98);
	nand (gm_n405, gm_n404, gm_n402, gm_n401);
	nand (gm_n406, gm_n295, gm_n233, gm_n43, gm_n392);
	nand (gm_n407, gm_n81, gm_n80, in_8, gm_n168, gm_n131);
	and (gm_n408, gm_n66, in_12, in_8, gm_n183, gm_n131);
	nand (gm_n409, gm_n408, gm_n69, gm_n62);
	nand (gm_n410, gm_n409, gm_n407, gm_n406);
	nor (gm_n411, gm_n400, gm_n242, gm_n238, gm_n410, gm_n405);
	and (gm_n412, gm_n349, gm_n109, gm_n45, gm_n295, gm_n255);
	and (gm_n413, gm_n126, gm_n65, gm_n45, gm_n224, gm_n170);
	or (gm_n414, gm_n89, gm_n57, gm_n45);
	nor (gm_n415, in_14, gm_n62, gm_n41, gm_n414, gm_n327);
	nor (gm_n416, gm_n415, gm_n413, gm_n412);
	nand (gm_n417, gm_n62, in_12, gm_n43);
	not (gm_n418, gm_n139);
	or (gm_n419, in_5, gm_n56, gm_n55, gm_n120, gm_n79);
	nor (gm_n420, gm_n417, in_14, in_10, gm_n419, gm_n418);
	and (gm_n421, gm_n73, gm_n44, gm_n45, gm_n88, gm_n243);
	and (gm_n422, gm_n136, in_14, gm_n42, gm_n258, gm_n144);
	nor (gm_n423, gm_n422, gm_n421, gm_n420);
	nand (gm_n424, gm_n411, gm_n236, gm_n234, gm_n423, gm_n416);
	nand (gm_n425, gm_n117, gm_n72, in_8, gm_n246, gm_n131);
	nor (gm_n426, gm_n208, gm_n147, gm_n45);
	nand (gm_n427, in_14, in_13, in_12, gm_n426, gm_n53);
	nor (gm_n428, gm_n208, gm_n95, gm_n45);
	nand (gm_n429, in_14, gm_n62, in_12, gm_n428, gm_n191);
	nand (gm_n430, gm_n429, gm_n427, gm_n425);
	or (gm_n431, gm_n143, in_14, gm_n42, gm_n302, gm_n177);
	and (gm_n432, gm_n161, gm_n81, gm_n45);
	nand (gm_n433, gm_n69, in_13, in_12, gm_n432, gm_n349);
	nand (gm_n434, gm_n109, gm_n370, gm_n45);
	or (gm_n435, in_14, in_10, gm_n70, gm_n434, gm_n119);
	nand (gm_n436, gm_n435, gm_n433, gm_n431);
	nor (gm_n437, gm_n424, gm_n232, gm_n228, gm_n436, gm_n430);
	nand (gm_n438, gm_n277, gm_n183, gm_n45);
	nor (gm_n439, gm_n69, in_13, in_12, gm_n438, gm_n327);
	nor (gm_n440, gm_n71, gm_n41, in_8, gm_n193, gm_n208);
	and (gm_n441, gm_n440, in_14, in_13);
	nand (gm_n442, gm_n88, gm_n44, in_8, gm_n133);
	nor (gm_n443, in_14, gm_n62, in_12, gm_n442);
	nor (gm_n444, gm_n443, gm_n441, gm_n439);
	nand (gm_n445, gm_n86, gm_n69, in_10, gm_n289, gm_n211);
	nand (gm_n446, gm_n105, gm_n88, in_8);
	or (gm_n447, gm_n69, gm_n62, in_12, gm_n446, gm_n63);
	nand (gm_n448, gm_n345, gm_n102, gm_n69);
	and (gm_n449, gm_n448, gm_n447, gm_n445);
	nand (gm_n450, gm_n437, gm_n223, gm_n221, gm_n449, gm_n444);
	and (gm_n451, gm_n42, gm_n70, gm_n45, gm_n199, gm_n161);
	nand (gm_n452, gm_n451, gm_n300, in_14);
	nand (gm_n453, gm_n73, gm_n65, gm_n43, gm_n295, gm_n284);
	not (gm_n454, gm_n305);
	nand (gm_n455, gm_n139, in_14, in_10, gm_n454, gm_n178);
	nand (gm_n456, gm_n455, gm_n453, gm_n452);
	nand (gm_n457, gm_n136, gm_n109, in_14, gm_n266, gm_n170);
	nand (gm_n458, gm_n81, gm_n65, gm_n43, gm_n284, gm_n104);
	nor (gm_n459, gm_n201, gm_n208, gm_n45);
	nand (gm_n460, gm_n69, gm_n62, gm_n41, gm_n459, gm_n98);
	nand (gm_n461, gm_n460, gm_n458, gm_n457);
	nor (out_1, gm_n456, gm_n450, gm_n218, gm_n461);
	and (gm_n463, in_14, in_13, gm_n41, gm_n379, gm_n53);
	or (gm_n464, gm_n90, gm_n385, gm_n43, gm_n225, gm_n156);
	and (gm_n465, gm_n66, gm_n41, gm_n45, gm_n126, gm_n161);
	nand (gm_n466, gm_n465, in_14, gm_n62);
	not (gm_n467, gm_n212);
	nor (gm_n468, gm_n119, in_14, in_10, gm_n419, gm_n467);
	nand (gm_n469, gm_n42, gm_n70, gm_n45, gm_n274, gm_n161);
	nor (gm_n470, gm_n469, gm_n108, in_14);
	and (gm_n471, gm_n255, gm_n72, in_8);
	nand (gm_n472, gm_n69, in_13, gm_n41, gm_n471, gm_n53);
	or (gm_n473, gm_n108, gm_n69, in_10, gm_n237, gm_n467);
	nand (gm_n474, gm_n80, gm_n66, gm_n45);
	nor (gm_n475, gm_n69, in_13, gm_n41, gm_n474, gm_n342);
	nor (gm_n476, gm_n69, in_10, gm_n70, gm_n446, gm_n84);
	nand (gm_n477, gm_n116, gm_n83, in_14, gm_n199, gm_n183);
	nor (gm_n478, gm_n208, gm_n396, in_8);
	nand (gm_n479, gm_n69, in_13, gm_n41, gm_n478, gm_n131);
	and (gm_n480, gm_n199, gm_n109, in_8);
	and (gm_n481, gm_n69, in_13, gm_n41, gm_n480, gm_n98);
	and (gm_n482, gm_n161, gm_n93, gm_n45, gm_n246, gm_n168);
	or (gm_n483, in_14, gm_n62, in_12, gm_n282, gm_n76);
	and (gm_n484, gm_n109, in_12, gm_n45, gm_n255, gm_n93);
	nand (gm_n485, gm_n484, gm_n69, in_13);
	and (gm_n486, gm_n124, gm_n88, gm_n45);
	and (gm_n487, gm_n69, gm_n62, in_12, gm_n486, gm_n131);
	and (gm_n488, gm_n73, gm_n46, gm_n45);
	and (gm_n489, in_14, gm_n62, in_12, gm_n488, gm_n93);
	nor (gm_n490, gm_n42, in_9, in_8, gm_n193, gm_n150);
	nand (gm_n491, gm_n490, gm_n245, in_14);
	and (gm_n492, gm_n124, gm_n46, in_8);
	nand (gm_n493, gm_n69, gm_n62, gm_n41, gm_n492, gm_n93);
	nor (gm_n494, gm_n69, in_13, in_12, gm_n366, gm_n230);
	and (gm_n495, gm_n116, gm_n161, gm_n43, gm_n124, gm_n117);
	nand (gm_n496, gm_n69, gm_n62, in_12, gm_n148, gm_n44);
	nand (gm_n497, gm_n126, gm_n104, gm_n60);
	nand (gm_n498, gm_n88, in_12, in_8, gm_n274, gm_n126);
	nor (gm_n499, gm_n498, gm_n69, gm_n62);
	nand (gm_n500, gm_n381, gm_n183, in_8);
	nor (gm_n501, gm_n69, gm_n62, gm_n41, gm_n500, gm_n76);
	nor (gm_n502, in_14, in_13, in_12, gm_n262, gm_n216);
	nand (gm_n503, gm_n79, in_5, in_4, gm_n114, gm_n58);
	nor (gm_n504, gm_n177, gm_n249, in_14, gm_n503);
	nor (gm_n505, gm_n57, gm_n47, in_8);
	and (gm_n506, in_14, gm_n62, gm_n41, gm_n505, gm_n349);
	nor (gm_n507, gm_n502, gm_n501, gm_n499, gm_n506, gm_n504);
	nor (gm_n508, gm_n145, in_14, in_10, gm_n287, gm_n271);
	nand (gm_n509, gm_n349, in_12, gm_n45, gm_n274, gm_n80);
	nor (gm_n510, gm_n509, gm_n69, gm_n62);
	or (gm_n511, gm_n42, in_9, gm_n45, gm_n193, gm_n351);
	nor (gm_n512, gm_n511, gm_n417, gm_n69);
	nor (gm_n513, gm_n512, gm_n510, gm_n508);
	nand (gm_n514, gm_n320, gm_n65, in_8);
	nor (gm_n515, gm_n69, gm_n62, in_12, gm_n514, gm_n63);
	nand (gm_n516, gm_n69, in_13, gm_n41);
	nor (gm_n517, gm_n94, gm_n90, in_11, gm_n516, gm_n226);
	nor (gm_n518, in_14, gm_n62, gm_n41, gm_n414, gm_n216);
	nor (gm_n519, gm_n518, gm_n517, gm_n515);
	nand (gm_n520, gm_n507, gm_n497, gm_n496, gm_n519, gm_n513);
	nand (gm_n521, gm_n184, gm_n161, in_8);
	or (gm_n522, in_14, gm_n42, in_9, gm_n521, gm_n177);
	nand (gm_n523, gm_n69, gm_n62, in_12, gm_n196, gm_n53);
	nand (gm_n524, in_14, gm_n62, gm_n41, gm_n264, gm_n44);
	nand (gm_n525, gm_n524, gm_n523, gm_n522);
	nand (gm_n526, gm_n69, in_13, in_12, gm_n397, gm_n98);
	and (gm_n527, gm_n255, gm_n72, gm_n45);
	nand (gm_n528, gm_n69, gm_n62, in_12, gm_n527, gm_n191);
	or (gm_n529, gm_n193, gm_n47, gm_n45);
	or (gm_n530, in_14, gm_n62, gm_n41, gm_n529, gm_n327);
	nand (gm_n531, gm_n530, gm_n528, gm_n526);
	nor (gm_n532, gm_n520, gm_n495, gm_n494, gm_n531, gm_n525);
	nand (gm_n533, gm_n79, gm_n64, in_4, gm_n114, in_7);
	nor (gm_n534, gm_n162, gm_n87, in_14, gm_n533);
	and (gm_n535, gm_n69, in_10, in_9, gm_n202, gm_n86);
	or (gm_n536, gm_n64, in_4, in_3, gm_n137, in_6);
	nor (gm_n537, gm_n119, in_14, gm_n42, gm_n536, gm_n418);
	nor (gm_n538, gm_n537, gm_n535, gm_n534);
	nor (gm_n539, gm_n69, in_13, gm_n41, gm_n434, gm_n216);
	nand (gm_n540, gm_n381, gm_n65, in_8);
	nor (gm_n541, in_14, gm_n42, in_9, gm_n540, gm_n271);
	nand (gm_n542, gm_n255, gm_n183, in_8);
	nor (gm_n543, gm_n69, gm_n42, in_9, gm_n542, gm_n108);
	nor (gm_n544, gm_n543, gm_n541, gm_n539);
	nand (gm_n545, gm_n532, gm_n493, gm_n491, gm_n544, gm_n538);
	nand (gm_n546, gm_n83, in_14, in_10, gm_n303);
	nor (gm_n547, gm_n150, gm_n41, gm_n45, gm_n261, gm_n95);
	nand (gm_n548, gm_n547, gm_n69, in_13);
	and (gm_n549, gm_n199, gm_n88, in_8);
	nand (gm_n550, in_14, in_13, in_12, gm_n549, gm_n349);
	nand (gm_n551, gm_n550, gm_n548, gm_n546);
	nand (gm_n552, gm_n101, in_14, in_10, gm_n138, gm_n322);
	nor (gm_n553, gm_n59, gm_n41, gm_n45, gm_n201, gm_n327);
	nand (gm_n554, gm_n553, in_14, in_13);
	and (gm_n555, gm_n246, gm_n183, in_8);
	nand (gm_n556, gm_n69, gm_n62, gm_n41, gm_n555, gm_n53);
	nand (gm_n557, gm_n556, gm_n554, gm_n552);
	nor (gm_n558, gm_n545, gm_n489, gm_n487, gm_n557, gm_n551);
	not (gm_n559, gm_n156);
	and (gm_n560, gm_n559, gm_n243, gm_n43, gm_n268, gm_n183);
	nor (gm_n561, in_14, in_10, gm_n70, gm_n434, gm_n84);
	not (gm_n562, gm_n116);
	nand (gm_n563, gm_n79, in_5, gm_n56, gm_n240, in_7);
	nor (gm_n564, gm_n562, gm_n77, gm_n43, gm_n563);
	nor (gm_n565, gm_n564, gm_n561, gm_n560);
	not (gm_n566, gm_n266);
	nor (gm_n567, gm_n241, gm_n229, gm_n43, gm_n566);
	nor (gm_n568, in_14, in_13, gm_n41, gm_n388, gm_n230);
	and (gm_n569, gm_n73, gm_n65, in_11, gm_n224, gm_n559);
	nor (gm_n570, gm_n569, gm_n568, gm_n567);
	nand (gm_n571, gm_n558, gm_n485, gm_n483, gm_n570, gm_n565);
	and (gm_n572, gm_n133, gm_n72, in_8);
	nand (gm_n573, in_14, in_13, gm_n41, gm_n572, gm_n93);
	nand (gm_n574, gm_n69, in_13, in_12, gm_n492, gm_n44);
	nor (gm_n575, gm_n90, gm_n150, gm_n45);
	nand (gm_n576, gm_n69, gm_n42, gm_n70, gm_n575, gm_n178);
	nand (gm_n577, gm_n576, gm_n574, gm_n573);
	nand (gm_n578, gm_n349, gm_n46, gm_n45, gm_n255, gm_n168);
	and (gm_n579, gm_n183, gm_n129, gm_n45);
	nand (gm_n580, in_14, gm_n62, in_12, gm_n579, gm_n93);
	nor (gm_n581, gm_n208, gm_n90, gm_n45);
	nand (gm_n582, gm_n69, in_13, in_12, gm_n581, gm_n93);
	nand (gm_n583, gm_n582, gm_n580, gm_n578);
	nor (gm_n584, gm_n571, gm_n482, gm_n481, gm_n583, gm_n577);
	and (gm_n585, gm_n164, gm_n88, in_11, gm_n233, gm_n170);
	and (gm_n586, gm_n161, gm_n73, gm_n45);
	and (gm_n587, in_14, gm_n42, in_9, gm_n586, gm_n178);
	nor (gm_n588, gm_n219, gm_n59, in_8);
	and (gm_n589, gm_n69, in_13, in_12, gm_n588, gm_n93);
	nor (gm_n590, gm_n589, gm_n587, gm_n585);
	nand (gm_n591, gm_n246, gm_n80, in_8);
	nor (gm_n592, in_14, gm_n62, in_12, gm_n591, gm_n71);
	nand (gm_n593, gm_n79, in_5, in_4, gm_n114, in_7);
	nor (gm_n594, gm_n516, gm_n249, gm_n43, gm_n593);
	nand (gm_n595, gm_n170, gm_n161, in_8);
	nor (gm_n596, gm_n69, in_10, in_9, gm_n595, gm_n271);
	nor (gm_n597, gm_n596, gm_n594, gm_n592);
	nand (gm_n598, gm_n584, gm_n479, gm_n477, gm_n597, gm_n590);
	nor (gm_n599, gm_n301, gm_n89, in_8);
	nand (gm_n600, in_14, gm_n62, gm_n41, gm_n599, gm_n126);
	nor (gm_n601, gm_n147, gm_n59, in_8);
	nand (gm_n602, in_14, in_13, gm_n41, gm_n601, gm_n126);
	nand (gm_n603, gm_n88, gm_n66, gm_n43, gm_n117, gm_n116);
	nand (gm_n604, gm_n603, gm_n602, gm_n600);
	nor (gm_n605, gm_n42, gm_n70, in_8, gm_n208, gm_n95);
	nand (gm_n606, gm_n605, gm_n245, gm_n69);
	and (gm_n607, gm_n170, gm_n41, in_8, gm_n191, gm_n183);
	nand (gm_n608, gm_n607, in_14, gm_n62);
	nand (gm_n609, gm_n80, gm_n370, gm_n45);
	or (gm_n610, in_14, in_13, in_12, gm_n609, gm_n76);
	nand (gm_n611, gm_n610, gm_n608, gm_n606);
	nor (gm_n612, gm_n598, gm_n476, gm_n475, gm_n611, gm_n604);
	and (gm_n613, gm_n83, gm_n65, gm_n69, gm_n266, gm_n381);
	nor (gm_n614, gm_n119, in_14, in_10, gm_n287, gm_n145);
	nand (gm_n615, gm_n129, gm_n79, in_5);
	nor (gm_n616, gm_n84, in_14, in_10, gm_n615, gm_n307);
	nor (gm_n617, gm_n616, gm_n614, gm_n613);
	and (gm_n618, in_14, in_10, in_9, gm_n527, gm_n345);
	nor (gm_n619, in_14, in_13, gm_n41, gm_n366, gm_n63);
	and (gm_n620, gm_n268, gm_n109, gm_n45);
	and (gm_n621, gm_n69, in_13, in_12, gm_n620, gm_n53);
	nor (gm_n622, gm_n621, gm_n619, gm_n618);
	nand (gm_n623, gm_n612, gm_n473, gm_n472, gm_n622, gm_n617);
	and (gm_n624, gm_n277, gm_n80, in_8);
	nand (gm_n625, gm_n69, in_13, gm_n41, gm_n624, gm_n349);
	nand (gm_n626, gm_n110, gm_n72, in_8);
	or (gm_n627, gm_n69, gm_n62, gm_n41, gm_n626, gm_n76);
	or (gm_n628, gm_n58, in_6, gm_n64, gm_n189, gm_n45);
	or (gm_n629, gm_n69, in_13, gm_n41, gm_n628, gm_n327);
	nand (gm_n630, gm_n629, gm_n627, gm_n625);
	and (gm_n631, in_6, in_5, gm_n56, gm_n240, in_7);
	nand (gm_n632, gm_n233, gm_n224, gm_n43, gm_n631);
	nand (gm_n633, gm_n161, gm_n243, in_11, gm_n129, gm_n116);
	nand (gm_n634, in_14, gm_n62, in_12, gm_n397, gm_n131);
	nand (gm_n635, gm_n634, gm_n633, gm_n632);
	nor (gm_n636, gm_n623, gm_n470, gm_n468, gm_n635, gm_n630);
	or (gm_n637, gm_n193, gm_n150, gm_n45);
	or (gm_n638, in_14, gm_n42, gm_n70, gm_n637, gm_n108);
	or (gm_n639, in_7, gm_n79, gm_n64, gm_n189, gm_n45);
	or (gm_n640, gm_n69, gm_n42, gm_n70, gm_n639, gm_n108);
	and (gm_n641, gm_n640, gm_n638, t_4);
	nand (gm_n642, gm_n66, gm_n109, in_8);
	nor (gm_n643, in_14, gm_n62, gm_n41, gm_n642, gm_n327);
	or (gm_n644, gm_n227, gm_n351, in_8);
	nor (gm_n645, gm_n69, gm_n62, in_12, gm_n644, gm_n216);
	nand (gm_n646, gm_n42, in_9, in_8);
	nor (gm_n647, gm_n646, gm_n77, gm_n43, gm_n593);
	nor (gm_n648, gm_n647, gm_n645, gm_n643);
	nand (gm_n649, gm_n636, gm_n466, gm_n464, gm_n648, gm_n641);
	nand (gm_n650, gm_n88, gm_n243, in_8, gm_n246, gm_n98);
	and (gm_n651, gm_n80, gm_n73, in_8);
	nand (gm_n652, gm_n69, gm_n62, in_12, gm_n651, gm_n191);
	nand (gm_n653, gm_n349, gm_n109, gm_n45, gm_n255, gm_n168);
	nand (gm_n654, gm_n653, gm_n652, gm_n650);
	and (gm_n655, gm_n79, gm_n64, gm_n56, gm_n240, gm_n58);
	nand (gm_n656, gm_n295, gm_n116, gm_n43, gm_n655);
	nor (gm_n657, gm_n90, in_12, in_8, gm_n208, gm_n342);
	nand (gm_n658, gm_n657, in_14, gm_n62);
	or (gm_n659, gm_n69, gm_n62, gm_n41, gm_n628, gm_n230);
	nand (gm_n660, gm_n659, gm_n658, gm_n656);
	nor (out_2, gm_n654, gm_n649, gm_n463, gm_n660);
	nor (gm_n662, gm_n69, in_10, gm_n70, gm_n446, gm_n119);
	nor (gm_n663, in_14, in_13, gm_n41, gm_n474, gm_n216);
	nor (gm_n664, gm_n90, gm_n89, in_8);
	nand (gm_n665, in_14, gm_n62, gm_n41, gm_n664, gm_n191);
	and (gm_n666, gm_n93, gm_n88, gm_n45, gm_n174, gm_n170);
	nor (gm_n667, gm_n122, in_14, in_10, gm_n305, gm_n271);
	nor (gm_n668, gm_n351, gm_n57, in_8);
	nand (gm_n669, gm_n69, in_13, gm_n41, gm_n668, gm_n349);
	nor (gm_n670, gm_n227, gm_n150, gm_n45);
	nand (gm_n671, in_14, gm_n62, gm_n41, gm_n670, gm_n53);
	and (gm_n672, in_14, in_13, in_12, gm_n579, gm_n53);
	and (gm_n673, gm_n69, in_13, in_12, gm_n394, gm_n349);
	nand (gm_n674, gm_n245, gm_n116, in_14, gm_n199, gm_n183);
	or (gm_n675, gm_n327, gm_n385, in_8, gm_n229, gm_n147);
	nand (gm_n676, gm_n69, in_13, in_12, gm_n575, gm_n349);
	nor (gm_n677, gm_n95, gm_n150, in_8);
	nand (gm_n678, in_14, gm_n62, in_12, gm_n677, gm_n191);
	nor (gm_n679, in_10, gm_n70, in_8, gm_n193, gm_n150);
	nand (gm_n680, gm_n679, gm_n345, in_14);
	and (gm_n681, gm_n199, gm_n65, in_8);
	nand (gm_n682, in_14, in_13, in_12, gm_n681, gm_n126);
	and (gm_n683, gm_n678, gm_n676, t_3, gm_n682, gm_n680);
	nor (gm_n684, gm_n122, gm_n69, gm_n42, gm_n287, gm_n177);
	nand (gm_n685, gm_n80, in_12, gm_n45, gm_n129, gm_n98);
	nor (gm_n686, gm_n685, in_14, in_13);
	nand (gm_n687, gm_n199, gm_n46, gm_n45);
	nor (gm_n688, in_14, gm_n62, gm_n41, gm_n687, gm_n216);
	nor (gm_n689, gm_n688, gm_n686, gm_n684);
	and (gm_n690, in_14, in_10, in_9, gm_n345, gm_n130);
	nor (gm_n691, gm_n396, gm_n385, gm_n45);
	and (gm_n692, gm_n69, gm_n62, gm_n41, gm_n691, gm_n93);
	nand (gm_n693, gm_n105, gm_n109, in_8);
	nor (gm_n694, gm_n69, gm_n62, gm_n41, gm_n693, gm_n327);
	nor (gm_n695, gm_n694, gm_n692, gm_n690);
	nand (gm_n696, gm_n683, gm_n675, gm_n674, gm_n695, gm_n689);
	and (gm_n697, gm_n174, gm_n109, gm_n45, gm_n381, gm_n191);
	and (gm_n698, gm_n178, gm_n69, gm_n42, gm_n323, gm_n289);
	or (gm_n699, gm_n698, gm_n697, t_0);
	nand (gm_n700, gm_n93, gm_n109, in_8, gm_n295, gm_n255);
	nand (gm_n701, gm_n183, gm_n158, gm_n45);
	or (gm_n702, in_14, gm_n62, in_12, gm_n701, gm_n76);
	or (gm_n703, gm_n95, gm_n351, gm_n69, gm_n417, gm_n249);
	nand (gm_n704, gm_n703, gm_n702, gm_n700);
	nor (gm_n705, gm_n696, gm_n673, gm_n672, gm_n704, gm_n699);
	nand (gm_n706, gm_n88, gm_n41, gm_n45, gm_n184, gm_n93);
	nor (gm_n707, gm_n706, in_14, gm_n62);
	nand (gm_n708, in_6, in_5, in_4, gm_n114, in_7);
	nor (gm_n709, gm_n229, gm_n156, in_11, gm_n708);
	or (gm_n710, gm_n385, in_12, in_8, gm_n227, gm_n216);
	nor (gm_n711, gm_n710, in_14, in_13);
	nor (gm_n712, gm_n711, gm_n709, gm_n707);
	nor (gm_n713, gm_n145, gm_n69, gm_n42, gm_n536, gm_n177);
	nor (gm_n714, in_14, gm_n42, gm_n70, gm_n87, gm_n82);
	nand (gm_n715, gm_n199, gm_n80, gm_n45);
	nor (gm_n716, gm_n69, in_10, gm_n70, gm_n715, gm_n271);
	nor (gm_n717, gm_n716, gm_n714, gm_n713);
	nand (gm_n718, gm_n705, gm_n671, gm_n669, gm_n717, gm_n712);
	or (gm_n719, in_14, in_10, in_9, gm_n119, gm_n67);
	nor (gm_n720, gm_n54, in_1, gm_n48, in_4, gm_n55);
	nand (gm_n721, gm_n720, gm_n72, in_8);
	or (gm_n722, in_14, gm_n62, in_12, gm_n721, gm_n76);
	nand (gm_n723, gm_n126, gm_n161, in_8, gm_n295, gm_n268);
	nand (gm_n724, gm_n723, gm_n722, gm_n719);
	nor (gm_n725, gm_n231, gm_n94, in_8);
	nand (gm_n726, in_14, in_13, gm_n41, gm_n725, gm_n126);
	nand (gm_n727, gm_n83, gm_n65, gm_n69, gm_n246, gm_n559);
	or (gm_n728, gm_n239, gm_n69, gm_n42, gm_n536, gm_n286);
	nand (gm_n729, gm_n728, gm_n727, gm_n726);
	nor (gm_n730, gm_n718, gm_n667, gm_n666, gm_n729, gm_n724);
	nand (gm_n731, gm_n69, gm_n62, in_12, gm_n488, gm_n349);
	and (gm_n732, gm_n246, gm_n80, gm_n45);
	nand (gm_n733, in_14, in_13, gm_n41, gm_n732, gm_n191);
	or (gm_n734, gm_n122, in_14, in_10, gm_n419, gm_n177);
	nand (gm_n735, gm_n731, gm_n730, gm_n665, gm_n734, gm_n733);
	nand (gm_n736, gm_n80, gm_n44, in_8, gm_n174, gm_n81);
	nand (gm_n737, gm_n116, gm_n109, gm_n43, gm_n295, gm_n124);
	nor (gm_n738, gm_n71, gm_n41, gm_n45, gm_n351, gm_n57);
	nand (gm_n739, gm_n738, gm_n69, in_13);
	nand (gm_n740, gm_n739, gm_n737, gm_n736);
	nor (gm_n741, in_9, in_8, gm_n58);
	and (gm_n742, gm_n83, gm_n69, gm_n42, gm_n741, gm_n258);
	nor (out_3, gm_n735, gm_n663, gm_n662, gm_n742, gm_n740);
	nor (gm_n744, gm_n69, in_10, gm_n70, gm_n591, gm_n239);
	or (gm_n745, gm_n150, gm_n57, gm_n69, gm_n646, gm_n87);
	nor (gm_n746, gm_n95, gm_n385, in_8);
	nand (gm_n747, in_14, gm_n62, gm_n41, gm_n746, gm_n191);
	and (gm_n748, gm_n58, gm_n79, in_5, gm_n124, gm_n45);
	and (gm_n749, in_14, gm_n62, in_12, gm_n748, gm_n191);
	and (gm_n750, in_14, gm_n62, in_12, gm_n204, gm_n349);
	or (gm_n751, gm_n280, gm_n94, gm_n69, gm_n156, gm_n119);
	nand (gm_n752, in_14, gm_n62, gm_n41, gm_n572, gm_n44);
	and (gm_n753, gm_n129, gm_n161, gm_n43, gm_n224, gm_n169);
	and (gm_n754, gm_n93, gm_n243, gm_n45, gm_n255, gm_n161);
	not (gm_n755, t_2);
	nand (gm_n756, gm_n136, in_14, in_10, gm_n329, gm_n212);
	nor (gm_n757, in_7, in_6, gm_n64, gm_n189, in_8);
	nor (gm_n758, in_12, in_11, gm_n42);
	nand (gm_n759, in_14, in_13, in_9, gm_n758, gm_n757);
	and (gm_n760, gm_n277, gm_n65, gm_n45);
	nand (gm_n761, in_14, in_13, gm_n41, gm_n760, gm_n191);
	nor (gm_n762, gm_n396, gm_n150, in_8);
	nand (gm_n763, in_14, in_13, gm_n41, gm_n762, gm_n349);
	nand (gm_n764, gm_n759, gm_n756, gm_n755, gm_n763, gm_n761);
	nand (gm_n765, in_14, in_13, in_12, gm_n624, gm_n44);
	or (gm_n766, gm_n177, in_14, gm_n42, gm_n615, gm_n307);
	and (gm_n767, gm_n183, gm_n133, gm_n45);
	nand (gm_n768, in_14, in_13, in_12, gm_n767, gm_n53);
	nand (gm_n769, gm_n768, gm_n766, gm_n765);
	nand (gm_n770, gm_n255, gm_n80, gm_n45);
	or (gm_n771, gm_n69, in_13, gm_n41, gm_n770, gm_n342);
	nand (gm_n772, in_14, in_13, in_12, gm_n488, gm_n349);
	nor (gm_n773, gm_n94, gm_n50, gm_n45);
	nand (gm_n774, gm_n69, in_13, in_12, gm_n773, gm_n53);
	nand (gm_n775, gm_n774, gm_n772, gm_n771);
	nor (gm_n776, gm_n764, gm_n754, gm_n753, gm_n775, gm_n769);
	and (gm_n777, gm_n116, gm_n86, in_14, gm_n631);
	and (gm_n778, gm_n86, gm_n69, in_10, gm_n323, gm_n289);
	and (gm_n779, gm_n136, in_14, gm_n42, gm_n346, gm_n289);
	nor (gm_n780, gm_n779, gm_n778, gm_n777);
	nor (gm_n781, gm_n90, gm_n385, gm_n43, gm_n226, gm_n225);
	not (gm_n782, gm_n233);
	nor (gm_n783, gm_n150, gm_n57, gm_n69, gm_n782, gm_n177);
	and (gm_n784, in_10, in_9, in_8, gm_n88, gm_n370);
	and (gm_n785, gm_n784, gm_n178, in_14);
	nor (gm_n786, gm_n785, gm_n783, gm_n781);
	nand (gm_n787, gm_n776, gm_n752, gm_n751, gm_n786, gm_n780);
	nand (gm_n788, gm_n183, gm_n169, gm_n69, gm_n345, gm_n199);
	nand (gm_n789, gm_n106, gm_n88, gm_n43, gm_n246, gm_n224);
	or (gm_n790, in_5, in_4, in_3, gm_n137, in_6);
	or (gm_n791, gm_n417, gm_n69, in_10, gm_n790, gm_n145);
	nand (gm_n792, gm_n791, gm_n789, gm_n788);
	nand (gm_n793, gm_n98, gm_n46, in_8, gm_n295, gm_n184);
	and (gm_n794, gm_n44, gm_n41, in_8, gm_n170, gm_n65);
	nand (gm_n795, gm_n794, in_14, in_13);
	nand (gm_n796, gm_n284, gm_n46, in_11, gm_n295, gm_n268);
	nand (gm_n797, gm_n796, gm_n795, gm_n793);
	nor (gm_n798, gm_n787, gm_n750, gm_n749, gm_n797, gm_n792);
	nor (gm_n799, in_7, in_6, in_5, gm_n189, in_8);
	and (gm_n800, gm_n799, gm_n174, gm_n53);
	nor (gm_n801, in_14, in_13, gm_n41, gm_n591, gm_n63);
	nor (gm_n802, gm_n516, gm_n156, gm_n43, gm_n563);
	nor (gm_n803, gm_n802, gm_n801, gm_n800);
	and (gm_n804, gm_n69, gm_n62, in_12, gm_n194, gm_n44);
	nor (gm_n805, gm_n122, gm_n69, in_10, gm_n790, gm_n417);
	nand (gm_n806, gm_n199, gm_n72, in_8);
	nor (gm_n807, in_14, in_13, in_12, gm_n806, gm_n76);
	nor (gm_n808, gm_n807, gm_n805, gm_n804);
	nand (gm_n809, gm_n798, gm_n747, gm_n745, gm_n808, gm_n803);
	not (gm_n810, gm_n503);
	nand (gm_n811, gm_n233, gm_n104, in_11, gm_n810);
	nand (gm_n812, in_14, gm_n62, in_12, gm_n459, gm_n126);
	nand (gm_n813, gm_n88, gm_n81, gm_n69, gm_n163, gm_n245);
	nand (gm_n814, gm_n813, gm_n812, gm_n811);
	and (gm_n815, in_14, in_13, gm_n41, gm_n732, gm_n131);
	nor (gm_n816, gm_n193, gm_n385, in_8);
	and (gm_n817, gm_n69, in_13, in_12, gm_n816, gm_n98);
	or (gm_n818, gm_n817, gm_n815, t_9);
	nor (out_4, gm_n814, gm_n809, gm_n744, gm_n818);
	nand (gm_n820, gm_n184, gm_n183, in_8);
	nor (gm_n821, gm_n69, in_13, gm_n41, gm_n820, gm_n342);
	nand (gm_n822, gm_n340, gm_n117, gm_n93);
	nor (gm_n823, in_7, in_6, in_5, gm_n189, gm_n45);
	nand (gm_n824, gm_n69, in_13, gm_n41, gm_n823, gm_n44);
	and (gm_n825, gm_n83, gm_n69, in_10, gm_n741, gm_n323);
	nor (gm_n826, gm_n108, in_14, gm_n42, gm_n305, gm_n302);
	not (gm_n827, gm_n174);
	nor (gm_n828, gm_n827, gm_n646, in_11, gm_n533);
	nor (gm_n829, gm_n231, gm_n89, in_8);
	and (gm_n830, in_14, gm_n62, in_12, gm_n829, gm_n44);
	nor (gm_n831, in_7, gm_n79, in_5, gm_n189, in_8);
	and (gm_n832, gm_n69, gm_n62, in_12, gm_n831, gm_n131);
	nor (gm_n833, gm_n271, gm_n69, gm_n42, gm_n302, gm_n287);
	or (gm_n834, gm_n830, gm_n828, t_7, gm_n833, gm_n832);
	nand (gm_n835, gm_n277, gm_n65, in_8);
	or (gm_n836, gm_n69, gm_n42, gm_n70, gm_n835, gm_n417);
	nand (gm_n837, gm_n83, in_14, gm_n42, gm_n741, gm_n258);
	nand (gm_n838, gm_n69, in_13, gm_n41, gm_n185, gm_n126);
	nand (gm_n839, gm_n838, gm_n837, gm_n836);
	nor (gm_n840, in_5, in_4, gm_n55, gm_n120, gm_n79);
	nand (gm_n841, gm_n178, in_14, in_10, gm_n840, gm_n212);
	and (gm_n842, gm_n161, in_12, in_8, gm_n274, gm_n191);
	nand (gm_n843, gm_n842, in_14, in_13);
	nand (gm_n844, in_7, in_6, gm_n64, gm_n124, in_8);
	or (gm_n845, in_14, gm_n62, gm_n41, gm_n844, gm_n342);
	nand (gm_n846, gm_n845, gm_n843, gm_n841);
	nor (gm_n847, gm_n834, gm_n826, gm_n825, gm_n846, gm_n839);
	and (gm_n848, gm_n106, gm_n109, gm_n43, gm_n164, gm_n124);
	and (gm_n849, gm_n168, gm_n133, in_8, gm_n191, gm_n183);
	nor (gm_n850, gm_n69, gm_n42, in_9, gm_n820, gm_n417);
	nor (gm_n851, gm_n850, gm_n849, gm_n848);
	and (gm_n852, gm_n243, gm_n65, in_11, gm_n559, gm_n81);
	and (gm_n853, gm_n174, gm_n559, gm_n43, gm_n253);
	and (gm_n854, gm_n116, gm_n161, gm_n43, gm_n295, gm_n158);
	nor (gm_n855, gm_n854, gm_n853, gm_n852);
	nand (gm_n856, gm_n847, gm_n824, gm_n822, gm_n855, gm_n851);
	nand (gm_n857, in_14, in_13, in_12, gm_n748, gm_n53);
	nand (gm_n858, gm_n110, gm_n46, gm_n45, gm_n224, gm_n126);
	nand (gm_n859, gm_n80, gm_n53, gm_n45, gm_n224, gm_n133);
	nand (gm_n860, gm_n859, gm_n858, gm_n857);
	nand (gm_n861, gm_n133, gm_n65, in_11, gm_n266, gm_n224);
	nand (gm_n862, gm_n93, gm_n88, gm_n45, gm_n170, gm_n117);
	and (gm_n863, gm_n46, gm_n41, gm_n45, gm_n131, gm_n81);
	nand (gm_n864, gm_n863, gm_n69, gm_n62);
	nand (gm_n865, gm_n864, gm_n862, gm_n861);
	nor (out_5, gm_n860, gm_n856, gm_n821, gm_n865);
	nand (gm_n867, gm_n274, gm_n80, in_8);
	nor (gm_n868, gm_n69, in_13, gm_n41, gm_n867, gm_n71);
	nand (gm_n869, in_14, in_13, in_12, gm_n278, gm_n53);
	or (gm_n870, gm_n467, gm_n69, gm_n42, gm_n305, gm_n239);
	or (gm_n871, gm_n227, gm_n47, in_8);
	nor (gm_n872, gm_n69, in_13, gm_n41, gm_n871, gm_n327);
	and (gm_n873, gm_n163, gm_n243, in_11, gm_n373);
	or (gm_n874, gm_n269, gm_n417, gm_n69);
	nand (gm_n875, gm_n83, in_14, gm_n42, gm_n329, gm_n289);
	nor (gm_n876, gm_n229, gm_n351, gm_n43, gm_n782, gm_n201);
	and (gm_n877, gm_n105, gm_n104, in_11, gm_n266, gm_n183);
	nand (gm_n878, gm_n93, gm_n46, gm_n45, gm_n274, gm_n224);
	nand (gm_n879, gm_n69, gm_n62, in_12, gm_n664, gm_n44);
	and (gm_n880, gm_n69, gm_n62, gm_n41, gm_n403, gm_n44);
	nor (gm_n881, gm_n119, in_14, gm_n42, gm_n536, gm_n467);
	not (gm_n882, gm_n168);
	or (gm_n883, gm_n882, gm_n156, in_11, gm_n593);
	and (gm_n884, gm_n81, gm_n46, in_8);
	nand (gm_n885, in_14, gm_n62, gm_n41, gm_n884, gm_n191);
	nor (gm_n886, gm_n511, gm_n239, gm_n69);
	nor (gm_n887, in_14, in_13, in_12, gm_n111, gm_n76);
	nand (gm_n888, gm_n83, in_14, gm_n42, gm_n741, gm_n323);
	nand (gm_n889, in_14, gm_n62, gm_n41, gm_n588, gm_n98);
	nor (gm_n890, in_14, in_13, gm_n41, gm_n529, gm_n63);
	and (gm_n891, gm_n126, gm_n72, in_8, gm_n164, gm_n133);
	nand (gm_n892, gm_n164, gm_n80, gm_n43, gm_n255, gm_n169);
	nand (gm_n893, gm_n320, gm_n65, gm_n45, gm_n295, gm_n98);
	nor (gm_n894, gm_n108, gm_n69, gm_n42, gm_n237, gm_n467);
	nor (gm_n895, gm_n385, gm_n76, in_8, gm_n95, gm_n77);
	and (gm_n896, gm_n93, gm_n80, in_8, gm_n199, gm_n174);
	nor (gm_n897, in_14, in_10, gm_n70, gm_n521, gm_n108);
	and (gm_n898, gm_n80, gm_n44, gm_n45, gm_n164, gm_n133);
	nor (gm_n899, gm_n896, gm_n895, gm_n894, gm_n898, gm_n897);
	nor (gm_n900, in_14, in_10, gm_n70, gm_n500, gm_n108);
	nand (gm_n901, gm_n158, gm_n80, in_8);
	nor (gm_n902, in_14, gm_n62, gm_n41, gm_n901, gm_n216);
	nand (gm_n903, gm_n80, gm_n41, gm_n45, gm_n191, gm_n105);
	nor (gm_n904, gm_n903, gm_n69, in_13);
	nor (gm_n905, gm_n904, gm_n902, gm_n900);
	or (gm_n906, in_10, gm_n70, gm_n45, gm_n189, gm_n150);
	nor (gm_n907, gm_n906, gm_n108, in_14);
	or (gm_n908, gm_n227, gm_n351, gm_n45);
	nor (gm_n909, in_14, in_13, gm_n41, gm_n908, gm_n342);
	and (gm_n910, gm_n199, gm_n88, gm_n45);
	and (gm_n911, gm_n69, in_13, in_12, gm_n910, gm_n53);
	nor (gm_n912, gm_n911, gm_n909, gm_n907);
	nand (gm_n913, gm_n899, gm_n893, gm_n892, gm_n912, gm_n905);
	nand (gm_n914, gm_n136, in_14, in_10, gm_n346, gm_n139);
	nor (gm_n915, gm_n89, gm_n41, in_8, gm_n227, gm_n216);
	nand (gm_n916, gm_n915, gm_n69, in_13);
	not (gm_n917, gm_n302);
	nand (gm_n918, gm_n101, in_14, gm_n42, gm_n329, gm_n917);
	nand (gm_n919, gm_n918, gm_n916, gm_n914);
	nand (gm_n920, gm_n69, gm_n62, in_12, gm_n98, gm_n60);
	nand (gm_n921, gm_n170, gm_n109, in_14, gm_n266, gm_n300);
	and (gm_n922, gm_n184, gm_n65, in_8);
	nand (gm_n923, gm_n69, gm_n62, gm_n41, gm_n922, gm_n191);
	nand (gm_n924, gm_n923, gm_n921, gm_n920);
	nor (gm_n925, gm_n913, gm_n891, gm_n890, gm_n924, gm_n919);
	nand (gm_n926, gm_n183, gm_n110, in_8);
	nor (gm_n927, gm_n69, gm_n62, gm_n41, gm_n926, gm_n63);
	and (gm_n928, in_14, gm_n62, in_12, gm_n278, gm_n44);
	and (gm_n929, gm_n233, gm_n117, gm_n43, gm_n631);
	nor (gm_n930, gm_n929, gm_n928, gm_n927);
	nor (gm_n931, gm_n69, gm_n62, in_12, gm_n542, gm_n230);
	nor (gm_n932, gm_n69, gm_n62, in_12, gm_n364, gm_n216);
	nand (gm_n933, gm_n81, gm_n41, in_8, gm_n183, gm_n126);
	nor (gm_n934, gm_n933, in_14, gm_n62);
	nor (gm_n935, gm_n934, gm_n932, gm_n931);
	nand (gm_n936, gm_n925, gm_n889, gm_n888, gm_n935, gm_n930);
	and (gm_n937, in_6, gm_n64, gm_n56, gm_n240);
	nand (gm_n938, gm_n117, in_11, gm_n58, gm_n937, gm_n559);
	or (gm_n939, gm_n108, in_14, in_10, gm_n286, gm_n121);
	nand (gm_n940, gm_n349, gm_n46, gm_n45, gm_n255, gm_n243);
	nand (gm_n941, gm_n940, gm_n939, gm_n938);
	or (gm_n942, gm_n69, gm_n62, gm_n41, gm_n591, gm_n63);
	not (gm_n943, gm_n307);
	nand (gm_n944, gm_n245, in_14, gm_n42, gm_n943, gm_n258);
	nand (gm_n945, gm_n131, gm_n243, in_8, gm_n246, gm_n183);
	nand (gm_n946, gm_n945, gm_n944, gm_n942);
	nor (gm_n947, gm_n936, gm_n887, gm_n886, gm_n946, gm_n941);
	and (gm_n948, gm_n104, gm_n109, gm_n43, gm_n246, gm_n116);
	and (gm_n949, in_14, in_10, in_9, gm_n101, gm_n99);
	nor (gm_n950, gm_n949, gm_n948, gm_n504);
	nor (gm_n951, gm_n69, in_13, in_12, gm_n835, gm_n71);
	nor (gm_n952, in_14, gm_n62, gm_n41, gm_n595, gm_n76);
	and (gm_n953, gm_n170, gm_n98, gm_n45, gm_n295, gm_n183);
	nor (gm_n954, gm_n953, gm_n952, gm_n951);
	nand (gm_n955, gm_n947, gm_n885, gm_n883, gm_n954, gm_n950);
	nand (gm_n956, gm_n133, gm_n161, gm_n43, gm_n174, gm_n163);
	nand (gm_n957, in_14, in_13, in_12, gm_n130, gm_n93);
	nand (gm_n958, in_14, gm_n62, in_12, gm_n191, gm_n179);
	nand (gm_n959, gm_n958, gm_n957, gm_n956);
	nor (gm_n960, gm_n76, gm_n41, in_8, gm_n90, gm_n150);
	nand (gm_n961, gm_n960, gm_n69, in_13);
	nand (gm_n962, gm_n69, gm_n42, gm_n70, gm_n125, gm_n245);
	not (gm_n963, gm_n117);
	or (gm_n964, gm_n226, gm_n963, gm_n43, gm_n533);
	nand (gm_n965, gm_n964, gm_n962, gm_n961);
	nor (gm_n966, gm_n955, gm_n881, gm_n880, gm_n965, gm_n959);
	nor (gm_n967, in_14, in_13, gm_n41, gm_n67, gm_n63);
	nand (gm_n968, in_7, gm_n79, in_5, gm_n124, in_8);
	nor (gm_n969, gm_n69, in_13, in_12, gm_n968, gm_n63);
	nor (gm_n970, gm_n150, gm_n57, in_11, gm_n566, gm_n827);
	nor (gm_n971, gm_n970, gm_n969, gm_n967);
	nor (gm_n972, gm_n84, gm_n69, in_10, gm_n307, gm_n237);
	and (gm_n973, gm_n105, gm_n46, in_8);
	and (gm_n974, gm_n69, gm_n62, gm_n41, gm_n973, gm_n98);
	and (gm_n975, gm_n320, gm_n109, gm_n43, gm_n168, gm_n116);
	nor (gm_n976, gm_n975, gm_n974, gm_n972);
	nand (gm_n977, gm_n966, gm_n879, gm_n878, gm_n976, gm_n971);
	nand (gm_n978, in_14, gm_n62, in_12, gm_n829, gm_n349);
	nand (gm_n979, gm_n106, gm_n65, gm_n43, gm_n295, gm_n255);
	nand (gm_n980, in_14, in_13, in_12, gm_n394, gm_n93);
	nand (gm_n981, gm_n980, gm_n979, gm_n978);
	nand (gm_n982, in_14, gm_n42, gm_n70, gm_n575, gm_n345);
	nand (gm_n983, in_14, in_10, gm_n70, gm_n586, gm_n345);
	nand (gm_n984, gm_n109, gm_n44, gm_n45, gm_n199, gm_n117);
	nand (gm_n985, gm_n984, gm_n983, gm_n982);
	nor (gm_n986, gm_n977, gm_n877, gm_n876, gm_n985, gm_n981);
	nand (gm_n987, gm_n110, gm_n80, in_8);
	nor (gm_n988, gm_n69, in_13, in_12, gm_n987, gm_n76);
	and (gm_n989, gm_n174, gm_n80, gm_n43, gm_n266, gm_n381);
	or (gm_n990, gm_n219, in_6, in_5, gm_n122);
	nor (gm_n991, gm_n239, in_14, in_10, gm_n990);
	nor (gm_n992, gm_n991, gm_n989, gm_n988);
	and (gm_n993, gm_n115, gm_n106, in_11, gm_n174);
	nor (gm_n994, gm_n119, gm_n69, in_10, gm_n302, gm_n143);
	or (gm_n995, gm_n59, gm_n41, gm_n45, gm_n227, gm_n327);
	nor (gm_n996, gm_n995, gm_n69, in_13);
	nor (gm_n997, gm_n996, gm_n994, gm_n993);
	nand (gm_n998, gm_n986, gm_n875, gm_n874, gm_n997, gm_n992);
	nand (gm_n999, gm_n69, gm_n62, gm_n41, gm_n471, gm_n53);
	and (gm_n1000, gm_n246, gm_n65, gm_n45);
	nand (gm_n1001, gm_n69, gm_n62, gm_n41, gm_n1000, gm_n93);
	and (gm_n1002, gm_n80, gm_n41, gm_n45, gm_n191, gm_n81);
	nand (gm_n1003, gm_n1002, gm_n69, in_13);
	nand (gm_n1004, gm_n1003, gm_n1001, gm_n999);
	nand (gm_n1005, gm_n101, in_14, gm_n42, gm_n346, gm_n144);
	nand (gm_n1006, in_14, in_13, in_12, gm_n96, gm_n53);
	and (gm_n1007, gm_n349, in_12, gm_n45, gm_n133, gm_n72);
	nand (gm_n1008, gm_n1007, in_14, gm_n62);
	nand (gm_n1009, gm_n1008, gm_n1006, gm_n1005);
	nor (gm_n1010, gm_n998, gm_n873, gm_n872, gm_n1009, gm_n1004);
	nor (gm_n1011, gm_n417, in_14, in_10, gm_n419, gm_n145);
	nor (gm_n1012, gm_n827, gm_n562, in_11, gm_n708);
	and (gm_n1013, gm_n93, gm_n109, in_8, gm_n255, gm_n117);
	nor (gm_n1014, gm_n1013, gm_n1012, gm_n1011);
	nor (gm_n1015, gm_n229, gm_n342, in_8, gm_n208, gm_n396);
	nor (gm_n1016, in_14, gm_n62, gm_n41, gm_n926, gm_n261);
	nor (gm_n1017, gm_n69, gm_n42, gm_n70, gm_n835, gm_n119);
	nor (gm_n1018, gm_n1017, gm_n1016, gm_n1015);
	nand (gm_n1019, gm_n1010, gm_n870, gm_n869, gm_n1018, gm_n1014);
	or (gm_n1020, in_14, in_10, in_9, gm_n871, gm_n87);
	nor (gm_n1021, gm_n208, gm_n280, in_8);
	nand (gm_n1022, gm_n69, in_13, in_12, gm_n1021, gm_n93);
	or (gm_n1023, gm_n261, gm_n150, gm_n45, gm_n193, gm_n882);
	nand (gm_n1024, gm_n1023, gm_n1022, gm_n1020);
	or (gm_n1025, gm_n119, gm_n69, in_10, gm_n467, gm_n121);
	or (gm_n1026, gm_n90, gm_n385, in_14, gm_n119, gm_n249);
	and (gm_n1027, gm_n46, gm_n41, gm_n45, gm_n274, gm_n98);
	nand (gm_n1028, gm_n1027, in_14, gm_n62);
	nand (gm_n1029, gm_n1028, gm_n1026, gm_n1025);
	nor (out_6, gm_n1024, gm_n1019, gm_n868, gm_n1029);
	nor (gm_n1031, gm_n69, in_13, gm_n41, gm_n693, gm_n261);
	nand (gm_n1032, gm_n101, gm_n69, in_10, gm_n741, gm_n138);
	nor (gm_n1033, gm_n69, in_13, gm_n41, gm_n446, gm_n216);
	and (gm_n1034, in_10, in_9, in_8, gm_n274, gm_n80);
	and (gm_n1035, gm_n1034, gm_n83, gm_n69);
	nor (gm_n1036, gm_n57, in_12, in_8, gm_n230, gm_n94);
	nand (gm_n1037, gm_n1036, gm_n69, gm_n62);
	and (gm_n1038, gm_n183, gm_n105, in_8);
	nand (gm_n1039, gm_n69, in_13, gm_n41, gm_n1038, gm_n126);
	and (gm_n1040, gm_n247, gm_n101, in_14);
	nor (gm_n1041, gm_n119, gm_n59, in_14, gm_n566, gm_n227);
	nand (gm_n1042, in_14, gm_n62, gm_n41, gm_n1021, gm_n126);
	or (gm_n1043, gm_n193, gm_n351, in_8);
	or (gm_n1044, gm_n69, gm_n62, in_12, gm_n1043, gm_n71);
	nor (gm_n1045, gm_n469, gm_n87, gm_n69);
	nor (gm_n1046, gm_n208, gm_n57, in_8);
	and (gm_n1047, gm_n69, in_13, in_12, gm_n1046, gm_n131);
	nand (gm_n1048, gm_n86, gm_n66, in_14, gm_n106, gm_n88);
	nand (gm_n1049, gm_n246, gm_n183, gm_n45);
	or (gm_n1050, in_14, gm_n62, in_12, gm_n1049, gm_n71);
	nor (gm_n1051, gm_n342, gm_n150, gm_n45, gm_n516, gm_n193);
	nor (gm_n1052, gm_n145, gm_n69, in_10, gm_n287, gm_n239);
	and (gm_n1053, gm_n109, in_12, in_8, gm_n274, gm_n126);
	nand (gm_n1054, gm_n1053, gm_n69, in_13);
	nand (gm_n1055, gm_n320, gm_n109, gm_n43, gm_n117, gm_n106);
	and (gm_n1056, gm_n104, gm_n46, in_11, gm_n381, gm_n169);
	nor (gm_n1057, gm_n231, gm_n385, gm_n45);
	and (gm_n1058, gm_n69, gm_n42, in_9, gm_n1057, gm_n300);
	and (gm_n1059, gm_n349, in_12, gm_n45, gm_n129, gm_n72);
	nand (gm_n1060, gm_n1059, gm_n69, gm_n62);
	or (gm_n1061, gm_n90, gm_n351, in_8, gm_n882, gm_n342);
	nand (gm_n1062, gm_n245, in_14, in_10, gm_n741, gm_n454);
	nand (gm_n1063, in_14, gm_n62, gm_n41, gm_n829, gm_n93);
	nand (gm_n1064, gm_n1061, gm_n1060, t_8, gm_n1063, gm_n1062);
	nand (gm_n1065, in_14, in_13, gm_n41, gm_n670, gm_n131);
	nand (gm_n1066, in_14, gm_n62, gm_n41, gm_n922, gm_n349);
	nand (gm_n1067, gm_n129, gm_n161, in_11, gm_n233, gm_n174);
	nand (gm_n1068, gm_n1067, gm_n1066, gm_n1065);
	nand (gm_n1069, gm_n88, gm_n73, in_8, gm_n117, gm_n93);
	nand (gm_n1070, gm_n243, gm_n65, in_11, gm_n163, gm_n133);
	nand (gm_n1071, gm_n72, gm_n370, in_8, gm_n224, gm_n126);
	nand (gm_n1072, gm_n1071, gm_n1070, gm_n1069);
	nor (gm_n1073, gm_n1064, gm_n1058, gm_n1056, gm_n1072, gm_n1068);
	nor (gm_n1074, in_14, gm_n62, in_12, gm_n926, gm_n230);
	nor (gm_n1075, gm_n108, gm_n69, in_10, gm_n307, gm_n287);
	nor (gm_n1076, gm_n906, gm_n119, in_14);
	nor (gm_n1077, gm_n1076, gm_n1075, gm_n1074);
	nor (gm_n1078, gm_n69, in_13, gm_n41, gm_n474, gm_n76);
	nor (gm_n1079, gm_n351, gm_n57, gm_n45, gm_n261, gm_n154);
	nor (gm_n1080, in_14, gm_n42, in_9, gm_n521, gm_n119);
	nor (gm_n1081, gm_n1080, gm_n1079, gm_n1078);
	nand (gm_n1082, gm_n1073, gm_n1055, gm_n1054, gm_n1081, gm_n1077);
	nand (gm_n1083, gm_n322, in_14, gm_n42, gm_n329, gm_n178);
	nand (gm_n1084, gm_n799, gm_n164, gm_n53);
	nor (gm_n1085, gm_n42, gm_n70, in_8, gm_n189, gm_n385);
	nand (gm_n1086, gm_n1085, gm_n178, gm_n69);
	nand (gm_n1087, gm_n1086, gm_n1084, gm_n1083);
	nand (gm_n1088, gm_n69, gm_n42, in_9, gm_n1057, gm_n101);
	nand (gm_n1089, gm_n440, gm_n69, gm_n62);
	nand (gm_n1090, gm_n93, gm_n88, in_8, gm_n277, gm_n117);
	nand (gm_n1091, gm_n1090, gm_n1089, gm_n1088);
	nor (gm_n1092, gm_n1082, gm_n1052, gm_n1051, gm_n1091, gm_n1087);
	nor (gm_n1093, gm_n155, in_11, gm_n58, gm_n882, gm_n156);
	nor (gm_n1094, in_14, in_13, gm_n41, gm_n926, gm_n261);
	nand (gm_n1095, gm_n268, gm_n46, gm_n45);
	nor (gm_n1096, gm_n69, in_13, in_12, gm_n1095, gm_n76);
	nor (gm_n1097, gm_n1096, gm_n1094, gm_n1093);
	and (gm_n1098, gm_n106, gm_n72, gm_n43, gm_n381, gm_n174);
	nand (gm_n1099, in_7, gm_n79, gm_n64, gm_n124, in_8);
	nor (gm_n1100, gm_n69, gm_n62, in_12, gm_n1099, gm_n71);
	and (gm_n1101, gm_n133, gm_n65, in_8);
	and (gm_n1102, gm_n69, in_13, gm_n41, gm_n1101, gm_n191);
	nor (gm_n1103, gm_n1102, gm_n1100, gm_n1098);
	nand (gm_n1104, gm_n1092, gm_n1050, gm_n1048, gm_n1103, gm_n1097);
	and (gm_n1105, gm_n58, in_6, gm_n64, gm_n124, in_8);
	nand (gm_n1106, in_14, gm_n42, gm_n70, gm_n1105, gm_n83);
	nor (gm_n1107, gm_n147, gm_n385, in_8);
	nand (gm_n1108, gm_n69, gm_n62, gm_n41, gm_n1107, gm_n349);
	and (gm_n1109, gm_n277, gm_n88, gm_n45);
	nand (gm_n1110, in_14, in_13, in_12, gm_n1109, gm_n191);
	nand (gm_n1111, gm_n1110, gm_n1108, gm_n1106);
	or (gm_n1112, gm_n108, in_14, in_10, gm_n307, gm_n305);
	nand (gm_n1113, gm_n322, in_14, gm_n42, gm_n329, gm_n300);
	nand (gm_n1114, gm_n93, gm_n46, gm_n45, gm_n274, gm_n168);
	nand (gm_n1115, gm_n1114, gm_n1113, gm_n1112);
	nor (gm_n1116, gm_n1104, gm_n1047, gm_n1045, gm_n1115, gm_n1111);
	and (gm_n1117, gm_n69, in_13, in_12, gm_n767, gm_n131);
	nor (gm_n1118, gm_n108, in_14, gm_n42, gm_n290);
	and (gm_n1119, gm_n105, gm_n72, gm_n45, gm_n191, gm_n174);
	nor (gm_n1120, gm_n1119, gm_n1118, gm_n1117);
	and (gm_n1121, gm_n93, gm_n46, in_8, gm_n168, gm_n110);
	nor (gm_n1122, gm_n87, gm_n385, in_14, gm_n249, gm_n90);
	nor (gm_n1123, gm_n562, gm_n77, gm_n43, gm_n593);
	nor (gm_n1124, gm_n1123, gm_n1122, gm_n1121);
	nand (gm_n1125, gm_n1116, gm_n1044, gm_n1042, gm_n1124, gm_n1120);
	nand (gm_n1126, gm_n86, gm_n69, in_10, gm_n211, gm_n144);
	or (gm_n1127, gm_n69, gm_n62, in_12, gm_n644, gm_n261);
	nand (gm_n1128, in_14, gm_n42, gm_n70, gm_n799, gm_n101);
	nand (gm_n1129, gm_n1128, gm_n1127, gm_n1126);
	nor (gm_n1130, gm_n64, in_4, gm_n55, gm_n120, gm_n79);
	nand (gm_n1131, gm_n322, in_14, in_10, gm_n1130, gm_n300);
	nand (gm_n1132, gm_n161, gm_n93, gm_n45, gm_n295, gm_n246);
	nand (gm_n1133, gm_n126, gm_n65, gm_n45, gm_n170, gm_n164);
	nand (gm_n1134, gm_n1133, gm_n1132, gm_n1131);
	nor (gm_n1135, gm_n1125, gm_n1041, gm_n1040, gm_n1134, gm_n1129);
	nor (gm_n1136, in_14, in_13, gm_n41, gm_n217, gm_n216);
	and (gm_n1137, gm_n69, in_13, in_12, gm_n278, gm_n44);
	nand (gm_n1138, gm_n42, gm_n70, gm_n45, gm_n274, gm_n88);
	nor (gm_n1139, gm_n1138, gm_n84, in_14);
	nor (gm_n1140, gm_n1139, gm_n1137, gm_n1136);
	and (gm_n1141, gm_n69, in_13, in_12, gm_n668, gm_n191);
	nor (gm_n1142, gm_n84, in_14, in_10, gm_n155, gm_n122);
	nor (gm_n1143, gm_n1142, gm_n1141, gm_n135);
	nand (gm_n1144, gm_n1135, gm_n1039, gm_n1037, gm_n1143, gm_n1140);
	nand (gm_n1145, gm_n69, gm_n62, in_12, gm_n581, gm_n349);
	nand (gm_n1146, gm_n69, in_13, in_9, gm_n758, gm_n757);
	nand (gm_n1147, gm_n720, gm_n46, in_11, gm_n233, gm_n117);
	nand (gm_n1148, gm_n1147, gm_n1146, gm_n1145);
	nor (gm_n1149, gm_n147, gm_n351, gm_n45);
	nand (gm_n1150, in_14, in_13, gm_n41, gm_n1149, gm_n349);
	nand (gm_n1151, gm_n110, gm_n161, gm_n43, gm_n284, gm_n117);
	nor (gm_n1152, gm_n227, gm_n208, in_8);
	nand (gm_n1153, gm_n69, gm_n62, gm_n41, gm_n1152, gm_n349);
	nand (gm_n1154, gm_n1153, gm_n1151, gm_n1150);
	nor (gm_n1155, gm_n1144, gm_n1035, gm_n1033, gm_n1154, gm_n1148);
	nand (gm_n1156, in_14, gm_n62, gm_n41, gm_n459, gm_n191);
	nand (gm_n1157, gm_n104, gm_n46, gm_n43, gm_n170, gm_n163);
	nand (gm_n1158, gm_n69, in_13, in_12, gm_n98, gm_n60);
	nand (gm_n1159, gm_n1156, gm_n1155, gm_n1032, gm_n1158, gm_n1157);
	nor (gm_n1160, gm_n351, in_12, gm_n45, gm_n193, gm_n261);
	and (gm_n1161, gm_n1160, gm_n69, gm_n62);
	nor (gm_n1162, in_14, in_10, in_9, gm_n119, gm_n82);
	and (gm_n1163, gm_n104, gm_n161, gm_n43, gm_n266, gm_n133);
	or (gm_n1164, gm_n1163, gm_n1162, gm_n1161);
	or (gm_n1165, in_14, gm_n62, in_12, gm_n637, gm_n327);
	nand (gm_n1166, gm_n69, gm_n62, gm_n41, gm_n691, gm_n53);
	and (gm_n1167, gm_n184, gm_n88, in_8);
	nand (gm_n1168, gm_n69, gm_n62, gm_n41, gm_n1167, gm_n53);
	nand (gm_n1169, gm_n1168, gm_n1166, gm_n1165);
	nor (out_7, gm_n1164, gm_n1159, gm_n1031, gm_n1169);
	and (gm_n1171, gm_n69, gm_n42, gm_n70, gm_n125, gm_n101);
	nand (gm_n1172, gm_n144, gm_n69, in_10, gm_n300, gm_n211);
	nand (gm_n1173, gm_n300, gm_n69, gm_n42, gm_n323, gm_n289);
	and (gm_n1174, gm_n69, gm_n62, in_12, gm_n725, gm_n126);
	nor (gm_n1175, gm_n280, gm_n47, in_8);
	and (gm_n1176, gm_n69, in_10, gm_n70, gm_n1175, gm_n345);
	nand (gm_n1177, in_14, gm_n62, in_12, gm_n677, gm_n44);
	nand (gm_n1178, in_14, in_13, in_12, gm_n222, gm_n53);
	and (gm_n1179, gm_n245, gm_n69, gm_n42, gm_n329, gm_n943);
	or (gm_n1180, gm_n89, gm_n41, gm_n45, gm_n201, gm_n261);
	nor (gm_n1181, gm_n1180, gm_n69, gm_n62);
	nand (gm_n1182, gm_n86, in_14, gm_n42, gm_n346, gm_n943);
	and (gm_n1183, gm_n161, in_12, gm_n45, gm_n126, gm_n105);
	nand (gm_n1184, gm_n1183, in_14, in_13);
	or (gm_n1185, gm_n42, in_6, gm_n64, gm_n307, gm_n301);
	nor (gm_n1186, gm_n1185, gm_n271, gm_n69);
	nor (gm_n1187, gm_n226, gm_n229, gm_n43, gm_n241);
	nand (gm_n1188, gm_n42, gm_n70, in_8, gm_n133, gm_n80);
	or (gm_n1189, gm_n1188, gm_n87, in_14);
	nand (gm_n1190, gm_n69, in_10, gm_n70, gm_n394, gm_n178);
	nor (gm_n1191, in_14, in_10, in_9, gm_n134, gm_n119);
	and (gm_n1192, gm_n163, gm_n115, in_11, gm_n174);
	nand (gm_n1193, gm_n86, in_14, in_10, gm_n211, gm_n144);
	nand (gm_n1194, in_14, gm_n62, in_12, gm_n131, gm_n60);
	and (gm_n1195, gm_n243, gm_n46, gm_n45, gm_n126, gm_n110);
	and (gm_n1196, gm_n349, gm_n370, gm_n45, gm_n174, gm_n80);
	and (gm_n1197, gm_n349, in_12, gm_n45, gm_n129, gm_n88);
	nand (gm_n1198, gm_n1197, gm_n69, gm_n62);
	nand (gm_n1199, gm_n131, gm_n161, in_8, gm_n246, gm_n224);
	and (gm_n1200, gm_n72, gm_n53, in_8, gm_n274, gm_n117);
	and (gm_n1201, gm_n109, gm_n44, gm_n45, gm_n199, gm_n174);
	nand (gm_n1202, gm_n105, gm_n88, gm_n45);
	nor (gm_n1203, in_14, gm_n62, gm_n41, gm_n1202, gm_n342);
	and (gm_n1204, in_14, in_13, in_12, gm_n670, gm_n126);
	nor (gm_n1205, in_14, gm_n42, gm_n70, gm_n637, gm_n119);
	nor (gm_n1206, gm_n1203, gm_n1201, gm_n1200, gm_n1205, gm_n1204);
	and (gm_n1207, gm_n69, gm_n62, in_12, gm_n471, gm_n349);
	nand (gm_n1208, gm_n53, in_12, in_8, gm_n105, gm_n161);
	nor (gm_n1209, gm_n1208, in_14, in_13);
	and (gm_n1210, gm_n69, gm_n62, in_12, gm_n428, gm_n98);
	nor (gm_n1211, gm_n1210, gm_n1209, gm_n1207);
	nor (gm_n1212, gm_n417, in_14, in_10, gm_n302, gm_n287);
	nor (gm_n1213, gm_n177, gm_n151, gm_n69);
	and (gm_n1214, gm_n88, gm_n66, gm_n69, gm_n136, gm_n106);
	nor (gm_n1215, gm_n1214, gm_n1213, gm_n1212);
	nand (gm_n1216, gm_n1206, gm_n1199, gm_n1198, gm_n1215, gm_n1211);
	or (gm_n1217, gm_n119, in_14, gm_n42, gm_n287, gm_n467);
	nand (gm_n1218, in_14, gm_n62, in_12, gm_n1107, gm_n44);
	nor (gm_n1219, gm_n50, gm_n41, gm_n45, gm_n208, gm_n63);
	nand (gm_n1220, gm_n1219, gm_n69, gm_n62);
	nand (gm_n1221, gm_n1220, gm_n1218, gm_n1217);
	nand (gm_n1222, gm_n295, gm_n169, gm_n43, gm_n655);
	nand (gm_n1223, gm_n1034, gm_n86, gm_n69);
	nand (gm_n1224, gm_n1223, gm_n1222, gm_n763);
	nor (gm_n1225, gm_n1216, gm_n1196, gm_n1195, gm_n1224, gm_n1221);
	not (gm_n1226, gm_n741);
	nor (gm_n1227, gm_n121, in_14, in_10, gm_n1226, gm_n271);
	nand (gm_n1228, gm_n109, gm_n41, in_8, gm_n277, gm_n131);
	nor (gm_n1229, gm_n1228, in_14, in_13);
	nor (gm_n1230, gm_n69, in_10, gm_n70, gm_n500, gm_n119);
	nor (gm_n1231, gm_n1230, gm_n1229, gm_n1227);
	nor (gm_n1232, gm_n94, gm_n76, gm_n45, gm_n516, gm_n231);
	nor (gm_n1233, gm_n69, gm_n42, in_9, gm_n987, gm_n108);
	nand (gm_n1234, gm_n42, gm_n70, in_8, gm_n105, gm_n65);
	nor (gm_n1235, gm_n1234, gm_n239, in_14);
	nor (gm_n1236, gm_n1235, gm_n1233, gm_n1232);
	nand (gm_n1237, gm_n1225, gm_n1194, gm_n1193, gm_n1236, gm_n1231);
	nand (gm_n1238, gm_n178, gm_n116, in_14, gm_n631);
	nand (gm_n1239, gm_n69, gm_n62, gm_n41, gm_n668, gm_n53);
	nand (gm_n1240, gm_n129, gm_n161, in_11, gm_n233, gm_n168);
	nand (gm_n1241, gm_n1240, gm_n1239, gm_n1238);
	nand (gm_n1242, in_14, gm_n62, in_12, gm_n760, gm_n126);
	and (gm_n1243, in_6, gm_n64, in_4, gm_n114);
	nand (gm_n1244, gm_n144, in_14, in_10, gm_n1243, gm_n300);
	nand (gm_n1245, gm_n233, gm_n104, in_11, gm_n655);
	nand (gm_n1246, gm_n1245, gm_n1244, gm_n1242);
	nor (gm_n1247, gm_n1237, gm_n1192, gm_n1191, gm_n1246, gm_n1241);
	nand (gm_n1248, gm_n72, gm_n41, gm_n45, gm_n191, gm_n110);
	nor (gm_n1249, gm_n1248, in_14, in_13);
	nor (gm_n1250, gm_n119, gm_n249, in_14, gm_n503);
	nand (gm_n1251, gm_n42, in_9, in_8, gm_n268, gm_n65);
	nor (gm_n1252, gm_n1251, gm_n417, gm_n69);
	nor (gm_n1253, gm_n1252, gm_n1250, gm_n1249);
	nand (gm_n1254, gm_n349, in_12, in_8, gm_n277, gm_n88);
	nor (gm_n1255, gm_n1254, in_14, gm_n62);
	nor (gm_n1256, gm_n69, in_13, gm_n41, gm_n770, gm_n216);
	nor (gm_n1257, gm_n108, in_14, in_10, gm_n305, gm_n145);
	nor (gm_n1258, gm_n1257, gm_n1256, gm_n1255);
	nand (gm_n1259, gm_n1247, gm_n1190, gm_n1189, gm_n1258, gm_n1253);
	nand (gm_n1260, gm_n233, gm_n104, in_11, gm_n253);
	nand (gm_n1261, in_14, gm_n62, gm_n41, gm_n222, gm_n126);
	or (gm_n1262, in_14, in_13, gm_n41, gm_n770, gm_n327);
	nand (gm_n1263, gm_n1262, gm_n1261, gm_n1260);
	nand (gm_n1264, in_14, gm_n42, in_9, gm_n278, gm_n345);
	or (gm_n1265, gm_n417, gm_n69, in_10, gm_n1226, gm_n287);
	or (gm_n1266, in_14, gm_n62, in_12, gm_n901, gm_n342);
	nand (gm_n1267, gm_n1266, gm_n1265, gm_n1264);
	nor (gm_n1268, gm_n1259, gm_n1187, gm_n1186, gm_n1267, gm_n1263);
	and (gm_n1269, in_14, in_13, gm_n41, gm_n624, gm_n191);
	and (gm_n1270, gm_n80, gm_n44, gm_n45, gm_n199, gm_n117);
	nand (gm_n1271, gm_n268, gm_n72, in_8);
	nor (gm_n1272, in_14, gm_n62, gm_n41, gm_n1271, gm_n327);
	nor (gm_n1273, gm_n1272, gm_n1270, gm_n1269);
	nand (gm_n1274, gm_n720, gm_n109, gm_n45);
	nor (gm_n1275, in_14, in_13, in_12, gm_n1274, gm_n216);
	nor (gm_n1276, gm_n119, gm_n69, gm_n42, gm_n330, gm_n418);
	and (gm_n1277, gm_n164, gm_n65, in_11, gm_n246, gm_n284);
	nor (gm_n1278, gm_n1277, gm_n1276, gm_n1275);
	nand (gm_n1279, gm_n1268, gm_n1184, gm_n1182, gm_n1278, gm_n1273);
	nand (gm_n1280, gm_n69, gm_n42, in_9, gm_n492, gm_n83);
	nand (gm_n1281, in_14, in_13, gm_n41, gm_n480, gm_n191);
	nand (gm_n1282, in_14, gm_n62, gm_n41, gm_n492, gm_n191);
	nand (gm_n1283, gm_n1282, gm_n1281, gm_n1280);
	and (gm_n1284, in_7, gm_n79, gm_n64, gm_n124, gm_n45);
	nand (gm_n1285, gm_n69, gm_n62, gm_n41, gm_n1284, gm_n126);
	nand (gm_n1286, gm_n86, in_14, gm_n42, gm_n1130, gm_n139);
	nand (gm_n1287, gm_n243, gm_n46, gm_n43, gm_n169, gm_n133);
	nand (gm_n1288, gm_n1287, gm_n1286, gm_n1285);
	nor (gm_n1289, gm_n1279, gm_n1181, gm_n1179, gm_n1288, gm_n1283);
	nor (gm_n1290, gm_n162, gm_n89, in_11, gm_n201, gm_n229);
	nor (gm_n1291, in_14, in_13, in_12, gm_n438, gm_n327);
	nor (gm_n1292, gm_n69, in_13, gm_n41, gm_n687, gm_n76);
	nor (gm_n1293, gm_n1292, gm_n1291, gm_n1290);
	nor (gm_n1294, gm_n69, gm_n62, in_12, gm_n342, gm_n67);
	and (gm_n1295, gm_n104, gm_n505, gm_n53);
	nor (gm_n1296, in_14, in_10, in_9, gm_n108, gm_n67);
	nor (gm_n1297, gm_n1296, gm_n1295, gm_n1294);
	nand (gm_n1298, gm_n1289, gm_n1178, gm_n1177, gm_n1297, gm_n1293);
	or (gm_n1299, gm_n69, in_13, gm_n41, gm_n1202, gm_n327);
	nand (gm_n1300, gm_n69, in_13, gm_n41, gm_n691, gm_n349);
	nand (gm_n1301, in_14, gm_n62, in_12, gm_n725, gm_n93);
	nand (gm_n1302, gm_n1301, gm_n1300, gm_n1299);
	nand (gm_n1303, in_14, gm_n62, in_12, gm_n386, gm_n191);
	nand (gm_n1304, gm_n69, gm_n62, gm_n41, gm_n823, gm_n44);
	nand (gm_n1305, gm_n69, in_13, gm_n41, gm_n973, gm_n98);
	nand (gm_n1306, gm_n1305, gm_n1304, gm_n1303);
	nor (gm_n1307, gm_n1298, gm_n1176, gm_n1174, gm_n1306, gm_n1302);
	nor (gm_n1308, gm_n154, gm_n89, in_11, gm_n566, gm_n201);
	nor (gm_n1309, gm_n69, gm_n62, gm_n41, gm_n256, gm_n261);
	nor (gm_n1310, gm_n69, gm_n62, gm_n41, gm_n514, gm_n230);
	nor (gm_n1311, gm_n1310, gm_n1309, gm_n1308);
	and (gm_n1312, gm_n245, gm_n65, gm_n69, gm_n246, gm_n559);
	nand (gm_n1313, gm_n129, gm_n109, in_8);
	nor (gm_n1314, in_14, gm_n62, in_12, gm_n1313, gm_n342);
	and (gm_n1315, in_14, in_13, gm_n41, gm_n459, gm_n126);
	nor (gm_n1316, gm_n1315, gm_n1314, gm_n1312);
	nand (gm_n1317, gm_n1307, gm_n1173, gm_n1172, gm_n1316, gm_n1311);
	nor (gm_n1318, in_10, gm_n70, gm_n45, gm_n231, gm_n89);
	nand (gm_n1319, gm_n1318, gm_n178, in_14);
	or (gm_n1320, gm_n201, gm_n385, gm_n45);
	or (gm_n1321, in_14, in_13, gm_n41, gm_n1320, gm_n63);
	and (gm_n1322, gm_n53, in_12, in_8, gm_n199, gm_n161);
	nand (gm_n1323, gm_n1322, gm_n69, in_13);
	nand (gm_n1324, gm_n1323, gm_n1321, gm_n1319);
	or (gm_n1325, gm_n249, gm_n351, in_14, gm_n239, gm_n201);
	or (gm_n1326, gm_n150, gm_n77, gm_n45, gm_n193, gm_n342);
	nand (gm_n1327, gm_n69, gm_n62, in_12, gm_n394, gm_n93);
	nand (gm_n1328, gm_n1327, gm_n1326, gm_n1325);
	nor (out_8, gm_n1324, gm_n1317, gm_n1171, gm_n1328);
	nand (gm_n1330, gm_n46, in_12, in_8, gm_n199, gm_n98);
	nor (gm_n1331, gm_n1330, gm_n69, gm_n62);
	nand (gm_n1332, gm_n104, gm_n46, gm_n43, gm_n381, gm_n116);
	nand (gm_n1333, gm_n73, gm_n41, gm_n45, gm_n98, gm_n88);
	nor (gm_n1334, gm_n1333, in_14, gm_n62);
	nor (gm_n1335, gm_n108, gm_n69, in_10, gm_n305, gm_n286);
	nand (gm_n1336, gm_n136, gm_n69, in_10, gm_n329, gm_n943);
	nand (gm_n1337, gm_n69, gm_n62, in_12, gm_n555, gm_n44);
	and (gm_n1338, in_14, in_10, in_9, gm_n178, gm_n130);
	or (gm_n1339, gm_n227, gm_n47, gm_n45);
	nor (gm_n1340, in_14, in_13, in_12, gm_n1339, gm_n76);
	nand (gm_n1341, in_14, in_13, in_12, gm_n194, gm_n349);
	and (gm_n1342, gm_n370, gm_n41, gm_n45, gm_n191, gm_n88);
	nand (gm_n1343, gm_n1342, gm_n69, gm_n62);
	nor (gm_n1344, in_14, gm_n62, in_12, gm_n1274, gm_n261);
	and (gm_n1345, gm_n69, gm_n62, in_12, gm_n922, gm_n126);
	nor (gm_n1346, gm_n95, gm_n59, gm_n45);
	nand (gm_n1347, gm_n69, gm_n62, gm_n41, gm_n1346, gm_n191);
	or (gm_n1348, gm_n1138, gm_n87, in_14);
	nand (gm_n1349, gm_n106, gm_n88, in_11, gm_n168, gm_n110);
	or (gm_n1350, gm_n69, in_13, gm_n41, gm_n626, gm_n216);
	nand (gm_n1351, gm_n80, gm_n44, gm_n45, gm_n224, gm_n133);
	or (gm_n1352, gm_n352, gm_n84, gm_n69);
	and (gm_n1353, gm_n1350, gm_n1349, t_6, gm_n1352, gm_n1351);
	and (gm_n1354, gm_n124, gm_n46, gm_n45);
	and (gm_n1355, gm_n69, in_13, in_12, gm_n1354, gm_n349);
	nand (gm_n1356, gm_n161, in_12, in_8, gm_n255, gm_n98);
	nor (gm_n1357, gm_n1356, in_14, in_13);
	and (gm_n1358, gm_n69, in_13, gm_n41, gm_n1346, gm_n98);
	nor (gm_n1359, gm_n1358, gm_n1357, gm_n1355);
	or (gm_n1360, gm_n385, gm_n57, in_8);
	nor (gm_n1361, in_14, gm_n42, gm_n70, gm_n1360, gm_n177);
	and (gm_n1362, gm_n233, gm_n174, in_11, gm_n655);
	and (gm_n1363, gm_n168, gm_n559, in_11, gm_n392);
	nor (gm_n1364, gm_n1363, gm_n1362, gm_n1361);
	nand (gm_n1365, gm_n1353, gm_n1348, gm_n1347, gm_n1364, gm_n1359);
	nor (gm_n1366, gm_n69, gm_n62, in_12, gm_n1313, gm_n71);
	and (gm_n1367, in_14, gm_n62, in_12, gm_n220, gm_n98);
	or (gm_n1368, gm_n1367, gm_n1366, gm_n1296);
	or (gm_n1369, gm_n69, gm_n62, in_12, gm_n67, gm_n76);
	and (gm_n1370, gm_n44, gm_n41, gm_n45, gm_n183, gm_n81);
	nand (gm_n1371, gm_n1370, gm_n69, in_13);
	or (gm_n1372, in_14, in_13, gm_n41, gm_n1320, gm_n327);
	nand (gm_n1373, gm_n1372, gm_n1371, gm_n1369);
	nor (gm_n1374, gm_n1365, gm_n1345, gm_n1344, gm_n1373, gm_n1368);
	and (gm_n1375, gm_n69, gm_n42, in_9, gm_n829, gm_n136);
	nand (gm_n1376, gm_n109, gm_n41, gm_n45, gm_n129, gm_n93);
	nor (gm_n1377, gm_n1376, gm_n69, in_13);
	and (gm_n1378, in_14, in_13, gm_n41, gm_n816, gm_n131);
	nor (gm_n1379, gm_n1378, gm_n1377, gm_n1375);
	and (gm_n1380, gm_n131, gm_n161, gm_n45, gm_n268, gm_n174);
	and (gm_n1381, gm_n69, gm_n62, in_12, gm_n394, gm_n126);
	nor (gm_n1382, gm_n63, gm_n50, in_8, gm_n150, gm_n77);
	nor (gm_n1383, gm_n1382, gm_n1381, gm_n1380);
	nand (gm_n1384, gm_n1374, gm_n1343, gm_n1341, gm_n1383, gm_n1379);
	nand (gm_n1385, in_14, in_13, gm_n41, gm_n1109, gm_n98);
	nand (gm_n1386, gm_n104, gm_n161, gm_n43, gm_n124, gm_n106);
	nand (gm_n1387, gm_n184, gm_n183, gm_n45, gm_n295, gm_n191);
	nand (gm_n1388, gm_n1387, gm_n1386, gm_n1385);
	nand (gm_n1389, gm_n131, gm_n161, in_8, gm_n246, gm_n168);
	or (gm_n1390, gm_n177, gm_n69, in_10, gm_n302, gm_n287);
	nand (gm_n1391, gm_n109, gm_n370, gm_n43, gm_n559, gm_n104);
	nand (gm_n1392, gm_n1391, gm_n1390, gm_n1389);
	nor (gm_n1393, gm_n1384, gm_n1340, gm_n1338, gm_n1392, gm_n1388);
	nand (gm_n1394, gm_n161, gm_n81, in_8);
	nor (gm_n1395, in_14, in_10, gm_n70, gm_n1394, gm_n239);
	nor (gm_n1396, gm_n59, gm_n57, gm_n45, gm_n882, gm_n261);
	nand (gm_n1397, gm_n73, in_12, in_8, gm_n131, gm_n88);
	nor (gm_n1398, gm_n1397, gm_n69, gm_n62);
	nor (gm_n1399, gm_n1398, gm_n1396, gm_n1395);
	nand (gm_n1400, gm_n268, gm_n161, in_8);
	nor (gm_n1401, in_14, gm_n42, gm_n70, gm_n1400, gm_n417);
	nor (gm_n1402, in_14, gm_n62, in_12, gm_n1095, gm_n216);
	and (gm_n1403, in_14, gm_n62, in_12, gm_n1167, gm_n98);
	nor (gm_n1404, gm_n1403, gm_n1402, gm_n1401);
	nand (gm_n1405, gm_n1393, gm_n1337, gm_n1336, gm_n1404, gm_n1399);
	nand (gm_n1406, gm_n559, gm_n117, gm_n43, gm_n311);
	nand (gm_n1407, gm_n101, in_14, in_10, gm_n258, gm_n139);
	and (gm_n1408, gm_n72, gm_n41, gm_n45, gm_n98, gm_n81);
	nand (gm_n1409, gm_n1408, gm_n69, gm_n62);
	nand (gm_n1410, gm_n1409, gm_n1407, gm_n1406);
	nand (gm_n1411, gm_n69, in_13, in_12, gm_n973, gm_n191);
	nand (gm_n1412, gm_n116, gm_n161, gm_n43, gm_n224, gm_n124);
	not (gm_n1413, gm_n237);
	nand (gm_n1414, gm_n139, in_14, in_10, gm_n300, gm_n1413);
	nand (gm_n1415, gm_n1414, gm_n1412, gm_n1411);
	nor (gm_n1416, gm_n1405, gm_n1335, gm_n1334, gm_n1415, gm_n1410);
	nand (gm_n1417, in_14, in_13, in_12, gm_n1149, gm_n44);
	nand (gm_n1418, gm_n93, gm_n46, in_8, gm_n110, gm_n104);
	nand (gm_n1419, gm_n69, gm_n62, in_12, gm_n148, gm_n93);
	nand (gm_n1420, gm_n1417, gm_n1416, gm_n1332, gm_n1419, gm_n1418);
	or (gm_n1421, gm_n143, in_14, in_10, gm_n307, gm_n177);
	or (gm_n1422, gm_n69, in_13, gm_n41, gm_n987, gm_n342);
	nor (gm_n1423, gm_n57, gm_n41, gm_n45, gm_n230, gm_n385);
	nand (gm_n1424, gm_n1423, gm_n69, in_13);
	nand (gm_n1425, gm_n1424, gm_n1422, gm_n1421);
	or (gm_n1426, gm_n566, gm_n882, in_11, gm_n593);
	nand (gm_n1427, gm_n86, in_14, in_10, gm_n346, gm_n943);
	nand (gm_n1428, gm_n69, gm_n42, in_9, gm_n426, gm_n245);
	nand (gm_n1429, gm_n1428, gm_n1427, gm_n1426);
	nor (out_9, gm_n1425, gm_n1420, gm_n1331, gm_n1429);
	and (gm_n1431, gm_n69, in_10, in_9, gm_n486, gm_n83);
	nand (gm_n1432, gm_n381, gm_n46, in_11, gm_n295, gm_n233);
	nor (gm_n1433, gm_n71, in_12, in_8, gm_n201, gm_n94);
	nand (gm_n1434, gm_n1433, gm_n69, gm_n62);
	nand (gm_n1435, gm_n42, in_9, in_8, gm_n183, gm_n133);
	nor (gm_n1436, gm_n1435, gm_n119, in_14);
	and (gm_n1437, gm_n320, gm_n109, in_11, gm_n224, gm_n116);
	nor (gm_n1438, gm_n385, in_12, in_8, gm_n201, gm_n230);
	nand (gm_n1439, gm_n1438, in_14, in_13);
	or (gm_n1440, in_14, gm_n62, in_12, gm_n438, gm_n63);
	or (gm_n1441, gm_n150, gm_n41, in_8, gm_n227, gm_n216);
	nor (gm_n1442, gm_n1441, in_14, in_13);
	and (gm_n1443, in_14, gm_n62, in_12, gm_n586, gm_n349);
	nand (gm_n1444, in_14, gm_n62, gm_n41, gm_n762, gm_n349);
	nand (gm_n1445, gm_n69, in_13, gm_n41, gm_n1000, gm_n53);
	nor (gm_n1446, gm_n637, gm_n261, gm_n154);
	nor (gm_n1447, gm_n351, gm_n50, gm_n45);
	and (gm_n1448, gm_n69, in_13, in_12, gm_n1447, gm_n93);
	nand (gm_n1449, gm_n124, gm_n88, in_11, gm_n224, gm_n169);
	or (gm_n1450, gm_n87, gm_n69, in_10, gm_n237, gm_n145);
	nor (gm_n1451, in_14, gm_n62, in_12, gm_n806, gm_n76);
	and (gm_n1452, gm_n69, gm_n62, in_12, gm_n488, gm_n93);
	nand (gm_n1453, in_14, gm_n62, in_12, gm_n620, gm_n131);
	nand (gm_n1454, in_14, in_13, gm_n41, gm_n1346, gm_n44);
	nor (gm_n1455, in_14, in_13, gm_n41, gm_n844, gm_n71);
	not (gm_n1456, gm_n840);
	nor (gm_n1457, gm_n418, gm_n69, gm_n42, gm_n1456, gm_n177);
	nand (gm_n1458, gm_n69, gm_n42, in_9, gm_n829, gm_n86);
	nand (gm_n1459, gm_n69, in_13, gm_n41, gm_n358, gm_n53);
	nor (gm_n1460, gm_n69, gm_n62, gm_n41, gm_n134, gm_n63);
	nor (gm_n1461, gm_n69, in_13, in_12, gm_n1049, gm_n342);
	nand (gm_n1462, gm_n73, gm_n41, in_8, gm_n183, gm_n126);
	nor (gm_n1463, gm_n1462, in_14, in_13);
	nor (gm_n1464, in_14, in_13, gm_n41, gm_n343, gm_n327);
	and (gm_n1465, gm_n720, gm_n46, in_11, gm_n224, gm_n106);
	nor (gm_n1466, gm_n1463, gm_n1461, gm_n1460, gm_n1465, gm_n1464);
	nor (gm_n1467, gm_n121, gm_n69, gm_n42, gm_n307, gm_n177);
	nor (gm_n1468, gm_n108, gm_n69, gm_n42, gm_n287, gm_n145);
	nor (gm_n1469, gm_n69, gm_n42, in_9, gm_n377, gm_n108);
	nor (gm_n1470, gm_n1469, gm_n1468, gm_n1467);
	nand (gm_n1471, gm_n133, gm_n109, in_8);
	nor (gm_n1472, in_14, in_13, gm_n41, gm_n1471, gm_n63);
	nor (gm_n1473, gm_n69, gm_n62, in_12, gm_n867, gm_n71);
	nor (gm_n1474, gm_n69, gm_n62, gm_n41, gm_n806, gm_n230);
	nor (gm_n1475, gm_n1474, gm_n1473, gm_n1472);
	nand (gm_n1476, gm_n1466, gm_n1459, gm_n1458, gm_n1475, gm_n1470);
	nand (gm_n1477, gm_n101, gm_n69, in_10, gm_n139, gm_n138);
	nand (gm_n1478, gm_n69, gm_n62, gm_n41, gm_n53, gm_n51);
	nand (gm_n1479, gm_n109, gm_n370, gm_n45, gm_n224, gm_n349);
	nand (gm_n1480, gm_n1479, gm_n1478, gm_n1477);
	nand (gm_n1481, gm_n268, gm_n161, gm_n45);
	or (gm_n1482, in_14, gm_n62, gm_n41, gm_n1481, gm_n342);
	nor (gm_n1483, gm_n57, gm_n41, in_8, gm_n261, gm_n59);
	nand (gm_n1484, gm_n1483, gm_n69, in_13);
	nor (gm_n1485, gm_n219, gm_n351, gm_n45);
	nand (gm_n1486, gm_n69, gm_n62, in_12, gm_n1485, gm_n53);
	nand (gm_n1487, gm_n1486, gm_n1484, gm_n1482);
	nor (gm_n1488, gm_n1476, gm_n1457, gm_n1455, gm_n1487, gm_n1480);
	nor (gm_n1489, gm_n385, gm_n219, gm_n43, gm_n162, gm_n77);
	nor (gm_n1490, gm_n119, in_14, gm_n42, gm_n1226, gm_n143);
	nor (gm_n1491, in_14, gm_n42, in_9, gm_n366, gm_n108);
	nor (gm_n1492, gm_n1491, gm_n1490, gm_n1489);
	nor (gm_n1493, gm_n1138, gm_n84, gm_n69);
	nor (gm_n1494, gm_n177, in_14, gm_n42, gm_n419, gm_n302);
	nor (gm_n1495, gm_n69, gm_n42, gm_n70, gm_n177, gm_n82);
	nor (gm_n1496, gm_n1495, gm_n1494, gm_n1493);
	nand (gm_n1497, gm_n1488, gm_n1454, gm_n1453, gm_n1496, gm_n1492);
	or (gm_n1498, gm_n229, gm_n562, in_11, gm_n708);
	nand (gm_n1499, gm_n105, gm_n80, gm_n45, gm_n164, gm_n131);
	nand (gm_n1500, in_14, in_13, in_12, gm_n471, gm_n191);
	nand (gm_n1501, gm_n1500, gm_n1499, gm_n1498);
	or (gm_n1502, gm_n1360, gm_n261, gm_n154);
	nand (gm_n1503, in_14, gm_n62, in_12, gm_n651, gm_n98);
	nand (gm_n1504, in_14, gm_n42, in_9, gm_n586, gm_n345);
	nand (gm_n1505, gm_n1504, gm_n1503, gm_n1502);
	nor (gm_n1506, gm_n1497, gm_n1452, gm_n1451, gm_n1505, gm_n1501);
	nand (gm_n1507, gm_n255, gm_n183, gm_n45);
	nor (gm_n1508, gm_n69, in_13, gm_n41, gm_n1507, gm_n63);
	nand (gm_n1509, gm_n170, gm_n80, in_8);
	nor (gm_n1510, gm_n69, gm_n42, gm_n70, gm_n1509, gm_n108);
	nor (gm_n1511, in_14, in_13, gm_n41, gm_n256, gm_n71);
	nor (gm_n1512, gm_n1511, gm_n1510, gm_n1508);
	or (gm_n1513, gm_n216, gm_n41, in_8, gm_n201, gm_n208);
	nor (gm_n1514, gm_n1513, in_14, gm_n62);
	and (gm_n1515, gm_n133, gm_n104, in_8, gm_n191, gm_n183);
	and (gm_n1516, gm_n116, gm_n88, in_11, gm_n268, gm_n168);
	nor (gm_n1517, gm_n1516, gm_n1515, gm_n1514);
	nand (gm_n1518, gm_n1506, gm_n1450, gm_n1449, gm_n1517, gm_n1512);
	nand (gm_n1519, gm_n69, gm_n62, in_12, gm_n1057, gm_n349);
	or (gm_n1520, gm_n69, gm_n62, in_12, gm_n908, gm_n230);
	or (gm_n1521, gm_n782, gm_n882, gm_n43, gm_n563);
	nand (gm_n1522, gm_n1521, gm_n1520, gm_n1519);
	nand (gm_n1523, gm_n69, in_13, gm_n41, gm_n486, gm_n93);
	nand (gm_n1524, in_14, in_13, gm_n41, gm_n202, gm_n191);
	nand (gm_n1525, gm_n69, gm_n62, gm_n41, gm_n581, gm_n349);
	nand (gm_n1526, gm_n1525, gm_n1524, gm_n1523);
	nor (gm_n1527, gm_n1518, gm_n1448, gm_n1446, gm_n1526, gm_n1522);
	nor (gm_n1528, in_14, in_13, gm_n41, gm_n721, gm_n342);
	nor (gm_n1529, gm_n231, gm_n59, in_8);
	and (gm_n1530, gm_n69, gm_n62, gm_n41, gm_n1529, gm_n93);
	and (gm_n1531, gm_n559, gm_n129, gm_n43, gm_n295, gm_n183);
	nor (gm_n1532, gm_n1531, gm_n1530, gm_n1528);
	and (gm_n1533, gm_n199, gm_n65, gm_n45);
	and (gm_n1534, in_14, in_13, in_12, gm_n1533, gm_n131);
	nor (gm_n1535, gm_n562, gm_n154, in_11, gm_n241);
	nor (gm_n1536, gm_n69, gm_n62, gm_n41, gm_n715, gm_n63);
	nor (gm_n1537, gm_n1536, gm_n1535, gm_n1534);
	nand (gm_n1538, gm_n1527, gm_n1445, gm_n1444, gm_n1537, gm_n1532);
	nand (gm_n1539, gm_n174, gm_n169, gm_n43, gm_n311);
	nand (gm_n1540, gm_n178, gm_n172, in_14);
	nand (gm_n1541, gm_n1318, gm_n300, gm_n69);
	nand (gm_n1542, gm_n1541, gm_n1540, gm_n1539);
	nand (gm_n1543, in_14, in_13, gm_n41, gm_n459, gm_n98);
	nand (gm_n1544, gm_n69, gm_n42, in_9, gm_n426, gm_n83);
	or (gm_n1545, in_14, in_13, in_12, gm_n637, gm_n216);
	nand (gm_n1546, gm_n1545, gm_n1544, gm_n1543);
	nor (gm_n1547, gm_n1538, gm_n1443, gm_n1442, gm_n1546, gm_n1542);
	and (gm_n1548, in_14, in_13, gm_n41, gm_n478, gm_n131);
	nor (gm_n1549, in_14, in_13, in_12, gm_n414, gm_n71);
	nor (gm_n1550, in_14, gm_n42, in_9, gm_n1274, gm_n119);
	nor (gm_n1551, gm_n1550, gm_n1549, gm_n1548);
	nand (gm_n1552, gm_n53, gm_n41, in_8, gm_n81, gm_n72);
	nor (gm_n1553, gm_n1552, gm_n69, gm_n62);
	nor (gm_n1554, gm_n229, gm_n94, in_11, gm_n566, gm_n227);
	nor (gm_n1555, gm_n69, gm_n42, in_9, gm_n542, gm_n87);
	nor (gm_n1556, gm_n1555, gm_n1554, gm_n1553);
	nand (gm_n1557, gm_n1547, gm_n1440, gm_n1439, gm_n1556, gm_n1551);
	nor (gm_n1558, gm_n301, gm_n385, gm_n45);
	nand (gm_n1559, in_14, in_13, gm_n41, gm_n1558, gm_n98);
	or (gm_n1560, gm_n94, gm_n77, in_11, gm_n227, gm_n156);
	nand (gm_n1561, gm_n72, gm_n66, in_11, gm_n284, gm_n164);
	nand (gm_n1562, gm_n1561, gm_n1560, gm_n1559);
	or (gm_n1563, gm_n69, gm_n62, gm_n41, gm_n926, gm_n342);
	nand (gm_n1564, in_14, in_13, gm_n41, gm_n884, gm_n349);
	nand (gm_n1565, gm_n451, gm_n83, in_14);
	nand (gm_n1566, gm_n1565, gm_n1564, gm_n1563);
	nor (gm_n1567, gm_n1557, gm_n1437, gm_n1436, gm_n1566, gm_n1562);
	nor (gm_n1568, in_14, gm_n62, gm_n41, gm_n591, gm_n230);
	nor (gm_n1569, gm_n94, gm_n90, in_11, gm_n226, gm_n882);
	nor (gm_n1570, gm_n69, in_13, gm_n41, gm_n343, gm_n63);
	nor (gm_n1571, gm_n1570, gm_n1569, gm_n1568);
	and (gm_n1572, in_14, in_13, gm_n41, gm_n691, gm_n131);
	and (gm_n1573, in_14, in_13, gm_n41, gm_n599, gm_n126);
	and (gm_n1574, gm_n81, gm_n109, in_8);
	and (gm_n1575, gm_n69, gm_n62, gm_n41, gm_n1574, gm_n53);
	nor (gm_n1576, gm_n1575, gm_n1573, gm_n1572);
	nand (gm_n1577, gm_n1567, gm_n1434, gm_n1432, gm_n1576, gm_n1571);
	nand (gm_n1578, gm_n117, gm_n65, gm_n43, gm_n266, gm_n184);
	nand (gm_n1579, gm_n69, in_13, gm_n41, gm_n1574, gm_n44);
	or (gm_n1580, in_14, in_13, gm_n41, gm_n1360, gm_n71);
	nand (gm_n1581, gm_n1580, gm_n1579, gm_n1578);
	or (gm_n1582, gm_n84, gm_n69, gm_n42, gm_n145, gm_n121);
	and (gm_n1583, gm_n44, in_12, gm_n45, gm_n80, gm_n73);
	nand (gm_n1584, gm_n1583, in_14, gm_n62);
	and (gm_n1585, gm_n53, in_12, in_8, gm_n255, gm_n109);
	nand (gm_n1586, gm_n1585, gm_n69, gm_n62);
	nand (gm_n1587, gm_n1586, gm_n1584, gm_n1582);
	nor (out_10, gm_n1581, gm_n1577, gm_n1431, gm_n1587);
	and (gm_n1589, in_14, gm_n62, in_12, gm_n1000, gm_n98);
	nand (gm_n1590, gm_n69, in_13, gm_n41, gm_n1529, gm_n53);
	and (gm_n1591, gm_n80, in_12, in_8, gm_n268, gm_n191);
	nand (gm_n1592, gm_n1591, in_14, in_13);
	or (gm_n1593, gm_n47, in_12, gm_n45, gm_n201, gm_n216);
	nor (gm_n1594, gm_n1593, in_14, gm_n62);
	nor (gm_n1595, in_14, gm_n42, gm_n70, gm_n1313, gm_n119);
	nand (gm_n1596, gm_n345, in_14, in_10, gm_n1130, gm_n289);
	nand (gm_n1597, gm_n88, gm_n66, gm_n43, gm_n224, gm_n116);
	and (gm_n1598, in_14, in_10, in_9, gm_n340, gm_n101);
	and (gm_n1599, in_14, in_13, gm_n41, gm_n1057, gm_n44);
	or (gm_n1600, in_14, in_13, in_12, gm_n642, gm_n261);
	nand (gm_n1601, gm_n161, gm_n243, gm_n43, gm_n233, gm_n720);
	and (gm_n1602, in_14, in_13, in_12, gm_n459, gm_n126);
	nor (gm_n1603, gm_n84, in_14, in_10, gm_n307, gm_n305);
	nand (gm_n1604, gm_n69, gm_n62, gm_n41, gm_n664, gm_n126);
	nand (gm_n1605, gm_n69, gm_n42, gm_n70, gm_n1533, gm_n178);
	and (gm_n1606, gm_n86, in_14, in_10, gm_n840, gm_n741);
	nand (gm_n1607, gm_n42, gm_n70, gm_n45, gm_n129, gm_n72);
	nor (gm_n1608, gm_n1607, gm_n119, gm_n69);
	nand (gm_n1609, gm_n66, gm_n65, in_8, gm_n168, gm_n93);
	nand (gm_n1610, gm_n105, gm_n72, gm_n45, gm_n295, gm_n191);
	nand (gm_n1611, gm_n46, in_12, in_8, gm_n129, gm_n53);
	nor (gm_n1612, gm_n1611, gm_n69, in_13);
	nor (gm_n1613, gm_n177, in_14, gm_n42, gm_n287, gm_n286);
	nand (gm_n1614, gm_n105, gm_n109, gm_n45);
	or (gm_n1615, in_14, in_13, in_12, gm_n1614, gm_n216);
	or (gm_n1616, gm_n69, gm_n62, in_12, gm_n1339, gm_n76);
	nand (gm_n1617, gm_n46, gm_n41, in_8, gm_n277, gm_n93);
	nor (gm_n1618, gm_n1617, in_14, gm_n62);
	nor (gm_n1619, in_14, gm_n62, gm_n41, gm_n628, gm_n76);
	nor (gm_n1620, gm_n122, gm_n69, gm_n42, gm_n790, gm_n177);
	nor (gm_n1621, gm_n69, in_13, in_12, gm_n1202, gm_n63);
	and (gm_n1622, gm_n370, gm_n46, gm_n43, gm_n106, gm_n243);
	nor (gm_n1623, gm_n1620, gm_n1619, gm_n1618, gm_n1622, gm_n1621);
	nor (gm_n1624, in_14, in_10, gm_n70, gm_n521, gm_n119);
	and (gm_n1625, gm_n69, gm_n62, in_12, gm_n318, gm_n349);
	nor (gm_n1626, in_14, gm_n62, gm_n41, gm_n871, gm_n342);
	nor (gm_n1627, gm_n1626, gm_n1625, gm_n1624);
	and (gm_n1628, gm_n69, gm_n62, in_12, gm_n581, gm_n126);
	and (gm_n1629, in_14, in_13, gm_n41, gm_n1107, gm_n349);
	nor (gm_n1630, in_14, gm_n62, gm_n41, gm_n844, gm_n76);
	nor (gm_n1631, gm_n1630, gm_n1629, gm_n1628);
	nand (gm_n1632, gm_n1623, gm_n1616, gm_n1615, gm_n1631, gm_n1627);
	nand (gm_n1633, gm_n115, gm_n104, in_11, gm_n266);
	or (gm_n1634, gm_n69, in_13, in_12, gm_n500, gm_n327);
	nand (gm_n1635, gm_n69, in_13, gm_n41, gm_n196, gm_n98);
	nand (gm_n1636, gm_n1635, gm_n1634, gm_n1633);
	nand (gm_n1637, gm_n86, gm_n69, gm_n42, gm_n840, gm_n212);
	nand (gm_n1638, gm_n69, gm_n62, in_12, gm_n202, gm_n131);
	nand (gm_n1639, gm_n69, in_13, in_12, gm_n126, gm_n505);
	nand (gm_n1640, gm_n1639, gm_n1638, gm_n1637);
	nor (gm_n1641, gm_n1632, gm_n1613, gm_n1612, gm_n1640, gm_n1636);
	nor (gm_n1642, in_14, gm_n62, in_12, gm_n414, gm_n71);
	nand (gm_n1643, gm_n133, gm_n161, in_8);
	nor (gm_n1644, in_14, in_13, in_12, gm_n1643, gm_n230);
	nor (gm_n1645, in_14, in_13, in_12, gm_n1274, gm_n63);
	nor (gm_n1646, gm_n1645, gm_n1644, gm_n1642);
	nor (gm_n1647, gm_n69, gm_n62, in_12, gm_n721, gm_n327);
	nor (gm_n1648, gm_n69, gm_n42, in_9, gm_n446, gm_n108);
	nor (gm_n1649, gm_n249, gm_n351, in_14, gm_n201, gm_n417);
	nor (gm_n1650, gm_n1649, gm_n1648, gm_n1647);
	nand (gm_n1651, gm_n1641, gm_n1610, gm_n1609, gm_n1650, gm_n1646);
	nand (gm_n1652, gm_n720, gm_n161, gm_n43, gm_n169, gm_n104);
	nand (gm_n1653, gm_n245, gm_n69, gm_n42, gm_n346, gm_n139);
	or (gm_n1654, gm_n145, gm_n69, in_10, gm_n305, gm_n271);
	nand (gm_n1655, gm_n1654, gm_n1653, gm_n1652);
	nand (gm_n1656, in_14, gm_n62, in_12, gm_n677, gm_n349);
	nand (gm_n1657, gm_n168, gm_n106, in_11, gm_n631);
	or (gm_n1658, gm_n156, gm_n77, in_11, gm_n503);
	nand (gm_n1659, gm_n1658, gm_n1657, gm_n1656);
	nor (gm_n1660, gm_n1651, gm_n1608, gm_n1606, gm_n1659, gm_n1655);
	nor (gm_n1661, in_14, in_13, in_12, gm_n1043, gm_n63);
	nor (gm_n1662, gm_n562, gm_n351, gm_n43, gm_n201, gm_n827);
	and (gm_n1663, gm_n81, gm_n80, in_8, gm_n131, gm_n104);
	nor (gm_n1664, gm_n1663, gm_n1662, gm_n1661);
	and (gm_n1665, gm_n88, gm_n83, in_14, gm_n255, gm_n116);
	and (gm_n1666, gm_n139, in_14, gm_n42, gm_n840, gm_n300);
	or (gm_n1667, in_10, in_9, in_8, gm_n59, gm_n57);
	nor (gm_n1668, gm_n1667, gm_n417, gm_n69);
	nor (gm_n1669, gm_n1668, gm_n1666, gm_n1665);
	nand (gm_n1670, gm_n1660, gm_n1605, gm_n1604, gm_n1669, gm_n1664);
	nand (gm_n1671, gm_n73, gm_n65, in_11, gm_n266, gm_n224);
	or (gm_n1672, gm_n417, in_14, in_10, gm_n1226, gm_n419);
	nand (gm_n1673, gm_n116, gm_n43, gm_n58, gm_n1243, gm_n224);
	nand (gm_n1674, gm_n1673, gm_n1672, gm_n1671);
	and (gm_n1675, gm_n69, gm_n62, in_12, gm_n318, gm_n44);
	and (gm_n1676, gm_n66, gm_n41, in_8, gm_n191, gm_n161);
	and (gm_n1677, gm_n1676, gm_n69, in_13);
	or (gm_n1678, gm_n1677, gm_n1675, gm_n1451);
	nor (gm_n1679, gm_n1670, gm_n1603, gm_n1602, gm_n1678, gm_n1674);
	nor (gm_n1680, in_14, gm_n42, gm_n70, gm_n1313, gm_n177);
	and (gm_n1681, gm_n106, gm_n161, gm_n43, gm_n174, gm_n129);
	nor (gm_n1682, gm_n84, gm_n69, in_10, gm_n307, gm_n143);
	nor (gm_n1683, gm_n1682, gm_n1681, gm_n1680);
	nor (gm_n1684, gm_n84, in_14, in_10, gm_n305, gm_n467);
	nor (gm_n1685, gm_n108, gm_n59, in_14, gm_n566, gm_n227);
	nand (gm_n1686, gm_n46, gm_n41, gm_n45, gm_n277, gm_n93);
	nor (gm_n1687, gm_n1686, in_14, in_13);
	nor (gm_n1688, gm_n1687, gm_n1685, gm_n1684);
	nand (gm_n1689, gm_n1679, gm_n1601, gm_n1600, gm_n1688, gm_n1683);
	nand (gm_n1690, gm_n69, gm_n62, in_12, gm_n681, gm_n93);
	nand (gm_n1691, gm_n83, in_14, in_10, gm_n323, gm_n144);
	nand (gm_n1692, in_14, gm_n62, in_12, gm_n681, gm_n349);
	nand (gm_n1693, gm_n1692, gm_n1691, gm_n1690);
	nand (gm_n1694, gm_n69, in_10, gm_n70, gm_n1175, gm_n101);
	nand (gm_n1695, gm_n69, in_13, in_12, gm_n1558, gm_n191);
	nand (gm_n1696, gm_n490, gm_n101, in_14);
	nand (gm_n1697, gm_n1696, gm_n1695, gm_n1694);
	nor (gm_n1698, gm_n1689, gm_n1599, gm_n1598, gm_n1697, gm_n1693);
	nor (gm_n1699, gm_n1435, gm_n84, gm_n69);
	nor (gm_n1700, gm_n69, gm_n62, gm_n41, gm_n1339, gm_n71);
	nor (gm_n1701, gm_n87, gm_n351, gm_n69, gm_n249, gm_n95);
	nor (gm_n1702, gm_n1701, gm_n1700, gm_n1699);
	and (gm_n1703, gm_n69, gm_n62, gm_n41, gm_n760, gm_n191);
	nor (gm_n1704, in_14, in_13, in_12, gm_n442);
	nor (gm_n1705, in_14, gm_n62, gm_n41, gm_n844, gm_n71);
	nor (gm_n1706, gm_n1705, gm_n1704, gm_n1703);
	nand (gm_n1707, gm_n1698, gm_n1597, gm_n1596, gm_n1706, gm_n1702);
	nand (gm_n1708, gm_n245, in_14, in_10, gm_n289, gm_n258);
	or (gm_n1709, in_14, in_10, gm_n70, gm_n609, gm_n108);
	nand (gm_n1710, gm_n73, gm_n109, in_8);
	or (gm_n1711, gm_n69, gm_n62, gm_n41, gm_n1710, gm_n342);
	nand (gm_n1712, gm_n1711, gm_n1709, gm_n1708);
	nand (gm_n1713, gm_n69, gm_n62, gm_n41, gm_n432, gm_n98);
	and (gm_n1714, gm_n42, gm_n79, gm_n64, gm_n277, gm_n144);
	nand (gm_n1715, gm_n1714, gm_n86, in_14);
	nand (gm_n1716, gm_n69, in_13, in_12, gm_n488, gm_n93);
	nand (gm_n1717, gm_n1716, gm_n1715, gm_n1713);
	nor (gm_n1718, gm_n1707, gm_n1595, gm_n1594, gm_n1717, gm_n1712);
	and (gm_n1719, gm_n277, gm_n80, gm_n45);
	and (gm_n1720, gm_n69, in_13, in_12, gm_n1719, gm_n44);
	and (gm_n1721, gm_n69, gm_n42, gm_n70, gm_n300, gm_n179);
	nor (gm_n1722, gm_n417, gm_n69, in_10, gm_n419, gm_n307);
	nor (gm_n1723, gm_n1722, gm_n1721, gm_n1720);
	nor (gm_n1724, gm_n84, gm_n69, in_10, gm_n467, gm_n121);
	and (gm_n1725, gm_n178, gm_n73, in_14, gm_n266, gm_n183);
	nand (gm_n1726, gm_n133, gm_n80, gm_n45);
	nor (gm_n1727, in_14, in_10, gm_n70, gm_n1726, gm_n108);
	nor (gm_n1728, gm_n1727, gm_n1725, gm_n1724);
	nand (gm_n1729, gm_n1718, gm_n1592, gm_n1590, gm_n1728, gm_n1723);
	nand (gm_n1730, gm_n69, in_13, gm_n41, gm_n1558, gm_n44);
	nor (gm_n1731, gm_n385, in_12, gm_n45, gm_n193, gm_n342);
	nand (gm_n1732, gm_n1731, gm_n69, gm_n62);
	nand (gm_n1733, gm_n1732, gm_n1730, gm_n409);
	nand (gm_n1734, gm_n183, gm_n168, gm_n43, gm_n268, gm_n284);
	nand (gm_n1735, gm_n66, gm_n65, in_8, gm_n224, gm_n93);
	or (gm_n1736, gm_n69, in_13, in_12, gm_n1313, gm_n71);
	nand (gm_n1737, gm_n1736, gm_n1735, gm_n1734);
	nor (out_11, gm_n1733, gm_n1729, gm_n1589, gm_n1737);
	nor (gm_n1739, gm_n1607, gm_n417, gm_n69);
	nor (gm_n1740, in_14, gm_n62, gm_n41, gm_n968, gm_n216);
	nand (gm_n1741, gm_n69, in_13, in_12, gm_n575, gm_n126);
	nand (gm_n1742, in_14, in_13, gm_n41, gm_n1485, gm_n131);
	nor (gm_n1743, gm_n122, gm_n69, in_10, gm_n287, gm_n239);
	nor (gm_n1744, gm_n108, gm_n351, in_14, gm_n201, gm_n646);
	or (gm_n1745, gm_n119, gm_n69, in_10, gm_n286, gm_n237);
	nor (gm_n1746, gm_n69, in_13, gm_n41, gm_n360, gm_n71);
	nor (gm_n1747, gm_n162, gm_n59, in_11, gm_n225, gm_n396);
	and (gm_n1748, gm_n243, gm_n65, gm_n43, gm_n106, gm_n105);
	and (gm_n1749, gm_n245, gm_n69, in_10, gm_n1130, gm_n212);
	or (gm_n1750, gm_n1747, gm_n1746, t_1, gm_n1749, gm_n1748);
	nand (gm_n1751, gm_n46, gm_n41, gm_n45, gm_n191, gm_n158);
	nor (gm_n1752, gm_n1751, gm_n69, gm_n62);
	and (gm_n1753, gm_n104, gm_n161, gm_n43, gm_n169, gm_n129);
	and (gm_n1754, gm_n69, in_13, in_12, gm_n185, gm_n131);
	nor (gm_n1755, gm_n1753, gm_n1752, gm_n1750, gm_n1754);
	nand (gm_n1756, gm_n138, in_14, gm_n42, gm_n345, gm_n144);
	nand (gm_n1757, in_14, in_13, in_12, gm_n209, gm_n349);
	nand (gm_n1758, gm_n243, gm_n109, in_11, gm_n246, gm_n284);
	nand (gm_n1759, gm_n1756, gm_n1755, gm_n1745, gm_n1758, gm_n1757);
	or (gm_n1760, gm_n69, gm_n62, in_12, gm_n1726, gm_n216);
	nor (gm_n1761, gm_n147, gm_n351, in_8);
	nand (gm_n1762, gm_n69, in_13, in_12, gm_n1761, gm_n131);
	or (gm_n1763, gm_n1234, gm_n417, in_14);
	nand (gm_n1764, gm_n1763, gm_n1762, gm_n1760);
	or (gm_n1765, in_14, gm_n62, gm_n41, gm_n388, gm_n63);
	or (gm_n1766, gm_n417, in_14, gm_n42, gm_n1226, gm_n536);
	nand (gm_n1767, gm_n559, gm_n117, in_11, gm_n655);
	nand (gm_n1768, gm_n1767, gm_n1766, gm_n1765);
	nor (gm_n1769, gm_n1759, gm_n1744, gm_n1743, gm_n1768, gm_n1764);
	nor (gm_n1770, gm_n87, in_14, gm_n42, gm_n305, gm_n418);
	nor (gm_n1771, gm_n646, gm_n963, in_11, gm_n708);
	and (gm_n1772, gm_n117, gm_n106, in_11, gm_n311);
	nor (gm_n1773, gm_n1772, gm_n1771, gm_n1770);
	and (gm_n1774, gm_n86, in_14, in_10, gm_n346, gm_n212);
	nand (gm_n1775, gm_n349, in_12, gm_n45, gm_n184, gm_n161);
	nor (gm_n1776, gm_n1775, gm_n69, gm_n62);
	and (gm_n1777, in_14, gm_n62, gm_n41, gm_n1105, gm_n126);
	nor (gm_n1778, gm_n1777, gm_n1776, gm_n1774);
	nand (gm_n1779, gm_n1769, gm_n1742, gm_n1741, gm_n1778, gm_n1773);
	nand (gm_n1780, in_14, gm_n62, in_12, gm_n480, gm_n191);
	nand (gm_n1781, gm_n605, gm_n83, gm_n69);
	nand (gm_n1782, gm_n93, gm_n72, in_8, gm_n246, gm_n164);
	nand (gm_n1783, gm_n1782, gm_n1781, gm_n1780);
	or (gm_n1784, in_14, in_10, gm_n70, gm_n540, gm_n84);
	nand (gm_n1785, gm_n1784, gm_n1601, gm_n1145);
	nor (out_12, gm_n1779, gm_n1740, gm_n1739, gm_n1785, gm_n1783);
	and (gm_n1787, gm_n131, gm_n117, gm_n45, gm_n381, gm_n183);
	or (gm_n1788, gm_n69, gm_n62, in_12, gm_n414, gm_n76);
	or (gm_n1789, in_14, gm_n42, gm_n70, gm_n1360, gm_n239);
	nand (gm_n1790, gm_n109, in_12, gm_n45, gm_n191, gm_n73);
	nor (gm_n1791, gm_n1790, in_14, gm_n62);
	and (gm_n1792, gm_n72, gm_n53, gm_n45, gm_n104, gm_n720);
	and (gm_n1793, gm_n349, gm_n41, gm_n45, gm_n246, gm_n161);
	nand (gm_n1794, gm_n1793, gm_n69, in_13);
	nand (gm_n1795, gm_n124, gm_n109, in_11, gm_n295, gm_n233);
	nor (gm_n1796, gm_n69, in_10, in_9, gm_n1394, gm_n119);
	nor (gm_n1797, in_7, gm_n79, gm_n64, gm_n189, in_8);
	and (gm_n1798, gm_n69, gm_n62, gm_n41, gm_n1797, gm_n44);
	nand (gm_n1799, gm_n69, gm_n62, in_12, gm_n1447, gm_n53);
	nand (gm_n1800, in_14, gm_n62, gm_n41, gm_n973, gm_n126);
	and (gm_n1801, gm_n178, gm_n72, gm_n69, gm_n266, gm_n199);
	nor (gm_n1802, gm_n69, in_10, in_9, gm_n417, gm_n134);
	or (gm_n1803, in_14, gm_n62, gm_n41, gm_n217, gm_n216);
	nand (gm_n1804, in_14, gm_n62, in_12, gm_n549, gm_n349);
	nor (gm_n1805, in_14, gm_n62, in_12, gm_n360, gm_n63);
	nor (gm_n1806, gm_n69, in_13, gm_n41, gm_n529, gm_n63);
	or (gm_n1807, gm_n145, in_14, gm_n42, gm_n237, gm_n177);
	nand (gm_n1808, gm_n69, in_10, in_9, gm_n340, gm_n345);
	and (gm_n1809, gm_n106, gm_n43, in_7, gm_n164, gm_n138);
	nor (gm_n1810, in_14, gm_n62, in_12, gm_n701, gm_n327);
	nand (gm_n1811, gm_n69, gm_n62, gm_n41, gm_n1354, gm_n191);
	nand (gm_n1812, in_14, gm_n62, in_12, gm_n757, gm_n191);
	nor (gm_n1813, in_14, gm_n62, gm_n41, gm_n642, gm_n342);
	nor (gm_n1814, in_14, gm_n62, gm_n41, gm_n442);
	nor (gm_n1815, gm_n225, gm_n162, in_11, gm_n563);
	and (gm_n1816, gm_n184, gm_n80, in_8);
	and (gm_n1817, gm_n69, in_13, in_12, gm_n1816, gm_n44);
	and (gm_n1818, gm_n93, gm_n72, in_8, gm_n246, gm_n104);
	nor (gm_n1819, gm_n1815, gm_n1814, gm_n1813, gm_n1818, gm_n1817);
	or (gm_n1820, gm_n58, in_6, in_5, gm_n189, gm_n45);
	nor (gm_n1821, gm_n69, gm_n62, in_12, gm_n1820, gm_n71);
	nor (gm_n1822, gm_n646, gm_n229, gm_n43, gm_n593);
	nor (gm_n1823, gm_n280, gm_n94, in_14, gm_n177, gm_n156);
	nor (gm_n1824, gm_n1823, gm_n1822, gm_n1821);
	nor (gm_n1825, gm_n1667, gm_n271, gm_n69);
	and (gm_n1826, gm_n117, gm_n72, in_8, gm_n246, gm_n126);
	nor (gm_n1827, in_14, in_13, in_12, gm_n644, gm_n261);
	nor (gm_n1828, gm_n1827, gm_n1826, gm_n1825);
	nand (gm_n1829, gm_n1819, gm_n1812, gm_n1811, gm_n1828, gm_n1824);
	nand (gm_n1830, gm_n42, in_9, gm_n45, gm_n274, gm_n72);
	or (gm_n1831, gm_n1830, gm_n119, in_14);
	nand (gm_n1832, gm_n164, gm_n88, in_11, gm_n268, gm_n233);
	or (gm_n1833, gm_n90, gm_n385, in_14, gm_n177, gm_n249);
	nand (gm_n1834, gm_n1833, gm_n1832, gm_n1831);
	nand (gm_n1835, gm_n83, gm_n69, in_10, gm_n258, gm_n144);
	nand (gm_n1836, in_14, in_13, in_12, gm_n1719, gm_n349);
	nand (gm_n1837, gm_n1836, gm_n1835, gm_n445);
	nor (gm_n1838, gm_n1829, gm_n1810, gm_n1809, gm_n1837, gm_n1834);
	nor (gm_n1839, gm_n69, in_13, gm_n41, gm_n806, gm_n342);
	nor (gm_n1840, in_14, gm_n62, gm_n41, gm_n1471, gm_n63);
	nand (gm_n1841, gm_n370, in_12, in_8, gm_n191, gm_n88);
	nor (gm_n1842, gm_n1841, gm_n69, gm_n62);
	nor (gm_n1843, gm_n1842, gm_n1840, gm_n1839);
	nor (gm_n1844, gm_n1188, gm_n108, gm_n69);
	nor (gm_n1845, gm_n119, in_14, gm_n42, gm_n287, gm_n418);
	nor (gm_n1846, gm_n119, gm_n69, gm_n42, gm_n419, gm_n302);
	nor (gm_n1847, gm_n1846, gm_n1845, gm_n1844);
	nand (gm_n1848, gm_n1838, gm_n1808, gm_n1807, gm_n1847, gm_n1843);
	or (gm_n1849, in_14, gm_n42, in_9, gm_n377, gm_n119);
	nand (gm_n1850, gm_n320, gm_n109, in_11, gm_n168, gm_n116);
	nand (gm_n1851, gm_n69, gm_n62, in_12, gm_n1046, gm_n131);
	nand (gm_n1852, gm_n1851, gm_n1850, gm_n1849);
	nor (gm_n1853, gm_n208, gm_n50, in_8);
	nand (gm_n1854, gm_n69, in_13, gm_n41, gm_n1853, gm_n53);
	nand (gm_n1855, gm_n69, in_13, in_12, gm_n588, gm_n53);
	nand (gm_n1856, gm_n1855, gm_n1854, gm_n363);
	nor (gm_n1857, gm_n1848, gm_n1806, gm_n1805, gm_n1856, gm_n1852);
	nor (gm_n1858, gm_n69, in_10, gm_n70, gm_n609, gm_n239);
	nor (gm_n1859, gm_n69, in_10, gm_n70, gm_n715, gm_n108);
	nor (gm_n1860, gm_n69, in_13, gm_n41, gm_n293, gm_n216);
	nor (gm_n1861, gm_n1860, gm_n1859, gm_n1858);
	nor (gm_n1862, gm_n69, gm_n62, in_12, gm_n1320, gm_n342);
	nor (gm_n1863, in_14, gm_n62, gm_n41, gm_n521, gm_n63);
	and (gm_n1864, gm_n69, in_13, in_12, gm_n831, gm_n53);
	nor (gm_n1865, gm_n1864, gm_n1863, gm_n1862);
	nand (gm_n1866, gm_n1857, gm_n1804, gm_n1803, gm_n1865, gm_n1861);
	or (gm_n1867, in_14, gm_n42, in_9, gm_n987, gm_n239);
	nand (gm_n1868, gm_n69, gm_n62, gm_n41, gm_n99, gm_n44);
	nand (gm_n1869, gm_n163, gm_n72, in_11, gm_n224, gm_n199);
	nand (gm_n1870, gm_n1869, gm_n1868, gm_n1867);
	or (gm_n1871, gm_n150, gm_n57, gm_n69, gm_n646, gm_n108);
	or (gm_n1872, in_14, in_13, gm_n41, gm_n542, gm_n342);
	nand (gm_n1873, gm_n69, in_13, in_12, gm_n202, gm_n98);
	nand (gm_n1874, gm_n1873, gm_n1872, gm_n1871);
	nor (gm_n1875, gm_n1866, gm_n1802, gm_n1801, gm_n1874, gm_n1870);
	nor (gm_n1876, in_14, gm_n62, in_12, gm_n1643, gm_n327);
	nor (gm_n1877, in_14, gm_n62, in_12, gm_n1043, gm_n71);
	nor (gm_n1878, gm_n827, gm_n249, gm_n43, gm_n593);
	nor (gm_n1879, gm_n1878, gm_n1877, gm_n1876);
	and (gm_n1880, in_14, gm_n62, in_12, gm_n426, gm_n191);
	and (gm_n1881, gm_n69, in_10, gm_n70, gm_n179, gm_n136);
	nor (gm_n1882, in_14, in_13, gm_n41, gm_n1509, gm_n71);
	nor (gm_n1883, gm_n1882, gm_n1881, gm_n1880);
	nand (gm_n1884, gm_n1875, gm_n1800, gm_n1799, gm_n1883, gm_n1879);
	nand (gm_n1885, gm_n101, gm_n88, gm_n69, gm_n169, gm_n110);
	nand (gm_n1886, gm_n163, gm_n104, in_11, gm_n631);
	and (gm_n1887, gm_n46, gm_n41, gm_n45, gm_n184, gm_n98);
	nand (gm_n1888, gm_n1887, in_14, in_13);
	nand (gm_n1889, gm_n1888, gm_n1886, gm_n1885);
	or (gm_n1890, gm_n87, in_14, gm_n42, gm_n790, gm_n467);
	nand (gm_n1891, in_14, in_13, in_12, gm_n773, gm_n126);
	nor (gm_n1892, gm_n47, in_12, gm_n45, gm_n216, gm_n57);
	nand (gm_n1893, gm_n1892, in_14, gm_n62);
	nand (gm_n1894, gm_n1893, gm_n1891, gm_n1890);
	nor (gm_n1895, gm_n1884, gm_n1798, gm_n1796, gm_n1894, gm_n1889);
	nor (gm_n1896, gm_n177, gm_n91, gm_n69);
	nor (gm_n1897, gm_n69, in_13, in_12, gm_n1271, gm_n216);
	or (gm_n1898, gm_n89, gm_n41, gm_n45, gm_n231, gm_n327);
	nor (gm_n1899, gm_n1898, gm_n69, gm_n62);
	nor (gm_n1900, gm_n1899, gm_n1897, gm_n1896);
	nor (gm_n1901, gm_n646, gm_n77, gm_n43, gm_n563);
	nor (gm_n1902, gm_n69, gm_n62, in_12, gm_n377, gm_n342);
	or (gm_n1903, gm_n201, gm_n94, gm_n45);
	nor (gm_n1904, gm_n69, gm_n62, in_12, gm_n1903, gm_n63);
	nor (gm_n1905, gm_n1904, gm_n1902, gm_n1901);
	nand (gm_n1906, gm_n1895, gm_n1795, gm_n1794, gm_n1905, gm_n1900);
	nand (gm_n1907, gm_n784, gm_n345, gm_n69);
	nand (gm_n1908, in_14, gm_n62, in_12, gm_n1105, gm_n53);
	or (gm_n1909, gm_n249, gm_n89, in_11, gm_n193, gm_n882);
	nand (gm_n1910, gm_n1909, gm_n1908, gm_n1907);
	nor (gm_n1911, gm_n239, gm_n69, in_10, gm_n330, gm_n307);
	and (gm_n1912, gm_n72, gm_n66, gm_n43, gm_n266, gm_n243);
	or (gm_n1913, gm_n1912, gm_n1911, gm_n1210);
	nor (gm_n1914, gm_n1906, gm_n1792, gm_n1791, gm_n1913, gm_n1910);
	nand (gm_n1915, gm_n370, gm_n41, gm_n45, gm_n98, gm_n72);
	nor (gm_n1916, gm_n1915, gm_n69, gm_n62);
	and (gm_n1917, gm_n136, gm_n80, gm_n69, gm_n255, gm_n233);
	nor (gm_n1918, gm_n782, gm_n77, in_11, gm_n708);
	nor (gm_n1919, gm_n1918, gm_n1917, gm_n1916);
	nor (gm_n1920, gm_n69, in_10, in_9, gm_n595, gm_n108);
	nand (gm_n1921, gm_n44, gm_n41, in_8, gm_n246, gm_n72);
	nor (gm_n1922, gm_n1921, gm_n69, in_13);
	nor (gm_n1923, gm_n69, gm_n62, gm_n41, gm_n1507, gm_n71);
	nor (gm_n1924, gm_n1923, gm_n1922, gm_n1920);
	nand (gm_n1925, gm_n1914, gm_n1789, gm_n1788, gm_n1924, gm_n1919);
	nand (gm_n1926, gm_n69, in_13, in_12, gm_n1038, gm_n191);
	nand (gm_n1927, gm_n170, gm_n109, in_14, gm_n345, gm_n266);
	nand (gm_n1928, gm_n178, gm_n69, in_10, gm_n840, gm_n943);
	nand (gm_n1929, gm_n1928, gm_n1927, gm_n1926);
	nand (gm_n1930, gm_n720, gm_n65, gm_n43, gm_n233, gm_n168);
	or (gm_n1931, gm_n1251, gm_n271, in_14);
	nand (gm_n1932, gm_n69, in_13, gm_n41, gm_n181, gm_n53);
	nand (gm_n1933, gm_n1932, gm_n1931, gm_n1930);
	nor (out_13, gm_n1929, gm_n1925, gm_n1787, gm_n1933);
	and (gm_n1935, gm_n93, gm_n66, in_8, gm_n168, gm_n161);
	nand (gm_n1936, gm_n245, in_14, in_10, gm_n329, gm_n144);
	nand (gm_n1937, gm_n183, gm_n73, gm_n69, gm_n266, gm_n300);
	nor (gm_n1938, in_14, in_10, gm_n70, gm_n1394, gm_n108);
	nand (gm_n1939, gm_n72, gm_n41, gm_n45, gm_n246, gm_n98);
	nor (gm_n1940, gm_n1939, in_14, gm_n62);
	nand (gm_n1941, gm_n345, in_14, in_10, gm_n741, gm_n329);
	nand (gm_n1942, in_14, in_13, gm_n41, gm_n1046, gm_n126);
	nand (gm_n1943, gm_n80, gm_n41, gm_n45, gm_n158, gm_n131);
	nor (gm_n1944, gm_n1943, in_14, in_13);
	and (gm_n1945, gm_n93, gm_n243, gm_n45, gm_n246, gm_n161);
	nand (gm_n1946, gm_n69, gm_n62, gm_n41, gm_n1797, gm_n53);
	or (gm_n1947, gm_n69, gm_n62, gm_n41, gm_n901, gm_n63);
	and (gm_n1948, gm_n69, gm_n62, in_12, gm_n1853, gm_n191);
	and (gm_n1949, gm_n243, gm_n72, gm_n43, gm_n184, gm_n163);
	nand (gm_n1950, in_14, in_13, in_12, gm_n397, gm_n53);
	nand (gm_n1951, gm_n69, in_10, in_9, gm_n345, gm_n99);
	nor (gm_n1952, gm_n69, gm_n62, gm_n41, gm_n1394, gm_n63);
	nor (gm_n1953, gm_n1830, gm_n108, in_14);
	nand (gm_n1954, in_14, in_13, in_12, gm_n823, gm_n53);
	nand (gm_n1955, gm_n69, gm_n62, gm_n41, gm_n1101, gm_n349);
	nor (gm_n1956, gm_n162, gm_n84, in_14, gm_n533);
	and (gm_n1957, gm_n136, in_14, in_10, gm_n258, gm_n144);
	nand (gm_n1958, gm_n116, in_11, gm_n58, gm_n937, gm_n164);
	nand (gm_n1959, gm_n136, in_14, in_10, gm_n289, gm_n258);
	and (gm_n1960, in_14, in_13, in_12, gm_n555, gm_n126);
	and (gm_n1961, gm_n98, gm_n72, gm_n45, gm_n224, gm_n170);
	nor (gm_n1962, in_14, gm_n62, in_12, gm_n1710, gm_n230);
	nor (gm_n1963, gm_n69, gm_n62, in_12, gm_n364, gm_n261);
	nor (gm_n1964, in_14, gm_n62, in_12, gm_n1614, gm_n63);
	nor (gm_n1965, gm_n1962, gm_n1961, gm_n1960, gm_n1964, gm_n1963);
	and (gm_n1966, gm_n88, gm_n81, in_11, gm_n169, gm_n117);
	nand (gm_n1967, gm_n58, gm_n79, in_5, gm_n124, in_8);
	nor (gm_n1968, gm_n69, gm_n62, gm_n41, gm_n1967, gm_n63);
	nor (gm_n1969, in_14, gm_n62, gm_n41, gm_n446, gm_n216);
	nor (gm_n1970, gm_n1969, gm_n1968, gm_n1966);
	nor (gm_n1971, in_14, in_13, in_12, gm_n820, gm_n76);
	nor (gm_n1972, gm_n385, gm_n57, in_8, gm_n229, gm_n261);
	nor (gm_n1973, gm_n69, in_10, gm_n70, gm_n1726, gm_n87);
	nor (gm_n1974, gm_n1973, gm_n1972, gm_n1971);
	nand (gm_n1975, gm_n1965, gm_n1959, gm_n1958, gm_n1974, gm_n1970);
	nand (gm_n1976, in_14, gm_n62, gm_n41, gm_n732, gm_n126);
	nand (gm_n1977, gm_n69, gm_n62, in_12, gm_n1485, gm_n126);
	nand (gm_n1978, gm_n169, gm_n243, in_11, gm_n631);
	nand (gm_n1979, gm_n1978, gm_n1977, gm_n1976);
	nand (gm_n1980, gm_n266, gm_n164, gm_n43, gm_n373);
	and (gm_n1981, gm_n88, in_12, gm_n45, gm_n158, gm_n93);
	nand (gm_n1982, gm_n1981, in_14, in_13);
	nand (gm_n1983, gm_n69, in_13, gm_n41, gm_n1816, gm_n349);
	nand (gm_n1984, gm_n1983, gm_n1982, gm_n1980);
	nor (gm_n1985, gm_n1975, gm_n1957, gm_n1956, gm_n1984, gm_n1979);
	nor (gm_n1986, gm_n84, gm_n69, gm_n42, gm_n615, gm_n307);
	and (gm_n1987, gm_n211, in_14, in_10, gm_n345, gm_n212);
	nor (gm_n1988, gm_n566, gm_n882, in_11, gm_n708);
	nor (gm_n1989, gm_n1988, gm_n1987, gm_n1986);
	nor (gm_n1990, gm_n385, gm_n219, in_11, gm_n827, gm_n156);
	nor (gm_n1991, gm_n271, in_14, gm_n42, gm_n990);
	and (gm_n1992, gm_n1322, gm_n69, gm_n62);
	nor (gm_n1993, gm_n1992, gm_n1991, gm_n1990);
	nand (gm_n1994, gm_n1985, gm_n1955, gm_n1954, gm_n1993, gm_n1989);
	nand (gm_n1995, gm_n110, gm_n109, in_11, gm_n284, gm_n164);
	nand (gm_n1996, gm_n131, gm_n72, gm_n45, gm_n224, gm_n158);
	nand (gm_n1997, gm_n69, gm_n62, in_12, gm_n910, gm_n131);
	nand (gm_n1998, gm_n1997, gm_n1996, gm_n1995);
	nand (gm_n1999, gm_n81, gm_n109, gm_n43, gm_n266, gm_n168);
	nand (gm_n2000, in_14, gm_n62, in_12, gm_n601, gm_n44);
	nand (gm_n2001, gm_n1085, gm_n300, in_14);
	nand (gm_n2002, gm_n2001, gm_n2000, gm_n1999);
	nor (gm_n2003, gm_n1994, gm_n1953, gm_n1952, gm_n2002, gm_n1998);
	and (gm_n2004, gm_n320, gm_n72, gm_n43, gm_n168, gm_n116);
	and (gm_n2005, gm_n116, gm_n161, gm_n43, gm_n164, gm_n158);
	nor (gm_n2006, in_14, in_13, gm_n41, gm_n1481, gm_n230);
	nor (gm_n2007, gm_n2006, gm_n2005, gm_n2004);
	and (gm_n2008, in_14, gm_n62, in_12, gm_n432, gm_n349);
	nor (gm_n2009, gm_n69, in_13, in_12, gm_n1400, gm_n216);
	nor (gm_n2010, gm_n2009, gm_n2008, gm_n475);
	nand (gm_n2011, gm_n2003, gm_n1951, gm_n1950, gm_n2010, gm_n2007);
	nand (gm_n2012, gm_n224, gm_n43, gm_n58, gm_n1243, gm_n284);
	nand (gm_n2013, gm_n104, gm_n72, gm_n43, gm_n268, gm_n266);
	nand (gm_n2014, gm_n69, gm_n62, gm_n41, gm_n823, gm_n126);
	nand (gm_n2015, gm_n2014, gm_n2013, gm_n2012);
	nand (gm_n2016, in_14, in_13, in_12, gm_n1533, gm_n349);
	nand (gm_n2017, gm_n126, gm_n72, in_8, gm_n174, gm_n133);
	nand (gm_n2018, gm_n164, gm_n559, gm_n43, gm_n253);
	nand (gm_n2019, gm_n2018, gm_n2017, gm_n2016);
	nor (gm_n2020, gm_n2011, gm_n1949, gm_n1948, gm_n2019, gm_n2015);
	nand (gm_n2021, gm_n44, in_12, in_8, gm_n73, gm_n72);
	nor (gm_n2022, gm_n2021, gm_n69, in_13);
	or (gm_n2023, gm_n50, in_12, gm_n45, gm_n216, gm_n385);
	nor (gm_n2024, gm_n2023, gm_n69, in_13);
	and (gm_n2025, gm_n106, gm_n161, in_11, gm_n158, gm_n117);
	nor (gm_n2026, gm_n2025, gm_n2024, gm_n2022);
	and (gm_n2027, gm_n69, gm_n62, gm_n41, gm_n691, gm_n349);
	and (gm_n2028, gm_n69, in_13, in_12, gm_n1152, gm_n191);
	nor (gm_n2029, gm_n57, gm_n76, gm_n45, gm_n225, gm_n94);
	nor (gm_n2030, gm_n2029, gm_n2028, gm_n2027);
	nand (gm_n2031, gm_n2020, gm_n1947, gm_n1946, gm_n2030, gm_n2026);
	or (gm_n2032, gm_n69, gm_n62, gm_n41, gm_n595, gm_n342);
	nand (gm_n2033, gm_n69, in_13, in_12, gm_n131, gm_n505);
	nand (gm_n2034, gm_n2033, gm_n2032, gm_n1504);
	nor (gm_n2035, gm_n41, gm_n43, in_10);
	nand (gm_n2036, in_14, gm_n62, in_9, gm_n2035, gm_n757);
	nand (gm_n2037, gm_n69, gm_n62, gm_n41, gm_n251, gm_n126);
	nand (gm_n2038, gm_n109, gm_n370, in_11, gm_n284, gm_n104);
	nand (gm_n2039, gm_n2038, gm_n2037, gm_n2036);
	nor (gm_n2040, gm_n2031, gm_n1945, gm_n1944, gm_n2039, gm_n2034);
	and (gm_n2041, gm_n381, gm_n65, gm_n69, gm_n266, gm_n300);
	nor (gm_n2042, gm_n385, gm_n50, gm_n45, gm_n229, gm_n261);
	and (gm_n2043, gm_n161, gm_n93, gm_n45, gm_n255, gm_n224);
	nor (gm_n2044, gm_n2043, gm_n2042, gm_n2041);
	nor (gm_n2045, in_14, gm_n62, in_12, gm_n74, gm_n63);
	nor (gm_n2046, gm_n108, in_14, gm_n42, gm_n286, gm_n143);
	nor (gm_n2047, gm_n84, gm_n69, gm_n42, gm_n287, gm_n467);
	nor (gm_n2048, gm_n2047, gm_n2046, gm_n2045);
	nand (gm_n2049, gm_n2040, gm_n1942, gm_n1941, gm_n2048, gm_n2044);
	nand (gm_n2050, gm_n174, gm_n131, gm_n45, gm_n381, gm_n183);
	nor (gm_n2051, gm_n94, in_12, gm_n45, gm_n193, gm_n342);
	nand (gm_n2052, gm_n2051, gm_n69, gm_n62);
	nand (gm_n2053, gm_n73, gm_n44, gm_n45, gm_n104, gm_n88);
	nand (gm_n2054, gm_n2053, gm_n2052, gm_n2050);
	nand (gm_n2055, gm_n88, gm_n66, in_8, gm_n191, gm_n168);
	or (gm_n2056, gm_n271, gm_n69, in_10, gm_n419, gm_n307);
	nor (gm_n2057, gm_n342, gm_n41, gm_n45, gm_n193, gm_n208);
	nand (gm_n2058, gm_n2057, in_14, in_13);
	nand (gm_n2059, gm_n2058, gm_n2056, gm_n2055);
	nor (gm_n2060, gm_n2049, gm_n1940, gm_n1938, gm_n2059, gm_n2054);
	nor (gm_n2061, gm_n229, gm_n89, gm_n43, gm_n193, gm_n646);
	and (gm_n2062, gm_n320, gm_n109, gm_n43, gm_n174, gm_n116);
	nor (gm_n2063, gm_n2062, gm_n2061, gm_n1163);
	and (gm_n2064, gm_n245, in_14, gm_n42, gm_n917, gm_n211);
	nor (gm_n2065, gm_n69, gm_n62, in_12, gm_n1903, gm_n71);
	nor (gm_n2066, in_14, gm_n42, in_9, gm_n1274, gm_n84);
	nor (gm_n2067, gm_n2066, gm_n2065, gm_n2064);
	nand (gm_n2068, gm_n2060, gm_n1937, gm_n1936, gm_n2067, gm_n2063);
	nand (gm_n2069, gm_n126, gm_n161, in_8, gm_n268, gm_n164);
	nand (gm_n2070, gm_n69, in_10, gm_n70, gm_n746, gm_n83);
	or (gm_n2071, gm_n566, gm_n827, in_11, gm_n593);
	nand (gm_n2072, gm_n2071, gm_n2070, gm_n2069);
	nand (gm_n2073, gm_n69, gm_n62, gm_n41, gm_n601, gm_n53);
	or (gm_n2074, in_14, in_13, gm_n41, gm_n262, gm_n327);
	nand (gm_n2075, gm_n69, gm_n62, gm_n41, gm_n1761, gm_n349);
	nand (gm_n2076, gm_n2075, gm_n2074, gm_n2073);
	nor (out_14, gm_n2072, gm_n2068, gm_n1935, gm_n2076);
endmodule
