module top ( g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 , g98 , g99 , g100 , g101 , g102 , g103 , g104 , g105 , g106 , g107 , g108 , g109 , g110 , g111 , g112 , g113 , g114 , g115 , g116 , g117 , g118 , g119 , g120 , g121 , g122 , g123 , g124 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g136 , g137 , g138 , g139 , g140 , g141 , g142 , g143 , g144 , g145 , g146 , g147 , g148 , g149 , g150 , g151 , g152 , g153 , g154 , g155 , g156 , g157 , g158 , g159 , g160 , g161 , g162 , g163 , g164 , g165 , g166 , g167 , g168 , g169 , g170 , g171 , g172 , g173 , g174 , g175 , g176 , g177 , g178 , g179 , g180 , g181 , g182 , g183 , g184 , g185 , g186 , g187 , g188 , g189 , g190 , g191 , g192 , g193 , g194 , g195 , g196 , g197 , g198 , g199 , g200 , g201 , g202 , g203 , g204 , g205 , g206 , g207 , g208 , g209 , g210 , g211 , g212 , g213 , g214 , g215 , g216 , g217 , g218 , g219 , g220 , g221 , g222 , g223 , g224 , g225 , g226 , g227 , g228 , g229 , g230 , g231 , g232 , g233 , g234 , g235 , g236 , g237 , g238 , g239 , g240 , g241 , g242 , g243 , g244 , g245 , g246 , g247 , g248 , g249 , g250 , g251 , g252 , g253 , g254 , g255 , g256 , g257 , g258 , g259 , g260 , g261 , g262 , g263 , g264 , g265 , g266 , g267 , g268 , g269 , g270 , g271 , g272 , g273 , g274 , g275 , g276 , g277 , g278 , g279 , g280 , g281 , g282 , g283 , g284 , g285 , g286 , g287 , g288 , g289 , g290 , g291 , g292 , g293 , g294 , g295 , g296 , g297 , g298 , g299 , g300 , g301 , g302 , g303 , g304 , g305 , g306 , g307 , g308 , g309 , g310 , g311 , g312 , g313 , g314 , g315 , g316 , g317 , g318 , g319 , g320 , g321 , g322 , g323 , g324 , g325 , g326 , g327 , g328 , g329 , g330 , g331 , g332 , g333 , g334 , g335 , g336 , g337 , g338 , g339 , g340 , g341 , g342 , g343 , g344 , g345 , g346 , g347 , g348 , g349 , g350 , g351 , g352 , g353 , g354 , g355 , g356 , g357 , g358 , g359 , g360 , g361 , g362 , g363 , g364 , g365 , g366 , g367 , g368 , g369 , g370 , g371 , g372 , g373 , g374 , g375 , g376 , g377 , g378 , g379 , g380 , g381 , g382 , g383 , g384 , g385 , g386 , g387 , g388 , g389 , g390 , g391 , g392 , g393 , g394 , g395 , g396 , g397 , g398 , g399 , g400 , g401 , g402 , g403 , g404 , g405 , g406 , g407 , g408 , g409 , g410 , g411 , g412 , g413 , g414 , g415 , g416 , g417 , g418 , g419 , g420 , g421 , g422 , g423 , g424 , g425 , g426 , g427 , g428 , g429 , g430 , g431 , g432 , g433 , g434 , g435 , g436 , g437 , g438 , g439 , g440 , g441 , g442 , g443 , g444 , g445 , g446 , g447 , g448 , g449 , g450 , g451 , g452 , g453 , g454 , g455 , g456 , g457 , g458 , g459 , g460 , g461 , g462 , g463 , g464 , g465 , g466 , g467 , g468 , g469 , g470 , g471 , g472 , g473 , g474 , g475 , g476 , g477 , g478 , g479 , g480 , g481 , g482 , g483 , g484 , g485 , g486 , g487 , g488 , g489 , g490 , g491 , g492 , g493 , g494 , g495 , g496 , g497 , g498 , g499 , g500 , g501 , g502 , g503 , g504 , g505 , g506 , g507 , g508 , g509 , g510 , g511 , g512 , g513 , g514 , g515 , g516 , g517 , g518 , g519 , g520 , g521 , g522 , g523 , g524 , g525 , g526 , g527 , g528 , g529 , g530 , g531 , g532 , g533 , g534 , g535 , g536 , g537 , g538 , g539 , g540 , g541 , g542 , g543 , g544 , g545 , g546 , g547 , g548 , g549 , g550 , g551 , g552 , g553 , g554 , g555 , g556 , g557 , g558 , g559 , g560 , g561 , g562 , g563 , g564 , g565 , g566 , g567 , g568 , g569 , g570 , g571 , g572 , g573 , g574 , g575 , g576 , g577 , g578 , g579 , g580 , g581 , g582 , g583 , g584 , g585 , g586 , g587 , g588 , g589 , g590 , g591 , g592 , g593 , g594 , g595 , g596 , g597 , g598 , g599 , g600 , g601 , g602 , g603 , g604 , g605 , g606 , g607 , g608 , g609 , g610 , g611 , g612 , g613 , g614 , g615 , g616 , g617 , g618 , g619 , g620 , g621 , g622 , g623 , g624 , g625 , g626 , g627 , g628 , g629 , g630 );
input g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 , g98 , g99 , g100 , g101 , g102 , g103 , g104 , g105 , g106 , g107 , g108 , g109 , g110 , g111 , g112 , g113 , g114 , g115 , g116 , g117 , g118 , g119 , g120 , g121 , g122 , g123 , g124 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g136 , g137 , g138 , g139 , g140 , g141 , g142 , g143 , g144 , g145 , g146 , g147 , g148 , g149 , g150 , g151 , g152 , g153 , g154 , g155 , g156 , g157 , g158 , g159 , g160 , g161 , g162 , g163 , g164 , g165 , g166 , g167 , g168 , g169 , g170 , g171 , g172 , g173 , g174 , g175 , g176 , g177 , g178 , g179 , g180 , g181 , g182 , g183 , g184 , g185 , g186 , g187 , g188 , g189 , g190 , g191 , g192 , g193 , g194 , g195 , g196 , g197 , g198 , g199 , g200 , g201 , g202 , g203 , g204 , g205 , g206 , g207 , g208 , g209 , g210 , g211 , g212 , g213 , g214 , g215 , g216 , g217 , g218 , g219 , g220 , g221 , g222 , g223 , g224 , g225 , g226 , g227 , g228 , g229 , g230 , g231 , g232 , g233 , g234 , g235 , g236 , g237 , g238 , g239 , g240 , g241 , g242 , g243 , g244 , g245 , g246 , g247 , g248 , g249 , g250 , g251 , g252 , g253 , g254 , g255 , g256 , g257 , g258 , g259 , g260 , g261 , g262 , g263 , g264 , g265 , g266 , g267 , g268 , g269 , g270 , g271 , g272 , g273 , g274 , g275 , g276 , g277 , g278 , g279 , g280 , g281 , g282 , g283 , g284 , g285 , g286 , g287 , g288 , g289 , g290 , g291 , g292 , g293 , g294 , g295 , g296 , g297 , g298 , g299 , g300 , g301 , g302 , g303 , g304 , g305 , g306 , g307 , g308 , g309 , g310 , g311 , g312 , g313 , g314 , g315 , g316 , g317 , g318 , g319 , g320 , g321 , g322 , g323 , g324 , g325 , g326 , g327 , g328 , g329 , g330 , g331 , g332 , g333 , g334 , g335 , g336 , g337 , g338 , g339 , g340 , g341 , g342 , g343 , g344 , g345 , g346 , g347 , g348 , g349 , g350 , g351 , g352 , g353 , g354 , g355 , g356 , g357 , g358 , g359 , g360 , g361 , g362 , g363 , g364 , g365 , g366 , g367 , g368 , g369 , g370 , g371 , g372 , g373 , g374 , g375 , g376 , g377 , g378 , g379 , g380 , g381 , g382 , g383 , g384 , g385 , g386 , g387 , g388 , g389 , g390 , g391 , g392 , g393 , g394 , g395 , g396 , g397 , g398 , g399 , g400 , g401 , g402 , g403 , g404 , g405 , g406 , g407 , g408 , g409 , g410 , g411 , g412 , g413 , g414 , g415 , g416 ;
output g417 , g418 , g419 , g420 , g421 , g422 , g423 , g424 , g425 , g426 , g427 , g428 , g429 , g430 , g431 , g432 , g433 , g434 , g435 , g436 , g437 , g438 , g439 , g440 , g441 , g442 , g443 , g444 , g445 , g446 , g447 , g448 , g449 , g450 , g451 , g452 , g453 , g454 , g455 , g456 , g457 , g458 , g459 , g460 , g461 , g462 , g463 , g464 , g465 , g466 , g467 , g468 , g469 , g470 , g471 , g472 , g473 , g474 , g475 , g476 , g477 , g478 , g479 , g480 , g481 , g482 , g483 , g484 , g485 , g486 , g487 , g488 , g489 , g490 , g491 , g492 , g493 , g494 , g495 , g496 , g497 , g498 , g499 , g500 , g501 , g502 , g503 , g504 , g505 , g506 , g507 , g508 , g509 , g510 , g511 , g512 , g513 , g514 , g515 , g516 , g517 , g518 , g519 , g520 , g521 , g522 , g523 , g524 , g525 , g526 , g527 , g528 , g529 , g530 , g531 , g532 , g533 , g534 , g535 , g536 , g537 , g538 , g539 , g540 , g541 , g542 , g543 , g544 , g545 , g546 , g547 , g548 , g549 , g550 , g551 , g552 , g553 , g554 , g555 , g556 , g557 , g558 , g559 , g560 , g561 , g562 , g563 , g564 , g565 , g566 , g567 , g568 , g569 , g570 , g571 , g572 , g573 , g574 , g575 , g576 , g577 , g578 , g579 , g580 , g581 , g582 , g583 , g584 , g585 , g586 , g587 , g588 , g589 , g590 , g591 , g592 , g593 , g594 , g595 , g596 , g597 , g598 , g599 , g600 , g601 , g602 , g603 , g604 , g605 , g606 , g607 , g608 , g609 , g610 , g611 , g612 , g613 , g614 , g615 , g616 , g617 , g618 , g619 , g620 , g621 , g622 , g623 , g624 , g625 , g626 , g627 , g628 , g629 , g630 ;

wire n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , 
     n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , 
     n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , 
     n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , 
     n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , 
     n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , 
     n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , 
     n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , 
     n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , 
     n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , 
     n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , 
     n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , 
     n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , 
     n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , 
     n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , 
     n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , 
     n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , 
     n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , 
     n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , 
     n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , 
     n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , 
     n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , 
     n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , 
     n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , 
     n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , 
     n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , 
     n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , 
     n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , 
     n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , 
     n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , 
     n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , 
     n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , 
     n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , 
     n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , 
     n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , 
     n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , 
     n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , 
     n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , 
     n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , 
     n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , 
     n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , 
     n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , 
     n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , 
     n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , 
     n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , 
     n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , 
     n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , 
     n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , 
     n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , 
     n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , 
     n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , 
     n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , 
     n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , 
     n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , 
     n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , 
     n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , 
     n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , 
     n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , 
     n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , 
     n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , 
     n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , 
     n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , 
     n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , 
     n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , 
     n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , 
     n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , 
     n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , 
     n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , 
     n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , 
     n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , 
     n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , 
     n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , 
     n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , 
     n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , 
     n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , 
     n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , 
     n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , 
     n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , 
     n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , 
     n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , 
     n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , 
     n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , 
     n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , 
     n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , 
     n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , 
     n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , 
     n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , 
     n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , 
     n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , 
     n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , 
     n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , 
     n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , 
     n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , 
     n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , 
     n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , 
     n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , 
     n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , 
     n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , 
     n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , 
     n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , 
     n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , 
     n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , 
     n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , 
     n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , 
     n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , 
     n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , 
     n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , 
     n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , 
     n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , 
     n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , 
     n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , 
     n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , 
     n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , 
     n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , 
     n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , 
     n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , 
     n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , 
     n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , 
     n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , 
     n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , 
     n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , 
     n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , 
     n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , 
     n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , 
     n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , 
     n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , 
     n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , 
     n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , 
     n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , 
     n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , 
     n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , 
     n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , 
     n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , 
     n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , 
     n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , 
     n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , 
     n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , 
     n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , 
     n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , 
     n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , 
     n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , 
     n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , 
     n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , 
     n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , 
     n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , 
     n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , 
     n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , 
     n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , 
     n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , 
     n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , 
     n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , 
     n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , 
     n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , 
     n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , 
     n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , 
     n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , 
     n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , 
     n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , 
     n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , 
     n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , 
     n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , 
     n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , 
     n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , 
     n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , 
     n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , 
     n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , 
     n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , 
     n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , 
     n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , 
     n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , 
     n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , 
     n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , 
     n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , 
     n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , 
     n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , 
     n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , 
     n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , 
     n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , 
     n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , 
     n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , 
     n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , 
     n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , 
     n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , 
     n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , 
     n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , 
     n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , 
     n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , 
     n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , 
     n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , 
     n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , 
     n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , 
     n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , 
     n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , 
     n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , 
     n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , 
     n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , 
     n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , 
     n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , 
     n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , 
     n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , 
     n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , 
     n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , 
     n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , 
     n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , 
     n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , 
     n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , 
     n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , 
     n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , 
     n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , 
     n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , 
     n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , 
     n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , 
     n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , 
     n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , 
     n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , 
     n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , 
     n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , 
     n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , 
     n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , 
     n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , 
     n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , 
     n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , 
     n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , 
     n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , 
     n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , 
     n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , 
     n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , 
     n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , 
     n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , 
     n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , 
     n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , 
     n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , 
     n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , 
     n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , 
     n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , 
     n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , 
     n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , 
     n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , 
     n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , 
     n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , 
     n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , 
     n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , 
     n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , 
     n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , 
     n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , 
     n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , 
     n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , 
     n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , 
     n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , 
     n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , 
     n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , 
     n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , 
     n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , 
     n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , 
     n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , 
     n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , 
     n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , 
     n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , 
     n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , 
     n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , 
     n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , 
     n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , 
     n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , 
     n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , 
     n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , 
     n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , 
     n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , 
     n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , 
     n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , 
     n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , 
     n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , 
     n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , 
     n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , 
     n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , 
     n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , 
     n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , 
     n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , 
     n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , 
     n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , 
     n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , 
     n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , 
     n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , 
     n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , 
     n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , 
     n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , 
     n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , 
     n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , 
     n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , 
     n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , 
     n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , 
     n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , 
     n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , 
     n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , 
     n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , 
     n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , 
     n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , 
     n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , 
     n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , 
     n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , 
     n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , 
     n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , 
     n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , 
     n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , 
     n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , 
     n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , 
     n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , 
     n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , 
     n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , 
     n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , 
     n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , 
     n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , 
     n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , 
     n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , 
     n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , 
     n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , 
     n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , 
     n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , 
     n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , 
     n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , 
     n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , 
     n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , 
     n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , 
     n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , 
     n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , 
     n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , 
     n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , 
     n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , 
     n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , 
     n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , 
     n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , 
     n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , 
     n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , 
     n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , 
     n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , 
     n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , 
     n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , 
     n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , 
     n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , 
     n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , 
     n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , 
     n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , 
     n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , 
     n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , 
     n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , 
     n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , 
     n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , 
     n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , 
     n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , 
     n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , 
     n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , 
     n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , 
     n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , 
     n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , 
     n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , 
     n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , 
     n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , 
     n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , 
     n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , 
     n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , 
     n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , 
     n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , 
     n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , 
     n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , 
     n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , 
     n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , 
     n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , 
     n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , 
     n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , 
     n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , 
     n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , 
     n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , 
     n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , 
     n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , 
     n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , 
     n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , 
     n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , 
     n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , 
     n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , 
     n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , 
     n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , 
     n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , 
     n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , 
     n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , 
     n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , 
     n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , 
     n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , 
     n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , 
     n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , 
     n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , 
     n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , 
     n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , 
     n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , 
     n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , 
     n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , 
     n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , 
     n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , 
     n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , 
     n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , 
     n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , 
     n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , 
     n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , 
     n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , 
     n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , 
     n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , 
     n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , 
     n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , 
     n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , 
     n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , 
     n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , 
     n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , 
     n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , 
     n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , 
     n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , 
     n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , 
     n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , 
     n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , 
     n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , 
     n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , 
     n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , 
     n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , 
     n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , 
     n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , 
     n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , 
     n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , 
     n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , 
     n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , 
     n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , 
     n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , 
     n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , 
     n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , 
     n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , 
     n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , 
     n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , 
     n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , 
     n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , 
     n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , 
     n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , 
     n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , 
     n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , 
     n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , 
     n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , 
     n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , 
     n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , 
     n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , 
     n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , 
     n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , 
     n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , 
     n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , 
     n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , 
     n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , 
     n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , 
     n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , 
     n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , 
     n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , 
     n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , 
     n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , 
     n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , 
     n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , 
     n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , 
     n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , 
     n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , 
     n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , 
     n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , 
     n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , 
     n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , 
     n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , 
     n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , 
     n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , 
     n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , 
     n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , 
     n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , 
     n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , 
     n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , 
     n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , 
     n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , 
     n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , 
     n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , 
     n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , 
     n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , 
     n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , 
     n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , 
     n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , 
     n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , 
     n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , 
     n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , 
     n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , 
     n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , 
     n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , 
     n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , 
     n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , 
     n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , 
     n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , 
     n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , 
     n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , 
     n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , 
     n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , 
     n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , 
     n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , 
     n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , 
     n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , 
     n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , 
     n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , 
     n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , 
     n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , 
     n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , 
     n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , 
     n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , 
     n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , 
     n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , 
     n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , 
     n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , 
     n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , 
     n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , 
     n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , 
     n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , 
     n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , 
     n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , 
     n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , 
     n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , 
     n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , 
     n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , 
     n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , 
     n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , 
     n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , 
     n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , 
     n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , 
     n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , 
     n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , 
     n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , 
     n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , 
     n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , 
     n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , 
     n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , 
     n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , 
     n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , 
     n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , 
     n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , 
     n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , 
     n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , 
     n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , 
     n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , 
     n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , 
     n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , 
     n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , 
     n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , 
     n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , 
     n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , 
     n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , 
     n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , 
     n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , 
     n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , 
     n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , 
     n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , 
     n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , 
     n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , 
     n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , 
     n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , 
     n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , 
     n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , 
     n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , 
     n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , 
     n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , 
     n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , 
     n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , 
     n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , 
     n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , 
     n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , 
     n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , 
     n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , 
     n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , 
     n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , 
     n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , 
     n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , 
     n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , 
     n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , 
     n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , 
     n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , 
     n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , 
     n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , 
     n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , 
     n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , 
     n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , 
     n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , 
     n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , 
     n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , 
     n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , 
     n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , 
     n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , 
     n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , 
     n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , 
     n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , 
     n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , 
     n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , 
     n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , 
     n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , 
     n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , 
     n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , 
     n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , 
     n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , 
     n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , 
     n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , 
     n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , 
     n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , 
     n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , 
     n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , 
     n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , 
     n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , 
     n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , 
     n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , 
     n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , 
     n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , 
     n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , 
     n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , 
     n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , 
     n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , 
     n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , 
     n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , 
     n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , 
     n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , 
     n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , 
     n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , 
     n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , 
     n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , 
     n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , 
     n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , 
     n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , 
     n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , 
     n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , 
     n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , 
     n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , 
     n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , 
     n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , 
     n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , 
     n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , 
     n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , 
     n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , 
     n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , 
     n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , 
     n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , 
     n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , 
     n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , 
     n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , 
     n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , 
     n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , 
     n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , 
     n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , 
     n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , 
     n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , 
     n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , 
     n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , 
     n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , 
     n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , 
     n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , 
     n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , 
     n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , 
     n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , 
     n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , 
     n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , 
     n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , 
     n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , 
     n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , 
     n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , 
     n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , 
     n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , 
     n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , 
     n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , 
     n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , 
     n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , 
     n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , 
     n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , 
     n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , 
     n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , 
     n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , 
     n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , 
     n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , 
     n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , 
     n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , 
     n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , 
     n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , 
     n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , 
     n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , 
     n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , 
     n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , 
     n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , 
     n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , 
     n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , 
     n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , 
     n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , 
     n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , 
     n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , 
     n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , 
     n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , 
     n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , 
     n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , 
     n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , 
     n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , 
     n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , 
     n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , 
     n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , 
     n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , 
     n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , 
     n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , 
     n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , 
     n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , 
     n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , 
     n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , 
     n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , 
     n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , 
     n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , 
     n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , 
     n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , 
     n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , 
     n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , 
     n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , 
     n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , 
     n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , 
     n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , 
     n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , 
     n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , 
     n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , 
     n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , 
     n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , 
     n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , 
     n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , 
     n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , 
     n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , 
     n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , 
     n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , 
     n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , 
     n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , 
     n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , 
     n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , 
     n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , 
     n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , 
     n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , 
     n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , 
     n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , 
     n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , 
     n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , 
     n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , 
     n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , 
     n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , 
     n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , 
     n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , 
     n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , 
     n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , 
     n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , 
     n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , 
     n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , 
     n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , 
     n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , 
     n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , 
     n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , 
     n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , 
     n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , 
     n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , 
     n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , 
     n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , 
     n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , 
     n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , 
     n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , 
     n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , 
     n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , 
     n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , 
     n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , 
     n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , 
     n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , 
     n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , 
     n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , 
     n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , 
     n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , 
     n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , 
     n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , 
     n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , 
     n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , 
     n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , 
     n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , 
     n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , 
     n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , 
     n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , 
     n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , 
     n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , 
     n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , 
     n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , 
     n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , 
     n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , 
     n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , 
     n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , 
     n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , 
     n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , 
     n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , 
     n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , 
     n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , 
     n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , 
     n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , 
     n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , 
     n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , 
     n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , 
     n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , 
     n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , 
     n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , 
     n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , 
     n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , 
     n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , 
     n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , 
     n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , 
     n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , 
     n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , 
     n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , 
     n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , 
     n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , 
     n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , 
     n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , 
     n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , 
     n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , 
     n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , 
     n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , 
     n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , 
     n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , 
     n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , 
     n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , 
     n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , 
     n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , 
     n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , 
     n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , 
     n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , 
     n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , 
     n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , 
     n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , 
     n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , 
     n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , 
     n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , 
     n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , 
     n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , 
     n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , 
     n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , 
     n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , 
     n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , 
     n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , 
     n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , 
     n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , 
     n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , 
     n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , 
     n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , 
     n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , 
     n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , 
     n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , 
     n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , 
     n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , 
     n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , 
     n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , 
     n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , 
     n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , 
     n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , 
     n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , 
     n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , 
     n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , 
     n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , 
     n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , 
     n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , 
     n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , 
     n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , 
     n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , 
     n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , 
     n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , 
     n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , 
     n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , 
     n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , 
     n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , 
     n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , 
     n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , 
     n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , 
     n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , 
     n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , 
     n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , 
     n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , 
     n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , 
     n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , 
     n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , 
     n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , 
     n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , 
     n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , 
     n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , 
     n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , 
     n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , 
     n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , 
     n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , 
     n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , 
     n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , 
     n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , 
     n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , 
     n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , 
     n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , 
     n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , 
     n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , 
     n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , 
     n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , 
     n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , 
     n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , 
     n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , 
     n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , 
     n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , 
     n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , 
     n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , 
     n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , 
     n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , 
     n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , 
     n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , 
     n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , 
     n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , 
     n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , 
     n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , 
     n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , 
     n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , 
     n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , 
     n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , 
     n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , 
     n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , 
     n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , 
     n9190 , n9191 ;
buf ( n1 , g0 );
buf ( n2 , g1 );
buf ( n3 , g2 );
buf ( n4 , g3 );
buf ( n5 , g4 );
buf ( n6 , g5 );
buf ( n7 , g6 );
buf ( n8 , g7 );
buf ( n9 , g8 );
buf ( n10 , g9 );
buf ( n11 , g10 );
buf ( n12 , g11 );
buf ( n13 , g12 );
buf ( n14 , g13 );
buf ( n15 , g14 );
buf ( n16 , g15 );
buf ( n17 , g16 );
buf ( n18 , g17 );
buf ( n19 , g18 );
buf ( n20 , g19 );
buf ( n21 , g20 );
buf ( n22 , g21 );
buf ( n23 , g22 );
buf ( n24 , g23 );
buf ( n25 , g24 );
buf ( n26 , g25 );
buf ( n27 , g26 );
buf ( n28 , g27 );
buf ( n29 , g28 );
buf ( n30 , g29 );
buf ( n31 , g30 );
buf ( n32 , g31 );
buf ( n33 , g32 );
buf ( n34 , g33 );
buf ( n35 , g34 );
buf ( n36 , g35 );
buf ( n37 , g36 );
buf ( n38 , g37 );
buf ( n39 , g38 );
buf ( n40 , g39 );
buf ( n41 , g40 );
buf ( n42 , g41 );
buf ( n43 , g42 );
buf ( n44 , g43 );
buf ( n45 , g44 );
buf ( n46 , g45 );
buf ( n47 , g46 );
buf ( n48 , g47 );
buf ( n49 , g48 );
buf ( n50 , g49 );
buf ( n51 , g50 );
buf ( n52 , g51 );
buf ( n53 , g52 );
buf ( n54 , g53 );
buf ( n55 , g54 );
buf ( n56 , g55 );
buf ( n57 , g56 );
buf ( n58 , g57 );
buf ( n59 , g58 );
buf ( n60 , g59 );
buf ( n61 , g60 );
buf ( n62 , g61 );
buf ( n63 , g62 );
buf ( n64 , g63 );
buf ( n65 , g64 );
buf ( n66 , g65 );
buf ( n67 , g66 );
buf ( n68 , g67 );
buf ( n69 , g68 );
buf ( n70 , g69 );
buf ( n71 , g70 );
buf ( n72 , g71 );
buf ( n73 , g72 );
buf ( n74 , g73 );
buf ( n75 , g74 );
buf ( n76 , g75 );
buf ( n77 , g76 );
buf ( n78 , g77 );
buf ( n79 , g78 );
buf ( n80 , g79 );
buf ( n81 , g80 );
buf ( n82 , g81 );
buf ( n83 , g82 );
buf ( n84 , g83 );
buf ( n85 , g84 );
buf ( n86 , g85 );
buf ( n87 , g86 );
buf ( n88 , g87 );
buf ( n89 , g88 );
buf ( n90 , g89 );
buf ( n91 , g90 );
buf ( n92 , g91 );
buf ( n93 , g92 );
buf ( n94 , g93 );
buf ( n95 , g94 );
buf ( n96 , g95 );
buf ( n97 , g96 );
buf ( n98 , g97 );
buf ( n99 , g98 );
buf ( n100 , g99 );
buf ( n101 , g100 );
buf ( n102 , g101 );
buf ( n103 , g102 );
buf ( n104 , g103 );
buf ( n105 , g104 );
buf ( n106 , g105 );
buf ( n107 , g106 );
buf ( n108 , g107 );
buf ( n109 , g108 );
buf ( n110 , g109 );
buf ( n111 , g110 );
buf ( n112 , g111 );
buf ( n113 , g112 );
buf ( n114 , g113 );
buf ( n115 , g114 );
buf ( n116 , g115 );
buf ( n117 , g116 );
buf ( n118 , g117 );
buf ( n119 , g118 );
buf ( n120 , g119 );
buf ( n121 , g120 );
buf ( n122 , g121 );
buf ( n123 , g122 );
buf ( n124 , g123 );
buf ( n125 , g124 );
buf ( n126 , g125 );
buf ( n127 , g126 );
buf ( n128 , g127 );
buf ( n129 , g128 );
buf ( n130 , g129 );
buf ( n131 , g130 );
buf ( n132 , g131 );
buf ( n133 , g132 );
buf ( n134 , g133 );
buf ( n135 , g134 );
buf ( n136 , g135 );
buf ( n137 , g136 );
buf ( n138 , g137 );
buf ( n139 , g138 );
buf ( n140 , g139 );
buf ( n141 , g140 );
buf ( n142 , g141 );
buf ( n143 , g142 );
buf ( n144 , g143 );
buf ( n145 , g144 );
buf ( n146 , g145 );
buf ( n147 , g146 );
buf ( n148 , g147 );
buf ( n149 , g148 );
buf ( n150 , g149 );
buf ( n151 , g150 );
buf ( n152 , g151 );
buf ( n153 , g152 );
buf ( n154 , g153 );
buf ( n155 , g154 );
buf ( n156 , g155 );
buf ( n157 , g156 );
buf ( n158 , g157 );
buf ( n159 , g158 );
buf ( n160 , g159 );
buf ( n161 , g160 );
buf ( n162 , g161 );
buf ( n163 , g162 );
buf ( n164 , g163 );
buf ( n165 , g164 );
buf ( n166 , g165 );
buf ( n167 , g166 );
buf ( n168 , g167 );
buf ( n169 , g168 );
buf ( n170 , g169 );
buf ( n171 , g170 );
buf ( n172 , g171 );
buf ( n173 , g172 );
buf ( n174 , g173 );
buf ( n175 , g174 );
buf ( n176 , g175 );
buf ( n177 , g176 );
buf ( n178 , g177 );
buf ( n179 , g178 );
buf ( n180 , g179 );
buf ( n181 , g180 );
buf ( n182 , g181 );
buf ( n183 , g182 );
buf ( n184 , g183 );
buf ( n185 , g184 );
buf ( n186 , g185 );
buf ( n187 , g186 );
buf ( n188 , g187 );
buf ( n189 , g188 );
buf ( n190 , g189 );
buf ( n191 , g190 );
buf ( n192 , g191 );
buf ( n193 , g192 );
buf ( n194 , g193 );
buf ( n195 , g194 );
buf ( n196 , g195 );
buf ( n197 , g196 );
buf ( n198 , g197 );
buf ( n199 , g198 );
buf ( n200 , g199 );
buf ( n201 , g200 );
buf ( n202 , g201 );
buf ( n203 , g202 );
buf ( n204 , g203 );
buf ( n205 , g204 );
buf ( n206 , g205 );
buf ( n207 , g206 );
buf ( n208 , g207 );
buf ( n209 , g208 );
buf ( n210 , g209 );
buf ( n211 , g210 );
buf ( n212 , g211 );
buf ( n213 , g212 );
buf ( n214 , g213 );
buf ( n215 , g214 );
buf ( n216 , g215 );
buf ( n217 , g216 );
buf ( n218 , g217 );
buf ( n219 , g218 );
buf ( n220 , g219 );
buf ( n221 , g220 );
buf ( n222 , g221 );
buf ( n223 , g222 );
buf ( n224 , g223 );
buf ( n225 , g224 );
buf ( n226 , g225 );
buf ( n227 , g226 );
buf ( n228 , g227 );
buf ( n229 , g228 );
buf ( n230 , g229 );
buf ( n231 , g230 );
buf ( n232 , g231 );
buf ( n233 , g232 );
buf ( n234 , g233 );
buf ( n235 , g234 );
buf ( n236 , g235 );
buf ( n237 , g236 );
buf ( n238 , g237 );
buf ( n239 , g238 );
buf ( n240 , g239 );
buf ( n241 , g240 );
buf ( n242 , g241 );
buf ( n243 , g242 );
buf ( n244 , g243 );
buf ( n245 , g244 );
buf ( n246 , g245 );
buf ( n247 , g246 );
buf ( n248 , g247 );
buf ( n249 , g248 );
buf ( n250 , g249 );
buf ( n251 , g250 );
buf ( n252 , g251 );
buf ( n253 , g252 );
buf ( n254 , g253 );
buf ( n255 , g254 );
buf ( n256 , g255 );
buf ( n257 , g256 );
buf ( n258 , g257 );
buf ( n259 , g258 );
buf ( n260 , g259 );
buf ( n261 , g260 );
buf ( n262 , g261 );
buf ( n263 , g262 );
buf ( n264 , g263 );
buf ( n265 , g264 );
buf ( n266 , g265 );
buf ( n267 , g266 );
buf ( n268 , g267 );
buf ( n269 , g268 );
buf ( n270 , g269 );
buf ( n271 , g270 );
buf ( n272 , g271 );
buf ( n273 , g272 );
buf ( n274 , g273 );
buf ( n275 , g274 );
buf ( n276 , g275 );
buf ( n277 , g276 );
buf ( n278 , g277 );
buf ( n279 , g278 );
buf ( n280 , g279 );
buf ( n281 , g280 );
buf ( n282 , g281 );
buf ( n283 , g282 );
buf ( n284 , g283 );
buf ( n285 , g284 );
buf ( n286 , g285 );
buf ( n287 , g286 );
buf ( n288 , g287 );
buf ( n289 , g288 );
buf ( n290 , g289 );
buf ( n291 , g290 );
buf ( n292 , g291 );
buf ( n293 , g292 );
buf ( n294 , g293 );
buf ( n295 , g294 );
buf ( n296 , g295 );
buf ( n297 , g296 );
buf ( n298 , g297 );
buf ( n299 , g298 );
buf ( n300 , g299 );
buf ( n301 , g300 );
buf ( n302 , g301 );
buf ( n303 , g302 );
buf ( n304 , g303 );
buf ( n305 , g304 );
buf ( n306 , g305 );
buf ( n307 , g306 );
buf ( n308 , g307 );
buf ( n309 , g308 );
buf ( n310 , g309 );
buf ( n311 , g310 );
buf ( n312 , g311 );
buf ( n313 , g312 );
buf ( n314 , g313 );
buf ( n315 , g314 );
buf ( n316 , g315 );
buf ( n317 , g316 );
buf ( n318 , g317 );
buf ( n319 , g318 );
buf ( n320 , g319 );
buf ( n321 , g320 );
buf ( n322 , g321 );
buf ( n323 , g322 );
buf ( n324 , g323 );
buf ( n325 , g324 );
buf ( n326 , g325 );
buf ( n327 , g326 );
buf ( n328 , g327 );
buf ( n329 , g328 );
buf ( n330 , g329 );
buf ( n331 , g330 );
buf ( n332 , g331 );
buf ( n333 , g332 );
buf ( n334 , g333 );
buf ( n335 , g334 );
buf ( n336 , g335 );
buf ( n337 , g336 );
buf ( n338 , g337 );
buf ( n339 , g338 );
buf ( n340 , g339 );
buf ( n341 , g340 );
buf ( n342 , g341 );
buf ( n343 , g342 );
buf ( n344 , g343 );
buf ( n345 , g344 );
buf ( n346 , g345 );
buf ( n347 , g346 );
buf ( n348 , g347 );
buf ( n349 , g348 );
buf ( n350 , g349 );
buf ( n351 , g350 );
buf ( n352 , g351 );
buf ( n353 , g352 );
buf ( n354 , g353 );
buf ( n355 , g354 );
buf ( n356 , g355 );
buf ( n357 , g356 );
buf ( n358 , g357 );
buf ( n359 , g358 );
buf ( n360 , g359 );
buf ( n361 , g360 );
buf ( n362 , g361 );
buf ( n363 , g362 );
buf ( n364 , g363 );
buf ( n365 , g364 );
buf ( n366 , g365 );
buf ( n367 , g366 );
buf ( n368 , g367 );
buf ( n369 , g368 );
buf ( n370 , g369 );
buf ( n371 , g370 );
buf ( n372 , g371 );
buf ( n373 , g372 );
buf ( n374 , g373 );
buf ( n375 , g374 );
buf ( n376 , g375 );
buf ( n377 , g376 );
buf ( n378 , g377 );
buf ( n379 , g378 );
buf ( n380 , g379 );
buf ( n381 , g380 );
buf ( n382 , g381 );
buf ( n383 , g382 );
buf ( n384 , g383 );
buf ( n385 , g384 );
buf ( n386 , g385 );
buf ( n387 , g386 );
buf ( n388 , g387 );
buf ( n389 , g388 );
buf ( n390 , g389 );
buf ( n391 , g390 );
buf ( n392 , g391 );
buf ( n393 , g392 );
buf ( n394 , g393 );
buf ( n395 , g394 );
buf ( n396 , g395 );
buf ( n397 , g396 );
buf ( n398 , g397 );
buf ( n399 , g398 );
buf ( n400 , g399 );
buf ( n401 , g400 );
buf ( n402 , g401 );
buf ( n403 , g402 );
buf ( n404 , g403 );
buf ( n405 , g404 );
buf ( n406 , g405 );
buf ( n407 , g406 );
buf ( n408 , g407 );
buf ( n409 , g408 );
buf ( n410 , g409 );
buf ( n411 , g410 );
buf ( n412 , g411 );
buf ( n413 , g412 );
buf ( n414 , g413 );
buf ( n415 , g414 );
buf ( n416 , g415 );
buf ( n417 , g416 );
buf ( g417 , n418 );
buf ( g418 , n419 );
buf ( g419 , n420 );
buf ( g420 , n421 );
buf ( g421 , n422 );
buf ( g422 , n423 );
buf ( g423 , n424 );
buf ( g424 , n425 );
buf ( g425 , n426 );
buf ( g426 , n427 );
buf ( g427 , n428 );
buf ( g428 , n429 );
buf ( g429 , n430 );
buf ( g430 , n431 );
buf ( g431 , n432 );
buf ( g432 , n433 );
buf ( g433 , n434 );
buf ( g434 , n435 );
buf ( g435 , n436 );
buf ( g436 , n437 );
buf ( g437 , n438 );
buf ( g438 , n439 );
buf ( g439 , n440 );
buf ( g440 , n441 );
buf ( g441 , n442 );
buf ( g442 , n443 );
buf ( g443 , n444 );
buf ( g444 , n445 );
buf ( g445 , n446 );
buf ( g446 , n447 );
buf ( g447 , n448 );
buf ( g448 , n449 );
buf ( g449 , n450 );
buf ( g450 , n451 );
buf ( g451 , n452 );
buf ( g452 , n453 );
buf ( g453 , n454 );
buf ( g454 , n455 );
buf ( g455 , n456 );
buf ( g456 , n457 );
buf ( g457 , n458 );
buf ( g458 , n459 );
buf ( g459 , n460 );
buf ( g460 , n461 );
buf ( g461 , n462 );
buf ( g462 , n463 );
buf ( g463 , n464 );
buf ( g464 , n465 );
buf ( g465 , n466 );
buf ( g466 , n467 );
buf ( g467 , n468 );
buf ( g468 , n469 );
buf ( g469 , n470 );
buf ( g470 , n471 );
buf ( g471 , n472 );
buf ( g472 , n473 );
buf ( g473 , n474 );
buf ( g474 , n475 );
buf ( g475 , n476 );
buf ( g476 , n477 );
buf ( g477 , n478 );
buf ( g478 , n479 );
buf ( g479 , n480 );
buf ( g480 , n481 );
buf ( g481 , n482 );
buf ( g482 , n483 );
buf ( g483 , n484 );
buf ( g484 , n485 );
buf ( g485 , n486 );
buf ( g486 , n487 );
buf ( g487 , n488 );
buf ( g488 , n489 );
buf ( g489 , n490 );
buf ( g490 , n491 );
buf ( g491 , n492 );
buf ( g492 , n493 );
buf ( g493 , n494 );
buf ( g494 , n495 );
buf ( g495 , n496 );
buf ( g496 , n497 );
buf ( g497 , n498 );
buf ( g498 , n499 );
buf ( g499 , n500 );
buf ( g500 , n501 );
buf ( g501 , n502 );
buf ( g502 , n503 );
buf ( g503 , n504 );
buf ( g504 , n505 );
buf ( g505 , n506 );
buf ( g506 , n507 );
buf ( g507 , n508 );
buf ( g508 , n509 );
buf ( g509 , n510 );
buf ( g510 , n511 );
buf ( g511 , n512 );
buf ( g512 , n513 );
buf ( g513 , n514 );
buf ( g514 , n515 );
buf ( g515 , n516 );
buf ( g516 , n517 );
buf ( g517 , n518 );
buf ( g518 , n519 );
buf ( g519 , n520 );
buf ( g520 , n521 );
buf ( g521 , n522 );
buf ( g522 , n523 );
buf ( g523 , n524 );
buf ( g524 , n525 );
buf ( g525 , n526 );
buf ( g526 , n527 );
buf ( g527 , n528 );
buf ( g528 , n529 );
buf ( g529 , n530 );
buf ( g530 , n531 );
buf ( g531 , n532 );
buf ( g532 , n533 );
buf ( g533 , n534 );
buf ( g534 , n535 );
buf ( g535 , n536 );
buf ( g536 , n537 );
buf ( g537 , n538 );
buf ( g538 , n539 );
buf ( g539 , n540 );
buf ( g540 , n541 );
buf ( g541 , n542 );
buf ( g542 , n543 );
buf ( g543 , n544 );
buf ( g544 , n545 );
buf ( g545 , n546 );
buf ( g546 , n547 );
buf ( g547 , n548 );
buf ( g548 , n549 );
buf ( g549 , n550 );
buf ( g550 , n551 );
buf ( g551 , n552 );
buf ( g552 , n553 );
buf ( g553 , n554 );
buf ( g554 , n555 );
buf ( g555 , n556 );
buf ( g556 , n557 );
buf ( g557 , n558 );
buf ( g558 , n559 );
buf ( g559 , n560 );
buf ( g560 , n561 );
buf ( g561 , n562 );
buf ( g562 , n563 );
buf ( g563 , n564 );
buf ( g564 , n565 );
buf ( g565 , n566 );
buf ( g566 , n567 );
buf ( g567 , n568 );
buf ( g568 , n569 );
buf ( g569 , n570 );
buf ( g570 , n571 );
buf ( g571 , n572 );
buf ( g572 , n573 );
buf ( g573 , n574 );
buf ( g574 , n575 );
buf ( g575 , n576 );
buf ( g576 , n577 );
buf ( g577 , n578 );
buf ( g578 , n579 );
buf ( g579 , n580 );
buf ( g580 , n581 );
buf ( g581 , n582 );
buf ( g582 , n583 );
buf ( g583 , n584 );
buf ( g584 , n585 );
buf ( g585 , n586 );
buf ( g586 , n587 );
buf ( g587 , n588 );
buf ( g588 , n589 );
buf ( g589 , n590 );
buf ( g590 , n591 );
buf ( g591 , n592 );
buf ( g592 , n593 );
buf ( g593 , n594 );
buf ( g594 , n595 );
buf ( g595 , n596 );
buf ( g596 , n597 );
buf ( g597 , n598 );
buf ( g598 , n599 );
buf ( g599 , n600 );
buf ( g600 , n601 );
buf ( g601 , n602 );
buf ( g602 , n603 );
buf ( g603 , n604 );
buf ( g604 , n605 );
buf ( g605 , n606 );
buf ( g606 , n607 );
buf ( g607 , n608 );
buf ( g608 , n609 );
buf ( g609 , n610 );
buf ( g610 , n611 );
buf ( g611 , n612 );
buf ( g612 , n613 );
buf ( g613 , n614 );
buf ( g614 , n615 );
buf ( g615 , n616 );
buf ( g616 , n617 );
buf ( g617 , n618 );
buf ( g618 , n619 );
buf ( g619 , n620 );
buf ( g620 , n621 );
buf ( g621 , n622 );
buf ( g622 , n623 );
buf ( g623 , n624 );
buf ( g624 , n625 );
buf ( g625 , n626 );
buf ( g626 , n627 );
buf ( g627 , n628 );
buf ( g628 , n629 );
buf ( g629 , n630 );
buf ( g630 , n631 );
buf ( n418 , 1'b0 );
buf ( n419 , n9144 );
buf ( n420 , 1'b0 );
buf ( n421 , n9187 );
buf ( n422 , 1'b0 );
buf ( n423 , n9134 );
buf ( n424 , 1'b0 );
buf ( n425 , 1'b0 );
buf ( n426 , n9135 );
buf ( n427 , 1'b0 );
buf ( n428 , n9164 );
buf ( n429 , n9138 );
buf ( n430 , 1'b0 );
buf ( n431 , n9159 );
buf ( n432 , n8861 );
buf ( n433 , n9098 );
buf ( n434 , n9165 );
buf ( n435 , n9161 );
buf ( n436 , n2986 );
buf ( n437 , n8850 );
buf ( n438 , n9095 );
buf ( n439 , n9156 );
buf ( n440 , n9158 );
buf ( n441 , n2986 );
buf ( n442 , n9094 );
buf ( n443 , n9140 );
buf ( n444 , n9147 );
buf ( n445 , n9149 );
buf ( n446 , n9182 );
buf ( n447 , n9155 );
buf ( n448 , n9116 );
buf ( n449 , n9121 );
buf ( n450 , n9143 );
buf ( n451 , n9160 );
buf ( n452 , n9163 );
buf ( n453 , 1'b0 );
buf ( n454 , n8874 );
buf ( n455 , n9174 );
buf ( n456 , n9054 );
buf ( n457 , n9146 );
buf ( n458 , n9122 );
buf ( n459 , n9162 );
buf ( n460 , n9031 );
buf ( n461 , n9184 );
buf ( n462 , n9168 );
buf ( n463 , n9167 );
buf ( n464 , n9142 );
buf ( n465 , n9124 );
buf ( n466 , n9120 );
buf ( n467 , n9125 );
buf ( n468 , n4144 );
buf ( n469 , n9117 );
buf ( n470 , n8020 );
buf ( n471 , n9123 );
buf ( n472 , n9145 );
buf ( n473 , n9152 );
buf ( n474 , n9185 );
buf ( n475 , 1'b0 );
buf ( n476 , n9097 );
buf ( n477 , n9148 );
buf ( n478 , n9151 );
buf ( n479 , n9157 );
buf ( n480 , 1'b0 );
buf ( n481 , n9189 );
buf ( n482 , n9136 );
buf ( n483 , n9153 );
buf ( n484 , n9183 );
buf ( n485 , 1'b0 );
buf ( n486 , n9133 );
buf ( n487 , n9154 );
buf ( n488 , n9166 );
buf ( n489 , 1'b0 );
buf ( n490 , n9141 );
buf ( n491 , n9181 );
buf ( n492 , n9118 );
buf ( n493 , n9173 );
buf ( n494 , n9139 );
buf ( n495 , 1'b0 );
buf ( n496 , n9175 );
buf ( n497 , n9137 );
buf ( n498 , 1'b0 );
buf ( n499 , n9186 );
buf ( n500 , 1'b0 );
buf ( n501 , 1'b0 );
buf ( n502 , n1 );
buf ( n503 , n8674 );
buf ( n504 , 1'b0 );
buf ( n505 , 1'b0 );
buf ( n506 , n1 );
buf ( n507 , n6223 );
buf ( n508 , 1'b0 );
buf ( n509 , 1'b0 );
buf ( n510 , n1 );
buf ( n511 , n8798 );
buf ( n512 , 1'b0 );
buf ( n513 , 1'b0 );
buf ( n514 , n1 );
buf ( n515 , n3017 );
buf ( n516 , 1'b0 );
buf ( n517 , 1'b0 );
buf ( n518 , n1 );
buf ( n519 , n9024 );
buf ( n520 , 1'b0 );
buf ( n521 , 1'b0 );
buf ( n522 , n1 );
buf ( n523 , n8894 );
buf ( n524 , 1'b0 );
buf ( n525 , 1'b0 );
buf ( n526 , n1 );
buf ( n527 , n9091 );
buf ( n528 , 1'b0 );
buf ( n529 , 1'b0 );
buf ( n530 , n1 );
buf ( n531 , n4912 );
buf ( n532 , 1'b0 );
buf ( n533 , 1'b0 );
buf ( n534 , n1 );
buf ( n535 , n8990 );
buf ( n536 , 1'b0 );
buf ( n537 , 1'b0 );
buf ( n538 , n1 );
buf ( n539 , n7644 );
buf ( n540 , 1'b0 );
buf ( n541 , 1'b0 );
buf ( n542 , n1 );
buf ( n543 , n9084 );
buf ( n544 , 1'b0 );
buf ( n545 , 1'b0 );
buf ( n546 , n1 );
buf ( n547 , n8542 );
buf ( n548 , 1'b0 );
buf ( n549 , 1'b0 );
buf ( n550 , n1 );
buf ( n551 , n2986 );
buf ( n552 , 1'b0 );
buf ( n553 , 1'b0 );
buf ( n554 , n1 );
buf ( n555 , n9101 );
buf ( n556 , 1'b0 );
buf ( n557 , 1'b0 );
buf ( n558 , n1 );
buf ( n559 , n8967 );
buf ( n560 , 1'b0 );
buf ( n561 , 1'b0 );
buf ( n562 , n1 );
buf ( n563 , n8776 );
buf ( n564 , 1'b0 );
buf ( n565 , 1'b0 );
buf ( n566 , n1 );
buf ( n567 , n9052 );
buf ( n568 , 1'b0 );
buf ( n569 , 1'b0 );
buf ( n570 , n1 );
buf ( n571 , n8917 );
buf ( n572 , 1'b0 );
buf ( n573 , 1'b0 );
buf ( n574 , n1 );
buf ( n575 , n8980 );
buf ( n576 , 1'b0 );
buf ( n577 , 1'b0 );
buf ( n578 , n1 );
buf ( n579 , n9046 );
buf ( n580 , 1'b0 );
buf ( n581 , 1'b0 );
buf ( n582 , n1 );
buf ( n583 , n9127 );
buf ( n584 , 1'b0 );
buf ( n585 , 1'b0 );
buf ( n586 , n1 );
buf ( n587 , n9003 );
buf ( n588 , 1'b0 );
buf ( n589 , 1'b0 );
buf ( n590 , n1 );
buf ( n591 , n8947 );
buf ( n592 , 1'b0 );
buf ( n593 , 1'b0 );
buf ( n594 , n1 );
buf ( n595 , n9115 );
buf ( n596 , 1'b0 );
buf ( n597 , 1'b0 );
buf ( n598 , n1 );
buf ( n599 , n9172 );
buf ( n600 , 1'b0 );
buf ( n601 , 1'b0 );
buf ( n602 , n1 );
buf ( n603 , n9180 );
buf ( n604 , 1'b0 );
buf ( n605 , 1'b0 );
buf ( n606 , n1 );
buf ( n607 , n9108 );
buf ( n608 , 1'b0 );
buf ( n609 , 1'b0 );
buf ( n610 , n1 );
buf ( n611 , n9132 );
buf ( n612 , 1'b0 );
buf ( n613 , 1'b0 );
buf ( n614 , n1 );
buf ( n615 , n8885 );
buf ( n616 , 1'b0 );
buf ( n617 , 1'b0 );
buf ( n618 , n1 );
buf ( n619 , n8835 );
buf ( n620 , 1'b0 );
buf ( n621 , 1'b0 );
buf ( n622 , n1 );
buf ( n623 , n9076 );
buf ( n624 , 1'b0 );
buf ( n625 , 1'b0 );
buf ( n626 , n1 );
buf ( n627 , n9020 );
buf ( n628 , 1'b0 );
buf ( n629 , 1'b0 );
buf ( n630 , n1 );
buf ( n631 , n9191 );
not ( n714 , n391 );
nor ( n715 , n389 , n395 );
and ( n716 , n393 , n715 );
nand ( n717 , n265 , n281 );
not ( n718 , n717 );
nor ( n719 , n24 , n64 );
nand ( n720 , n718 , n719 );
nand ( n721 , n386 , n394 );
not ( n722 , n721 );
not ( n723 , n722 );
not ( n724 , n723 );
not ( n725 , n416 );
nand ( n726 , n725 , n415 );
buf ( n727 , n726 );
not ( n728 , n727 );
not ( n729 , n728 );
not ( n730 , n404 );
nor ( n731 , n730 , n407 );
not ( n732 , n731 );
and ( n733 , n729 , n732 );
nor ( n734 , n410 , n412 );
buf ( n735 , n734 );
not ( n736 , n735 );
nor ( n737 , n733 , n736 );
not ( n738 , n737 );
and ( n739 , n724 , n738 );
not ( n740 , n402 );
nand ( n741 , n417 , n740 );
not ( n742 , n741 );
nand ( n743 , n730 , n742 );
not ( n744 , n734 );
not ( n745 , n744 );
not ( n746 , n407 );
nand ( n747 , n745 , n746 );
not ( n748 , n747 );
nand ( n749 , n743 , n748 );
not ( n750 , n415 );
and ( n751 , n414 , n750 );
not ( n752 , n751 );
not ( n753 , n416 );
nor ( n754 , n410 , n412 );
and ( n755 , n753 , n754 );
not ( n756 , n755 );
not ( n757 , n409 );
nor ( n758 , n757 , n414 );
nor ( n759 , n415 , n416 );
nand ( n760 , n758 , n759 );
not ( n761 , n760 );
nor ( n762 , n756 , n761 );
nand ( n763 , n752 , n762 );
buf ( n764 , n763 );
and ( n765 , n749 , n764 );
not ( n766 , n390 );
nor ( n767 , n388 , n392 );
and ( n768 , n766 , n767 );
not ( n769 , n768 );
not ( n770 , n769 );
not ( n771 , n770 );
nor ( n772 , n765 , n771 );
not ( n773 , n769 );
not ( n774 , n402 );
not ( n775 , n404 );
nor ( n776 , n775 , n407 );
nor ( n777 , n774 , n776 );
not ( n778 , n777 );
nand ( n779 , n402 , n404 );
not ( n780 , n779 );
not ( n781 , n735 );
nand ( n782 , n746 , n781 );
not ( n783 , n782 );
nand ( n784 , n780 , n783 );
nand ( n785 , n773 , n778 , n784 );
nand ( n786 , n764 , n785 );
nand ( n787 , n772 , n786 );
nor ( n788 , n739 , n787 );
not ( n789 , n788 );
not ( n790 , n388 );
not ( n791 , n392 );
and ( n792 , n394 , n791 );
not ( n793 , n386 );
nor ( n794 , n793 , n390 );
and ( n795 , n794 , n737 );
nand ( n796 , n792 , n795 );
and ( n797 , n790 , n796 );
nand ( n798 , n789 , n797 );
and ( n799 , n311 , n798 );
not ( n800 , n311 );
not ( n801 , n739 );
not ( n802 , n801 );
nor ( n803 , n409 , n414 );
nand ( n804 , n750 , n803 );
nor ( n805 , n756 , n751 );
nand ( n806 , n804 , n805 );
nand ( n807 , n806 , n785 );
not ( n808 , n807 );
not ( n809 , n746 );
nor ( n810 , n402 , n417 );
nand ( n811 , n730 , n810 );
not ( n812 , n811 );
or ( n813 , n809 , n812 );
nand ( n814 , n813 , n806 );
not ( n815 , n748 );
not ( n816 , n815 );
not ( n817 , n816 );
not ( n818 , n804 );
not ( n819 , n755 );
not ( n820 , n819 );
not ( n821 , n820 );
nor ( n822 , n818 , n821 );
not ( n823 , n822 );
and ( n824 , n817 , n823 );
buf ( n825 , n768 );
not ( n826 , n825 );
nor ( n827 , n824 , n826 );
nand ( n828 , n814 , n827 );
nor ( n829 , n808 , n828 );
not ( n830 , n829 );
or ( n831 , n802 , n830 );
nand ( n832 , n831 , n797 );
and ( n833 , n800 , n832 );
nor ( n834 , n799 , n833 );
nor ( n835 , n720 , n834 );
not ( n836 , n835 );
not ( n837 , n402 );
or ( n838 , n837 , n771 );
not ( n839 , n838 );
not ( n840 , n819 );
nand ( n841 , n840 , n752 );
nand ( n842 , n815 , n841 );
and ( n843 , n842 , n770 );
not ( n844 , n843 );
not ( n845 , n410 );
nand ( n846 , n726 , n845 );
not ( n847 , n846 );
not ( n848 , n416 );
nand ( n849 , n847 , n848 );
not ( n850 , n849 );
nor ( n851 , n409 , n414 );
not ( n852 , n851 );
nand ( n853 , n850 , n852 );
not ( n854 , n412 );
nand ( n855 , n726 , n854 );
not ( n856 , n855 );
nor ( n857 , n856 , n410 );
not ( n858 , n857 );
and ( n859 , n853 , n858 );
nand ( n860 , n407 , n413 );
not ( n861 , n416 );
not ( n862 , n412 );
not ( n863 , n862 );
or ( n864 , n861 , n863 );
not ( n865 , n410 );
nand ( n866 , n864 , n865 );
nand ( n867 , n407 , n866 );
nand ( n868 , n860 , n867 );
nand ( n869 , n859 , n868 );
not ( n870 , n736 );
buf ( n871 , n870 );
nand ( n872 , n869 , n871 );
not ( n873 , n872 );
not ( n874 , n873 );
or ( n875 , n844 , n874 );
nor ( n876 , n392 , n402 );
not ( n877 , n399 );
nor ( n878 , n388 , n390 );
not ( n879 , n878 );
nor ( n880 , n877 , n879 );
nand ( n881 , n876 , n880 );
nand ( n882 , n875 , n881 );
nor ( n883 , n839 , n882 );
not ( n884 , n883 );
not ( n885 , n842 );
not ( n886 , n872 );
not ( n887 , n886 );
or ( n888 , n885 , n887 );
nand ( n889 , n413 , n777 );
not ( n890 , n889 );
and ( n891 , n890 , n806 );
not ( n892 , n413 );
and ( n893 , n892 , n777 );
not ( n894 , n893 );
not ( n895 , n841 );
or ( n896 , n894 , n895 );
nand ( n897 , n896 , n784 );
nor ( n898 , n891 , n897 );
nand ( n899 , n888 , n898 );
not ( n900 , n899 );
and ( n901 , n900 , n404 );
not ( n902 , n743 );
not ( n903 , n902 );
not ( n904 , n783 );
not ( n905 , n904 );
not ( n906 , n905 );
or ( n907 , n903 , n906 );
not ( n908 , n402 );
nor ( n909 , n908 , n404 );
not ( n910 , n909 );
not ( n911 , n810 );
nand ( n912 , n911 , n730 );
not ( n913 , n912 );
nand ( n914 , n913 , n748 );
nand ( n915 , n910 , n914 );
nor ( n916 , n915 , n404 );
not ( n917 , n916 );
or ( n918 , n892 , n917 );
nand ( n919 , n907 , n918 );
nor ( n920 , n901 , n919 );
nand ( n921 , n851 , n759 );
or ( n922 , n920 , n921 );
not ( n923 , n917 );
not ( n924 , n899 );
or ( n925 , n923 , n924 );
buf ( n926 , n841 );
nand ( n927 , n925 , n926 );
nand ( n928 , n922 , n927 );
not ( n929 , n915 );
nand ( n930 , n399 , n929 );
not ( n931 , n930 );
nand ( n932 , n928 , n931 );
nand ( n933 , n884 , n932 , n898 );
not ( n934 , n933 );
not ( n935 , n739 );
not ( n936 , n935 );
not ( n937 , n936 );
not ( n938 , n937 );
not ( n939 , n938 );
buf ( n940 , n939 );
nand ( n941 , n934 , n940 );
not ( n942 , n797 );
not ( n943 , n942 );
buf ( n944 , n943 );
nand ( n945 , n941 , n944 );
not ( n946 , n24 );
nand ( n947 , n946 , n64 );
not ( n948 , n947 );
not ( n949 , n311 );
nand ( n950 , n949 , n718 );
not ( n951 , n950 );
nand ( n952 , n948 , n951 );
not ( n953 , n952 );
nand ( n954 , n945 , n953 );
not ( n955 , n843 );
not ( n956 , n414 );
nor ( n957 , n415 , n416 );
nand ( n958 , n957 , n754 );
nor ( n959 , n803 , n958 );
nand ( n960 , n956 , n959 );
not ( n961 , n866 );
nand ( n962 , n960 , n961 );
nand ( n963 , n868 , n962 );
nand ( n964 , n871 , n963 );
or ( n965 , n955 , n964 );
nand ( n966 , n965 , n881 );
not ( n967 , n966 );
nand ( n968 , n967 , n838 );
not ( n969 , n890 );
not ( n970 , n764 );
or ( n971 , n969 , n970 );
not ( n972 , n897 );
nand ( n973 , n971 , n972 );
not ( n974 , n973 );
not ( n975 , n842 );
not ( n976 , n975 );
not ( n977 , n974 );
or ( n978 , n976 , n977 );
and ( n979 , n974 , n964 );
not ( n980 , n402 );
nand ( n981 , n730 , n741 );
not ( n982 , n981 );
not ( n983 , n747 );
nand ( n984 , n982 , n983 );
nand ( n985 , n980 , n984 );
nor ( n986 , n985 , n404 );
not ( n987 , n986 );
not ( n988 , n764 );
nor ( n989 , n987 , n988 );
nor ( n990 , n979 , n989 );
nand ( n991 , n978 , n990 );
nand ( n992 , n730 , n985 );
and ( n993 , n399 , n992 );
nor ( n994 , n404 , n841 );
not ( n995 , n413 );
not ( n996 , n409 );
nor ( n997 , n996 , n414 );
nand ( n998 , n995 , n997 );
not ( n999 , n998 );
not ( n1000 , n999 );
not ( n1001 , n986 );
or ( n1002 , n1000 , n1001 );
not ( n1003 , n760 );
nand ( n1004 , n1002 , n1003 );
nand ( n1005 , n994 , n1004 );
nand ( n1006 , n991 , n993 , n1005 );
and ( n1007 , n968 , n974 , n1006 );
nand ( n1008 , n939 , n1007 );
and ( n1009 , n944 , n1008 );
and ( n1010 , n64 , n311 );
nor ( n1011 , n717 , n24 );
buf ( n1012 , n1011 );
and ( n1013 , n1010 , n1012 );
not ( n1014 , n1013 );
nor ( n1015 , n1009 , n1014 );
not ( n1016 , n1015 );
nand ( n1017 , n836 , n954 , n1016 );
not ( n1018 , n1017 );
not ( n1019 , n373 );
nand ( n1020 , n265 , n281 );
not ( n1021 , n1020 );
not ( n1022 , n1021 );
not ( n1023 , n1022 );
not ( n1024 , n1023 );
not ( n1025 , n1024 );
nand ( n1026 , n1019 , n1025 );
not ( n1027 , n24 );
and ( n1028 , n311 , n1027 );
nand ( n1029 , n64 , n1028 );
nor ( n1030 , n1026 , n1029 );
and ( n1031 , n359 , n1030 );
nor ( n1032 , n390 , n394 );
or ( n1033 , n790 , n1032 );
nand ( n1034 , n1033 , n796 );
not ( n1035 , n1034 );
nand ( n1036 , n1035 , n1008 );
nand ( n1037 , n1031 , n1036 );
and ( n1038 , n1018 , n1037 );
nor ( n1039 , n1038 , n358 );
not ( n1040 , n359 );
or ( n1041 , n1040 , n373 );
not ( n1042 , n1041 );
nor ( n1043 , n1039 , n1042 );
not ( n1044 , n1043 );
not ( n1045 , n936 );
not ( n1046 , n1045 );
not ( n1047 , n1046 );
not ( n1048 , n966 );
not ( n1049 , n783 );
and ( n1050 , n1049 , n768 );
not ( n1051 , n820 );
nor ( n1052 , n1051 , n1003 );
nand ( n1053 , n1050 , n1052 );
buf ( n1054 , n1053 );
nand ( n1055 , n1048 , n838 , n1054 );
not ( n1056 , n1052 );
nand ( n1057 , n1056 , n973 );
not ( n1058 , n990 );
not ( n1059 , n821 );
not ( n1060 , n1059 );
not ( n1061 , n1060 );
nand ( n1062 , n1061 , n1004 );
nand ( n1063 , n1058 , n993 , n1062 );
and ( n1064 , n1055 , n1057 , n1063 );
nand ( n1065 , n1047 , n1064 );
nand ( n1066 , n943 , n1065 );
not ( n1067 , n64 );
or ( n1068 , n1067 , n1020 );
not ( n1069 , n1068 );
and ( n1070 , n311 , n1069 );
and ( n1071 , n1066 , n1070 );
not ( n1072 , n942 );
not ( n1073 , n838 );
buf ( n1074 , n825 );
not ( n1075 , n1074 );
not ( n1076 , n1075 );
and ( n1077 , n873 , n1076 );
not ( n1078 , n881 );
nor ( n1079 , n1077 , n1078 );
not ( n1080 , n1079 );
or ( n1081 , n1073 , n1080 );
not ( n1082 , n804 );
nand ( n1083 , n413 , n1082 );
nand ( n1084 , n1059 , n1083 );
nand ( n1085 , n730 , n1084 );
and ( n1086 , n873 , n1085 );
nor ( n1087 , n1086 , n930 );
not ( n1088 , n959 );
not ( n1089 , n1088 );
not ( n1090 , n1089 );
not ( n1091 , n731 );
not ( n1092 , n1091 );
not ( n1093 , n1092 );
not ( n1094 , n1093 );
or ( n1095 , n1090 , n1094 );
nand ( n1096 , n1095 , n402 );
nor ( n1097 , n1096 , n898 );
nor ( n1098 , n1087 , n1097 );
nand ( n1099 , n1081 , n1098 );
not ( n1100 , n1099 );
nand ( n1101 , n937 , n1100 );
and ( n1102 , n1072 , n1101 );
not ( n1103 , n311 );
and ( n1104 , n1103 , n1069 );
not ( n1105 , n1104 );
nor ( n1106 , n1102 , n1105 );
nor ( n1107 , n1071 , n1106 );
or ( n1108 , n1107 , n24 );
not ( n1109 , n720 );
and ( n1110 , n1054 , n787 );
and ( n1111 , n311 , n1110 );
not ( n1112 , n311 );
nand ( n1113 , n1074 , n822 );
nor ( n1114 , n404 , n407 );
not ( n1115 , n1114 );
not ( n1116 , n1115 );
nand ( n1117 , n1116 , n870 );
not ( n1118 , n1117 );
nand ( n1119 , n1113 , n402 , n1118 );
not ( n1120 , n822 );
nand ( n1121 , n1120 , n916 );
and ( n1122 , n827 , n1121 );
nand ( n1123 , n1119 , n1122 );
and ( n1124 , n1112 , n1123 );
or ( n1125 , n1111 , n1124 );
or ( n1126 , n1046 , n1125 );
not ( n1127 , n942 );
nand ( n1128 , n1126 , n1127 );
nand ( n1129 , n1109 , n1128 );
nand ( n1130 , n1108 , n1129 );
nand ( n1131 , n358 , n1130 );
not ( n1132 , n1131 );
not ( n1133 , n358 );
not ( n1134 , n1133 );
nor ( n1135 , n1027 , n64 );
nand ( n1136 , n311 , n1135 );
not ( n1137 , n1136 );
and ( n1138 , n1023 , n1137 );
not ( n1139 , n1138 );
not ( n1140 , n1047 );
not ( n1141 , n843 );
and ( n1142 , n407 , n892 );
not ( n1143 , n1142 );
nand ( n1144 , n1143 , n867 );
nand ( n1145 , n1144 , n962 );
nand ( n1146 , n871 , n1145 );
not ( n1147 , n1146 );
not ( n1148 , n1147 );
or ( n1149 , n1141 , n1148 );
not ( n1150 , n399 );
not ( n1151 , n879 );
and ( n1152 , n1150 , n1151 );
nand ( n1153 , n876 , n1152 );
nand ( n1154 , n1149 , n1153 );
not ( n1155 , n1154 );
nand ( n1156 , n838 , n1155 );
not ( n1157 , n893 );
not ( n1158 , n763 );
or ( n1159 , n1157 , n1158 );
not ( n1160 , n889 );
not ( n1161 , n805 );
and ( n1162 , n1160 , n1161 );
nor ( n1163 , n779 , n782 );
nor ( n1164 , n1162 , n1163 );
nand ( n1165 , n1159 , n1164 );
not ( n1166 , n1165 );
and ( n1167 , n759 , n999 , n986 );
not ( n1168 , n1167 );
nand ( n1169 , n994 , n1168 );
not ( n1170 , n989 );
not ( n1171 , n842 );
not ( n1172 , n1147 );
or ( n1173 , n1171 , n1172 );
nand ( n1174 , n1173 , n1166 );
and ( n1175 , n1170 , n1174 );
not ( n1176 , n399 );
and ( n1177 , n1176 , n992 );
not ( n1178 , n1177 );
nor ( n1179 , n1175 , n1178 );
nand ( n1180 , n1169 , n1179 );
nand ( n1181 , n1156 , n1166 , n1180 );
not ( n1182 , n1181 );
not ( n1183 , n1182 );
or ( n1184 , n1140 , n1183 );
nand ( n1185 , n1184 , n943 );
not ( n1186 , n1185 );
or ( n1187 , n1139 , n1186 );
not ( n1188 , n938 );
not ( n1189 , n410 );
not ( n1190 , n416 );
nand ( n1191 , n1190 , n856 );
not ( n1192 , n1191 );
nor ( n1193 , n1192 , n746 );
not ( n1194 , n1114 );
not ( n1195 , n856 );
not ( n1196 , n1195 );
or ( n1197 , n1194 , n1196 );
nand ( n1198 , n1197 , n1091 );
nor ( n1199 , n1193 , n1198 );
nand ( n1200 , n1189 , n1199 );
not ( n1201 , n1200 );
and ( n1202 , n1201 , n1074 );
not ( n1203 , n1202 );
nand ( n1204 , n407 , n414 );
not ( n1205 , n1204 );
nor ( n1206 , n1203 , n1205 );
not ( n1207 , n958 );
not ( n1208 , n1207 );
nor ( n1209 , n414 , n1208 );
not ( n1210 , n1209 );
nand ( n1211 , n402 , n1210 );
nand ( n1212 , n1206 , n1211 );
nand ( n1213 , n770 , n737 );
nand ( n1214 , n1212 , n1213 );
not ( n1215 , n64 );
or ( n1216 , n1027 , n1020 );
or ( n1217 , n1215 , n1216 );
not ( n1218 , n1217 );
nand ( n1219 , n1214 , n1218 );
nand ( n1220 , n859 , n1144 );
nand ( n1221 , n1220 , n871 );
not ( n1222 , n1221 );
and ( n1223 , n843 , n1222 );
not ( n1224 , n1153 );
nor ( n1225 , n1223 , n1224 );
nand ( n1226 , n838 , n1225 );
nand ( n1227 , n893 , n806 );
and ( n1228 , n1227 , n1164 );
and ( n1229 , n929 , n806 );
or ( n1230 , n1221 , n975 );
nand ( n1231 , n1230 , n1228 );
and ( n1232 , n404 , n1231 );
not ( n1233 , n413 );
not ( n1234 , n994 );
or ( n1235 , n1233 , n1234 );
not ( n1236 , n399 );
nand ( n1237 , n1235 , n1236 );
nor ( n1238 , n1232 , n1237 );
nand ( n1239 , n1229 , n1238 );
nand ( n1240 , n1226 , n1228 , n1239 );
not ( n1241 , n1240 );
not ( n1242 , n64 );
not ( n1243 , n311 );
and ( n1244 , n1242 , n1243 );
not ( n1245 , n1216 );
and ( n1246 , n1244 , n1245 );
nand ( n1247 , n1241 , n1246 );
nand ( n1248 , n1219 , n1247 );
and ( n1249 , n1188 , n1248 );
not ( n1250 , n64 );
nand ( n1251 , n311 , n1250 );
not ( n1252 , n1251 );
nor ( n1253 , n1252 , n1216 );
nand ( n1254 , n1253 , n942 );
not ( n1255 , n1254 );
nor ( n1256 , n1249 , n1255 );
nand ( n1257 , n1187 , n1256 );
not ( n1258 , n1257 );
or ( n1259 , n1134 , n1258 );
and ( n1260 , n24 , n358 );
not ( n1261 , n1260 );
not ( n1262 , n1020 );
nand ( n1263 , n311 , n1262 );
or ( n1264 , n64 , n1263 );
nand ( n1265 , n1056 , n1165 );
not ( n1266 , n1265 );
not ( n1267 , n1266 );
and ( n1268 , n1146 , n1265 );
not ( n1269 , n1268 );
nand ( n1270 , n404 , n1269 );
not ( n1271 , n1003 );
nor ( n1272 , n782 , n811 );
not ( n1273 , n1272 );
or ( n1274 , n1271 , n1273 );
nand ( n1275 , n1274 , n730 );
not ( n1276 , n1275 );
not ( n1277 , n1268 );
or ( n1278 , n1276 , n1277 );
nor ( n1279 , n1060 , n1167 );
nand ( n1280 , n1278 , n1279 );
nand ( n1281 , n1270 , n1177 , n1280 );
not ( n1282 , n1154 );
buf ( n1283 , n1054 );
nand ( n1284 , n1282 , n1283 , n838 );
nand ( n1285 , n1267 , n1281 , n1284 );
or ( n1286 , n1264 , n1285 );
not ( n1287 , n1237 );
not ( n1288 , n1121 );
nand ( n1289 , n1287 , n1288 );
and ( n1290 , n1289 , n1076 , n1222 );
nor ( n1291 , n950 , n64 );
or ( n1292 , n1096 , n1228 );
nand ( n1293 , n1290 , n1291 , n1292 );
nand ( n1294 , n1286 , n1293 );
not ( n1295 , n1294 );
or ( n1296 , n1261 , n1295 );
not ( n1297 , n1260 );
or ( n1298 , n1068 , n1297 );
not ( n1299 , n416 );
and ( n1300 , n402 , n1114 );
not ( n1301 , n1300 );
or ( n1302 , n1299 , n1301 );
nand ( n1303 , n407 , n1060 );
and ( n1304 , n1303 , n1050 );
nand ( n1305 , n1302 , n1304 );
or ( n1306 , n1298 , n1305 );
nand ( n1307 , n1296 , n1306 );
and ( n1308 , n940 , n1307 );
not ( n1309 , n942 );
not ( n1310 , n1309 );
and ( n1311 , n358 , n1245 , n1310 );
nor ( n1312 , n1308 , n1311 );
nand ( n1313 , n1259 , n1312 );
nor ( n1314 , n1132 , n1313 );
not ( n1315 , n1314 );
or ( n1316 , n1044 , n1315 );
not ( n1317 , n358 );
not ( n1318 , n1035 );
not ( n1319 , n941 );
or ( n1320 , n1318 , n1319 );
nand ( n1321 , n1320 , n953 );
nand ( n1322 , n1317 , n1037 , n1321 );
nand ( n1323 , n390 , n394 );
not ( n1324 , n1323 );
nor ( n1325 , n1324 , n1032 );
nor ( n1326 , n790 , n1325 );
nand ( n1327 , n766 , n1326 );
not ( n1328 , n1327 );
not ( n1329 , n1027 );
not ( n1330 , n1106 );
or ( n1331 , n1329 , n1330 );
nand ( n1332 , n1331 , n1129 );
not ( n1333 , n1332 );
or ( n1334 , n1328 , n1333 );
not ( n1335 , n1101 );
and ( n1336 , n953 , n1335 );
nand ( n1337 , n1252 , n1011 );
not ( n1338 , n1337 );
not ( n1339 , n1338 );
nor ( n1340 , n1339 , n739 );
not ( n1341 , n1110 );
and ( n1342 , n1340 , n1341 );
not ( n1343 , n311 );
and ( n1344 , n1343 , n1109 );
not ( n1345 , n1344 );
nand ( n1346 , n935 , n1122 );
nor ( n1347 , n1345 , n1346 );
and ( n1348 , n1119 , n1347 );
nor ( n1349 , n1342 , n1348 );
not ( n1350 , n1010 );
nand ( n1351 , n1350 , n1012 );
or ( n1352 , n1033 , n1351 );
nand ( n1353 , n1349 , n358 , n1352 );
nor ( n1354 , n1336 , n1353 );
nand ( n1355 , n1334 , n1354 );
nand ( n1356 , n1322 , n1355 );
and ( n1357 , n1035 , n1065 );
nand ( n1358 , n358 , n1027 );
not ( n1359 , n1358 );
and ( n1360 , n1010 , n1359 );
and ( n1361 , n1023 , n1360 );
not ( n1362 , n1361 );
nor ( n1363 , n1357 , n1362 );
not ( n1364 , n1363 );
not ( n1365 , n1327 );
not ( n1366 , n1365 );
nand ( n1367 , n1366 , n1313 );
not ( n1368 , n940 );
not ( n1369 , n1368 );
not ( n1370 , n358 );
not ( n1371 , n1138 );
not ( n1372 , n1182 );
or ( n1373 , n1371 , n1372 );
nand ( n1374 , n1373 , n1219 );
nand ( n1375 , n1370 , n1374 );
not ( n1376 , n358 );
nand ( n1377 , n1376 , n1135 );
or ( n1378 , n311 , n1377 );
or ( n1379 , n1024 , n1378 );
not ( n1380 , n1379 );
nand ( n1381 , n1380 , n1241 );
not ( n1382 , n1307 );
nand ( n1383 , n1375 , n1381 , n1382 );
and ( n1384 , n1369 , n1383 );
nor ( n1385 , n1216 , n1033 );
nor ( n1386 , n1384 , n1385 );
nand ( n1387 , n1364 , n1367 , n1386 );
not ( n1388 , n1387 );
nand ( n1389 , n1356 , n1042 , n1388 );
nand ( n1390 , n1316 , n1389 );
not ( n1391 , n358 );
nand ( n1392 , n1391 , n1042 );
or ( n1393 , n1365 , n834 );
nand ( n1394 , n1393 , n1033 );
and ( n1395 , n1109 , n1394 );
not ( n1396 , n828 );
nand ( n1397 , n937 , n1396 );
nor ( n1398 , n1345 , n1397 );
and ( n1399 , n807 , n1398 );
not ( n1400 , n1339 );
not ( n1401 , n1400 );
not ( n1402 , n1401 );
not ( n1403 , n1402 );
not ( n1404 , n1403 );
and ( n1405 , n1404 , n788 );
nor ( n1406 , n1395 , n1399 , n1405 );
or ( n1407 , n1392 , n1406 );
nor ( n1408 , n394 , n1041 );
and ( n1409 , n766 , n1408 );
not ( n1410 , n1409 );
not ( n1411 , n1022 );
not ( n1412 , n1411 );
and ( n1413 , n388 , n1412 );
nand ( n1414 , n1410 , n1413 );
nand ( n1415 , n1390 , n1407 , n1414 );
nor ( n1416 , n398 , n406 );
nand ( n1417 , n403 , n1416 );
not ( n1418 , n1417 );
buf ( n1419 , n1418 );
not ( n1420 , n1419 );
nor ( n1421 , n372 , n1420 );
nand ( n1422 , n1415 , n1421 );
not ( n1423 , n398 );
not ( n1424 , n406 );
nand ( n1425 , n403 , n1424 );
nand ( n1426 , n1423 , n1425 );
buf ( n1427 , n1025 );
not ( n1428 , n1213 );
nand ( n1429 , n1427 , n1428 );
and ( n1430 , n790 , n1429 );
or ( n1431 , n1426 , n1430 );
not ( n1432 , n1431 );
nand ( n1433 , n388 , n1409 );
nand ( n1434 , n1432 , n1433 );
and ( n1435 , n358 , n372 );
nand ( n1436 , n1435 , n1419 );
not ( n1437 , n1436 );
not ( n1438 , n953 );
not ( n1439 , n942 );
nor ( n1440 , n1087 , n1079 );
nand ( n1441 , n1045 , n1440 );
nand ( n1442 , n1439 , n1441 );
not ( n1443 , n1442 );
or ( n1444 , n1438 , n1443 );
not ( n1445 , n797 );
not ( n1446 , n1346 );
or ( n1447 , n1445 , n1446 );
nand ( n1448 , n1447 , n1344 );
not ( n1449 , n797 );
not ( n1450 , n739 );
and ( n1451 , n749 , n764 );
nor ( n1452 , n1451 , n771 );
nand ( n1453 , n1450 , n1452 );
not ( n1454 , n1453 );
or ( n1455 , n1449 , n1454 );
nand ( n1456 , n1455 , n1400 );
not ( n1457 , n1452 );
nand ( n1458 , n1457 , n1054 );
nand ( n1459 , n1340 , n1458 );
and ( n1460 , n1448 , n1456 , n1459 );
nand ( n1461 , n1444 , n1460 );
and ( n1462 , n1437 , n1461 );
not ( n1463 , n1462 );
not ( n1464 , n372 );
or ( n1465 , n1464 , n358 );
not ( n1466 , n1419 );
nor ( n1467 , n1465 , n1466 );
buf ( n1468 , n1309 );
not ( n1469 , n1468 );
and ( n1470 , n966 , n1006 );
nand ( n1471 , n939 , n1470 );
not ( n1472 , n1471 );
or ( n1473 , n1469 , n1472 );
nand ( n1474 , n1473 , n1013 );
not ( n1475 , n1072 );
not ( n1476 , n1397 );
or ( n1477 , n1475 , n1476 );
nand ( n1478 , n1477 , n1344 );
nand ( n1479 , n1474 , n1456 , n1478 );
nand ( n1480 , n1467 , n1479 );
nand ( n1481 , n1463 , n1480 );
and ( n1482 , n1327 , n1481 );
not ( n1483 , n1467 );
not ( n1484 , n1471 );
and ( n1485 , n1013 , n1484 );
not ( n1486 , n1401 );
not ( n1487 , n1486 );
not ( n1488 , n1487 );
not ( n1489 , n1488 );
or ( n1490 , n1489 , n1453 );
not ( n1491 , n1025 );
not ( n1492 , n1491 );
not ( n1493 , n311 );
and ( n1494 , n64 , n1493 );
nor ( n1495 , n24 , n1494 );
nand ( n1496 , n1492 , n1495 );
or ( n1497 , n1033 , n1496 );
nand ( n1498 , n1490 , n1497 );
nor ( n1499 , n1485 , n1498 , n1398 );
or ( n1500 , n1483 , n1499 );
not ( n1501 , n1441 );
and ( n1502 , n953 , n1501 );
nand ( n1503 , n1352 , n1459 );
nor ( n1504 , n1502 , n1503 , n1347 );
or ( n1505 , n1436 , n1504 );
nand ( n1506 , n1500 , n1505 );
nor ( n1507 , n1482 , n1506 );
not ( n1508 , n1507 );
not ( n1509 , n358 );
not ( n1510 , n938 );
not ( n1511 , n1510 );
nand ( n1512 , n1218 , n843 );
and ( n1513 , n1238 , n1229 );
nor ( n1514 , n1513 , n1225 );
nand ( n1515 , n1246 , n1514 );
nand ( n1516 , n1512 , n1515 );
not ( n1517 , n1516 );
or ( n1518 , n1511 , n1517 );
nand ( n1519 , n1518 , n1254 );
and ( n1520 , n1169 , n1179 );
nor ( n1521 , n1520 , n1155 );
nand ( n1522 , n1047 , n1521 );
and ( n1523 , n1522 , n1468 );
not ( n1524 , n1138 );
nor ( n1525 , n1523 , n1524 );
nor ( n1526 , n1519 , n1525 );
or ( n1527 , n1365 , n1526 );
not ( n1528 , n1138 );
not ( n1529 , n1521 );
or ( n1530 , n1528 , n1529 );
not ( n1531 , n1516 );
nand ( n1532 , n1530 , n1531 );
not ( n1533 , n1532 );
or ( n1534 , n1533 , n1368 );
not ( n1535 , n1385 );
nand ( n1536 , n1527 , n1534 , n1535 );
nand ( n1537 , n1509 , n1536 );
not ( n1538 , n1298 );
nand ( n1539 , n1045 , n1304 );
not ( n1540 , n1539 );
and ( n1541 , n1538 , n1540 );
and ( n1542 , n358 , n1385 );
nor ( n1543 , n1541 , n1542 );
not ( n1544 , n1543 );
or ( n1545 , n64 , n1297 );
nor ( n1546 , n1263 , n1545 );
not ( n1547 , n1546 );
nand ( n1548 , n1283 , n1155 );
nand ( n1549 , n1281 , n1548 );
nor ( n1550 , n1549 , n938 );
not ( n1551 , n1550 );
or ( n1552 , n1547 , n1551 );
and ( n1553 , n1260 , n1291 );
not ( n1554 , n1553 );
not ( n1555 , n936 );
nand ( n1556 , n1290 , n1555 );
or ( n1557 , n1554 , n1556 );
nand ( n1558 , n1552 , n1557 );
nor ( n1559 , n1544 , n1558 );
nand ( n1560 , n1264 , n1556 );
not ( n1561 , n1560 );
not ( n1562 , n1550 );
or ( n1563 , n1561 , n1562 );
nand ( n1564 , n1563 , n1468 );
not ( n1565 , n1291 );
nor ( n1566 , n1565 , n1556 );
or ( n1567 , n1564 , n1566 );
nand ( n1568 , n1264 , n1565 );
nand ( n1569 , n1567 , n1568 );
nand ( n1570 , n1072 , n1539 );
nand ( n1571 , n1069 , n1570 );
and ( n1572 , n1569 , n1571 );
nor ( n1573 , n1572 , n1297 );
nand ( n1574 , n1327 , n1573 );
nand ( n1575 , n1537 , n1559 , n1574 );
not ( n1576 , n966 );
nand ( n1577 , n1576 , n1054 );
nand ( n1578 , n1577 , n1063 );
not ( n1579 , n1578 );
nand ( n1580 , n1047 , n1579 );
and ( n1581 , n1035 , n1580 );
nor ( n1582 , n1581 , n1362 );
or ( n1583 , n1575 , n1582 );
and ( n1584 , n372 , n403 );
nand ( n1585 , n1584 , n1416 );
not ( n1586 , n1585 );
nand ( n1587 , n1583 , n1586 );
not ( n1588 , n1587 );
or ( n1589 , n1508 , n1588 );
nand ( n1590 , n1589 , n1042 );
not ( n1591 , n358 );
nand ( n1592 , n932 , n882 );
not ( n1593 , n1592 );
nand ( n1594 , n1593 , n1188 );
not ( n1595 , n1594 );
nor ( n1596 , n1595 , n1034 );
or ( n1597 , n1596 , n952 , n1392 );
nand ( n1598 , n944 , n1594 );
and ( n1599 , n1598 , n953 );
nor ( n1600 , n1599 , n1479 );
or ( n1601 , n1600 , n1042 );
nand ( n1602 , n1597 , n1601 );
and ( n1603 , n1591 , n1602 );
not ( n1604 , n1414 );
nor ( n1605 , n1603 , n1604 );
nor ( n1606 , n1585 , n1605 );
nor ( n1607 , n1014 , n1436 );
nand ( n1608 , n1468 , n1580 );
nand ( n1609 , n1607 , n1608 );
not ( n1610 , n358 );
not ( n1611 , n1526 );
nand ( n1612 , n1610 , n1611 );
not ( n1613 , n1573 );
nand ( n1614 , n1612 , n1613 );
and ( n1615 , n1586 , n1614 );
nor ( n1616 , n1615 , n1462 );
and ( n1617 , n1609 , n1616 );
nor ( n1618 , n1617 , n1042 );
nor ( n1619 , n1606 , n1618 );
nand ( n1620 , n1422 , n1434 , n1590 , n1619 );
not ( n1621 , n401 );
nand ( n1622 , n1620 , n1621 );
nor ( n1623 , n1423 , n401 );
nand ( n1624 , n406 , n1623 );
not ( n1625 , n401 );
or ( n1626 , n1625 , n1418 );
nand ( n1627 , n1624 , n1626 );
not ( n1628 , n1627 );
nor ( n1629 , n1628 , n1430 );
nand ( n1630 , n1433 , n1629 );
not ( n1631 , n1492 );
not ( n1632 , n401 );
or ( n1633 , n1632 , n1417 );
not ( n1634 , n1633 );
nand ( n1635 , n1631 , n1634 );
not ( n1636 , n1326 );
or ( n1637 , n1019 , n1636 );
nand ( n1638 , n388 , n390 );
or ( n1639 , n373 , n1638 );
nand ( n1640 , n1637 , n1639 );
not ( n1641 , n1640 );
nand ( n1642 , n44 , n344 );
not ( n1643 , n44 );
not ( n1644 , n344 );
nand ( n1645 , n1643 , n1644 );
nand ( n1646 , n1642 , n1645 );
nand ( n1647 , n388 , n1325 );
not ( n1648 , n1647 );
nand ( n1649 , n1646 , n1648 );
nand ( n1650 , n1641 , n1649 );
not ( n1651 , n1650 );
or ( n1652 , n1635 , n1651 );
nand ( n1653 , n1652 , n359 );
not ( n1654 , n1492 );
not ( n1655 , n1623 );
or ( n1656 , n1655 , n1425 );
nor ( n1657 , n1654 , n1656 );
not ( n1658 , n1657 );
not ( n1659 , n1492 );
not ( n1660 , n1659 );
nor ( n1661 , n403 , n406 );
nand ( n1662 , n1623 , n1661 );
nor ( n1663 , n1660 , n1662 );
not ( n1664 , n1663 );
and ( n1665 , n1658 , n1664 );
not ( n1666 , n1645 );
not ( n1667 , n1666 );
not ( n1668 , n1667 );
not ( n1669 , n1668 );
buf ( n1670 , n1648 );
nand ( n1671 , n1669 , n1670 );
not ( n1672 , n1671 );
and ( n1673 , n1663 , n1672 );
not ( n1674 , n1657 );
not ( n1675 , n1672 );
and ( n1676 , n1674 , n1675 );
nand ( n1677 , n1643 , n1648 );
not ( n1678 , n1677 );
nor ( n1679 , n1678 , n1428 );
nor ( n1680 , n1676 , n1679 );
nor ( n1681 , n1673 , n1640 , n1680 );
nor ( n1682 , n1665 , n1681 );
nor ( n1683 , n1631 , n1662 );
not ( n1684 , n1325 );
or ( n1685 , n1667 , n1684 );
nand ( n1686 , n388 , n1685 );
nand ( n1687 , n1686 , n1213 );
and ( n1688 , n1683 , n1687 );
nand ( n1689 , n1636 , n1677 );
and ( n1690 , n1491 , n1689 );
not ( n1691 , n1690 );
nor ( n1692 , n1691 , n1656 );
nor ( n1693 , n1688 , n1692 );
not ( n1694 , n1693 );
not ( n1695 , n1631 );
nand ( n1696 , n1695 , n1634 );
nand ( n1697 , n1636 , n1649 );
nor ( n1698 , n1428 , n1697 );
nor ( n1699 , n1696 , n1698 );
nor ( n1700 , n1694 , n1699 );
and ( n1701 , n373 , n1700 );
and ( n1702 , n1649 , n1638 , n1213 );
nor ( n1703 , n1702 , n1696 );
not ( n1704 , n1703 );
nand ( n1705 , n394 , n1643 );
not ( n1706 , n388 );
nor ( n1707 , n1706 , n390 );
nand ( n1708 , n1705 , n1707 );
not ( n1709 , n1708 );
nor ( n1710 , n1709 , n1656 );
and ( n1711 , n1413 , n1710 );
nand ( n1712 , n1638 , n1671 );
or ( n1713 , n1712 , n1428 );
nand ( n1714 , n1713 , n1683 );
not ( n1715 , n1714 );
nor ( n1716 , n1711 , n373 , n1715 );
and ( n1717 , n1704 , n1716 );
nor ( n1718 , n1701 , n1717 );
or ( n1719 , n1653 , n1682 , n1718 );
not ( n1720 , n1697 );
or ( n1721 , n1635 , n1720 );
not ( n1722 , n1664 );
not ( n1723 , n1686 );
and ( n1724 , n1722 , n1723 );
nand ( n1725 , n1636 , n1679 );
and ( n1726 , n1657 , n1725 );
nor ( n1727 , n1724 , n1726 );
nand ( n1728 , n1721 , n1727 );
not ( n1729 , n1700 );
or ( n1730 , n1728 , n359 , n1729 );
nand ( n1731 , n1719 , n1730 );
nand ( n1732 , n1622 , n1630 , n1731 );
and ( n1733 , n716 , n1732 );
not ( n1734 , n389 );
not ( n1735 , n395 );
nand ( n1736 , n393 , n1735 );
not ( n1737 , n401 );
not ( n1738 , n1586 );
not ( n1739 , n358 );
nand ( n1740 , n1739 , n948 );
not ( n1741 , n1740 );
nand ( n1742 , n951 , n1741 );
not ( n1743 , n1742 );
and ( n1744 , n1743 , n1598 );
not ( n1745 , n1744 );
nand ( n1746 , n1359 , n1494 );
or ( n1747 , n1024 , n1746 );
not ( n1748 , n1747 );
nand ( n1749 , n1748 , n1442 );
not ( n1750 , n64 );
nand ( n1751 , n1750 , n1413 );
and ( n1752 , n1751 , n1569 );
nor ( n1753 , n1752 , n1297 );
not ( n1754 , n1753 );
nand ( n1755 , n1745 , n1749 , n1754 );
not ( n1756 , n1755 );
or ( n1757 , n1738 , n1756 );
and ( n1758 , n1586 , n1538 , n1570 );
and ( n1759 , n358 , n1464 );
not ( n1760 , n1759 );
nor ( n1761 , n1760 , n1420 );
not ( n1762 , n1761 );
nor ( n1763 , n24 , n358 );
not ( n1764 , n1763 );
nor ( n1765 , n1464 , n1764 );
or ( n1766 , n1464 , n1297 );
nor ( n1767 , n64 , n1766 );
nor ( n1768 , n1464 , n1358 );
and ( n1769 , n64 , n1768 );
or ( n1770 , n1767 , n1769 );
nor ( n1771 , n1765 , n1770 );
nor ( n1772 , n1420 , n1771 );
not ( n1773 , n1772 );
and ( n1774 , n1762 , n1773 );
nand ( n1775 , n24 , n64 );
not ( n1776 , n719 );
nand ( n1777 , n1775 , n1776 );
nand ( n1778 , n358 , n1777 );
nand ( n1779 , n1413 , n1778 );
nor ( n1780 , n1774 , n1779 );
nor ( n1781 , n1758 , n1780 );
or ( n1782 , n1436 , n1460 );
not ( n1783 , n1129 );
nand ( n1784 , n1783 , n1761 );
and ( n1785 , n1781 , n1782 , n1431 , n1784 );
nand ( n1786 , n1757 , n1785 );
not ( n1787 , n1786 );
and ( n1788 , n1609 , n1480 );
not ( n1789 , n954 );
nand ( n1790 , n24 , n388 );
nor ( n1791 , n1492 , n1790 );
nor ( n1792 , n1015 , n1791 );
not ( n1793 , n1257 );
nand ( n1794 , n1792 , n1793 );
not ( n1795 , n1794 );
not ( n1796 , n1795 );
or ( n1797 , n1789 , n1796 );
not ( n1798 , n358 );
nand ( n1799 , n1797 , n1798 );
and ( n1800 , n1763 , n1291 );
and ( n1801 , n1800 , n832 );
and ( n1802 , n1764 , n1545 );
not ( n1803 , n1413 );
nor ( n1804 , n1802 , n1803 );
nor ( n1805 , n1801 , n1804 );
not ( n1806 , n1264 );
and ( n1807 , n1806 , n1763 );
nand ( n1808 , n1807 , n798 );
nand ( n1809 , n1805 , n1808 , n1312 );
not ( n1810 , n1809 );
and ( n1811 , n1799 , n1810 );
nor ( n1812 , n1811 , n372 );
nor ( n1813 , n24 , n1760 );
not ( n1814 , n1813 );
or ( n1815 , n1814 , n1107 );
not ( n1816 , n1791 );
and ( n1817 , n1526 , n1816 );
or ( n1818 , n1465 , n1817 );
nand ( n1819 , n1815 , n1818 );
or ( n1820 , n1812 , n1819 );
not ( n1821 , n1420 );
not ( n1822 , n1821 );
not ( n1823 , n1822 );
not ( n1824 , n1823 );
not ( n1825 , n1824 );
nand ( n1826 , n1820 , n1825 );
nand ( n1827 , n1787 , n1788 , n1826 );
nand ( n1828 , n1737 , n1827 );
or ( n1829 , n44 , n1670 );
not ( n1830 , n1646 );
nand ( n1831 , n1829 , n1830 );
nand ( n1832 , n388 , n1831 );
nor ( n1833 , n1635 , n1832 );
nor ( n1834 , n1833 , n1629 );
nand ( n1835 , n1828 , n1700 , n1727 , n1834 );
and ( n1836 , n1734 , n1736 , n1835 );
nor ( n1837 , n1733 , n1836 );
or ( n1838 , n714 , n1837 );
nand ( n1839 , n358 , n1643 );
nor ( n1840 , n344 , n1839 );
not ( n1841 , n1670 );
not ( n1842 , n1841 );
not ( n1843 , n1842 );
not ( n1844 , n1843 );
not ( n1845 , n1844 );
not ( n1846 , n1109 );
not ( n1847 , n394 );
nand ( n1848 , n386 , n1847 );
or ( n1849 , n737 , n1848 );
buf ( n1850 , n1849 );
buf ( n1851 , n1850 );
not ( n1852 , n1851 );
buf ( n1853 , n1852 );
or ( n1854 , n1125 , n1853 );
nor ( n1855 , n392 , n394 );
nand ( n1856 , n737 , n794 , n1855 );
and ( n1857 , n790 , n1856 );
not ( n1858 , n1857 );
not ( n1859 , n1858 );
not ( n1860 , n1859 );
not ( n1861 , n1860 );
nand ( n1862 , n1854 , n1861 );
not ( n1863 , n1862 );
or ( n1864 , n1846 , n1863 );
not ( n1865 , n1860 );
not ( n1866 , n1865 );
not ( n1867 , n1852 );
nand ( n1868 , n1867 , n1100 );
not ( n1869 , n1868 );
or ( n1870 , n1866 , n1869 );
nand ( n1871 , n1870 , n953 );
nand ( n1872 , n1864 , n1871 );
and ( n1873 , n1845 , n1872 );
nand ( n1874 , n1400 , n1851 );
or ( n1875 , n1874 , n1110 );
not ( n1876 , n1119 );
nand ( n1877 , n1851 , n1122 );
not ( n1878 , n1877 );
nand ( n1879 , n1878 , n1344 );
or ( n1880 , n1876 , n1879 );
not ( n1881 , n1868 );
and ( n1882 , n953 , n1881 );
nor ( n1883 , n1636 , n1351 );
nor ( n1884 , n1882 , n1883 );
nand ( n1885 , n1875 , n1880 , n1884 );
nor ( n1886 , n1873 , n1885 );
not ( n1887 , n1886 );
and ( n1888 , n1840 , n1887 );
not ( n1889 , n1669 );
not ( n1890 , n1889 );
not ( n1891 , n1890 );
nor ( n1892 , n358 , n1891 );
not ( n1893 , n1865 );
not ( n1894 , n1893 );
not ( n1895 , n1894 );
not ( n1896 , n1895 );
buf ( n1897 , n1867 );
not ( n1898 , n1897 );
nor ( n1899 , n1898 , n933 );
not ( n1900 , n1899 );
nand ( n1901 , n1896 , n1900 );
not ( n1902 , n1901 );
or ( n1903 , n1902 , n952 );
not ( n1904 , n787 );
nand ( n1905 , n1849 , n1904 );
nand ( n1906 , n1857 , n1905 );
not ( n1907 , n1906 );
nand ( n1908 , n1907 , n311 );
not ( n1909 , n311 );
not ( n1910 , n1850 );
not ( n1911 , n829 );
nor ( n1912 , n1910 , n1911 );
nor ( n1913 , n1858 , n1912 );
nand ( n1914 , n1909 , n1913 );
nand ( n1915 , n1908 , n1109 , n1914 );
nand ( n1916 , n1903 , n1915 );
and ( n1917 , n1892 , n1916 );
nor ( n1918 , n1888 , n1917 );
not ( n1919 , n1891 );
not ( n1920 , n1919 );
not ( n1921 , n1920 );
nand ( n1922 , n1897 , n1007 );
nand ( n1923 , n1894 , n1922 );
or ( n1924 , n1263 , n1740 );
not ( n1925 , n1924 );
nand ( n1926 , n1923 , n1925 );
buf ( n1927 , n1865 );
not ( n1928 , n1927 );
nand ( n1929 , n1897 , n1064 );
not ( n1930 , n1929 );
or ( n1931 , n1928 , n1930 );
nand ( n1932 , n1931 , n1361 );
nand ( n1933 , n1872 , n358 );
nand ( n1934 , n1932 , n1933 );
not ( n1935 , n1852 );
nand ( n1936 , n1935 , n1290 );
not ( n1937 , n1292 );
or ( n1938 , n1936 , n1937 );
nand ( n1939 , n1938 , n1861 );
and ( n1940 , n1553 , n1939 );
not ( n1941 , n1867 );
not ( n1942 , n1214 );
or ( n1943 , n1941 , n1942 );
nand ( n1944 , n1943 , n1861 );
or ( n1945 , n358 , n1775 );
or ( n1946 , n1412 , n1945 );
not ( n1947 , n1946 );
and ( n1948 , n1944 , n1947 );
nor ( n1949 , n1940 , n1948 );
and ( n1950 , n1861 , n1305 );
not ( n1951 , n1857 );
nand ( n1952 , n1850 , n1304 );
not ( n1953 , n1952 );
or ( n1954 , n1951 , n1953 );
nand ( n1955 , n1954 , n1538 );
nor ( n1956 , n1950 , n1955 );
nand ( n1957 , n1897 , n1182 );
and ( n1958 , n1894 , n1957 );
not ( n1959 , n1263 );
not ( n1960 , n1377 );
and ( n1961 , n1959 , n1960 );
not ( n1962 , n1961 );
nor ( n1963 , n1958 , n1962 );
nor ( n1964 , n1956 , n1963 );
not ( n1965 , n1897 );
or ( n1966 , n1965 , n1285 );
not ( n1967 , n1861 );
not ( n1968 , n1967 );
nand ( n1969 , n1966 , n1968 );
and ( n1970 , n1969 , n1546 );
nand ( n1971 , n1897 , n1241 );
and ( n1972 , n1927 , n1971 );
nor ( n1973 , n1972 , n1379 );
nor ( n1974 , n1970 , n1973 );
nand ( n1975 , n1949 , n1964 , n1974 );
nor ( n1976 , n1934 , n1975 );
nand ( n1977 , n1926 , n1976 );
and ( n1978 , n1921 , n1977 );
not ( n1979 , n1921 );
not ( n1980 , n358 );
nand ( n1981 , n1636 , n1856 );
not ( n1982 , n1981 );
and ( n1983 , n1982 , n1929 );
nor ( n1984 , n1983 , n1014 );
not ( n1985 , n1984 );
or ( n1986 , n1980 , n1985 );
not ( n1987 , n1922 );
or ( n1988 , n1987 , n1981 );
nand ( n1989 , n1988 , n1013 );
not ( n1990 , n1989 );
nand ( n1991 , n1850 , n1396 );
nor ( n1992 , n1345 , n1991 );
and ( n1993 , n807 , n1992 );
not ( n1994 , n1905 );
and ( n1995 , n1488 , n1994 );
or ( n1996 , n1915 , n1844 );
nand ( n1997 , n1109 , n1326 );
nand ( n1998 , n1996 , n1997 );
nor ( n1999 , n1993 , n1995 , n1998 );
not ( n2000 , n1999 );
or ( n2001 , n1990 , n2000 );
not ( n2002 , n358 );
nand ( n2003 , n2001 , n2002 );
not ( n2004 , n1845 );
not ( n2005 , n2004 );
and ( n2006 , n1975 , n2005 );
nor ( n2007 , n1216 , n1636 );
nor ( n2008 , n2006 , n2007 );
not ( n2009 , n1898 );
and ( n2010 , n2009 , n1383 );
not ( n2011 , n1899 );
not ( n2012 , n1981 );
and ( n2013 , n2011 , n2012 );
nor ( n2014 , n2013 , n1742 );
nor ( n2015 , n2010 , n2014 );
nand ( n2016 , n2003 , n2008 , n2015 );
not ( n2017 , n2016 );
nand ( n2018 , n1986 , n2017 );
and ( n2019 , n1979 , n2018 );
nor ( n2020 , n1978 , n2019 );
nand ( n2021 , n1413 , n1685 );
and ( n2022 , n1918 , n2020 , n2021 );
nor ( n2023 , n372 , n403 );
nand ( n2024 , n398 , n1424 );
nor ( n2025 , n401 , n2024 );
nand ( n2026 , n2023 , n2025 );
nor ( n2027 , n2022 , n2026 );
not ( n2028 , n403 );
nor ( n2029 , n2028 , n372 );
not ( n2030 , n2029 );
not ( n2031 , n2025 );
nor ( n2032 , n2030 , n2031 );
not ( n2033 , n2032 );
not ( n2034 , n1984 );
nand ( n2035 , n2034 , n1886 );
nand ( n2036 , n358 , n2035 );
not ( n2037 , n2036 );
nor ( n2038 , n2037 , n2016 );
or ( n2039 , n2038 , n1643 );
not ( n2040 , n1976 );
and ( n2041 , n1643 , n2040 );
nor ( n2042 , n2041 , n1690 );
not ( n2043 , n1923 );
nor ( n2044 , n1014 , n2043 );
or ( n2045 , n1916 , n2044 );
nor ( n2046 , n44 , n358 );
nand ( n2047 , n2045 , n2046 );
nand ( n2048 , n2039 , n2042 , n2047 );
not ( n2049 , n2048 );
or ( n2050 , n2033 , n2049 );
nand ( n2051 , n953 , n1593 );
not ( n2052 , n1790 );
nor ( n2053 , n2052 , n1532 );
nand ( n2054 , n2051 , n2053 );
not ( n2055 , n2054 );
or ( n2056 , n2055 , n1465 );
not ( n2057 , n1747 );
not ( n2058 , n1099 );
and ( n2059 , n2057 , n2058 );
and ( n2060 , n1807 , n1904 );
nor ( n2061 , n2059 , n2060 );
nand ( n2062 , n1800 , n829 );
nand ( n2063 , n2061 , n1306 , n2062 );
and ( n2064 , n2063 , n1464 );
nor ( n2065 , n1760 , n1487 );
and ( n2066 , n2065 , n1341 );
not ( n2067 , n358 );
nor ( n2068 , n2067 , n64 );
nor ( n2069 , n24 , n311 );
nand ( n2070 , n2068 , n2069 );
not ( n2071 , n2070 );
nand ( n2072 , n1023 , n2071 );
nor ( n2073 , n372 , n2072 );
not ( n2074 , n1123 );
and ( n2075 , n2073 , n2074 );
nor ( n2076 , n2064 , n2066 , n2075 );
not ( n2077 , n1766 );
not ( n2078 , n64 );
nand ( n2079 , n388 , n2078 );
not ( n2080 , n2079 );
or ( n2081 , n1264 , n1549 );
nand ( n2082 , n1291 , n1290 );
nand ( n2083 , n2081 , n2082 );
nor ( n2084 , n2080 , n2083 );
not ( n2085 , n2084 );
and ( n2086 , n2077 , n2085 );
nor ( n2087 , n372 , n1740 );
nand ( n2088 , n1104 , n2087 );
nor ( n2089 , n2088 , n933 );
nor ( n2090 , n2086 , n2089 );
nand ( n2091 , n2056 , n2076 , n2090 );
not ( n2092 , n2091 );
nor ( n2093 , n64 , n1024 );
nand ( n2094 , n358 , n1028 );
not ( n2095 , n2094 );
nand ( n2096 , n2093 , n2095 );
nor ( n2097 , n1464 , n2096 );
and ( n2098 , n2097 , n1458 );
not ( n2099 , n358 );
nand ( n2100 , n24 , n2099 );
and ( n2101 , n1464 , n1778 );
nand ( n2102 , n2100 , n2101 );
nand ( n2103 , n2102 , n1771 );
and ( n2104 , n388 , n2103 );
nand ( n2105 , n1069 , n2077 );
not ( n2106 , n2105 );
and ( n2107 , n2106 , n1304 );
nor ( n2108 , n2098 , n2104 , n2107 );
nor ( n2109 , n372 , n1297 );
not ( n2110 , n1294 );
nand ( n2111 , n2079 , n2110 );
nand ( n2112 , n2109 , n2111 );
nand ( n2113 , n1013 , n1007 );
not ( n2114 , n1247 );
not ( n2115 , n2114 );
not ( n2116 , n1374 );
nand ( n2117 , n2115 , n2116 , n1790 );
not ( n2118 , n2117 );
and ( n2119 , n2113 , n2118 );
or ( n2120 , n358 , n372 );
nor ( n2121 , n2119 , n2120 );
buf ( n2122 , n1064 );
nand ( n2123 , n1013 , n1759 , n2122 );
not ( n2124 , n2123 );
nor ( n2125 , n2121 , n2124 );
nand ( n2126 , n2092 , n2108 , n2112 , n2125 );
not ( n2127 , n1824 );
nand ( n2128 , n2126 , n2127 );
and ( n2129 , n1768 , n1104 );
and ( n2130 , n1821 , n2129 );
and ( n2131 , n2130 , n1440 );
nor ( n2132 , n1585 , n2072 );
and ( n2133 , n2132 , n1122 );
nand ( n2134 , n1586 , n1800 );
or ( n2135 , n2134 , n828 );
not ( n2136 , n1489 );
nand ( n2137 , n2136 , n1467 );
not ( n2138 , n1457 );
not ( n2139 , n2138 );
or ( n2140 , n2137 , n2139 );
nand ( n2141 , n2135 , n2140 );
nor ( n2142 , n2131 , n2133 , n2141 );
nor ( n2143 , n1585 , n1924 );
and ( n2144 , n2143 , n1470 );
and ( n2145 , n1607 , n1579 );
nor ( n2146 , n2144 , n2145 );
nand ( n2147 , n2128 , n2142 , n2146 );
or ( n2148 , n1853 , n955 );
nand ( n2149 , n2148 , n1865 );
nand ( n2150 , n1947 , n2149 );
not ( n2151 , n2150 );
nor ( n2152 , n1298 , n1952 );
nor ( n2153 , n2151 , n2152 );
nand ( n2154 , n1897 , n1470 );
nand ( n2155 , n1927 , n2154 );
nand ( n2156 , n1925 , n2155 );
nor ( n2157 , n1853 , n1578 );
nor ( n2158 , n2157 , n1893 );
nor ( n2159 , n2158 , n1014 );
nand ( n2160 , n358 , n2159 );
not ( n2161 , n1861 );
not ( n2162 , n1936 );
or ( n2163 , n2161 , n2162 );
nand ( n2164 , n2163 , n1553 );
nand ( n2165 , n2156 , n2160 , n2164 );
not ( n2166 , n1800 );
not ( n2167 , n1858 );
and ( n2168 , n2167 , n1991 );
nor ( n2169 , n2166 , n2168 );
nor ( n2170 , n2165 , n2169 );
and ( n2171 , n2153 , n2170 );
nor ( n2172 , n2171 , n1464 );
not ( n2173 , n2172 );
not ( n2174 , n2088 );
nand ( n2175 , n2174 , n1901 );
not ( n2176 , n1765 );
nor ( n2177 , n2176 , n1105 );
nor ( n2178 , n1592 , n1898 );
nor ( n2179 , n2178 , n1895 );
not ( n2180 , n2179 );
nand ( n2181 , n2177 , n2180 );
nand ( n2182 , n1974 , n1932 , n1464 );
not ( n2183 , n1963 );
nand ( n2184 , n2183 , n1926 );
or ( n2185 , n2182 , n2184 );
not ( n2186 , n1860 );
not ( n2187 , n2186 );
not ( n2188 , n1852 );
nand ( n2189 , n2188 , n1440 );
not ( n2190 , n2189 );
or ( n2191 , n2187 , n2190 );
nand ( n2192 , n2191 , n953 );
not ( n2193 , n1874 );
nand ( n2194 , n2193 , n1458 );
nand ( n2195 , n1849 , n1452 );
and ( n2196 , n1857 , n2195 );
nor ( n2197 , n2196 , n1339 );
and ( n2198 , n1859 , n1877 );
nor ( n2199 , n2198 , n1345 );
nor ( n2200 , n2197 , n2199 );
nand ( n2201 , n2192 , n2194 , n2200 );
nand ( n2202 , n358 , n2201 );
not ( n2203 , n1853 );
and ( n2204 , n2203 , n1514 );
nor ( n2205 , n2204 , n1967 );
nor ( n2206 , n2205 , n1379 );
nand ( n2207 , n2203 , n1521 );
and ( n2208 , n2207 , n1927 );
nor ( n2209 , n2208 , n1962 );
nor ( n2210 , n2206 , n2209 );
not ( n2211 , n1968 );
not ( n2212 , n1549 );
nand ( n2213 , n2203 , n2212 );
not ( n2214 , n2213 );
or ( n2215 , n2211 , n2214 );
nand ( n2216 , n2215 , n1546 );
nand ( n2217 , n2202 , n2210 , n2216 , n372 );
nand ( n2218 , n2185 , n2217 );
nand ( n2219 , n2175 , n2181 , n2218 );
not ( n2220 , n2219 );
and ( n2221 , n1933 , n1949 );
nor ( n2222 , n2221 , n372 );
nor ( n2223 , n372 , n2166 );
not ( n2224 , n2223 );
or ( n2225 , n2224 , n1913 );
not ( n2226 , n1465 );
and ( n2227 , n2226 , n2197 );
nor ( n2228 , n2120 , n1487 );
and ( n2229 , n2228 , n1906 );
not ( n2230 , n1779 );
nor ( n2231 , n2227 , n2229 , n2230 );
not ( n2232 , n1956 );
nand ( n2233 , n2225 , n2231 , n2232 );
nor ( n2234 , n2222 , n2233 );
nand ( n2235 , n2173 , n2220 , n2234 );
not ( n2236 , n2235 );
nor ( n2237 , n2236 , n1426 );
or ( n2238 , n2147 , n2237 );
not ( n2239 , n401 );
nand ( n2240 , n2238 , n2239 );
nand ( n2241 , n2050 , n2240 );
nor ( n2242 , n2027 , n2241 );
nor ( n2243 , n1902 , n1742 );
or ( n2244 , n2243 , n1977 );
nand ( n2245 , n2244 , n1646 );
not ( n2246 , n358 );
or ( n2247 , n1830 , n1915 );
or ( n2248 , n1646 , n1989 );
not ( n2249 , n311 );
nand ( n2250 , n2249 , n948 );
not ( n2251 , n265 );
not ( n2252 , n311 );
nand ( n2253 , n2252 , n265 );
or ( n2254 , n281 , n2253 );
not ( n2255 , n2254 );
or ( n2256 , n2251 , n2255 );
nand ( n2257 , n2256 , n1697 );
or ( n2258 , n2250 , n2257 );
nand ( n2259 , n2247 , n2248 , n2258 );
nand ( n2260 , n2246 , n2259 );
nand ( n2261 , n344 , n2046 );
not ( n2262 , n2261 );
not ( n2263 , n1999 );
and ( n2264 , n2262 , n2263 );
nand ( n2265 , n1494 , n1763 );
nand ( n2266 , n1413 , n1831 );
not ( n2267 , n2266 );
and ( n2268 , n2265 , n2267 );
nor ( n2269 , n2264 , n2268 );
nand ( n2270 , n2245 , n2260 , n2269 );
and ( n2271 , n2008 , n2015 );
and ( n2272 , n2271 , n2036 );
or ( n2273 , n1644 , n44 );
nor ( n2274 , n2272 , n2273 );
or ( n2275 , n2270 , n2274 );
nor ( n2276 , n372 , n1633 );
nand ( n2277 , n2275 , n2276 );
not ( n2278 , n2004 );
nand ( n2279 , n2216 , n1955 , n2164 );
nand ( n2280 , n2278 , n2279 );
or ( n2281 , n1547 , n2213 );
not ( n2282 , n1246 );
or ( n2283 , n2282 , n1936 );
not ( n2284 , n2007 );
nand ( n2285 , n2283 , n2284 );
and ( n2286 , n358 , n2285 );
nor ( n2287 , n2286 , n2152 );
nand ( n2288 , n2280 , n2281 , n2287 );
and ( n2289 , n1845 , n2201 );
nor ( n2290 , n2289 , n1883 );
not ( n2291 , n2189 );
nand ( n2292 , n2291 , n953 );
and ( n2293 , n1879 , n2194 );
nand ( n2294 , n2290 , n2292 , n2293 );
not ( n2295 , n2294 );
not ( n2296 , n358 );
nor ( n2297 , n2295 , n2296 );
nor ( n2298 , n2288 , n2297 );
and ( n2299 , n44 , n2298 );
not ( n2300 , n44 );
not ( n2301 , n2279 );
and ( n2302 , n2300 , n2301 );
or ( n2303 , n2299 , n2302 );
not ( n2304 , n1013 );
nand ( n2305 , n1982 , n2154 );
not ( n2306 , n2305 );
or ( n2307 , n2304 , n2306 );
or ( n2308 , n2178 , n1981 );
nand ( n2309 , n2308 , n953 );
nand ( n2310 , n2307 , n2309 );
or ( n2311 , n1643 , n2310 );
not ( n2312 , n2179 );
not ( n2313 , n952 );
and ( n2314 , n2312 , n2313 );
not ( n2315 , n2155 );
nor ( n2316 , n2315 , n1014 );
nor ( n2317 , n2314 , n2316 );
and ( n2318 , n2317 , n1643 );
nor ( n2319 , n2318 , n358 );
and ( n2320 , n2311 , n2319 );
not ( n2321 , n2201 );
not ( n2322 , n2159 );
nand ( n2323 , n2321 , n2322 );
not ( n2324 , n2323 );
and ( n2325 , n2324 , n1643 );
not ( n2326 , n2157 );
nand ( n2327 , n1982 , n2326 );
nand ( n2328 , n1013 , n2327 );
and ( n2329 , n44 , n2328 );
nor ( n2330 , n2325 , n2329 );
not ( n2331 , n2330 );
not ( n2332 , n1690 );
and ( n2333 , n2331 , n2332 );
not ( n2334 , n358 );
nor ( n2335 , n2333 , n2334 );
nor ( n2336 , n2320 , n2335 );
and ( n2337 , n2303 , n2336 );
not ( n2338 , n1584 );
nor ( n2339 , n2338 , n2031 );
not ( n2340 , n2339 );
nor ( n2341 , n2337 , n2340 );
not ( n2342 , n2235 );
nor ( n2343 , n2342 , n1628 );
nor ( n2344 , n2341 , n2343 );
not ( n2345 , n358 );
or ( n2346 , n2168 , n1345 );
not ( n2347 , n2197 );
nand ( n2348 , n2346 , n2347 );
and ( n2349 , n2348 , n1845 );
not ( n2350 , n2195 );
and ( n2351 , n1404 , n2350 );
not ( n2352 , n1992 );
nand ( n2353 , n2352 , n1997 );
nor ( n2354 , n2349 , n2351 , n2353 );
not ( n2355 , n2354 );
nand ( n2356 , n2345 , n2355 );
nand ( n2357 , n2210 , n2150 );
and ( n2358 , n2005 , n2357 );
and ( n2359 , n2009 , n1532 );
nor ( n2360 , n2359 , n2007 );
nor ( n2361 , n2360 , n358 );
nor ( n2362 , n2358 , n2361 );
and ( n2363 , n2356 , n2362 );
nand ( n2364 , n44 , n2339 );
not ( n2365 , n2273 );
and ( n2366 , n401 , n1586 );
nand ( n2367 , n2365 , n2366 );
and ( n2368 , n2364 , n2367 );
nor ( n2369 , n2363 , n2368 );
and ( n2370 , n1643 , n2339 );
not ( n2371 , n2366 );
nor ( n2372 , n1830 , n2371 );
nor ( n2373 , n2370 , n2372 );
not ( n2374 , n358 );
and ( n2375 , n2374 , n2348 );
nor ( n2376 , n2375 , n2357 );
or ( n2377 , n2373 , n2376 );
nand ( n2378 , n2372 , n1743 , n2180 );
nor ( n2379 , n1924 , n2367 );
and ( n2380 , n2379 , n2305 );
and ( n2381 , n2226 , n1833 );
nor ( n2382 , n2380 , n2381 );
nand ( n2383 , n2377 , n2378 , n2382 );
nor ( n2384 , n2369 , n2383 );
not ( n2385 , n358 );
or ( n2386 , n2367 , n2309 );
and ( n2387 , n2372 , n2316 );
and ( n2388 , n372 , n1692 );
nor ( n2389 , n2387 , n2388 );
nand ( n2390 , n2386 , n2389 );
nand ( n2391 , n2385 , n2390 );
or ( n2392 , n2298 , n2273 );
nand ( n2393 , n358 , n2323 );
nand ( n2394 , n2301 , n2393 );
nand ( n2395 , n1646 , n2394 );
nand ( n2396 , n2392 , n2395 );
not ( n2397 , n1839 );
nand ( n2398 , n344 , n2397 );
or ( n2399 , n2398 , n2328 );
not ( n2400 , n358 );
or ( n2401 , n2400 , n2266 );
nand ( n2402 , n2399 , n2401 );
or ( n2403 , n2396 , n2402 );
nand ( n2404 , n2403 , n2366 );
nand ( n2405 , n2384 , n2391 , n2404 );
not ( n2406 , n2405 );
nor ( n2407 , n1464 , n403 );
not ( n2408 , n2407 );
nor ( n2409 , n2408 , n2031 );
nand ( n2410 , n1644 , n2046 );
not ( n2411 , n2410 );
not ( n2412 , n2310 );
nand ( n2413 , n2354 , n2412 );
nand ( n2414 , n2411 , n2413 );
and ( n2415 , n1840 , n2294 );
and ( n2416 , n1890 , n2158 );
nor ( n2417 , n2416 , n1362 );
and ( n2418 , n2327 , n2417 );
nor ( n2419 , n2415 , n2418 );
and ( n2420 , n2414 , n2021 , n2419 );
not ( n2421 , n2317 );
or ( n2422 , n2421 , n2348 );
nand ( n2423 , n2422 , n1892 );
not ( n2424 , n2357 );
nand ( n2425 , n2301 , n2202 , n2424 );
not ( n2426 , n1919 );
or ( n2427 , n2425 , n2426 , n2417 );
nand ( n2428 , n1920 , n2362 );
or ( n2429 , n2428 , n2288 );
nand ( n2430 , n2427 , n2429 );
nand ( n2431 , n2420 , n2423 , n2430 );
nand ( n2432 , n2409 , n2431 );
and ( n2433 , n2277 , n2344 , n2406 , n2432 );
and ( n2434 , n2242 , n2433 );
nor ( n2435 , n389 , n391 );
nand ( n2436 , n1735 , n2435 );
nor ( n2437 , n2434 , n2436 );
and ( n2438 , n393 , n2437 );
nand ( n2439 , n1693 , n1727 );
and ( n2440 , n359 , n2439 );
not ( n2441 , n1040 );
not ( n2442 , n1682 );
or ( n2443 , n2441 , n2442 );
nor ( n2444 , n359 , n373 );
not ( n2445 , n1032 );
not ( n2446 , n2445 );
nand ( n2447 , n2444 , n2446 );
and ( n2448 , n1707 , n2447 );
nand ( n2449 , n1033 , n1429 );
nor ( n2450 , n2448 , n2449 );
or ( n2451 , n1624 , n2450 );
nand ( n2452 , n2443 , n2451 );
not ( n2453 , n2444 );
and ( n2454 , n2453 , n1693 );
nor ( n2455 , n2454 , n1716 );
nor ( n2456 , n2440 , n2452 , n2455 );
not ( n2457 , n358 );
nand ( n2458 , n1017 , n2457 );
nand ( n2459 , n2458 , n1314 );
and ( n2460 , n2453 , n2459 );
not ( n2461 , n2453 );
and ( n2462 , n2461 , n1387 );
nor ( n2463 , n2460 , n2462 );
and ( n2464 , n1013 , n1036 );
nor ( n2465 , n2464 , n358 );
nand ( n2466 , n1321 , n2465 , n1406 );
nand ( n2467 , n2466 , n2444 , n1355 );
nand ( n2468 , n1413 , n2447 );
nand ( n2469 , n2463 , n2467 , n2468 );
nand ( n2470 , n2469 , n1421 );
not ( n2471 , n2450 );
not ( n2472 , n1426 );
nand ( n2473 , n2471 , n2472 );
not ( n2474 , n1596 );
nor ( n2475 , n952 , n1483 );
nand ( n2476 , n2474 , n2475 );
and ( n2477 , n2476 , n1507 );
and ( n2478 , n1586 , n1575 );
nor ( n2479 , n2478 , n2453 );
and ( n2480 , n2477 , n2479 );
nor ( n2481 , n2444 , n1481 );
or ( n2482 , n1614 , n1744 );
nand ( n2483 , n2482 , n1586 );
and ( n2484 , n2481 , n1609 , n2483 );
nor ( n2485 , n2480 , n2484 );
nand ( n2486 , n2444 , n1582 );
and ( n2487 , n2468 , n2486 );
nor ( n2488 , n2487 , n1585 );
nor ( n2489 , n2485 , n2488 );
nand ( n2490 , n2470 , n2473 , n2489 );
not ( n2491 , n401 );
nand ( n2492 , n2490 , n2491 );
and ( n2493 , n2456 , n2492 );
and ( n2494 , n389 , n714 );
nor ( n2495 , n393 , n395 );
nand ( n2496 , n2494 , n2495 );
nor ( n2497 , n2493 , n2496 );
nor ( n2498 , n2438 , n2497 );
not ( n2499 , n2494 );
nor ( n2500 , n2499 , n1736 );
not ( n2501 , n2477 );
not ( n2502 , n1587 );
or ( n2503 , n2501 , n2502 );
nand ( n2504 , n2503 , n373 );
or ( n2505 , n1483 , n1600 );
and ( n2506 , n2505 , n1616 );
nor ( n2507 , n2506 , n373 );
and ( n2508 , n1030 , n1437 , n1608 );
nand ( n2509 , n373 , n1847 );
and ( n2510 , n2509 , n1707 );
nor ( n2511 , n2510 , n2449 );
or ( n2512 , n1426 , n2511 );
not ( n2513 , n1823 );
not ( n2514 , n2445 );
nand ( n2515 , n373 , n2514 );
nand ( n2516 , n1413 , n2515 );
or ( n2517 , n2513 , n2516 );
nand ( n2518 , n2512 , n2517 );
nor ( n2519 , n2507 , n2508 , n2518 );
and ( n2520 , n1030 , n1066 );
or ( n2521 , n1355 , n2520 );
nand ( n2522 , n2521 , n2466 );
nand ( n2523 , n1388 , n373 , n2522 );
not ( n2524 , n1313 );
or ( n2525 , n2520 , n1332 );
and ( n2526 , n358 , n2525 );
nor ( n2527 , n2526 , n373 );
nand ( n2528 , n2524 , n2527 , n2458 );
nand ( n2529 , n2523 , n1421 , n2528 );
and ( n2530 , n2504 , n2519 , n2529 );
or ( n2531 , n2530 , n401 );
and ( n2532 , n1019 , n2439 );
or ( n2533 , n1624 , n2511 );
not ( n2534 , n1656 );
nand ( n2535 , n373 , n2534 );
not ( n2536 , n1638 );
nor ( n2537 , n2536 , n1678 );
or ( n2538 , n2535 , n2537 );
nand ( n2539 , n2533 , n2538 );
and ( n2540 , n1657 , n1428 );
and ( n2541 , n1663 , n1712 );
nor ( n2542 , n2540 , n2541 );
and ( n2543 , n1714 , n2542 );
nor ( n2544 , n2543 , n1019 );
nor ( n2545 , n2532 , n2539 , n2544 );
nand ( n2546 , n2531 , n2545 );
and ( n2547 , n2500 , n2546 );
not ( n2548 , n1695 );
not ( n2549 , n2548 );
buf ( n2550 , n2549 );
not ( n2551 , n2550 );
not ( n2552 , n2551 );
and ( n2553 , n2273 , n1670 );
or ( n2554 , n2536 , n2553 );
nand ( n2555 , n2554 , n2500 );
or ( n2556 , n1019 , n2555 );
or ( n2557 , n1040 , n2496 );
nand ( n2558 , n1019 , n2500 );
nand ( n2559 , n2557 , n2558 );
nand ( n2560 , n2559 , n1697 );
nand ( n2561 , n2556 , n2560 );
and ( n2562 , n1634 , n2561 );
not ( n2563 , n2496 );
nand ( n2564 , n401 , n2563 );
nor ( n2565 , n359 , n2564 );
and ( n2566 , n1419 , n2565 );
and ( n2567 , n2566 , n1650 );
nor ( n2568 , n2562 , n2567 );
or ( n2569 , n2552 , n2568 );
not ( n2570 , n1626 );
nand ( n2571 , n2570 , n2500 );
or ( n2572 , n2571 , n2511 );
not ( n2573 , n2444 );
not ( n2574 , n2495 );
or ( n2575 , n2573 , n2574 );
nor ( n2576 , n1734 , n1736 );
nand ( n2577 , n373 , n2576 );
nand ( n2578 , n2575 , n2577 );
and ( n2579 , n2494 , n2578 );
and ( n2580 , n2579 , n1703 );
nor ( n2581 , n1821 , n2564 );
not ( n2582 , n2581 );
or ( n2583 , n2582 , n2450 );
not ( n2584 , n2558 );
or ( n2585 , n2444 , n2564 );
not ( n2586 , n2585 );
or ( n2587 , n2584 , n2586 );
nand ( n2588 , n2587 , n1699 );
nand ( n2589 , n2583 , n2588 );
nor ( n2590 , n2580 , n2589 );
nand ( n2591 , n2569 , n2572 , n2590 );
nor ( n2592 , n2547 , n2591 );
nand ( n2593 , n2435 , n2495 );
not ( n2594 , n2593 );
not ( n2595 , n1628 );
not ( n2596 , n329 );
and ( n2597 , n2596 , n1021 );
not ( n2598 , n2597 );
nor ( n2599 , n2598 , n1430 );
and ( n2600 , n329 , n1344 );
and ( n2601 , n2600 , n829 );
not ( n2602 , n2601 );
nand ( n2603 , n281 , n329 );
or ( n2604 , n2251 , n1251 );
nor ( n2605 , n2603 , n2604 );
and ( n2606 , n2605 , n1027 );
nand ( n2607 , n2606 , n1904 );
nand ( n2608 , n2602 , n2607 );
not ( n2609 , n2608 );
nor ( n2610 , n790 , n2597 );
nand ( n2611 , n1495 , n2610 );
not ( n2612 , n1020 );
and ( n2613 , n329 , n2612 );
not ( n2614 , n2613 );
nor ( n2615 , n2614 , n1029 );
nand ( n2616 , n2615 , n1007 );
nand ( n2617 , n2609 , n2611 , n2616 );
nor ( n2618 , n2599 , n2617 );
nand ( n2619 , n2596 , n1803 );
and ( n2620 , n2619 , n2117 );
and ( n2621 , n934 , n2613 );
nor ( n2622 , n2621 , n2610 );
nor ( n2623 , n2622 , n2250 );
nor ( n2624 , n2620 , n2623 );
and ( n2625 , n2618 , n2624 );
nor ( n2626 , n2625 , n358 );
and ( n2627 , n329 , n1260 );
and ( n2628 , n2111 , n2627 );
and ( n2629 , n1069 , n2627 );
not ( n2630 , n2629 );
nor ( n2631 , n2630 , n1305 );
nor ( n2632 , n2628 , n2631 );
nand ( n2633 , n1464 , n2632 );
or ( n2634 , n2626 , n2633 );
not ( n2635 , n358 );
and ( n2636 , n2635 , n2619 );
not ( n2637 , n2636 );
not ( n2638 , n2053 );
not ( n2639 , n2638 );
or ( n2640 , n2637 , n2639 );
not ( n2641 , n2627 );
or ( n2642 , n2084 , n2641 );
not ( n2643 , n358 );
nand ( n2644 , n2643 , n2606 );
not ( n2645 , n2644 );
and ( n2646 , n2645 , n2138 );
not ( n2647 , n2629 );
not ( n2648 , n1304 );
or ( n2649 , n2647 , n2648 );
and ( n2650 , n329 , n1800 );
not ( n2651 , n2650 );
or ( n2652 , n2651 , n828 );
nand ( n2653 , n2649 , n2652 );
nor ( n2654 , n2646 , n2653 );
nand ( n2655 , n2642 , n2654 );
not ( n2656 , n2655 );
nand ( n2657 , n2640 , n2656 );
or ( n2658 , n1464 , n2657 );
nand ( n2659 , n2634 , n2658 );
not ( n2660 , n1435 );
not ( n2661 , n2660 );
not ( n2662 , n951 );
not ( n2663 , n2662 );
nor ( n2664 , n2596 , n24 );
and ( n2665 , n64 , n2664 );
and ( n2666 , n2663 , n2665 );
and ( n2667 , n2666 , n1440 );
not ( n2668 , n2606 );
not ( n2669 , n1458 );
or ( n2670 , n2668 , n2669 );
nand ( n2671 , n2600 , n1122 );
nand ( n2672 , n2670 , n2671 );
nor ( n2673 , n2667 , n2672 );
not ( n2674 , n2673 );
and ( n2675 , n2661 , n2674 );
not ( n2676 , n2666 );
not ( n2677 , n1100 );
or ( n2678 , n2676 , n2677 );
and ( n2679 , n2606 , n1341 );
nor ( n2680 , n1876 , n2671 );
nor ( n2681 , n2679 , n2680 );
nand ( n2682 , n2678 , n2681 );
and ( n2683 , n1759 , n2682 );
nor ( n2684 , n2675 , n2683 );
not ( n2685 , n2100 );
not ( n2686 , n2610 );
nor ( n2687 , n2685 , n2686 );
or ( n2688 , n2687 , n2599 );
nand ( n2689 , n2688 , n2120 );
and ( n2690 , n265 , n311 );
and ( n2691 , n64 , n1359 );
and ( n2692 , n2690 , n2691 );
not ( n2693 , n2603 );
and ( n2694 , n2692 , n2693 );
and ( n2695 , n2694 , n1579 );
nand ( n2696 , n1010 , n1763 );
nor ( n2697 , n2614 , n2696 );
not ( n2698 , n2697 );
not ( n2699 , n1470 );
nor ( n2700 , n2698 , n2699 );
nor ( n2701 , n2695 , n2700 );
not ( n2702 , n2701 );
nand ( n2703 , n2702 , n372 );
and ( n2704 , n2684 , n2689 , n2703 );
not ( n2705 , n2177 );
not ( n2706 , n1593 );
or ( n2707 , n2705 , n2706 );
nand ( n2708 , n2707 , n2123 );
nand ( n2709 , n329 , n2708 );
nand ( n2710 , n2659 , n2704 , n2709 );
not ( n2711 , n2710 );
not ( n2712 , n2711 );
and ( n2713 , n2595 , n2712 );
not ( n2714 , n1260 );
not ( n2715 , n1751 );
not ( n2716 , n2715 );
or ( n2717 , n2714 , n2716 );
or ( n2718 , n835 , n1794 );
not ( n2719 , n358 );
nand ( n2720 , n2718 , n2719 );
nand ( n2721 , n2717 , n2720 );
nand ( n2722 , n1312 , n1131 );
or ( n2723 , n2721 , n2722 );
nand ( n2724 , n2723 , n2596 );
not ( n2725 , n2663 );
buf ( n2726 , n2725 );
not ( n2727 , n2726 );
nand ( n2728 , n2596 , n2727 );
not ( n2729 , n945 );
or ( n2730 , n2728 , n2729 );
or ( n2731 , n311 , n2622 );
nand ( n2732 , n2730 , n2731 );
nand ( n2733 , n1741 , n2732 );
not ( n2734 , n2632 );
nand ( n2735 , n2615 , n2122 );
not ( n2736 , n2682 );
and ( n2737 , n2686 , n2735 , n2736 );
not ( n2738 , n358 );
nor ( n2739 , n2737 , n2738 );
nor ( n2740 , n2734 , n2739 );
nand ( n2741 , n2724 , n2733 , n2740 );
nand ( n2742 , n2741 , n1421 );
nand ( n2743 , n2472 , n2710 );
nand ( n2744 , n2596 , n1753 );
and ( n2745 , n1817 , n1600 );
not ( n2746 , n358 );
nand ( n2747 , n2596 , n2746 );
nor ( n2748 , n2745 , n2747 );
nor ( n2749 , n2700 , n2655 );
nand ( n2750 , n2636 , n2687 );
not ( n2751 , n358 );
and ( n2752 , n329 , n2751 );
nand ( n2753 , n2752 , n2054 );
nand ( n2754 , n2749 , n2750 , n2753 );
nor ( n2755 , n2748 , n2754 );
and ( n2756 , n2744 , n2755 );
nor ( n2757 , n2756 , n1585 );
not ( n2758 , n2690 );
nor ( n2759 , n2758 , n2603 );
not ( n2760 , n2759 );
not ( n2761 , n1579 );
or ( n2762 , n2760 , n2761 );
not ( n2763 , n281 );
nor ( n2764 , n2763 , n329 );
nand ( n2765 , n2764 , n2690 , n1608 );
nand ( n2766 , n2762 , n2765 );
and ( n2767 , n948 , n2766 );
nor ( n2768 , n329 , n1217 );
and ( n2769 , n2768 , n1570 );
nor ( n2770 , n2767 , n2769 );
not ( n2771 , n2687 );
and ( n2772 , n2770 , n2771 , n2673 );
nor ( n2773 , n2772 , n1436 );
and ( n2774 , n329 , n2117 );
nor ( n2775 , n2774 , n2617 );
or ( n2776 , n2775 , n2120 , n1822 );
not ( n2777 , n358 );
nor ( n2778 , n2777 , n329 );
nand ( n2779 , n1461 , n2778 , n1586 );
nand ( n2780 , n2776 , n2779 );
nor ( n2781 , n2757 , n2773 , n2780 );
and ( n2782 , n2742 , n2743 , n2781 );
nor ( n2783 , n2782 , n401 );
nor ( n2784 , n2713 , n2783 );
nand ( n2785 , n2694 , n2122 );
nand ( n2786 , n24 , n329 );
or ( n2787 , n2786 , n2110 );
nand ( n2788 , n2787 , n2681 );
and ( n2789 , n358 , n2788 );
not ( n2790 , n358 );
and ( n2791 , n2790 , n2608 );
nor ( n2792 , n2789 , n2791 );
not ( n2793 , n311 );
and ( n2794 , n2793 , n2613 );
nand ( n2795 , n2691 , n2794 );
not ( n2796 , n2795 );
not ( n2797 , n1099 );
and ( n2798 , n2796 , n2797 );
not ( n2799 , n358 );
nand ( n2800 , n2666 , n934 );
not ( n2801 , n1247 );
nand ( n2802 , n1138 , n1182 );
not ( n2803 , n2802 );
or ( n2804 , n2801 , n2803 );
nand ( n2805 , n2804 , n329 );
nand ( n2806 , n2800 , n2616 , n2805 );
and ( n2807 , n2799 , n2806 );
nor ( n2808 , n2798 , n2807 );
nand ( n2809 , n2785 , n2792 , n2808 );
nand ( n2810 , n2596 , n1428 );
or ( n2811 , n1491 , n2810 );
nand ( n2812 , n2811 , n790 );
and ( n2813 , n2812 , n1725 );
nor ( n2814 , n2614 , n1945 );
not ( n2815 , n2814 );
not ( n2816 , n1214 );
or ( n2817 , n2815 , n2816 );
not ( n2818 , n2631 );
nand ( n2819 , n2817 , n2818 );
or ( n2820 , n2809 , n2813 , n2819 );
nand ( n2821 , n2820 , n2032 );
or ( n2822 , n1775 , n2021 );
nand ( n2823 , n311 , n1775 );
not ( n2824 , n2823 );
and ( n2825 , n265 , n2812 );
nand ( n2826 , n1686 , n2810 );
and ( n2827 , n2824 , n2825 , n2826 );
nor ( n2828 , n2827 , n2680 );
nand ( n2829 , n2822 , n2828 , n2735 );
and ( n2830 , n358 , n2829 );
and ( n2831 , n1538 , n2826 );
nor ( n2832 , n2830 , n2831 );
or ( n2833 , n372 , n2832 );
not ( n2834 , n1293 );
and ( n2835 , n2627 , n2834 );
and ( n2836 , n1359 , n1252 );
nand ( n2837 , n2613 , n2836 );
or ( n2838 , n2837 , n1110 );
or ( n2839 , n358 , n2607 );
nand ( n2840 , n2838 , n2839 );
nor ( n2841 , n2835 , n2840 );
not ( n2842 , n2841 );
nand ( n2843 , n2690 , n948 );
nand ( n2844 , n2604 , n1775 , n2843 );
and ( n2845 , n2826 , n2844 , n2812 );
nor ( n2846 , n2845 , n2601 );
or ( n2847 , n358 , n2846 );
nand ( n2848 , n2847 , n1464 );
not ( n2849 , n1775 );
not ( n2850 , n2690 );
not ( n2851 , n1686 );
and ( n2852 , n2850 , n2851 );
nor ( n2853 , n2726 , n2810 );
nor ( n2854 , n2852 , n2853 );
nor ( n2855 , n2849 , n2854 );
nor ( n2856 , n2842 , n2848 , n2855 , n2819 );
nor ( n2857 , n2596 , n1547 );
not ( n2858 , n1285 );
nand ( n2859 , n2857 , n2858 );
and ( n2860 , n2859 , n2808 );
nand ( n2861 , n2833 , n2856 , n2860 );
nor ( n2862 , n948 , n2068 );
or ( n2863 , n281 , n1244 );
nand ( n2864 , n2863 , n265 );
and ( n2865 , n2862 , n2864 );
nor ( n2866 , n2865 , n2645 );
or ( n2867 , n1686 , n2866 );
not ( n2868 , n1244 );
and ( n2869 , n2868 , n2862 );
not ( n2870 , n358 );
nor ( n2871 , n2870 , n311 );
nor ( n2872 , n2869 , n2871 );
and ( n2873 , n2872 , n2250 , n2825 );
and ( n2874 , n1252 , n2597 );
not ( n2875 , n2874 );
nor ( n2876 , n1764 , n2875 );
nor ( n2877 , n2873 , n2876 );
nor ( n2878 , n1218 , n1961 );
nand ( n2879 , n2867 , n2877 , n2878 );
and ( n2880 , n2826 , n2879 );
nor ( n2881 , n2862 , n2854 );
not ( n2882 , n1515 );
not ( n2883 , n2051 );
or ( n2884 , n2882 , n2883 );
nand ( n2885 , n2884 , n2752 );
and ( n2886 , n1960 , n2759 );
and ( n2887 , n2886 , n1521 );
not ( n2888 , n2795 );
and ( n2889 , n2888 , n1440 );
nor ( n2890 , n2887 , n2889 );
nand ( n2891 , n2627 , n2083 );
nand ( n2892 , n2885 , n2890 , n2891 , n2701 );
nor ( n2893 , n2880 , n2881 , n2892 );
nor ( n2894 , n2596 , n2072 );
and ( n2895 , n2894 , n1122 );
not ( n2896 , n2837 );
and ( n2897 , n2896 , n1458 );
not ( n2898 , n2752 );
or ( n2899 , n2898 , n1512 );
nand ( n2900 , n2899 , n2654 );
nor ( n2901 , n2895 , n2897 , n2900 );
and ( n2902 , n2893 , n372 , n2901 );
nor ( n2903 , n2902 , n1662 );
and ( n2904 , n2861 , n2903 );
not ( n2905 , n2892 );
not ( n2906 , n1029 );
or ( n2907 , n2251 , n2764 , n1720 );
nor ( n2908 , n329 , n1698 );
nand ( n2909 , n1427 , n2908 );
nand ( n2910 , n2907 , n2909 );
and ( n2911 , n2906 , n2910 );
and ( n2912 , n1832 , n2909 );
nor ( n2913 , n2912 , n1775 );
not ( n2914 , n1776 );
not ( n2915 , n2914 );
not ( n2916 , n2915 );
not ( n2917 , n2908 );
and ( n2918 , n1832 , n2917 );
or ( n2919 , n2918 , n2726 );
nand ( n2920 , n2919 , n2257 );
and ( n2921 , n2916 , n2920 );
and ( n2922 , n1252 , n2910 );
nor ( n2923 , n2921 , n2922 );
not ( n2924 , n2923 );
nor ( n2925 , n2911 , n2913 , n2924 );
not ( n2926 , n1777 );
nand ( n2927 , n2926 , n2920 );
nand ( n2928 , n2905 , n2925 , n2927 , n2901 );
and ( n2929 , n2366 , n2928 );
nor ( n2930 , n2904 , n2929 );
nand ( n2931 , n1763 , n1068 , n2253 , n1697 );
not ( n2932 , n2931 );
not ( n2933 , n1360 );
not ( n2934 , n358 );
nand ( n2935 , n2934 , n1137 );
not ( n2936 , n358 );
not ( n2937 , n2069 );
nor ( n2938 , n64 , n2937 );
nand ( n2939 , n2936 , n2938 );
and ( n2940 , n2935 , n2939 );
and ( n2941 , n2265 , n2933 , n2940 );
not ( n2942 , n2910 );
nor ( n2943 , n2941 , n2942 );
or ( n2944 , n1924 , n2918 );
not ( n2945 , n1807 );
or ( n2946 , n2945 , n2810 );
not ( n2947 , n2596 );
not ( n2948 , n2062 );
and ( n2949 , n2947 , n2948 );
and ( n2950 , n2894 , n2074 );
nor ( n2951 , n2949 , n2950 );
nand ( n2952 , n2944 , n2946 , n2951 );
nor ( n2953 , n2932 , n2943 , n2952 , n2913 );
nand ( n2954 , n2923 , n2735 );
and ( n2955 , n358 , n2954 );
or ( n2956 , n1763 , n2927 );
nand ( n2957 , n2956 , n2841 );
nor ( n2958 , n2955 , n2957 , n2819 );
nand ( n2959 , n2860 , n2953 , n2958 );
and ( n2960 , n2276 , n2959 );
not ( n2961 , n358 );
not ( n2962 , n2672 );
or ( n2963 , n2961 , n2962 );
nor ( n2964 , n2813 , n2900 );
nand ( n2965 , n2963 , n2964 , n2905 );
and ( n2966 , n2339 , n2965 );
nor ( n2967 , n2960 , n2966 );
nand ( n2968 , n2784 , n2821 , n2930 , n2967 );
nand ( n2969 , n2594 , n2968 );
and ( n2970 , n2498 , n2592 , n2969 );
nand ( n2971 , n391 , n1734 );
nand ( n2972 , n714 , n1735 );
nand ( n2973 , n2971 , n2972 , n1835 );
nand ( n2974 , n1838 , n2970 , n2973 );
not ( n2975 , n397 );
not ( n2976 , n405 );
nand ( n2977 , n2975 , n2976 );
not ( n2978 , n387 );
nor ( n2979 , n385 , n400 );
and ( n2980 , n2978 , n2979 );
nor ( n2981 , n2977 , n2980 );
nand ( n2982 , n2974 , n2981 );
not ( n2983 , n401 );
and ( n2984 , n1423 , n2983 );
not ( n2985 , n2984 );
not ( n2986 , n2977 );
and ( n2987 , n2986 , n2436 );
and ( n2988 , n2980 , n2987 );
nand ( n2989 , n2985 , n2988 );
not ( n2990 , n2989 );
not ( n2991 , n1430 );
and ( n2992 , n2990 , n2991 );
and ( n2993 , n388 , n2977 );
nor ( n2994 , n2992 , n2993 );
nor ( n2995 , n2977 , n2593 );
nand ( n2996 , n2980 , n2995 );
not ( n2997 , n2996 );
not ( n2998 , n2783 );
not ( n2999 , n2998 );
and ( n3000 , n2997 , n2999 );
nand ( n3001 , n393 , n2986 );
nor ( n3002 , n395 , n3001 );
nand ( n3003 , n2435 , n3002 );
not ( n3004 , n3003 );
nand ( n3005 , n2980 , n3004 );
or ( n3006 , n3005 , n2240 );
nor ( n3007 , n2984 , n3005 );
not ( n3008 , n2342 );
and ( n3009 , n3007 , n3008 );
nor ( n3010 , n2984 , n2996 );
and ( n3011 , n3010 , n2710 );
nor ( n3012 , n3009 , n3011 );
not ( n3013 , n1828 );
nand ( n3014 , n2988 , n3013 );
nand ( n3015 , n3006 , n3012 , n3014 );
nor ( n3016 , n3000 , n3015 );
nand ( n3017 , n2982 , n2994 , n3016 );
not ( n3018 , n389 );
not ( n3019 , n1070 );
not ( n3020 , n399 );
nor ( n3021 , n3020 , n402 );
not ( n3022 , n3021 );
not ( n3023 , n3022 );
not ( n3024 , n3023 );
not ( n3025 , n963 );
and ( n3026 , n3024 , n3025 );
not ( n3027 , n3026 );
nand ( n3028 , n746 , n912 );
nor ( n3029 , n407 , n417 );
nor ( n3030 , n402 , n3029 );
nand ( n3031 , n3028 , n3030 );
not ( n3032 , n3031 );
not ( n3033 , n3032 );
buf ( n3034 , n962 );
not ( n3035 , n3034 );
or ( n3036 , n3033 , n3035 );
not ( n3037 , n410 );
nand ( n3038 , n3037 , n412 );
not ( n3039 , n3038 );
not ( n3040 , n3039 );
nand ( n3041 , n3040 , n776 );
nand ( n3042 , n3041 , n857 );
nand ( n3043 , n3042 , n746 );
not ( n3044 , n417 );
nor ( n3045 , n3044 , n407 );
and ( n3046 , n730 , n3045 );
nor ( n3047 , n3043 , n3046 );
not ( n3048 , n402 );
nand ( n3049 , n3047 , n3048 );
nand ( n3050 , n3036 , n3049 );
not ( n3051 , n3050 );
nor ( n3052 , n3046 , n3043 );
not ( n3053 , n3052 );
nand ( n3054 , n892 , n3053 );
not ( n3055 , n961 );
not ( n3056 , n3055 );
not ( n3057 , n3056 );
nor ( n3058 , n3054 , n3057 );
nor ( n3059 , n3051 , n3058 );
nand ( n3060 , n399 , n3059 );
not ( n3061 , n3043 );
nand ( n3062 , n3022 , n3061 );
not ( n3063 , n3062 );
not ( n3064 , n3063 );
nand ( n3065 , n3027 , n3060 , n3064 );
not ( n3066 , n879 );
not ( n3067 , n3066 );
not ( n3068 , n3067 );
buf ( n3069 , n3068 );
not ( n3070 , n3069 );
or ( n3071 , n3065 , n3070 );
nor ( n3072 , n791 , n388 );
not ( n3073 , n3072 );
not ( n3074 , n3073 );
not ( n3075 , n3074 );
not ( n3076 , n3075 );
not ( n3077 , n3076 );
buf ( n3078 , n3077 );
nand ( n3079 , n3071 , n3078 );
not ( n3080 , n3079 );
or ( n3081 , n3019 , n3080 );
not ( n3082 , n811 );
and ( n3083 , n892 , n3082 );
nand ( n3084 , n3057 , n3083 );
not ( n3085 , n3084 );
nor ( n3086 , n402 , n3045 );
and ( n3087 , n1093 , n3086 );
not ( n3088 , n3087 );
not ( n3089 , n859 );
not ( n3090 , n3089 );
not ( n3091 , n3090 );
or ( n3092 , n3088 , n3091 );
not ( n3093 , n985 );
not ( n3094 , n3041 );
not ( n3095 , n3045 );
not ( n3096 , n3095 );
nor ( n3097 , n3094 , n3096 );
not ( n3098 , n3042 );
nor ( n3099 , n3097 , n3098 );
nand ( n3100 , n3093 , n3099 );
nand ( n3101 , n3092 , n3100 );
not ( n3102 , n3099 );
nand ( n3103 , n3102 , n892 );
nand ( n3104 , n3101 , n3103 );
not ( n3105 , n3104 );
or ( n3106 , n3085 , n3105 );
nand ( n3107 , n3106 , n399 );
buf ( n3108 , n869 );
nand ( n3109 , n3107 , n3108 );
nand ( n3110 , n3068 , n3064 );
or ( n3111 , n3109 , n3110 );
nand ( n3112 , n3111 , n3078 );
nand ( n3113 , n1104 , n3112 );
nand ( n3114 , n3081 , n3113 );
nand ( n3115 , n3114 , n358 , n2664 );
not ( n3116 , n2886 );
not ( n3117 , n3061 );
not ( n3118 , n3117 );
not ( n3119 , n857 );
not ( n3120 , n866 );
nand ( n3121 , n956 , n3120 );
nand ( n3122 , n3119 , n3121 );
not ( n3123 , n3122 );
nand ( n3124 , n3123 , n407 );
nand ( n3125 , n3124 , n1145 );
not ( n3126 , n3125 );
not ( n3127 , n3126 );
or ( n3128 , n3118 , n3127 );
nor ( n3129 , n399 , n402 );
not ( n3130 , n3129 );
nand ( n3131 , n3128 , n3130 );
buf ( n3132 , n3131 );
nand ( n3133 , n413 , n902 );
not ( n3134 , n3133 );
not ( n3135 , n3122 );
not ( n3136 , n3135 );
not ( n3137 , n3136 );
not ( n3138 , n3137 );
not ( n3139 , n3138 );
nand ( n3140 , n3134 , n3139 );
not ( n3141 , n3140 );
nor ( n3142 , n3052 , n892 );
not ( n3143 , n3142 );
not ( n3144 , n3032 );
not ( n3145 , n3135 );
not ( n3146 , n960 );
not ( n3147 , n3146 );
nand ( n3148 , n3145 , n3147 );
not ( n3149 , n3148 );
or ( n3150 , n3144 , n3149 );
nand ( n3151 , n3150 , n3049 );
and ( n3152 , n3143 , n3151 );
not ( n3153 , n3125 );
nor ( n3154 , n3153 , n402 );
nor ( n3155 , n3152 , n3154 );
not ( n3156 , n3155 );
or ( n3157 , n3141 , n3156 );
not ( n3158 , n399 );
nand ( n3159 , n3157 , n3158 );
nand ( n3160 , n3132 , n3159 );
or ( n3161 , n3160 , n3070 );
nand ( n3162 , n3161 , n3078 );
not ( n3163 , n3162 );
or ( n3164 , n3116 , n3163 );
nor ( n3165 , n2596 , n1742 );
not ( n3166 , n3070 );
not ( n3167 , n3166 );
not ( n3168 , n402 );
not ( n3169 , n3168 );
buf ( n3170 , n3124 );
nand ( n3171 , n3170 , n869 );
not ( n3172 , n3171 );
or ( n3173 , n3169 , n3172 );
not ( n3174 , n3087 );
not ( n3175 , n410 );
nand ( n3176 , n1003 , n3175 );
nand ( n3177 , n3176 , n3119 );
not ( n3178 , n3177 );
not ( n3179 , n3178 );
or ( n3180 , n3174 , n3179 );
nand ( n3181 , n3180 , n3100 );
and ( n3182 , n3103 , n3181 );
not ( n3183 , n3083 );
nor ( n3184 , n3183 , n3136 );
nor ( n3185 , n3182 , n3184 );
nand ( n3186 , n3173 , n3185 );
and ( n3187 , n399 , n3186 );
or ( n3188 , n3063 , n3171 );
nor ( n3189 , n3187 , n3188 );
not ( n3190 , n3189 );
or ( n3191 , n3167 , n3190 );
nand ( n3192 , n3191 , n3078 );
nand ( n3193 , n3165 , n3192 );
nand ( n3194 , n3164 , n3193 );
and ( n3195 , n1960 , n2794 );
not ( n3196 , n3195 );
not ( n3197 , n3069 );
not ( n3198 , n399 );
nand ( n3199 , n413 , n3102 );
not ( n3200 , n3199 );
not ( n3201 , n3181 );
or ( n3202 , n3200 , n3201 );
not ( n3203 , n3030 );
nand ( n3204 , n413 , n3082 );
nand ( n3205 , n3203 , n3204 );
nand ( n3206 , n3205 , n3137 );
nand ( n3207 , n3202 , n3206 );
and ( n3208 , n3198 , n3207 );
nand ( n3209 , n3170 , n1220 );
nand ( n3210 , n3209 , n3130 );
nand ( n3211 , n3117 , n1220 );
nand ( n3212 , n3130 , n3211 );
nand ( n3213 , n3210 , n3212 );
nor ( n3214 , n3208 , n3213 );
not ( n3215 , n3214 );
or ( n3216 , n3197 , n3215 );
buf ( n3217 , n3077 );
nand ( n3218 , n3216 , n3217 );
not ( n3219 , n3218 );
or ( n3220 , n3196 , n3219 );
not ( n3221 , n3054 );
not ( n3222 , n3151 );
or ( n3223 , n3221 , n3222 );
not ( n3224 , n867 );
not ( n3225 , n402 );
nand ( n3226 , n3224 , n3225 );
and ( n3227 , n3226 , n3206 );
nand ( n3228 , n3223 , n3227 );
nand ( n3229 , n3228 , n399 );
not ( n3230 , n3023 );
nand ( n3231 , n3170 , n963 );
and ( n3232 , n3230 , n3231 );
nor ( n3233 , n3232 , n3063 );
nand ( n3234 , n3229 , n3233 , n3069 );
nand ( n3235 , n3234 , n3217 );
nand ( n3236 , n2613 , n3235 );
or ( n3237 , n2696 , n3236 );
nand ( n3238 , n3220 , n3237 );
nor ( n3239 , n3194 , n3238 );
and ( n3240 , n3115 , n3239 );
not ( n3241 , n951 );
nand ( n3242 , n388 , n392 );
not ( n3243 , n3242 );
and ( n3244 , n3243 , n1685 );
not ( n3245 , n3244 );
nand ( n3246 , n1668 , n1648 );
not ( n3247 , n3119 );
and ( n3248 , n878 , n3041 );
nand ( n3249 , n3247 , n3248 );
and ( n3250 , n791 , n3249 );
nor ( n3251 , n329 , n3250 );
nand ( n3252 , n3246 , n3251 );
nand ( n3253 , n3245 , n3252 );
not ( n3254 , n3253 );
or ( n3255 , n3241 , n3254 );
not ( n3256 , n311 );
nand ( n3257 , n392 , n2251 );
not ( n3258 , n3257 );
or ( n3259 , n3256 , n3258 );
not ( n3260 , n392 );
nand ( n3261 , n3260 , n388 );
or ( n3262 , n390 , n410 );
nand ( n3263 , n3262 , n791 );
nand ( n3264 , n2763 , n3261 , n3263 );
nor ( n3265 , n2251 , n3264 );
not ( n3266 , n3265 );
nand ( n3267 , n3257 , n3266 );
nand ( n3268 , n3246 , n3267 );
not ( n3269 , n3268 );
nand ( n3270 , n3259 , n3269 );
nand ( n3271 , n3255 , n3270 );
and ( n3272 , n1135 , n3271 );
not ( n3273 , n1025 );
not ( n3274 , n3253 );
or ( n3275 , n3273 , n3274 );
nand ( n3276 , n3275 , n3268 );
not ( n3277 , n3276 );
nor ( n3278 , n1775 , n3277 );
nor ( n3279 , n3272 , n358 , n3278 );
not ( n3280 , n3279 );
not ( n3281 , n2786 );
buf ( n3282 , n3077 );
nand ( n3283 , n3057 , n3205 );
not ( n3284 , n3283 );
nand ( n3285 , n3199 , n3101 );
not ( n3286 , n3285 );
or ( n3287 , n3284 , n3286 );
not ( n3288 , n399 );
nand ( n3289 , n3287 , n3288 );
nand ( n3290 , n3289 , n3212 , n3069 );
nand ( n3291 , n3282 , n3290 );
nand ( n3292 , n1291 , n3291 );
not ( n3293 , n3292 );
and ( n3294 , n3281 , n3293 );
not ( n3295 , n2606 );
not ( n3296 , n3039 );
and ( n3297 , n402 , n731 );
nand ( n3298 , n3296 , n3297 );
nand ( n3299 , n3066 , n3298 );
not ( n3300 , n3299 );
not ( n3301 , n3300 );
not ( n3302 , n3301 );
not ( n3303 , n778 );
not ( n3304 , n3303 );
nand ( n3305 , n3302 , n3304 , n3051 );
not ( n3306 , n3073 );
not ( n3307 , n3306 );
nand ( n3308 , n3248 , n3049 );
not ( n3309 , n3308 );
not ( n3310 , n3034 );
buf ( n3311 , n3310 );
nand ( n3312 , n3309 , n3311 );
nand ( n3313 , n3305 , n3307 , n3312 );
not ( n3314 , n3247 );
nand ( n3315 , n1300 , n3314 );
and ( n3316 , n3313 , n3315 );
not ( n3317 , n1115 );
not ( n3318 , n3249 );
nand ( n3319 , n3317 , n3318 );
not ( n3320 , n3319 );
not ( n3321 , n3320 );
not ( n3322 , n3051 );
or ( n3323 , n3321 , n3322 );
nand ( n3324 , n3323 , n3307 );
nor ( n3325 , n3316 , n3324 );
or ( n3326 , n3295 , n3325 );
not ( n3327 , n3101 );
buf ( n3328 , n3090 );
not ( n3329 , n3328 );
not ( n3330 , n3301 );
nand ( n3331 , n3327 , n3329 , n3330 );
not ( n3332 , n3315 );
or ( n3333 , n3331 , n3332 );
and ( n3334 , n3073 , n3319 );
nand ( n3335 , n3333 , n3334 );
nand ( n3336 , n2600 , n3335 );
nand ( n3337 , n3326 , n3336 );
not ( n3338 , n3337 );
nand ( n3339 , n1251 , n2250 );
nor ( n3340 , n3277 , n2251 );
and ( n3341 , n3339 , n3340 );
not ( n3342 , n358 );
nor ( n3343 , n3341 , n3342 );
nand ( n3344 , n1218 , n3253 );
not ( n3345 , n311 );
nand ( n3346 , n3345 , n3257 );
and ( n3347 , n3346 , n3276 );
and ( n3348 , n3347 , n948 );
not ( n3349 , n2662 );
not ( n3350 , n3252 );
and ( n3351 , n3349 , n3350 );
and ( n3352 , n2794 , n3244 );
nor ( n3353 , n3351 , n3352 );
and ( n3354 , n3270 , n3353 );
nor ( n3355 , n3354 , n1776 );
nor ( n3356 , n3348 , n3355 );
nand ( n3357 , n3338 , n3343 , n3344 , n3356 );
nor ( n3358 , n3294 , n3357 );
not ( n3359 , n3358 );
and ( n3360 , n3280 , n3359 );
not ( n3361 , n3069 );
not ( n3362 , n3061 );
and ( n3363 , n3362 , n3310 );
or ( n3364 , n3131 , n3363 );
not ( n3365 , n3056 );
not ( n3366 , n3142 );
or ( n3367 , n3365 , n3366 );
nand ( n3368 , n3367 , n3050 );
or ( n3369 , n3368 , n399 );
nand ( n3370 , n3364 , n3369 );
not ( n3371 , n3370 );
not ( n3372 , n3371 );
or ( n3373 , n3361 , n3372 );
nand ( n3374 , n3373 , n3282 );
nand ( n3375 , n3374 , n1806 );
not ( n3376 , n3375 );
and ( n3377 , n2627 , n3376 );
not ( n3378 , n2696 );
not ( n3379 , n2940 );
or ( n3380 , n3378 , n3379 );
nand ( n3381 , n3380 , n3340 );
and ( n3382 , n1807 , n3350 );
not ( n3383 , n3346 );
nor ( n3384 , n64 , n1764 );
not ( n3385 , n3384 );
or ( n3386 , n3383 , n3385 );
not ( n3387 , n358 );
nor ( n3388 , n3387 , n1775 );
not ( n3389 , n3388 );
nand ( n3390 , n3386 , n3389 );
and ( n3391 , n3390 , n3269 );
nor ( n3392 , n3382 , n3391 );
nor ( n3393 , n2068 , n1763 );
nand ( n3394 , n1776 , n3271 );
or ( n3395 , n3393 , n3394 );
not ( n3396 , n3315 );
and ( n3397 , n3300 , n3177 );
nand ( n3398 , n3397 , n3100 );
not ( n3399 , n3398 );
not ( n3400 , n3399 );
or ( n3401 , n3396 , n3400 );
nand ( n3402 , n3401 , n3334 );
nand ( n3403 , n2650 , n3402 );
nand ( n3404 , n2645 , n3244 );
nand ( n3405 , n3395 , n3403 , n3404 );
not ( n3406 , n3405 );
nand ( n3407 , n3381 , n3392 , n3406 );
nor ( n3408 , n3377 , n3407 );
nor ( n3409 , n3067 , n3061 );
nand ( n3410 , n867 , n3409 );
nand ( n3411 , n3075 , n3410 );
not ( n3412 , n3411 );
or ( n3413 , n2630 , n3412 );
and ( n3414 , n3170 , n3409 );
nor ( n3415 , n3414 , n3074 );
or ( n3416 , n1217 , n3415 );
not ( n3417 , n3416 );
nand ( n3418 , n3417 , n2752 );
nand ( n3419 , n3413 , n3418 );
not ( n3420 , n3419 );
not ( n3421 , n3308 );
not ( n3422 , n3148 );
and ( n3423 , n3421 , n3422 );
nor ( n3424 , n3423 , n3306 );
or ( n3425 , n3424 , n3332 );
not ( n3426 , n3151 );
not ( n3427 , n3319 );
and ( n3428 , n3426 , n3427 );
nor ( n3429 , n3428 , n3076 );
nand ( n3430 , n3425 , n3429 );
nand ( n3431 , n2645 , n3430 );
nand ( n3432 , n3408 , n3420 , n3431 );
nor ( n3433 , n3360 , n3432 );
and ( n3434 , n3240 , n3433 );
nor ( n3435 , n3434 , n2408 );
and ( n3436 , n3292 , n3375 );
not ( n3437 , n3436 );
nand ( n3438 , n2627 , n3437 );
nand ( n3439 , n3337 , n358 );
not ( n3440 , n3439 );
nand ( n3441 , n392 , n1689 );
not ( n3442 , n3072 );
and ( n3443 , n3442 , n3249 );
not ( n3444 , n3443 );
nand ( n3445 , n3444 , n2596 );
and ( n3446 , n3441 , n3445 );
or ( n3447 , n1631 , n3446 );
nand ( n3448 , n44 , n1842 );
not ( n3449 , n3267 );
not ( n3450 , n3449 );
nand ( n3451 , n3448 , n3450 );
nand ( n3452 , n3447 , n3451 );
and ( n3453 , n3403 , n3431 );
not ( n3454 , n3453 );
nor ( n3455 , n3440 , n3452 , n3419 , n3454 );
and ( n3456 , n3240 , n3438 , n3455 );
nor ( n3457 , n3456 , n2338 );
nor ( n3458 , n3435 , n3457 );
not ( n3459 , n3109 );
nand ( n3460 , n413 , n909 );
and ( n3461 , n779 , n3460 );
and ( n3462 , n3461 , n3068 , n3062 );
nand ( n3463 , n892 , n909 );
not ( n3464 , n3463 );
nand ( n3465 , n3055 , n3464 );
and ( n3466 , n3462 , n3465 , n3298 );
not ( n3467 , n3466 );
not ( n3468 , n399 );
nand ( n3469 , n3468 , n3461 );
not ( n3470 , n3469 );
not ( n3471 , n3460 );
nor ( n3472 , n3471 , n868 );
nor ( n3473 , n3472 , n3089 );
not ( n3474 , n3473 );
or ( n3475 , n3470 , n3474 );
and ( n3476 , n3465 , n3300 );
nand ( n3477 , n3475 , n3476 );
not ( n3478 , n3477 );
nand ( n3479 , n3064 , n3478 );
nand ( n3480 , n3467 , n3479 );
and ( n3481 , n3459 , n3480 );
not ( n3482 , n399 );
nand ( n3483 , n3482 , n3476 );
not ( n3484 , n3461 );
nand ( n3485 , n3484 , n3473 );
not ( n3486 , n3485 );
nor ( n3487 , n3483 , n3486 );
nor ( n3488 , n3487 , n3104 );
not ( n3489 , n402 );
or ( n3490 , n3488 , n3477 , n3489 );
nand ( n3491 , n3490 , n3077 );
nor ( n3492 , n3481 , n3491 );
not ( n3493 , n3492 );
not ( n3494 , n3493 );
or ( n3495 , n2795 , n3494 );
not ( n3496 , n3306 );
nand ( n3497 , n3496 , n3398 );
and ( n3498 , n2650 , n3497 );
not ( n3499 , n3057 );
and ( n3500 , n402 , n3248 );
nand ( n3501 , n3499 , n3500 );
nand ( n3502 , n3501 , n3412 );
and ( n3503 , n2629 , n3502 );
nor ( n3504 , n3498 , n3503 );
not ( n3505 , n3228 );
not ( n3506 , n3463 );
not ( n3507 , n3506 );
not ( n3508 , n3135 );
or ( n3509 , n3507 , n3508 );
nand ( n3510 , n3509 , n3300 );
or ( n3511 , n3471 , n3510 );
not ( n3512 , n3511 );
nor ( n3513 , n3301 , n3148 );
not ( n3514 , n3513 );
not ( n3515 , n3514 );
or ( n3516 , n3512 , n3515 );
nand ( n3517 , n3516 , n3233 );
nor ( n3518 , n3130 , n3117 );
not ( n3519 , n3518 );
not ( n3520 , n3514 );
and ( n3521 , n3519 , n3520 );
and ( n3522 , n779 , n3463 );
or ( n3523 , n3522 , n3510 );
nor ( n3524 , n3523 , n3231 );
nor ( n3525 , n3521 , n3524 );
nand ( n3526 , n3230 , n3231 );
not ( n3527 , n3462 );
nor ( n3528 , n3527 , n3510 );
and ( n3529 , n3526 , n3528 );
not ( n3530 , n3463 );
not ( n3531 , n3530 );
nor ( n3532 , n3531 , n3510 );
nor ( n3533 , n3529 , n3532 );
nand ( n3534 , n3517 , n3525 , n3533 );
nand ( n3535 , n3505 , n3534 );
not ( n3536 , n402 );
nand ( n3537 , n1152 , n3041 );
nor ( n3538 , n3536 , n3537 );
not ( n3539 , n3139 );
not ( n3540 , n3472 );
nand ( n3541 , n3540 , n3034 );
and ( n3542 , n3538 , n3539 , n3541 );
nor ( n3543 , n3542 , n3076 );
not ( n3544 , n910 );
nand ( n3545 , n3544 , n3513 );
not ( n3546 , n3517 );
nand ( n3547 , n3546 , n1152 );
nand ( n3548 , n3535 , n3543 , n3545 , n3547 );
and ( n3549 , n2697 , n3548 );
nor ( n3550 , n2644 , n3424 );
nor ( n3551 , n3549 , n3550 );
nand ( n3552 , n3495 , n3504 , n3551 );
nor ( n3553 , n3452 , n3552 );
not ( n3554 , n3121 );
nand ( n3555 , n3554 , n3500 );
and ( n3556 , n3555 , n3415 );
nor ( n3557 , n3556 , n1217 );
nand ( n3558 , n2752 , n3557 );
nand ( n3559 , n3305 , n3077 , n3312 );
not ( n3560 , n3559 );
or ( n3561 , n3295 , n3560 );
not ( n3562 , n2600 );
nand ( n3563 , n3307 , n3331 );
not ( n3564 , n3563 );
or ( n3565 , n3562 , n3564 );
nand ( n3566 , n3561 , n3565 );
nand ( n3567 , n358 , n3566 );
and ( n3568 , n3558 , n3567 );
nand ( n3569 , n3135 , n3471 );
nand ( n3570 , n402 , n880 , n3569 );
and ( n3571 , n3570 , n3160 );
nand ( n3572 , n3300 , n3569 );
nor ( n3573 , n3572 , n3530 );
not ( n3574 , n3573 );
not ( n3575 , n3574 );
and ( n3576 , n3575 , n3126 );
nor ( n3577 , n3576 , n3513 );
nor ( n3578 , n3571 , n3577 );
not ( n3579 , n3578 );
buf ( n3580 , n3155 );
and ( n3581 , n3140 , n3126 );
not ( n3582 , n3581 );
not ( n3583 , n3024 );
not ( n3584 , n3513 );
or ( n3585 , n3583 , n3584 );
not ( n3586 , n3023 );
not ( n3587 , n3117 );
not ( n3588 , n3587 );
or ( n3589 , n3586 , n3588 );
nand ( n3590 , n3589 , n3573 );
nand ( n3591 , n3585 , n3590 );
not ( n3592 , n3591 );
or ( n3593 , n3582 , n3592 );
nand ( n3594 , n3471 , n3068 , n3138 );
and ( n3595 , n3594 , n3545 );
nand ( n3596 , n3593 , n3595 );
nand ( n3597 , n3580 , n3596 );
not ( n3598 , n399 );
or ( n3599 , n3594 , n3598 );
nand ( n3600 , n3599 , n3496 );
not ( n3601 , n3600 );
nand ( n3602 , n3579 , n3597 , n3601 );
not ( n3603 , n3602 );
not ( n3604 , n3603 );
nand ( n3605 , n2886 , n3604 );
not ( n3606 , n3065 );
not ( n3607 , n3606 );
not ( n3608 , n3066 );
nor ( n3609 , n780 , n3608 );
not ( n3610 , n3609 );
buf ( n3611 , n3311 );
not ( n3612 , n3611 );
or ( n3613 , n3610 , n3612 );
not ( n3614 , n3541 );
nand ( n3615 , n3614 , n3469 );
nand ( n3616 , n3060 , n3476 , n3615 );
nand ( n3617 , n3613 , n3616 );
not ( n3618 , n3617 );
or ( n3619 , n3607 , n3618 );
not ( n3620 , n402 );
or ( n3621 , n3620 , n3616 );
not ( n3622 , n3312 );
nand ( n3623 , n3544 , n3622 );
nand ( n3624 , n3621 , n3623 );
not ( n3625 , n3059 );
and ( n3626 , n3625 , n3466 );
not ( n3627 , n3363 );
nor ( n3628 , n3627 , n3483 );
nor ( n3629 , n3626 , n3628 );
or ( n3630 , n3026 , n3629 );
nand ( n3631 , n3630 , n3078 );
nor ( n3632 , n3624 , n3631 );
nand ( n3633 , n3619 , n3632 );
nand ( n3634 , n2694 , n3633 );
not ( n3635 , n2596 );
not ( n3636 , n3230 );
and ( n3637 , n3636 , n3211 );
not ( n3638 , n3530 );
not ( n3639 , n1144 );
and ( n3640 , n3638 , n3639 );
nor ( n3641 , n3640 , n3522 );
and ( n3642 , n3328 , n3641 );
nor ( n3643 , n3637 , n3642 );
and ( n3644 , n3057 , n3471 );
nor ( n3645 , n3644 , n3301 );
nand ( n3646 , n3643 , n3645 , n3289 );
not ( n3647 , n3328 );
nand ( n3648 , n399 , n3647 , n3409 );
nand ( n3649 , n3646 , n3217 , n3648 );
nand ( n3650 , n1553 , n3649 );
not ( n3651 , n3650 );
and ( n3652 , n3635 , n3651 );
not ( n3653 , n3207 );
not ( n3654 , n3500 );
not ( n3655 , n3177 );
or ( n3656 , n3654 , n3655 );
not ( n3657 , n3210 );
or ( n3658 , n3657 , n3590 );
nand ( n3659 , n3656 , n3658 );
and ( n3660 , n3653 , n3659 );
nor ( n3661 , n3660 , n3600 );
nand ( n3662 , n3544 , n3397 );
not ( n3663 , n3662 );
nand ( n3664 , n399 , n3663 );
or ( n3665 , n3574 , n3209 );
nand ( n3666 , n3609 , n3177 );
nand ( n3667 , n3665 , n3666 );
not ( n3668 , n399 );
nor ( n3669 , n3522 , n3177 );
nor ( n3670 , n3668 , n3669 , n3572 );
nor ( n3671 , n3667 , n3670 );
not ( n3672 , n3671 );
nand ( n3673 , n3672 , n3214 );
nand ( n3674 , n3661 , n3664 , n3673 );
and ( n3675 , n3195 , n3674 );
nor ( n3676 , n3652 , n3675 );
not ( n3677 , n402 );
and ( n3678 , n3677 , n3370 );
not ( n3679 , n3611 );
and ( n3680 , n3679 , n3641 );
nor ( n3681 , n3678 , n3680 );
and ( n3682 , n3645 , n3681 );
not ( n3683 , n3282 );
nor ( n3684 , n3682 , n3683 );
or ( n3685 , n1264 , n3684 );
not ( n3686 , n3685 );
and ( n3687 , n2627 , n3686 );
nand ( n3688 , n3186 , n3537 );
not ( n3689 , n3523 );
and ( n3690 , n3688 , n3689 );
nor ( n3691 , n3537 , n3662 );
nor ( n3692 , n3690 , n3691 );
buf ( n3693 , n3171 );
or ( n3694 , n3692 , n3693 );
nand ( n3695 , n3694 , n3078 );
not ( n3696 , n3695 );
or ( n3697 , n3186 , n3666 );
not ( n3698 , n3691 );
nand ( n3699 , n3697 , n3511 , n3698 );
and ( n3700 , n3189 , n3699 );
not ( n3701 , n3518 );
nand ( n3702 , n3701 , n3397 );
not ( n3703 , n3230 );
nand ( n3704 , n1083 , n1209 );
nand ( n3705 , n407 , n3704 );
not ( n3706 , n3705 );
not ( n3707 , n3706 );
or ( n3708 , n3703 , n3707 );
nand ( n3709 , n3708 , n3528 );
not ( n3710 , n3532 );
and ( n3711 , n3702 , n3709 , n3710 );
nor ( n3712 , n3711 , n3186 );
nor ( n3713 , n3700 , n3712 );
nand ( n3714 , n3696 , n3713 );
not ( n3715 , n3714 );
not ( n3716 , n3165 );
nor ( n3717 , n3715 , n3716 );
nor ( n3718 , n3687 , n3717 );
and ( n3719 , n3605 , n3634 , n3676 , n3718 );
nand ( n3720 , n3553 , n3568 , n3719 );
nand ( n3721 , n2029 , n3720 );
not ( n3722 , n3552 );
not ( n3723 , n3560 );
and ( n3724 , n2896 , n3723 );
and ( n3725 , n2894 , n3563 );
nor ( n3726 , n3724 , n3725 );
nand ( n3727 , n3719 , n3722 , n3726 );
nand ( n3728 , n1358 , n2926 , n3347 );
nor ( n3729 , n1251 , n1764 );
not ( n3730 , n2265 );
not ( n3731 , n1378 );
nand ( n3732 , n1135 , n2871 );
nand ( n3733 , n2094 , n3732 );
or ( n3734 , n3729 , n3730 , n3731 , n3733 );
and ( n3735 , n3734 , n3340 );
nor ( n3736 , n3735 , n3355 );
and ( n3737 , n2691 , n3271 );
not ( n3738 , n3278 );
nand ( n3739 , n3738 , n3558 );
nor ( n3740 , n3737 , n3739 );
nand ( n3741 , n3728 , n3736 , n3740 );
or ( n3742 , n3727 , n3741 );
nand ( n3743 , n3742 , n2023 );
nand ( n3744 , n3458 , n3721 , n3743 );
and ( n3745 , n2025 , n3744 );
not ( n3746 , n64 );
nand ( n3747 , n392 , n1697 );
and ( n3748 , n3445 , n3747 );
not ( n3749 , n1427 );
or ( n3750 , n3748 , n3749 );
nand ( n3751 , n790 , n3263 );
not ( n3752 , n3751 );
not ( n3753 , n3747 );
or ( n3754 , n3752 , n3753 );
and ( n3755 , n265 , n2763 );
nand ( n3756 , n3754 , n3755 );
nand ( n3757 , n3750 , n3756 );
nand ( n3758 , n311 , n3757 );
or ( n3759 , n1297 , n3758 );
not ( n3760 , n311 );
not ( n3761 , n3756 );
nand ( n3762 , n3760 , n1297 , n3761 );
nand ( n3763 , n1670 , n1830 );
nand ( n3764 , n3258 , n3763 );
nand ( n3765 , n3759 , n3762 , n3764 );
and ( n3766 , n3746 , n3765 );
nand ( n3767 , n3258 , n1831 );
and ( n3768 , n3767 , n3756 );
or ( n3769 , n1775 , n3768 );
nor ( n3770 , n358 , n2849 );
nor ( n3771 , n2069 , n3770 );
or ( n3772 , n1244 , n3771 );
not ( n3773 , n3733 );
nand ( n3774 , n3772 , n3773 );
and ( n3775 , n3774 , n3757 );
and ( n3776 , n1344 , n3763 , n3251 );
nor ( n3777 , n3562 , n3747 );
nor ( n3778 , n3776 , n3777 );
not ( n3779 , n3764 );
nand ( n3780 , n948 , n3779 );
nand ( n3781 , n3778 , n3780 , n3418 );
and ( n3782 , n1217 , n1379 );
nor ( n3783 , n3782 , n3748 );
nor ( n3784 , n3775 , n3781 , n3783 );
nand ( n3785 , n3769 , n3784 );
nor ( n3786 , n3766 , n3785 , n3454 );
nand ( n3787 , n2888 , n3112 );
and ( n3788 , n3786 , n3787 , n3438 );
nand ( n3789 , n2694 , n3079 );
and ( n3790 , n3789 , n3413 , n3439 );
and ( n3791 , n3788 , n3239 , n3790 );
nor ( n3792 , n3791 , n2371 );
nor ( n3793 , n3745 , n3792 );
and ( n3794 , n3193 , n3453 );
nand ( n3795 , n3243 , n2093 );
not ( n3796 , n64 );
nand ( n3797 , n3796 , n3450 );
and ( n3798 , n3795 , n3797 );
nand ( n3799 , n3798 , n3436 );
nand ( n3800 , n2627 , n3799 );
nand ( n3801 , n3794 , n3800 , n3790 );
nand ( n3802 , n3801 , n372 );
not ( n3803 , n3715 );
nand ( n3804 , n3803 , n2794 , n2087 );
or ( n3805 , n1464 , n1924 );
or ( n3806 , n358 , n1216 );
nand ( n3807 , n3805 , n3806 );
nand ( n3808 , n3807 , n3251 );
nand ( n3809 , n329 , n2129 , n3112 );
and ( n3810 , n3808 , n3809 );
not ( n3811 , n2610 );
nor ( n3812 , n1435 , n2087 );
or ( n3813 , n1495 , n3812 );
nand ( n3814 , n1350 , n1765 );
nand ( n3815 , n3813 , n3814 );
not ( n3816 , n3815 );
and ( n3817 , n3811 , n3816 );
nand ( n3818 , n3243 , n2613 );
nor ( n3819 , n3817 , n3818 );
not ( n3820 , n3450 );
not ( n3821 , n3820 );
not ( n3822 , n3250 );
nand ( n3823 , n1411 , n3822 );
not ( n3824 , n3823 );
and ( n3825 , n2596 , n3824 );
or ( n3826 , n3819 , n3821 , n3825 );
and ( n3827 , n1760 , n1465 , n1495 );
or ( n3828 , n3827 , n3815 );
nand ( n3829 , n3826 , n3828 );
nand ( n3830 , n3818 , n3820 );
not ( n3831 , n3830 );
not ( n3832 , n3831 );
not ( n3833 , n3236 );
or ( n3834 , n3832 , n3833 );
nor ( n3835 , n1465 , n1029 );
nand ( n3836 , n3834 , n3835 );
and ( n3837 , n3804 , n3810 , n3829 , n3836 );
and ( n3838 , n3802 , n3837 );
not ( n3839 , n2596 );
not ( n3840 , n3264 );
nor ( n3841 , n3258 , n3840 );
not ( n3842 , n3841 );
or ( n3843 , n3839 , n3842 );
not ( n3844 , n1138 );
not ( n3845 , n3602 );
or ( n3846 , n3844 , n3845 );
not ( n3847 , n1246 );
not ( n3848 , n3674 );
or ( n3849 , n3847 , n3848 );
not ( n3850 , n3557 );
nand ( n3851 , n3849 , n3850 );
not ( n3852 , n3851 );
nand ( n3853 , n3846 , n3852 );
and ( n3854 , n3243 , n1245 );
and ( n3855 , n24 , n3450 );
nor ( n3856 , n3854 , n3855 );
not ( n3857 , n3856 );
nor ( n3858 , n3853 , n3857 );
or ( n3859 , n2120 , n3858 );
not ( n3860 , n1138 );
not ( n3861 , n3162 );
or ( n3862 , n3860 , n3861 );
not ( n3863 , n1246 );
not ( n3864 , n3218 );
or ( n3865 , n3863 , n3864 );
nand ( n3866 , n3865 , n3416 );
not ( n3867 , n3866 );
nand ( n3868 , n3862 , n3867 );
not ( n3869 , n3868 );
and ( n3870 , n3869 , n3856 );
nor ( n3871 , n3870 , n1465 );
not ( n3872 , n3871 );
nand ( n3873 , n3859 , n3872 );
nand ( n3874 , n3843 , n3873 );
or ( n3875 , n3830 , n3825 );
nand ( n3876 , n3875 , n358 );
nand ( n3877 , n1291 , n3649 );
nand ( n3878 , n3685 , n3798 , n3877 );
and ( n3879 , n3878 , n2627 );
not ( n3880 , n2694 );
not ( n3881 , n3633 );
or ( n3882 , n3880 , n3881 );
nand ( n3883 , n3882 , n3567 );
nor ( n3884 , n3879 , n3883 );
nand ( n3885 , n3722 , n3876 , n3884 );
nand ( n3886 , n3885 , n1464 );
nand ( n3887 , n3838 , n3874 , n3886 );
buf ( n3888 , n3887 );
nand ( n3889 , n1627 , n3888 );
nand ( n3890 , n3764 , n3758 );
and ( n3891 , n2926 , n3890 );
not ( n3892 , n2823 );
not ( n3893 , n3757 );
or ( n3894 , n3892 , n3893 );
or ( n3895 , n3295 , n3747 );
nand ( n3896 , n3894 , n3895 );
or ( n3897 , n1775 , n3767 );
not ( n3898 , n2916 );
not ( n3899 , n3898 );
not ( n3900 , n3899 );
not ( n3901 , n3763 );
not ( n3902 , n3825 );
or ( n3903 , n3901 , n3902 );
nand ( n3904 , n3903 , n3756 );
and ( n3905 , n311 , n3904 );
nor ( n3906 , n3905 , n3779 );
or ( n3907 , n3900 , n3906 );
nand ( n3908 , n3897 , n3907 , n3558 );
nor ( n3909 , n3891 , n3896 , n3908 );
not ( n3910 , n3727 );
nand ( n3911 , n3909 , n3910 );
nand ( n3912 , n2276 , n3911 );
not ( n3913 , n401 );
not ( n3914 , n1421 );
not ( n3915 , n3098 );
and ( n3916 , n722 , n3915 );
not ( n3917 , n3916 );
nand ( n3918 , n3803 , n3917 );
not ( n3919 , n724 );
not ( n3920 , n3318 );
or ( n3921 , n3919 , n3920 );
or ( n3922 , n386 , n388 );
nand ( n3923 , n3922 , n392 );
nand ( n3924 , n3921 , n3923 );
not ( n3925 , n3924 );
nand ( n3926 , n3918 , n3925 );
and ( n3927 , n3926 , n953 );
and ( n3928 , n3917 , n3497 );
nor ( n3929 , n3928 , n3924 );
or ( n3930 , n1345 , n3929 );
nor ( n3931 , n3916 , n3424 );
or ( n3932 , n3924 , n3931 );
nand ( n3933 , n3932 , n1488 );
nand ( n3934 , n3930 , n3933 );
nor ( n3935 , n3927 , n3934 );
not ( n3936 , n3917 );
not ( n3937 , n3602 );
or ( n3938 , n3936 , n3937 );
nand ( n3939 , n3938 , n3925 );
nand ( n3940 , n3939 , n1138 );
nand ( n3941 , n1253 , n3924 );
nand ( n3942 , n3851 , n3917 );
nand ( n3943 , n3940 , n3941 , n3942 );
nor ( n3944 , n3943 , n3855 );
and ( n3945 , n3935 , n3944 );
nor ( n3946 , n3945 , n2747 );
not ( n3947 , n3684 );
nand ( n3948 , n3947 , n3917 );
and ( n3949 , n3925 , n3948 );
nor ( n3950 , n3949 , n1264 );
nand ( n3951 , n3917 , n3649 );
and ( n3952 , n3951 , n3925 );
nor ( n3953 , n3952 , n1565 );
nor ( n3954 , n3950 , n3953 );
and ( n3955 , n3797 , n3954 );
nor ( n3956 , n3955 , n1027 );
or ( n3957 , n1496 , n3925 );
and ( n3958 , n1402 , n3559 );
and ( n3959 , n1344 , n3563 );
nor ( n3960 , n3958 , n3959 );
not ( n3961 , n3960 );
not ( n3962 , n3961 );
nand ( n3963 , n3633 , n1013 );
and ( n3964 , n3962 , n3963 );
nor ( n3965 , n3964 , n3916 );
not ( n3966 , n3965 );
nand ( n3967 , n3957 , n3966 );
or ( n3968 , n3956 , n3967 );
nand ( n3969 , n3968 , n2778 );
not ( n3970 , n3858 );
nand ( n3971 , n3970 , n2752 );
not ( n3972 , n2747 );
nand ( n3973 , n3917 , n3548 );
and ( n3974 , n3925 , n3973 );
nor ( n3975 , n3974 , n1014 );
nand ( n3976 , n3972 , n3975 );
nand ( n3977 , n3969 , n3971 , n3976 );
nand ( n3978 , n2100 , n3830 );
nand ( n3979 , n3502 , n1538 , n3917 );
not ( n3980 , n3925 );
nand ( n3981 , n3917 , n3411 );
not ( n3982 , n3981 );
or ( n3983 , n3980 , n3982 );
nand ( n3984 , n3983 , n1538 );
nand ( n3985 , n3979 , n3984 );
nand ( n3986 , n2596 , n3985 );
nand ( n3987 , n3978 , n3986 , n3884 );
not ( n3988 , n3987 );
nor ( n3989 , n3492 , n3916 );
nor ( n3990 , n3924 , n3989 );
nor ( n3991 , n2728 , n3990 );
and ( n3992 , n3991 , n2691 );
nor ( n3993 , n3992 , n3717 );
nand ( n3994 , n3988 , n3993 , n3722 );
nor ( n3995 , n3946 , n3977 , n3994 );
or ( n3996 , n3914 , n3995 );
and ( n3997 , n2472 , n3887 );
not ( n3998 , n1545 );
nand ( n3999 , n3998 , n3821 );
and ( n4000 , n3374 , n3917 );
nor ( n4001 , n4000 , n3924 );
or ( n4002 , n1547 , n4001 );
not ( n4003 , n3291 );
or ( n4004 , n4003 , n3916 );
nand ( n4005 , n4004 , n3925 );
nand ( n4006 , n1553 , n4005 );
nand ( n4007 , n4002 , n4006 , n3984 );
not ( n4008 , n4007 );
not ( n4009 , n3917 );
not ( n4010 , n3162 );
or ( n4011 , n4009 , n4010 );
nand ( n4012 , n4011 , n3925 );
nand ( n4013 , n1138 , n4012 );
nand ( n4014 , n3917 , n3866 );
nand ( n4015 , n4013 , n3941 , n4014 );
or ( n4016 , n4015 , n3855 );
not ( n4017 , n358 );
nand ( n4018 , n4016 , n4017 );
nand ( n4019 , n3999 , n4008 , n4018 );
not ( n4020 , n4019 );
not ( n4021 , n3925 );
nand ( n4022 , n3917 , n3192 );
not ( n4023 , n4022 );
or ( n4024 , n4021 , n4023 );
nand ( n4025 , n4024 , n953 );
not ( n4026 , n311 );
not ( n4027 , n3402 );
or ( n4028 , n4027 , n3916 );
nand ( n4029 , n4028 , n3925 );
nand ( n4030 , n4026 , n4029 );
not ( n4031 , n4030 );
nand ( n4032 , n3430 , n3917 );
nand ( n4033 , n3925 , n4032 );
nand ( n4034 , n311 , n4033 );
not ( n4035 , n4034 );
or ( n4036 , n4031 , n4035 );
nand ( n4037 , n4036 , n1109 );
not ( n4038 , n3925 );
nand ( n4039 , n3917 , n3235 );
not ( n4040 , n4039 );
or ( n4041 , n4038 , n4040 );
nand ( n4042 , n4041 , n1013 );
nand ( n4043 , n4037 , n4042 );
nor ( n4044 , n4043 , n4015 );
and ( n4045 , n4025 , n4044 );
nor ( n4046 , n4045 , n358 );
not ( n4047 , n358 );
nor ( n4048 , n3080 , n3916 );
nand ( n4049 , n1013 , n4048 );
or ( n4050 , n1109 , n1013 );
nand ( n4051 , n4050 , n3924 );
or ( n4052 , n1403 , n3325 );
nand ( n4053 , n1344 , n3335 );
nand ( n4054 , n4052 , n4053 );
nand ( n4055 , n3917 , n4054 );
nand ( n4056 , n4049 , n4051 , n4055 );
not ( n4057 , n4056 );
or ( n4058 , n4047 , n4057 );
nand ( n4059 , n3917 , n3112 );
and ( n4060 , n3925 , n4059 );
nor ( n4061 , n4060 , n1747 );
nor ( n4062 , n4061 , n4007 );
nand ( n4063 , n4058 , n4062 );
nor ( n4064 , n4046 , n4063 );
and ( n4065 , n4020 , n4064 );
nand ( n4066 , n2596 , n1586 );
nor ( n4067 , n4065 , n4066 );
nor ( n4068 , n3997 , n4067 );
and ( n4069 , n3809 , n3836 );
and ( n4070 , n329 , n3871 );
and ( n4071 , n2660 , n3814 );
nor ( n4072 , n4071 , n3831 );
nor ( n4073 , n4070 , n4072 );
nand ( n4074 , n4069 , n4073 , n3802 );
nand ( n4075 , n2127 , n4074 );
nand ( n4076 , n3996 , n4068 , n4075 );
nand ( n4077 , n3913 , n4076 );
nand ( n4078 , n3793 , n3889 , n3912 , n4077 );
nand ( n4079 , n3018 , n4078 , n2495 );
not ( n4080 , n3975 );
not ( n4081 , n4080 );
not ( n4082 , n3944 );
or ( n4083 , n4081 , n4082 );
not ( n4084 , n2120 );
nand ( n4085 , n4083 , n4084 );
or ( n4086 , n2166 , n3929 );
or ( n4087 , n358 , n3933 );
not ( n4088 , n3985 );
nand ( n4089 , n4086 , n4087 , n4088 );
nand ( n4090 , n1464 , n4089 );
not ( n4091 , n2102 );
not ( n4092 , n3821 );
not ( n4093 , n4092 );
and ( n4094 , n4091 , n4093 );
and ( n4095 , n3926 , n2174 );
nor ( n4096 , n4094 , n4095 );
nand ( n4097 , n4085 , n4090 , n4096 );
not ( n4098 , n3956 );
nor ( n4099 , n952 , n3990 );
nor ( n4100 , n4099 , n3967 );
and ( n4101 , n4098 , n4100 );
nor ( n4102 , n4101 , n1760 );
or ( n4103 , n4097 , n4102 );
nand ( n4104 , n4103 , n1825 );
not ( n4105 , n358 );
nand ( n4106 , n4042 , n4025 );
and ( n4107 , n4105 , n4106 );
nor ( n4108 , n4107 , n4061 );
not ( n4109 , n4108 );
not ( n4110 , n4020 );
or ( n4111 , n4109 , n4110 );
nand ( n4112 , n4111 , n1586 );
not ( n4113 , n4092 );
nand ( n4114 , n4113 , n1772 );
nand ( n4115 , n4104 , n4112 , n4114 );
not ( n4116 , n4056 );
or ( n4117 , n1436 , n4116 );
not ( n4118 , n4033 );
or ( n4119 , n2137 , n4118 );
not ( n4120 , n2134 );
and ( n4121 , n4120 , n4029 );
nand ( n4122 , n3449 , n3823 );
and ( n4123 , n2472 , n4122 );
nor ( n4124 , n4121 , n4123 );
nand ( n4125 , n4117 , n4119 , n4124 );
or ( n4126 , n4115 , n4125 );
not ( n4127 , n401 );
nand ( n4128 , n4126 , n4127 );
and ( n4129 , n3441 , n3443 );
nor ( n4130 , n4129 , n1658 );
or ( n4131 , n1425 , n3451 );
nand ( n4132 , n1661 , n3246 , n4122 );
nand ( n4133 , n4131 , n4132 );
not ( n4134 , n4133 );
nor ( n4135 , n4134 , n1655 );
nor ( n4136 , n4130 , n4135 );
and ( n4137 , n1627 , n4122 );
nand ( n4138 , n3763 , n3824 );
and ( n4139 , n4138 , n3768 );
nor ( n4140 , n4139 , n1633 );
nor ( n4141 , n4137 , n4140 );
nand ( n4142 , n4128 , n4136 , n4141 );
nand ( n4143 , n4142 , n1734 , n395 );
not ( n4144 , n1848 );
and ( n4145 , n4144 , n3915 );
buf ( n4146 , n4145 );
or ( n4147 , n4146 , n3424 );
not ( n4148 , n4144 );
not ( n4149 , n3318 );
or ( n4150 , n4148 , n4149 );
nand ( n4151 , n4150 , n3923 );
not ( n4152 , n4151 );
not ( n4153 , n4152 );
not ( n4154 , n4153 );
nand ( n4155 , n4147 , n4154 );
nand ( n4156 , n1807 , n4155 );
or ( n4157 , n720 , n4152 );
buf ( n4158 , n4146 );
or ( n4159 , n4158 , n3960 );
nand ( n4160 , n4157 , n4159 );
nand ( n4161 , n4160 , n358 );
and ( n4162 , n4156 , n4161 );
nor ( n4163 , n358 , n4145 );
nand ( n4164 , n4163 , n3557 );
not ( n4165 , n4145 );
nand ( n4166 , n1538 , n4165 );
not ( n4167 , n4166 );
nand ( n4168 , n4167 , n3502 );
not ( n4169 , n4145 );
not ( n4170 , n3415 );
and ( n4171 , n4169 , n4170 );
nor ( n4172 , n4171 , n4153 );
not ( n4173 , n4172 );
not ( n4174 , n1946 );
and ( n4175 , n4173 , n4174 );
or ( n4176 , n4145 , n3412 );
not ( n4177 , n4153 );
nand ( n4178 , n4176 , n4177 );
and ( n4179 , n1538 , n4178 );
nor ( n4180 , n4175 , n4179 );
and ( n4181 , n4164 , n4168 , n4180 );
not ( n4182 , n1961 );
buf ( n4183 , n4158 );
or ( n4184 , n3603 , n4183 );
buf ( n4185 , n4154 );
buf ( n4186 , n4185 );
nand ( n4187 , n4184 , n4186 );
not ( n4188 , n4187 );
or ( n4189 , n4182 , n4188 );
not ( n4190 , n4146 );
nand ( n4191 , n4190 , n3674 );
and ( n4192 , n4186 , n4191 );
nor ( n4193 , n4192 , n1379 );
or ( n4194 , n4158 , n3684 );
and ( n4195 , n4186 , n4194 );
nor ( n4196 , n4195 , n1547 );
nor ( n4197 , n4193 , n4196 );
nand ( n4198 , n4189 , n4197 );
not ( n4199 , n4198 );
nand ( n4200 , n4162 , n4181 , n4199 );
nand ( n4201 , n4200 , n1464 );
not ( n4202 , n4185 );
nand ( n4203 , n4190 , n3649 );
not ( n4204 , n4203 );
or ( n4205 , n4202 , n4204 );
nand ( n4206 , n4205 , n1553 );
not ( n4207 , n358 );
buf ( n4208 , n4186 );
not ( n4209 , n4183 );
nand ( n4210 , n4209 , n3548 );
and ( n4211 , n4208 , n4210 );
nor ( n4212 , n4211 , n1014 );
nand ( n4213 , n4207 , n4212 );
and ( n4214 , n4206 , n4213 );
nor ( n4215 , n4214 , n372 );
not ( n4216 , n1925 );
buf ( n4217 , n4146 );
not ( n4218 , n3235 );
or ( n4219 , n4217 , n4218 );
nand ( n4220 , n4219 , n4186 );
not ( n4221 , n4220 );
or ( n4222 , n4216 , n4221 );
nand ( n4223 , n3112 , n4190 );
and ( n4224 , n4186 , n4223 );
nor ( n4225 , n4224 , n1747 );
not ( n4226 , n4225 );
nand ( n4227 , n4222 , n4226 );
and ( n4228 , n4227 , n372 );
nand ( n4229 , n2226 , n1404 );
not ( n4230 , n4146 );
not ( n4231 , n4230 );
not ( n4232 , n3430 );
or ( n4233 , n4231 , n4232 );
nand ( n4234 , n4233 , n4185 );
not ( n4235 , n4234 );
or ( n4236 , n4229 , n4235 );
nand ( n4237 , n4165 , n3497 );
nand ( n4238 , n4154 , n4237 );
and ( n4239 , n2223 , n4238 );
and ( n4240 , n1778 , n3821 );
nor ( n4241 , n4239 , n4240 );
nor ( n4242 , n1464 , n2166 );
nand ( n4243 , n4165 , n3402 );
nand ( n4244 , n4154 , n4243 );
nand ( n4245 , n4242 , n4244 );
nand ( n4246 , n4236 , n4241 , n4245 );
nor ( n4247 , n4228 , n4246 );
not ( n4248 , n4217 );
nand ( n4249 , n3714 , n4248 );
nand ( n4250 , n4186 , n4249 );
and ( n4251 , n2174 , n4250 );
not ( n4252 , n2177 );
nand ( n4253 , n4248 , n3192 );
nand ( n4254 , n4186 , n4253 );
not ( n4255 , n4254 );
nor ( n4256 , n4252 , n4255 );
nor ( n4257 , n4251 , n4256 );
nand ( n4258 , n4247 , n4257 );
nor ( n4259 , n4215 , n4258 );
not ( n4260 , n4157 );
nand ( n4261 , n3079 , n4190 );
and ( n4262 , n4185 , n4261 );
nor ( n4263 , n4262 , n1014 );
not ( n4264 , n4054 );
nor ( n4265 , n4217 , n4264 );
nor ( n4266 , n4263 , n4265 );
not ( n4267 , n4266 );
or ( n4268 , n4260 , n4267 );
nand ( n4269 , n4268 , n358 );
not ( n4270 , n3162 );
or ( n4271 , n4270 , n4183 );
nand ( n4272 , n4271 , n4186 );
nand ( n4273 , n1961 , n4272 );
not ( n4274 , n4230 );
not ( n4275 , n3218 );
or ( n4276 , n4274 , n4275 );
nand ( n4277 , n4276 , n4185 );
and ( n4278 , n1380 , n4277 );
not ( n4279 , n4146 );
nand ( n4280 , n4279 , n3291 );
and ( n4281 , n4185 , n4280 );
nor ( n4282 , n4281 , n1554 );
nor ( n4283 , n4278 , n4282 );
not ( n4284 , n4185 );
nand ( n4285 , n4279 , n3374 );
not ( n4286 , n4285 );
or ( n4287 , n4284 , n4286 );
nand ( n4288 , n4287 , n1546 );
and ( n4289 , n4283 , n4180 , n4288 );
nand ( n4290 , n4269 , n4273 , n4289 );
and ( n4291 , n372 , n4290 );
not ( n4292 , n372 );
not ( n4293 , n4186 );
not ( n4294 , n4158 );
nand ( n4295 , n3493 , n4294 );
not ( n4296 , n4295 );
or ( n4297 , n4293 , n4296 );
nand ( n4298 , n4297 , n953 );
not ( n4299 , n4183 );
not ( n4300 , n4299 );
not ( n4301 , n3633 );
or ( n4302 , n4300 , n4301 );
nand ( n4303 , n4302 , n4208 );
nand ( n4304 , n4303 , n1013 );
and ( n4305 , n4298 , n4304 );
not ( n4306 , n358 );
nor ( n4307 , n4305 , n4306 );
and ( n4308 , n4292 , n4307 );
nor ( n4309 , n4291 , n4308 );
nand ( n4310 , n4201 , n4259 , n4309 );
nand ( n4311 , n4310 , n2472 );
and ( n4312 , n2143 , n3235 );
not ( n4313 , n3080 );
and ( n4314 , n1607 , n4313 );
nor ( n4315 , n4312 , n4314 );
and ( n4316 , n2130 , n3112 );
and ( n4317 , n2475 , n3192 );
not ( n4318 , n2132 );
not ( n4319 , n3335 );
or ( n4320 , n4318 , n4319 );
or ( n4321 , n2134 , n4027 );
nand ( n4322 , n4320 , n4321 );
nor ( n4323 , n4316 , n4317 , n4322 );
not ( n4324 , n1760 );
not ( n4325 , n3963 );
and ( n4326 , n4324 , n4325 );
nor ( n4327 , n4326 , n3873 );
and ( n4328 , n2077 , n3799 );
not ( n4329 , n2174 );
not ( n4330 , n3803 );
or ( n4331 , n4329 , n4330 );
and ( n4332 , n358 , n3961 );
nand ( n4333 , n791 , n3410 );
not ( n4334 , n4333 );
nand ( n4335 , n4334 , n3501 );
and ( n4336 , n1538 , n4335 );
not ( n4337 , n3424 );
and ( n4338 , n1807 , n4337 );
nor ( n4339 , n4332 , n4336 , n4338 );
or ( n4340 , n372 , n4339 );
nand ( n4341 , n4331 , n4340 );
nor ( n4342 , n4328 , n4341 );
nand ( n4343 , n2109 , n3878 );
and ( n4344 , n64 , n2100 , n3821 );
or ( n4345 , n3242 , n1068 );
nand ( n4346 , n4345 , n3798 );
and ( n4347 , n1027 , n4346 );
nor ( n4348 , n4344 , n4347 );
and ( n4349 , n2223 , n3497 );
and ( n4350 , n2106 , n4333 );
nor ( n4351 , n4349 , n4350 );
not ( n4352 , n3325 );
and ( n4353 , n2097 , n4352 );
not ( n4354 , n4229 );
and ( n4355 , n4354 , n3430 );
nor ( n4356 , n4353 , n4355 );
and ( n4357 , n1464 , n1925 , n3548 );
nor ( n4358 , n3494 , n1760 , n952 );
nor ( n4359 , n4357 , n4358 );
and ( n4360 , n4348 , n4351 , n4356 , n4359 );
nand ( n4361 , n4327 , n4342 , n4343 , n4360 );
nand ( n4362 , n1825 , n4361 );
nand ( n4363 , n4311 , n4315 , n4323 , n4362 );
not ( n4364 , n401 );
nand ( n4365 , n4363 , n4364 );
and ( n4366 , n1841 , n4153 );
not ( n4367 , n4366 );
nand ( n4368 , n4299 , n3633 );
nand ( n4369 , n4367 , n4368 );
nand ( n4370 , n1361 , n4369 );
not ( n4371 , n4370 );
nand ( n4372 , n4206 , n4181 );
nor ( n4373 , n4198 , n4372 );
and ( n4374 , n1643 , n4373 );
not ( n4375 , n4208 );
nand ( n4376 , n1361 , n4375 );
not ( n4377 , n358 );
not ( n4378 , n3451 );
not ( n4379 , n4160 );
nand ( n4380 , n4379 , n4298 );
nor ( n4381 , n4378 , n4380 );
not ( n4382 , n4381 );
or ( n4383 , n4377 , n4382 );
not ( n4384 , n4212 );
not ( n4385 , n358 );
nand ( n4386 , n4250 , n953 );
and ( n4387 , n1344 , n4238 );
and ( n4388 , n1404 , n4155 );
nor ( n4389 , n4387 , n4388 );
nand ( n4390 , n4386 , n4389 );
and ( n4391 , n1643 , n4390 );
nor ( n4392 , n4391 , n4378 );
nand ( n4393 , n4384 , n4385 , n4392 );
nand ( n4394 , n4383 , n4393 );
nand ( n4395 , n4374 , n4376 , n4394 );
nand ( n4396 , n1245 , n4366 );
not ( n4397 , n4396 );
nand ( n4398 , n3853 , n4299 );
not ( n4399 , n4398 );
or ( n4400 , n4397 , n4399 );
not ( n4401 , n358 );
nand ( n4402 , n4400 , n4401 );
not ( n4403 , n4183 );
not ( n4404 , n3650 );
and ( n4405 , n4403 , n4404 );
not ( n4406 , n4396 );
and ( n4407 , n358 , n4406 );
nor ( n4408 , n4405 , n4407 );
not ( n4409 , n4194 );
nand ( n4410 , n1546 , n4409 );
and ( n4411 , n4408 , n4168 , n4410 );
nand ( n4412 , n4367 , n4210 );
nand ( n4413 , n1925 , n4412 );
nand ( n4414 , n4402 , n4411 , n4413 );
not ( n4415 , n4414 );
or ( n4416 , n1345 , n4237 );
nor ( n4417 , n1403 , n4146 );
nand ( n4418 , n4417 , n4337 );
or ( n4419 , n1842 , n4157 );
nand ( n4420 , n4416 , n4418 , n4419 );
and ( n4421 , n4367 , n4249 );
nor ( n4422 , n4421 , n952 );
nor ( n4423 , n4420 , n4422 );
not ( n4424 , n4423 );
not ( n4425 , n4392 );
or ( n4426 , n4424 , n4425 );
not ( n4427 , n358 );
nand ( n4428 , n4426 , n4427 );
and ( n4429 , n4419 , n4159 );
nand ( n4430 , n4295 , n4367 );
nand ( n4431 , n953 , n4430 );
and ( n4432 , n4429 , n4431 );
nand ( n4433 , n3451 , n4432 );
and ( n4434 , n4433 , n358 );
nor ( n4435 , n4434 , n1643 );
nand ( n4436 , n4415 , n4428 , n4435 );
nand ( n4437 , n4395 , n4436 );
not ( n4438 , n4437 );
or ( n4439 , n4371 , n4438 );
nand ( n4440 , n4439 , n2032 );
nand ( n4441 , n4367 , n4219 );
and ( n4442 , n1925 , n4441 );
and ( n4443 , n4417 , n3430 );
or ( n4444 , n1345 , n4243 );
nand ( n4445 , n4444 , n4419 );
nor ( n4446 , n4443 , n4445 );
nor ( n4447 , n358 , n4446 );
nor ( n4448 , n4442 , n4447 );
not ( n4449 , n4448 );
not ( n4450 , n4163 );
not ( n4451 , n3868 );
or ( n4452 , n4450 , n4451 );
or ( n4453 , n4285 , n1547 );
nand ( n4454 , n4453 , n4396 );
or ( n4455 , n4280 , n1554 );
or ( n4456 , n4166 , n3412 );
nand ( n4457 , n4455 , n4456 );
nor ( n4458 , n4454 , n4457 );
nand ( n4459 , n4452 , n4458 );
not ( n4460 , n4459 );
and ( n4461 , n4367 , n4261 );
nor ( n4462 , n4461 , n1014 );
not ( n4463 , n4265 );
nand ( n4464 , n4419 , n4463 );
or ( n4465 , n4462 , n4464 );
nand ( n4466 , n4465 , n358 );
nand ( n4467 , n4460 , n4466 );
nor ( n4468 , n1643 , n4467 );
not ( n4469 , n4468 );
or ( n4470 , n4449 , n4469 );
not ( n4471 , n358 );
and ( n4472 , n4220 , n1013 );
not ( n4473 , n311 );
and ( n4474 , n4473 , n4244 );
not ( n4475 , n4473 );
and ( n4476 , n4475 , n4234 );
nor ( n4477 , n4474 , n4476 );
nor ( n4478 , n720 , n4477 );
nor ( n4479 , n4472 , n4478 );
not ( n4480 , n4479 );
nand ( n4481 , n4471 , n4480 );
not ( n4482 , n4290 );
nand ( n4483 , n1643 , n4481 , n4482 );
nand ( n4484 , n4470 , n4483 );
and ( n4485 , n3448 , n4375 );
not ( n4486 , n358 );
not ( n4487 , n3192 );
and ( n4488 , n4486 , n4487 );
not ( n4489 , n4163 );
and ( n4490 , n4489 , n4223 );
nor ( n4491 , n4488 , n4490 );
nor ( n4492 , n4485 , n4491 );
or ( n4493 , n952 , n4492 );
nand ( n4494 , n4484 , n4493 , n3451 );
nand ( n4495 , n4494 , n2339 );
nand ( n4496 , n4365 , n4440 , n4495 );
nand ( n4497 , n1627 , n4310 );
not ( n4498 , n358 );
not ( n4499 , n4498 );
nand ( n4500 , n953 , n4254 );
and ( n4501 , n4500 , n4479 );
or ( n4502 , n1830 , n4501 );
or ( n4503 , n2906 , n3768 );
nor ( n4504 , n3779 , n3761 );
not ( n4505 , n4504 );
nand ( n4506 , n2906 , n4505 );
nand ( n4507 , n4502 , n4503 , n4506 );
not ( n4508 , n4507 );
or ( n4509 , n4499 , n4508 );
not ( n4510 , n358 );
not ( n4511 , n4510 );
not ( n4512 , n4503 );
and ( n4513 , n4511 , n4512 );
nor ( n4514 , n2933 , n4504 );
nor ( n4515 , n4513 , n4514 );
nand ( n4516 , n4509 , n4515 );
nor ( n4517 , n4290 , n4225 );
or ( n4518 , n1830 , n4517 );
not ( n4519 , n4367 );
not ( n4520 , n4253 );
or ( n4521 , n4519 , n4520 );
nand ( n4522 , n4521 , n953 );
and ( n4523 , n4446 , n4522 );
nor ( n4524 , n4523 , n358 );
or ( n4525 , n4467 , n4524 );
nand ( n4526 , n4525 , n2365 );
nor ( n4527 , n1646 , n1747 );
nand ( n4528 , n4367 , n4223 );
nand ( n4529 , n4527 , n4528 );
nand ( n4530 , n4518 , n4526 , n4529 );
or ( n4531 , n4516 , n4530 );
nand ( n4532 , n4531 , n2366 );
not ( n4533 , n2026 );
nand ( n4534 , n1013 , n4369 );
and ( n4535 , n4534 , n4432 );
not ( n4536 , n1840 );
nor ( n4537 , n4535 , n4536 );
nand ( n4538 , n358 , n1919 , n4303 );
not ( n4539 , n2410 );
nand ( n4540 , n4539 , n4412 );
and ( n4541 , n4538 , n4540 );
nor ( n4542 , n4541 , n1014 );
or ( n4543 , n4423 , n2410 );
nand ( n4544 , n4543 , n3268 );
nor ( n4545 , n4537 , n4542 , n4544 );
or ( n4546 , n4390 , n4212 );
nand ( n4547 , n4546 , n1892 );
nand ( n4548 , n4402 , n4411 , n1920 );
nand ( n4549 , n358 , n4380 );
not ( n4550 , n2426 );
nand ( n4551 , n4549 , n4550 , n4373 );
nand ( n4552 , n4548 , n4551 );
nand ( n4553 , n4545 , n4547 , n4552 );
nand ( n4554 , n4533 , n4553 );
and ( n4555 , n4497 , n4532 , n4554 );
nand ( n4556 , n2379 , n4441 );
not ( n4557 , n4528 );
or ( n4558 , n952 , n4557 );
not ( n4559 , n4464 );
nand ( n4560 , n4558 , n4559 );
and ( n4561 , n1840 , n4560 );
not ( n4562 , n358 );
not ( n4563 , n4562 );
not ( n4564 , n4218 );
or ( n4565 , n4563 , n4564 );
nand ( n4566 , n4489 , n4261 );
nand ( n4567 , n4565 , n4566 );
and ( n4568 , n4367 , n4567 );
nor ( n4569 , n4568 , n1014 );
and ( n4570 , n2426 , n4569 );
nor ( n4571 , n4561 , n4570 );
or ( n4572 , n4524 , n4459 );
nand ( n4573 , n4572 , n1920 );
nand ( n4574 , n4571 , n3268 , n4573 );
not ( n4575 , n358 );
not ( n4576 , n4501 );
nand ( n4577 , n4575 , n4576 );
and ( n4578 , n4577 , n4517 );
not ( n4579 , n1921 );
nor ( n4580 , n4578 , n4579 );
or ( n4581 , n4574 , n4580 );
nand ( n4582 , n4581 , n2409 );
nor ( n4583 , n4414 , n1646 );
not ( n4584 , n4307 );
or ( n4585 , n358 , n4389 );
nand ( n4586 , n4584 , n4585 , n4161 );
nand ( n4587 , n1646 , n4373 );
nor ( n4588 , n4586 , n4587 );
or ( n4589 , n4583 , n4588 );
and ( n4590 , n4384 , n4386 );
nor ( n4591 , n4590 , n1830 );
not ( n4592 , n4422 );
nor ( n4593 , n2273 , n4592 );
or ( n4594 , n4591 , n4593 );
not ( n4595 , n358 );
nand ( n4596 , n4594 , n4595 );
nand ( n4597 , n4589 , n4515 , n4596 );
not ( n4598 , n2261 );
and ( n4599 , n4598 , n4420 );
not ( n4600 , n358 );
or ( n4601 , n311 , n3780 );
nand ( n4602 , n4601 , n3768 );
and ( n4603 , n4600 , n4602 );
nor ( n4604 , n4599 , n4603 );
nand ( n4605 , n4527 , n4430 );
not ( n4606 , n4429 );
not ( n4607 , n4534 );
or ( n4608 , n4606 , n4607 );
not ( n4609 , n2398 );
nand ( n4610 , n4608 , n4609 );
nand ( n4611 , n4604 , n4605 , n4610 );
or ( n4612 , n4597 , n4611 );
nand ( n4613 , n4612 , n2276 );
nand ( n4614 , n4555 , n4556 , n4582 , n4613 );
or ( n4615 , n4496 , n4614 );
nand ( n4616 , n4615 , n716 );
nand ( n4617 , n4079 , n4143 , n4616 );
nand ( n4618 , n4617 , n714 );
and ( n4619 , n391 , n716 );
not ( n4620 , n3917 );
not ( n4621 , n358 );
not ( n4622 , n4621 );
not ( n4623 , n3853 );
or ( n4624 , n4622 , n4623 );
nand ( n4625 , n4624 , n3650 );
not ( n4626 , n4625 );
or ( n4627 , n4620 , n4626 );
nor ( n4628 , n791 , n1033 );
not ( n4629 , n4628 );
nand ( n4630 , n4629 , n3443 );
nand ( n4631 , n4630 , n3924 );
or ( n4632 , n1496 , n4631 );
nand ( n4633 , n4632 , n358 , n3966 );
or ( n4634 , n952 , n3918 );
not ( n4635 , n4631 );
not ( n4636 , n3973 );
or ( n4637 , n4635 , n4636 );
nand ( n4638 , n4637 , n1013 );
and ( n4639 , n2136 , n3931 );
nand ( n4640 , n1344 , n3917 );
not ( n4641 , n3497 );
or ( n4642 , n4640 , n4641 );
or ( n4643 , n1351 , n4631 );
nand ( n4644 , n4642 , n4643 );
nor ( n4645 , n4639 , n4644 , n358 );
nand ( n4646 , n4634 , n4638 , n4645 );
and ( n4647 , n4633 , n4646 );
not ( n4648 , n4631 );
nand ( n4649 , n1245 , n4648 );
not ( n4650 , n3948 );
nand ( n4651 , n4650 , n1546 );
or ( n4652 , n4648 , n3989 );
nand ( n4653 , n4652 , n1748 );
nand ( n4654 , n4649 , n4651 , n3979 , n4653 );
nor ( n4655 , n4647 , n4654 );
nand ( n4656 , n4627 , n4655 );
and ( n4657 , n1042 , n4656 );
not ( n4658 , n1042 );
not ( n4659 , n3954 );
nand ( n4660 , n4659 , n24 );
not ( n4661 , n4660 );
not ( n4662 , n4100 );
or ( n4663 , n4661 , n4662 );
nand ( n4664 , n4663 , n358 );
not ( n4665 , n358 );
not ( n4666 , n3943 );
nand ( n4667 , n4666 , n3935 , n4080 );
and ( n4668 , n4665 , n4667 );
nor ( n4669 , n4668 , n3985 );
nand ( n4670 , n4664 , n4669 );
and ( n4671 , n4658 , n4670 );
nor ( n4672 , n4657 , n4671 );
or ( n4673 , n791 , n1414 );
and ( n4674 , n3258 , n1327 );
not ( n4675 , n4628 );
and ( n4676 , n4675 , n3751 );
not ( n4677 , n3755 );
nor ( n4678 , n4676 , n4677 );
nor ( n4679 , n4674 , n4678 );
nand ( n4680 , n4673 , n4679 );
not ( n4681 , n4680 );
and ( n4682 , n4672 , n4681 );
not ( n4683 , n401 );
nand ( n4684 , n4683 , n1416 );
nor ( n4685 , n2030 , n4684 );
not ( n4686 , n4685 );
nor ( n4687 , n4682 , n4686 );
not ( n4688 , n4687 );
nor ( n4689 , n401 , n1483 );
or ( n4690 , n1042 , n4044 );
not ( n4691 , n1031 );
and ( n4692 , n4631 , n4039 );
or ( n4693 , n4691 , n4692 );
nand ( n4694 , n4690 , n4693 );
and ( n4695 , n4689 , n4694 );
or ( n4696 , n359 , n4135 , n4140 );
and ( n4697 , n373 , n4133 );
nand ( n4698 , n2537 , n3443 );
and ( n4699 , n4122 , n4698 );
and ( n4700 , n1708 , n3265 );
nor ( n4701 , n4699 , n4700 );
not ( n4702 , n4701 );
not ( n4703 , n1425 );
nand ( n4704 , n4702 , n4703 );
nand ( n4705 , n1427 , n4630 );
nand ( n4706 , n4679 , n4705 );
or ( n4707 , n1644 , n4706 );
or ( n4708 , n4701 , n388 );
nand ( n4709 , n766 , n1689 );
nand ( n4710 , n4628 , n4709 );
nand ( n4711 , n4708 , n4710 );
or ( n4712 , n344 , n4711 );
nand ( n4713 , n4707 , n4712 , n1661 );
and ( n4714 , n4704 , n4713 );
nor ( n4715 , n4714 , n373 );
nor ( n4716 , n4697 , n4715 );
or ( n4717 , n1655 , n4716 );
nor ( n4718 , n1644 , n373 );
and ( n4719 , n4718 , n4711 );
nand ( n4720 , n4138 , n4504 );
and ( n4721 , n373 , n4720 );
nor ( n4722 , n344 , n373 );
and ( n4723 , n4722 , n4706 );
nor ( n4724 , n4719 , n4721 , n4723 );
or ( n4725 , n1633 , n4724 );
nand ( n4726 , n4717 , n4725 , n359 );
and ( n4727 , n4696 , n4726 );
nor ( n4728 , n4695 , n4727 );
not ( n4729 , n1041 );
not ( n4730 , n4025 );
or ( n4731 , n4729 , n4730 );
or ( n4732 , n1489 , n4032 );
or ( n4733 , n4640 , n4027 );
nand ( n4734 , n1109 , n4648 );
nand ( n4735 , n4732 , n4733 , n4734 );
or ( n4736 , n1041 , n4735 );
nand ( n4737 , n4731 , n4736 );
nand ( n4738 , n4681 , n4737 );
and ( n4739 , n4689 , n4738 );
nand ( n4740 , n392 , n1707 );
nor ( n4741 , n394 , n4740 );
or ( n4742 , n4741 , n4130 );
nand ( n4743 , n4742 , n1041 );
not ( n4744 , n4706 );
and ( n4745 , n4743 , n4744 );
and ( n4746 , n1041 , n4130 );
nor ( n4747 , n398 , n403 );
or ( n4748 , n406 , n4747 );
not ( n4749 , n401 );
nand ( n4750 , n4748 , n4749 );
nand ( n4751 , n1626 , n4750 );
nor ( n4752 , n4746 , n4751 );
nor ( n4753 , n4745 , n4752 );
nor ( n4754 , n4739 , n4753 );
nor ( n4755 , n401 , n1425 );
nand ( n4756 , n1423 , n4755 );
not ( n4757 , n4756 );
nand ( n4758 , n372 , n4757 );
not ( n4759 , n4758 );
not ( n4760 , n358 );
not ( n4761 , n4048 );
nand ( n4762 , n4631 , n4761 );
and ( n4763 , n1031 , n4762 );
nor ( n4764 , n4763 , n4680 );
or ( n4765 , n4760 , n4764 );
not ( n4766 , n4631 );
not ( n4767 , n4059 );
or ( n4768 , n4766 , n4767 );
nand ( n4769 , n4768 , n953 );
nand ( n4770 , n4055 , n4734 , n4769 );
nand ( n4771 , n358 , n4770 );
and ( n4772 , n4649 , n4771 );
not ( n4773 , n358 );
not ( n4774 , n4773 );
not ( n4775 , n3868 );
or ( n4776 , n4774 , n4775 );
nand ( n4777 , n1260 , n3437 );
nand ( n4778 , n4776 , n4777 );
and ( n4779 , n3917 , n4778 );
nor ( n4780 , n1298 , n3981 );
nor ( n4781 , n4779 , n4780 );
nand ( n4782 , n4772 , n4781 );
not ( n4783 , n4782 );
not ( n4784 , n4631 );
not ( n4785 , n4022 );
or ( n4786 , n4784 , n4785 );
nand ( n4787 , n4786 , n1743 );
nand ( n4788 , n4783 , n4787 );
and ( n4789 , n4788 , n1042 );
and ( n4790 , n1041 , n4063 );
nor ( n4791 , n4789 , n4790 );
nand ( n4792 , n4765 , n4791 );
nand ( n4793 , n4759 , n4792 );
nand ( n4794 , n4688 , n4728 , n4754 , n4793 );
nand ( n4795 , n4619 , n4794 );
not ( n4796 , n2500 );
or ( n4797 , n1656 , n4701 );
not ( n4798 , n1662 );
and ( n4799 , n344 , n4798 );
and ( n4800 , n1644 , n1634 );
nor ( n4801 , n4799 , n4800 );
or ( n4802 , n4801 , n4744 );
nand ( n4803 , n344 , n1634 );
not ( n4804 , n4803 );
nor ( n4805 , n344 , n1662 );
or ( n4806 , n4804 , n4805 );
nand ( n4807 , n4806 , n4711 );
nand ( n4808 , n4797 , n4802 , n4807 );
and ( n4809 , n373 , n4808 );
or ( n4810 , n1026 , n3250 );
not ( n4811 , n4705 );
or ( n4812 , n791 , n2516 );
nand ( n4813 , n4812 , n4679 );
nor ( n4814 , n4811 , n4813 );
nand ( n4815 , n4810 , n4814 );
and ( n4816 , n4751 , n4815 );
nor ( n4817 , n4809 , n4816 );
or ( n4818 , n4796 , n4817 );
and ( n4819 , n2559 , n4140 );
not ( n4820 , n2566 );
nor ( n4821 , n4820 , n4724 );
nor ( n4822 , n2558 , n4136 );
nor ( n4823 , n4819 , n4821 , n4822 );
nand ( n4824 , n4618 , n4795 , n4818 , n4823 );
and ( n4825 , n373 , n4656 );
not ( n4826 , n373 );
and ( n4827 , n4826 , n4670 );
nor ( n4828 , n4825 , n4827 );
and ( n4829 , n1464 , n4828 );
or ( n4830 , n373 , n4064 );
nand ( n4831 , n4830 , n372 );
not ( n4832 , n4692 );
nand ( n4833 , n4832 , n1925 );
and ( n4834 , n1361 , n4762 );
not ( n4835 , n4735 );
and ( n4836 , n4787 , n4835 );
nor ( n4837 , n4836 , n358 );
nor ( n4838 , n4834 , n4782 , n4837 );
and ( n4839 , n4833 , n4838 );
nor ( n4840 , n4839 , n1019 );
nor ( n4841 , n4831 , n4840 );
nor ( n4842 , n4829 , n4841 );
or ( n4843 , n4842 , n4813 );
nand ( n4844 , n4843 , n4757 );
not ( n4845 , n4844 );
not ( n4846 , n4796 );
and ( n4847 , n4845 , n4846 );
not ( n4848 , n791 );
not ( n4849 , n2468 );
and ( n4850 , n4848 , n4849 );
not ( n4851 , n4679 );
nor ( n4852 , n4850 , n4851 );
or ( n4853 , n2453 , n4630 );
nand ( n4854 , n4853 , n3824 );
nand ( n4855 , n4852 , n4854 );
and ( n4856 , n2581 , n4855 );
nor ( n4857 , n4847 , n4856 );
nand ( n4858 , n389 , n395 );
not ( n4859 , n4858 );
nor ( n4860 , n714 , n716 );
not ( n4861 , n4860 );
not ( n4862 , n4861 );
or ( n4863 , n4859 , n4862 );
nand ( n4864 , n4863 , n4142 );
not ( n4865 , n4852 );
and ( n4866 , n2444 , n4656 );
not ( n4867 , n2444 );
and ( n4868 , n4867 , n4670 );
nor ( n4869 , n4866 , n4868 );
not ( n4870 , n4869 );
or ( n4871 , n4865 , n4870 );
nand ( n4872 , n4871 , n4685 );
not ( n4873 , n4852 );
nand ( n4874 , n4873 , n4689 );
or ( n4875 , n4838 , n2453 );
or ( n4876 , n2444 , n4064 );
not ( n4877 , n358 );
or ( n4878 , n4877 , n4852 );
nand ( n4879 , n4875 , n4876 , n4878 );
nand ( n4880 , n4759 , n4879 );
and ( n4881 , n2453 , n4130 );
or ( n4882 , n4758 , n2453 , n4833 );
and ( n4883 , n1040 , n4715 );
and ( n4884 , n2453 , n4133 );
nor ( n4885 , n4883 , n4884 );
or ( n4886 , n1655 , n4885 );
nand ( n4887 , n4882 , n4886 );
not ( n4888 , n4855 );
nor ( n4889 , n4888 , n4750 );
nor ( n4890 , n4881 , n4887 , n4889 );
nand ( n4891 , n4872 , n4874 , n4880 , n4890 );
nand ( n4892 , n2563 , n4891 );
nand ( n4893 , n4857 , n4864 , n4892 );
or ( n4894 , n4824 , n4893 );
nand ( n4895 , n4894 , n2981 );
not ( n4896 , n2996 );
not ( n4897 , n4077 );
nand ( n4898 , n4896 , n4897 );
not ( n4899 , n3005 );
not ( n4900 , n4365 );
and ( n4901 , n4899 , n4900 );
not ( n4902 , n4128 );
and ( n4903 , n2988 , n4902 );
nor ( n4904 , n4901 , n4903 );
and ( n4905 , n3007 , n4310 );
and ( n4906 , n3010 , n3888 );
not ( n4907 , n4122 );
or ( n4908 , n2989 , n4907 );
or ( n4909 , n791 , n2986 );
nand ( n4910 , n4908 , n4909 );
nor ( n4911 , n4905 , n4906 , n4910 );
nand ( n4912 , n4895 , n4898 , n4904 , n4911 );
nor ( n4913 , n4677 , n1029 );
nand ( n4914 , n413 , n997 );
not ( n4915 , n4914 );
not ( n4916 , n849 );
not ( n4917 , n4916 );
nor ( n4918 , n4915 , n4917 );
nor ( n4919 , n791 , n4918 );
nand ( n4920 , n402 , n4919 );
not ( n4921 , n392 );
not ( n4922 , n388 );
nand ( n4923 , n4922 , n390 , n386 );
nor ( n4924 , n4921 , n4923 );
not ( n4925 , n4924 );
not ( n4926 , n3029 );
and ( n4927 , n3021 , n4926 );
nand ( n4928 , n4927 , n4919 );
nand ( n4929 , n730 , n746 );
nand ( n4930 , n392 , n4929 );
or ( n4931 , n4914 , n4930 );
not ( n4932 , n407 );
not ( n4933 , n4916 );
not ( n4934 , n4933 );
or ( n4935 , n4932 , n4934 );
nand ( n4936 , n730 , n847 );
nand ( n4937 , n746 , n4936 );
nand ( n4938 , n4935 , n4937 );
nand ( n4939 , n392 , n4938 );
nand ( n4940 , n4928 , n4931 , n4939 );
nor ( n4941 , n4925 , n4940 );
nand ( n4942 , n4920 , n4941 );
and ( n4943 , n4913 , n4942 );
nand ( n4944 , n790 , n794 );
not ( n4945 , n4944 );
nand ( n4946 , n893 , n1056 );
not ( n4947 , n3297 );
not ( n4948 , n1207 );
nand ( n4949 , n402 , n4948 );
and ( n4950 , n4947 , n4949 );
not ( n4951 , n998 );
not ( n4952 , n4951 );
nand ( n4953 , n4952 , n1192 );
nand ( n4954 , n3030 , n4953 );
not ( n4955 , n4954 );
not ( n4956 , n847 );
not ( n4957 , n4956 );
nor ( n4958 , n407 , n417 );
not ( n4959 , n4958 );
nor ( n4960 , n4959 , n402 );
not ( n4961 , n4960 );
or ( n4962 , n4957 , n4961 );
not ( n4963 , n402 );
nand ( n4964 , n4963 , n731 );
nand ( n4965 , n4962 , n4964 );
nor ( n4966 , n1272 , n4965 );
not ( n4967 , n4966 );
or ( n4968 , n4955 , n4967 );
not ( n4969 , n399 );
nand ( n4970 , n4968 , n4969 );
not ( n4971 , n410 );
not ( n4972 , n1198 );
nand ( n4973 , n407 , n4953 );
nand ( n4974 , n4972 , n4973 );
not ( n4975 , n4974 );
and ( n4976 , n4970 , n4971 , n4975 );
nand ( n4977 , n4946 , n4950 , n4976 );
not ( n4978 , n4977 );
not ( n4979 , n4978 );
and ( n4980 , n4945 , n4979 );
nand ( n4981 , n392 , n402 );
not ( n4982 , n4981 );
nor ( n4983 , n999 , n4917 );
not ( n4984 , n4983 );
and ( n4985 , n4982 , n4984 );
not ( n4986 , n4983 );
not ( n4987 , n4986 );
nor ( n4988 , n791 , n399 );
not ( n4989 , n4988 );
not ( n4990 , n3030 );
or ( n4991 , n4989 , n4990 );
not ( n4992 , n407 );
nor ( n4993 , n4992 , n3129 );
nand ( n4994 , n392 , n4993 );
nand ( n4995 , n4991 , n4994 );
not ( n4996 , n4995 );
or ( n4997 , n4987 , n4996 );
nand ( n4998 , n4997 , n4939 );
nor ( n4999 , n4985 , n4998 );
not ( n5000 , n1093 );
not ( n5001 , n5000 );
not ( n5002 , n5001 );
not ( n5003 , n5002 );
not ( n5004 , n4953 );
and ( n5005 , n5003 , n5004 );
nand ( n5006 , n402 , n791 );
nor ( n5007 , n5005 , n5006 );
nand ( n5008 , n791 , n3130 , n4974 );
not ( n5009 , n1195 );
not ( n5010 , n4960 );
or ( n5011 , n5009 , n5010 );
nand ( n5012 , n5011 , n4964 );
not ( n5013 , n5012 );
not ( n5014 , n5013 );
not ( n5015 , n4954 );
or ( n5016 , n5014 , n5015 );
nor ( n5017 , n392 , n399 );
nand ( n5018 , n5016 , n5017 );
nand ( n5019 , n5008 , n5018 );
nor ( n5020 , n5007 , n5019 );
and ( n5021 , n4999 , n5020 );
not ( n5022 , n4923 );
not ( n5023 , n5022 );
not ( n5024 , n5023 );
buf ( n5025 , n5024 );
not ( n5026 , n5025 );
nor ( n5027 , n5021 , n5026 );
nor ( n5028 , n4980 , n5027 );
nor ( n5029 , n793 , n3242 );
nand ( n5030 , n402 , n5029 );
buf ( n5031 , n997 );
nor ( n5032 , n5031 , n4948 );
not ( n5033 , n5032 );
not ( n5034 , n388 );
nor ( n5035 , n5034 , n392 );
nand ( n5036 , n386 , n5035 );
nand ( n5037 , n956 , n5004 );
nor ( n5038 , n410 , n5037 );
nor ( n5039 , n5036 , n5038 );
and ( n5040 , n5033 , n5039 );
nand ( n5041 , n5029 , n984 );
or ( n5042 , n399 , n5041 );
nand ( n5043 , n5029 , n1117 );
nand ( n5044 , n5042 , n5043 );
nor ( n5045 , n5040 , n5044 );
nand ( n5046 , n5028 , n5030 , n5045 );
and ( n5047 , n1138 , n5046 );
not ( n5048 , n5003 );
nand ( n5049 , n4914 , n1192 );
nor ( n5050 , n410 , n5049 );
not ( n5051 , n5050 );
or ( n5052 , n5048 , n5051 );
nand ( n5053 , n5052 , n402 );
not ( n5054 , n410 );
not ( n5055 , n5049 );
or ( n5056 , n746 , n5055 );
nand ( n5057 , n5056 , n4972 );
not ( n5058 , n5057 );
nor ( n5059 , n3203 , n5050 );
not ( n5060 , n4966 );
or ( n5061 , n5059 , n5060 );
nand ( n5062 , n5061 , n399 );
nand ( n5063 , n5054 , n5058 , n5062 );
not ( n5064 , n5063 );
nand ( n5065 , n5053 , n5064 );
not ( n5066 , n5065 );
or ( n5067 , n4944 , n5066 );
not ( n5068 , n5036 );
not ( n5069 , n5050 );
and ( n5070 , n5068 , n5069 );
not ( n5071 , n399 );
or ( n5072 , n5071 , n5041 );
nand ( n5073 , n5072 , n5043 );
nor ( n5074 , n5070 , n5073 );
and ( n5075 , n5030 , n5074 );
nand ( n5076 , n5067 , n5075 );
not ( n5077 , n5002 );
not ( n5078 , n5077 );
not ( n5079 , n5055 );
or ( n5080 , n5078 , n5079 );
not ( n5081 , n5006 );
nand ( n5082 , n5080 , n5081 );
not ( n5083 , n399 );
and ( n5084 , n3030 , n5049 );
nor ( n5085 , n5084 , n5012 );
or ( n5086 , n5083 , n392 , n5085 );
nor ( n5087 , n392 , n3021 );
nand ( n5088 , n5087 , n5057 );
nand ( n5089 , n5086 , n5088 );
nor ( n5090 , n4940 , n5089 );
and ( n5091 , n4920 , n5082 , n5090 );
nor ( n5092 , n5091 , n5026 );
nor ( n5093 , n5076 , n5092 );
or ( n5094 , n1014 , n5093 );
and ( n5095 , n416 , n5081 );
not ( n5096 , n1199 );
nand ( n5097 , n791 , n5096 );
not ( n5098 , n5097 );
nor ( n5099 , n5095 , n5098 );
or ( n5100 , n265 , n5099 );
not ( n5101 , n416 );
nor ( n5102 , n5101 , n4981 );
not ( n5103 , n4939 );
nor ( n5104 , n5102 , n5103 );
or ( n5105 , n4677 , n5104 );
nand ( n5106 , n390 , n767 );
nor ( n5107 , n793 , n5106 );
nand ( n5108 , n281 , n5107 );
or ( n5109 , n281 , n4924 );
nand ( n5110 , n5109 , n265 );
nand ( n5111 , n5108 , n5110 );
nand ( n5112 , n5100 , n5105 , n5111 );
nand ( n5113 , n2849 , n5112 );
not ( n5114 , n4925 );
not ( n5115 , n5114 );
not ( n5116 , n4999 );
or ( n5117 , n5115 , n5116 );
nor ( n5118 , n4677 , n1136 );
nand ( n5119 , n5117 , n5118 );
not ( n5120 , n5108 );
not ( n5121 , n5120 );
not ( n5122 , n5121 );
not ( n5123 , n5122 );
not ( n5124 , n5020 );
or ( n5125 , n5123 , n5124 );
nor ( n5126 , n265 , n1136 );
nand ( n5127 , n5125 , n5126 );
and ( n5128 , n5113 , n5119 , n5127 );
nand ( n5129 , n5094 , n5128 );
nor ( n5130 , n4943 , n5047 , n5129 );
or ( n5131 , n1760 , n5130 );
not ( n5132 , n358 );
and ( n5133 , n793 , n1021 );
not ( n5134 , n5120 );
not ( n5135 , n5134 );
not ( n5136 , n5135 );
not ( n5137 , n5136 );
not ( n5138 , n5031 );
not ( n5139 , n5138 );
nor ( n5140 , n3095 , n402 );
nor ( n5141 , n392 , n5140 );
not ( n5142 , n5141 );
or ( n5143 , n5139 , n5142 );
not ( n5144 , n851 );
and ( n5145 , n5144 , n1192 );
not ( n5146 , n5141 );
nor ( n5147 , n5145 , n5146 );
nor ( n5148 , n5147 , n5098 );
nand ( n5149 , n5143 , n5148 );
not ( n5150 , n5149 );
and ( n5151 , n5137 , n5150 );
nor ( n5152 , n265 , n311 );
not ( n5153 , n5152 );
nor ( n5154 , n5151 , n5153 );
or ( n5155 , n5133 , n5154 );
nand ( n5156 , n2916 , n5155 );
not ( n5157 , n5137 );
not ( n5158 , n5007 );
not ( n5159 , n5000 );
not ( n5160 , n5159 );
nand ( n5161 , n956 , n1192 );
not ( n5162 , n5161 );
not ( n5163 , n5162 );
or ( n5164 , n5160 , n5163 );
nand ( n5165 , n5164 , n5081 );
not ( n5166 , n742 );
not ( n5167 , n5017 );
or ( n5168 , n5166 , n5167 );
not ( n5169 , n407 );
nor ( n5170 , n5169 , n392 );
not ( n5171 , n5170 );
nand ( n5172 , n5168 , n5171 );
nand ( n5173 , n5172 , n5037 );
and ( n5174 , n5097 , n5173 );
nand ( n5175 , n5158 , n5165 , n5174 );
or ( n5176 , n5157 , n5175 );
nand ( n5177 , n5176 , n5126 );
not ( n5178 , n4960 );
not ( n5179 , n5178 );
not ( n5180 , n921 );
nand ( n5181 , n5180 , n870 );
not ( n5182 , n5181 );
or ( n5183 , n5179 , n5182 );
or ( n5184 , n5031 , n4917 );
nand ( n5185 , n5184 , n5178 );
nand ( n5186 , n4937 , n5185 );
nor ( n5187 , n905 , n5186 );
nand ( n5188 , n5183 , n5187 );
not ( n5189 , n5188 );
or ( n5190 , n4944 , n5189 );
not ( n5191 , n4965 );
or ( n5192 , n410 , n3297 , n921 );
or ( n5193 , n402 , n3030 );
nand ( n5194 , n5192 , n5193 );
and ( n5195 , n5191 , n5194 );
nor ( n5196 , n5195 , n791 );
not ( n5197 , n414 );
and ( n5198 , n791 , n5178 );
not ( n5199 , n5198 );
or ( n5200 , n5197 , n5199 );
and ( n5201 , n5138 , n1192 );
not ( n5202 , n5198 );
nor ( n5203 , n5201 , n5202 );
nor ( n5204 , n5203 , n5098 );
nand ( n5205 , n5200 , n5204 );
or ( n5206 , n5196 , n5205 );
not ( n5207 , n5023 );
nand ( n5208 , n5206 , n5207 );
nand ( n5209 , n5190 , n5208 );
and ( n5210 , n5068 , n5181 );
not ( n5211 , n5030 );
not ( n5212 , n5041 );
nor ( n5213 , n5211 , n5212 );
not ( n5214 , n5213 );
or ( n5215 , n5209 , n5210 , n5214 );
nand ( n5216 , n5215 , n1404 );
nand ( n5217 , n5177 , n5216 );
not ( n5218 , n5217 );
nand ( n5219 , n5068 , n1210 );
and ( n5220 , n5219 , n5075 );
not ( n5221 , n4944 );
nand ( n5222 , n1211 , n5062 );
not ( n5223 , n5222 );
not ( n5224 , n402 );
not ( n5225 , n5224 );
and ( n5226 , n4914 , n5162 );
nor ( n5227 , n407 , n4927 );
nor ( n5228 , n5226 , n5227 );
not ( n5229 , n5228 );
not ( n5230 , n5063 );
nand ( n5231 , n5229 , n5230 );
not ( n5232 , n5231 );
or ( n5233 , n5225 , n5232 );
nand ( n5234 , n5233 , n5053 );
not ( n5235 , n5234 );
nand ( n5236 , n5223 , n5235 );
and ( n5237 , n5221 , n5236 );
and ( n5238 , n956 , n4918 );
not ( n5239 , n402 );
and ( n5240 , n5239 , n5227 );
nor ( n5241 , n5238 , n5240 );
and ( n5242 , n392 , n5241 );
nor ( n5243 , n5242 , n5103 );
nand ( n5244 , n5198 , n5228 );
not ( n5245 , n5096 );
nand ( n5246 , n1204 , n5245 );
nand ( n5247 , n876 , n5246 );
and ( n5248 , n5165 , n5247 );
and ( n5249 , n5082 , n5244 , n5248 );
and ( n5250 , n5243 , n5249 );
not ( n5251 , n5025 );
nor ( n5252 , n5250 , n5251 );
nor ( n5253 , n5237 , n5252 );
and ( n5254 , n5220 , n5253 );
nor ( n5255 , n5254 , n1014 );
not ( n5256 , n5114 );
not ( n5257 , n5256 );
and ( n5258 , n5257 , n5243 );
not ( n5259 , n4913 );
nor ( n5260 , n5258 , n5259 );
and ( n5261 , n5137 , n5249 );
or ( n5262 , n24 , n265 );
or ( n5263 , n1350 , n5262 );
nor ( n5264 , n5261 , n5263 );
nor ( n5265 , n5260 , n5264 );
not ( n5266 , n5257 );
nand ( n5267 , n414 , n4995 );
nand ( n5268 , n392 , n414 );
not ( n5269 , n5268 );
not ( n5270 , n5104 );
or ( n5271 , n5269 , n5270 );
nand ( n5272 , n5271 , n402 );
nand ( n5273 , n4999 , n5267 , n5272 );
not ( n5274 , n5273 );
not ( n5275 , n5274 );
or ( n5276 , n5266 , n5275 );
nand ( n5277 , n5276 , n5118 );
nor ( n5278 , n5039 , n5044 );
and ( n5279 , n5030 , n5278 );
not ( n5280 , n402 );
not ( n5281 , n5037 );
nor ( n5282 , n5280 , n5281 );
not ( n5283 , n5282 );
buf ( n5284 , n1200 );
not ( n5285 , n5284 );
and ( n5286 , n1204 , n5285 );
not ( n5287 , n399 );
or ( n5288 , n3203 , n5038 );
not ( n5289 , n5060 );
nand ( n5290 , n5288 , n5289 );
and ( n5291 , n5287 , n5290 );
not ( n5292 , n4973 );
nor ( n5293 , n5291 , n5292 );
nand ( n5294 , n5286 , n5293 );
not ( n5295 , n5294 );
nand ( n5296 , n5283 , n5295 );
nand ( n5297 , n5221 , n5296 );
or ( n5298 , n5175 , n5273 );
not ( n5299 , n5024 );
not ( n5300 , n5299 );
nand ( n5301 , n5298 , n5300 );
nand ( n5302 , n5279 , n5297 , n5301 );
nand ( n5303 , n1138 , n5302 );
nand ( n5304 , n5265 , n5277 , n5303 );
nor ( n5305 , n5255 , n5304 );
and ( n5306 , n5156 , n5218 , n5305 );
nand ( n5307 , n5133 , n2844 );
not ( n5308 , n311 );
nand ( n5309 , n1192 , n1083 );
not ( n5310 , n5309 );
nand ( n5311 , n5001 , n5310 );
nand ( n5312 , n5081 , n5311 );
not ( n5313 , n956 );
not ( n5314 , n5310 );
or ( n5315 , n5313 , n5314 );
not ( n5316 , n399 );
not ( n5317 , n810 );
or ( n5318 , n5316 , n5317 );
nand ( n5319 , n5318 , n746 );
nand ( n5320 , n5315 , n5319 );
nand ( n5321 , n5245 , n5320 );
nand ( n5322 , n791 , n5321 );
nand ( n5323 , n5312 , n5165 , n5322 );
not ( n5324 , n5323 );
and ( n5325 , n5137 , n5324 );
nor ( n5326 , n5325 , n265 );
and ( n5327 , n5308 , n5326 );
not ( n5328 , n4917 );
nand ( n5329 , n5328 , n1083 );
not ( n5330 , n5329 );
nand ( n5331 , n956 , n5330 );
not ( n5332 , n5331 );
or ( n5333 , n4981 , n5332 );
and ( n5334 , n392 , n5319 );
nand ( n5335 , n5334 , n5331 );
and ( n5336 , n4939 , n5335 );
nand ( n5337 , n5333 , n5336 );
and ( n5338 , n2255 , n5337 );
nor ( n5339 , n5327 , n5338 );
not ( n5340 , n793 );
nand ( n5341 , n390 , n3072 );
and ( n5342 , n2763 , n5341 );
not ( n5343 , n5342 );
and ( n5344 , n5340 , n5343 );
nor ( n5345 , n5344 , n2253 );
not ( n5346 , n5345 );
nand ( n5347 , n5029 , n914 );
not ( n5348 , n5347 );
and ( n5349 , n399 , n5348 );
not ( n5350 , n3704 );
nand ( n5351 , n5068 , n1088 );
or ( n5352 , n5350 , n5351 );
nand ( n5353 , n5352 , n5043 );
nor ( n5354 , n5349 , n5353 );
and ( n5355 , n5030 , n5354 );
or ( n5356 , n5337 , n5323 );
nand ( n5357 , n5356 , n5025 );
and ( n5358 , n5355 , n5357 );
not ( n5359 , n3086 );
not ( n5360 , n3704 );
or ( n5361 , n5359 , n5360 );
nand ( n5362 , n5284 , n3093 );
nand ( n5363 , n5361 , n5362 );
and ( n5364 , n399 , n5363 );
nand ( n5365 , n904 , n4937 );
not ( n5366 , n5365 );
and ( n5367 , n5366 , n3705 );
nor ( n5368 , n5367 , n3023 );
nor ( n5369 , n5364 , n5368 );
or ( n5370 , n402 , n5369 );
nand ( n5371 , n4950 , n3485 );
not ( n5372 , n5371 );
and ( n5373 , n1211 , n5372 );
nand ( n5374 , n5370 , n5373 );
nand ( n5375 , n5221 , n5374 );
nand ( n5376 , n5358 , n5219 , n5375 );
nand ( n5377 , n2727 , n5376 );
nand ( n5378 , n5339 , n5346 , n5377 );
nand ( n5379 , n948 , n5378 );
nand ( n5380 , n5306 , n5307 , n5379 );
nand ( n5381 , n5132 , n5380 );
not ( n5382 , n5346 );
not ( n5383 , n2254 );
not ( n5384 , n413 );
nand ( n5385 , n5384 , n803 );
nand ( n5386 , n5385 , n4916 );
or ( n5387 , n5000 , n5386 );
not ( n5388 , n4981 );
nand ( n5389 , n5387 , n5388 );
not ( n5390 , n5389 );
not ( n5391 , n5386 );
not ( n5392 , n4988 );
not ( n5393 , n3086 );
or ( n5394 , n5392 , n5393 );
nand ( n5395 , n5394 , n4994 );
not ( n5396 , n5395 );
or ( n5397 , n5391 , n5396 );
nand ( n5398 , n5397 , n4939 );
nor ( n5399 , n5390 , n5398 );
not ( n5400 , n5399 );
and ( n5401 , n5383 , n5400 );
not ( n5402 , n311 );
not ( n5403 , n1695 );
not ( n5404 , n3086 );
not ( n5405 , n1089 );
not ( n5406 , n5405 );
or ( n5407 , n5404 , n5406 );
nand ( n5408 , n5407 , n5362 );
not ( n5409 , n5408 );
not ( n5410 , n5386 );
nor ( n5411 , n409 , n413 );
nor ( n5412 , n5411 , n5161 );
nand ( n5413 , n5410 , n5412 );
nand ( n5414 , n3086 , n5413 );
not ( n5415 , n5414 );
not ( n5416 , n5362 );
or ( n5417 , n5415 , n5416 );
not ( n5418 , n399 );
nand ( n5419 , n5417 , n5418 );
not ( n5420 , n5419 );
not ( n5421 , n5420 );
or ( n5422 , n5409 , n5421 );
not ( n5423 , n4993 );
not ( n5424 , n410 );
not ( n5425 , n5385 );
nor ( n5426 , n5425 , n1191 );
and ( n5427 , n5424 , n5426 );
or ( n5428 , n5423 , n5427 );
nand ( n5429 , n3130 , n5365 );
nand ( n5430 , n5428 , n5429 );
not ( n5431 , n5430 );
nand ( n5432 , n5422 , n5431 );
nor ( n5433 , n1937 , n5432 );
or ( n5434 , n4944 , n5433 );
or ( n5435 , n5036 , n5427 );
or ( n5436 , n399 , n5347 );
nand ( n5437 , n5436 , n5043 );
not ( n5438 , n5437 );
nand ( n5439 , n5435 , n5438 );
or ( n5440 , n5006 , n5426 );
not ( n5441 , n5440 );
and ( n5442 , n5017 , n810 );
nor ( n5443 , n5442 , n5170 );
or ( n5444 , n5443 , n5426 );
nand ( n5445 , n5444 , n5097 );
nor ( n5446 , n5441 , n5445 );
and ( n5447 , n5446 , n5399 );
nor ( n5448 , n5447 , n5299 );
nor ( n5449 , n5439 , n5448 );
nand ( n5450 , n5434 , n5449 , n5030 );
not ( n5451 , n5450 );
or ( n5452 , n5403 , n5451 );
not ( n5453 , n5157 );
not ( n5454 , n5453 );
not ( n5455 , n5446 );
or ( n5456 , n5454 , n5455 );
nand ( n5457 , n5456 , n2251 );
nand ( n5458 , n5452 , n5457 );
and ( n5459 , n5402 , n5458 );
nor ( n5460 , n5401 , n5459 );
not ( n5461 , n5460 );
or ( n5462 , n5382 , n5461 );
nand ( n5463 , n5462 , n3998 );
not ( n5464 , n3729 );
not ( n5465 , n4956 );
nand ( n5466 , n5465 , n1300 );
nand ( n5467 , n392 , n5466 );
and ( n5468 , n921 , n5467 );
nand ( n5469 , n5466 , n5196 );
nand ( n5470 , n5114 , n5469 );
nor ( n5471 , n5468 , n5470 );
or ( n5472 , n4677 , n5471 );
not ( n5473 , n5121 );
not ( n5474 , n5473 );
or ( n5475 , n5474 , n5205 );
nand ( n5476 , n5475 , n2251 );
nand ( n5477 , n5472 , n5476 );
not ( n5478 , n5477 );
or ( n5479 , n5464 , n5478 );
not ( n5480 , n1945 );
not ( n5481 , n4938 );
nand ( n5482 , n1204 , n5481 );
and ( n5483 , n392 , n5482 );
not ( n5484 , n5272 );
nor ( n5485 , n5483 , n5484 );
or ( n5486 , n4677 , n5485 );
or ( n5487 , n265 , n5248 );
nand ( n5488 , n5486 , n5487 , n5111 );
and ( n5489 , n5480 , n5488 );
nor ( n5490 , n5489 , n372 );
nand ( n5491 , n5479 , n5490 );
and ( n5492 , n413 , n956 );
nand ( n5493 , n5492 , n4918 );
and ( n5494 , n5395 , n3176 , n5493 );
nor ( n5495 , n5103 , n5494 );
not ( n5496 , n5495 );
nand ( n5497 , n5496 , n4981 );
nand ( n5498 , n5497 , n5389 , n5272 );
and ( n5499 , n2255 , n5498 );
not ( n5500 , n311 );
not ( n5501 , n5443 );
not ( n5502 , n5412 );
and ( n5503 , n5501 , n5502 );
nor ( n5504 , n5503 , n5098 );
and ( n5505 , n5165 , n5440 , n5504 );
and ( n5506 , n5137 , n5505 );
nor ( n5507 , n5506 , n265 );
and ( n5508 , n5500 , n5507 );
nor ( n5509 , n5499 , n5508 );
not ( n5510 , n2726 );
not ( n5511 , n5498 );
and ( n5512 , n5505 , n5511 );
nor ( n5513 , n5512 , n5026 );
nor ( n5514 , n5211 , n5513 );
and ( n5515 , n5068 , n5413 );
nor ( n5516 , n5515 , n5437 );
not ( n5517 , n5413 );
nor ( n5518 , n5423 , n5517 );
not ( n5519 , n5518 );
nand ( n5520 , n5519 , n5429 , n5419 );
not ( n5521 , n5520 );
nand ( n5522 , n402 , n5502 );
nand ( n5523 , n5521 , n5522 );
nand ( n5524 , n5221 , n5523 );
nand ( n5525 , n5514 , n5516 , n5524 );
and ( n5526 , n5510 , n5525 );
nor ( n5527 , n5526 , n5345 );
and ( n5528 , n5509 , n5527 );
nor ( n5529 , n5528 , n1377 );
nor ( n5530 , n5491 , n5529 );
and ( n5531 , n1211 , n5286 );
or ( n5532 , n4944 , n5531 );
nand ( n5533 , n5532 , n5030 );
nand ( n5534 , n5043 , n5219 );
and ( n5535 , n5248 , n5485 );
not ( n5536 , n5300 );
nor ( n5537 , n5535 , n5536 );
nor ( n5538 , n5533 , n5534 , n5537 );
nor ( n5539 , n1946 , n5538 );
not ( n5540 , n5221 );
not ( n5541 , n5187 );
nand ( n5542 , n1093 , n5032 );
not ( n5543 , n984 );
nand ( n5544 , n5465 , n5543 );
and ( n5545 , n5542 , n5544 );
or ( n5546 , n5541 , n5545 );
not ( n5547 , n5546 );
or ( n5548 , n5540 , n5547 );
nand ( n5549 , n5548 , n5213 );
and ( n5550 , n1486 , n5549 );
not ( n5551 , n64 );
nand ( n5552 , n5551 , n1028 );
not ( n5553 , n5552 );
nand ( n5554 , n3755 , n5553 );
nand ( n5555 , n5022 , n1338 );
and ( n5556 , n5554 , n5555 );
not ( n5557 , n5186 );
nor ( n5558 , n5556 , n5557 );
and ( n5559 , n392 , n5558 );
nor ( n5560 , n5550 , n5559 );
or ( n5561 , n5552 , n5111 );
nand ( n5562 , n5068 , n1338 , n5033 );
nand ( n5563 , n5561 , n5562 );
not ( n5564 , n5563 );
or ( n5565 , n1251 , n5262 );
nand ( n5566 , n5565 , n5555 );
not ( n5567 , n5204 );
nand ( n5568 , n5566 , n5567 );
nand ( n5569 , n5560 , n5564 , n5568 );
not ( n5570 , n5569 );
not ( n5571 , n1096 );
nor ( n5572 , n5571 , n5408 );
not ( n5573 , n5572 );
and ( n5574 , n5221 , n5573 );
and ( n5575 , n5347 , n5351 );
and ( n5576 , n5030 , n5575 );
not ( n5577 , n853 );
or ( n5578 , n5140 , n5577 );
nand ( n5579 , n5578 , n4937 );
nand ( n5580 , n392 , n5579 );
not ( n5581 , n5580 );
not ( n5582 , n5148 );
or ( n5583 , n5581 , n5582 );
not ( n5584 , n5023 );
nand ( n5585 , n5583 , n5584 );
nand ( n5586 , n5576 , n5585 );
nor ( n5587 , n5574 , n5586 );
or ( n5588 , n2725 , n5587 );
nor ( n5589 , n2254 , n5580 );
nor ( n5590 , n5345 , n5589 );
not ( n5591 , n5153 );
nand ( n5592 , n5135 , n5148 );
nand ( n5593 , n5591 , n5592 );
nand ( n5594 , n5588 , n5590 , n5593 );
nand ( n5595 , n2914 , n5594 );
not ( n5596 , n5355 );
nand ( n5597 , n5319 , n1084 );
not ( n5598 , n5284 );
nand ( n5599 , n5597 , n5598 );
nor ( n5600 , n5599 , n5371 );
nor ( n5601 , n4944 , n5600 );
nand ( n5602 , n5388 , n5329 );
nand ( n5603 , n5334 , n5329 );
and ( n5604 , n4939 , n5603 );
and ( n5605 , n5602 , n5604 );
not ( n5606 , n5312 );
not ( n5607 , n5087 );
not ( n5608 , n407 );
not ( n5609 , n5309 );
or ( n5610 , n5608 , n5609 );
nand ( n5611 , n5610 , n4972 );
not ( n5612 , n5611 );
or ( n5613 , n5607 , n5612 );
not ( n5614 , n1195 );
and ( n5615 , n5614 , n3046 );
not ( n5616 , n399 );
nor ( n5617 , n5615 , n5616 );
nand ( n5618 , n5617 , n876 , n5311 );
nand ( n5619 , n5613 , n5618 );
nor ( n5620 , n5606 , n5619 );
and ( n5621 , n5605 , n5620 );
nor ( n5622 , n5621 , n5299 );
nor ( n5623 , n5596 , n5601 , n5622 );
or ( n5624 , n2725 , n5623 );
not ( n5625 , n2254 );
not ( n5626 , n5605 );
and ( n5627 , n5625 , n5626 );
not ( n5628 , n311 );
and ( n5629 , n5620 , n5135 );
nor ( n5630 , n5629 , n265 );
and ( n5631 , n5628 , n5630 );
nor ( n5632 , n5627 , n5631 );
nand ( n5633 , n5624 , n5632 , n5346 );
nand ( n5634 , n948 , n5633 );
nand ( n5635 , n5570 , n5307 , n5595 , n5634 );
and ( n5636 , n358 , n5635 );
nor ( n5637 , n5121 , n5089 );
and ( n5638 , n5082 , n5637 );
nor ( n5639 , n5638 , n265 , n2933 );
nand ( n5640 , n5104 , n5099 );
and ( n5641 , n5025 , n5640 );
nand ( n5642 , n4949 , n5598 );
and ( n5643 , n5221 , n5642 );
nor ( n5644 , n5641 , n5643 );
and ( n5645 , n5068 , n4948 );
not ( n5646 , n5043 );
nor ( n5647 , n5645 , n5646 );
and ( n5648 , n5644 , n5030 , n5647 );
nor ( n5649 , n5648 , n1298 );
or ( n5650 , n5639 , n5649 );
nor ( n5651 , n5636 , n5650 );
or ( n5652 , n372 , n5651 );
not ( n5653 , n3176 );
and ( n5654 , n1093 , n5653 );
nor ( n5655 , n5654 , n791 );
nand ( n5656 , n402 , n5655 );
nand ( n5657 , n4924 , n5656 );
not ( n5658 , n5657 );
not ( n5659 , n3096 );
not ( n5660 , n4936 );
not ( n5661 , n5660 );
or ( n5662 , n5659 , n5661 );
nand ( n5663 , n5662 , n5655 );
and ( n5664 , n5658 , n5663 );
nor ( n5665 , n5664 , n2254 );
and ( n5666 , n5656 , n5150 );
nor ( n5667 , n5666 , n5299 );
or ( n5668 , n5657 , n5663 );
or ( n5669 , n5140 , n3146 );
nand ( n5670 , n5669 , n5285 );
not ( n5671 , n5670 );
or ( n5672 , n4944 , n5671 );
and ( n5673 , n5219 , n5576 );
nand ( n5674 , n5668 , n5672 , n5673 );
nor ( n5675 , n5667 , n5674 );
nor ( n5676 , n2726 , n5675 );
or ( n5677 , n5665 , n5676 );
nand ( n5678 , n5677 , n3384 );
nand ( n5679 , n5652 , n5678 );
nor ( n5680 , n5539 , n5679 );
nand ( n5681 , n5381 , n5463 , n5530 , n5680 );
not ( n5682 , n311 );
not ( n5683 , n1300 );
and ( n5684 , n5683 , n5149 );
nor ( n5685 , n4929 , n5614 );
nand ( n5686 , n5081 , n5685 );
not ( n5687 , n5686 );
nor ( n5688 , n5684 , n5687 );
and ( n5689 , n5688 , n5473 );
nor ( n5690 , n5689 , n265 );
and ( n5691 , n5682 , n5690 );
not ( n5692 , n5466 );
nor ( n5693 , n5692 , n5663 );
and ( n5694 , n2255 , n5693 );
nor ( n5695 , n5691 , n5694 );
and ( n5696 , n5219 , n5575 );
not ( n5697 , n5693 );
nand ( n5698 , n5697 , n5688 );
nand ( n5699 , n5300 , n5698 );
not ( n5700 , n5683 );
not ( n5701 , n5670 );
or ( n5702 , n5700 , n5701 );
not ( n5703 , n781 );
nand ( n5704 , n5703 , n727 );
buf ( n5705 , n5704 );
and ( n5706 , n1300 , n5705 );
nor ( n5707 , n5706 , n5408 );
nand ( n5708 , n5702 , n5707 );
nand ( n5709 , n5221 , n5708 );
nand ( n5710 , n5696 , n5699 , n5709 );
nand ( n5711 , n2727 , n5710 );
nand ( n5712 , n5695 , n5346 , n5711 );
and ( n5713 , n3384 , n5712 );
not ( n5714 , n5286 );
and ( n5715 , n5221 , n5714 );
nor ( n5716 , n5715 , n5534 );
and ( n5717 , n5107 , n5246 );
and ( n5718 , n5257 , n5482 );
nor ( n5719 , n5717 , n5718 );
nand ( n5720 , n5716 , n5719 );
and ( n5721 , n1947 , n5720 );
nor ( n5722 , n5713 , n5721 );
not ( n5723 , n2254 );
not ( n5724 , n5495 );
and ( n5725 , n5723 , n5724 );
not ( n5726 , n311 );
and ( n5727 , n5221 , n5520 );
not ( n5728 , n5504 );
not ( n5729 , n5495 );
or ( n5730 , n5728 , n5729 );
nand ( n5731 , n5730 , n5207 );
nand ( n5732 , n5516 , n5731 );
nor ( n5733 , n5727 , n5732 );
or ( n5734 , n5733 , n1631 );
and ( n5735 , n5473 , n5504 );
or ( n5736 , n265 , n5735 );
nand ( n5737 , n5734 , n5736 );
and ( n5738 , n5726 , n5737 );
nor ( n5739 , n5725 , n5738 );
and ( n5740 , n5346 , n5739 );
nor ( n5741 , n5740 , n1377 );
not ( n5742 , n5741 );
and ( n5743 , n5722 , n372 , n5742 );
not ( n5744 , n948 );
or ( n5745 , n2254 , n5604 );
not ( n5746 , n311 );
nand ( n5747 , n5221 , n5599 );
not ( n5748 , n5604 );
or ( n5749 , n5748 , n5619 );
nand ( n5750 , n5749 , n5584 );
and ( n5751 , n5747 , n5354 , n5750 );
or ( n5752 , n1659 , n5751 );
not ( n5753 , n5120 );
or ( n5754 , n5753 , n5619 );
nand ( n5755 , n5754 , n2251 );
nand ( n5756 , n5752 , n5755 );
and ( n5757 , n5746 , n5756 );
nor ( n5758 , n5757 , n5345 );
nand ( n5759 , n5745 , n5758 );
not ( n5760 , n5759 );
or ( n5761 , n5744 , n5760 );
not ( n5762 , n4929 );
not ( n5763 , n5762 );
not ( n5764 , n5763 );
not ( n5765 , n5571 );
or ( n5766 , n5764 , n5765 );
nand ( n5767 , n5766 , n5707 );
nand ( n5768 , n5221 , n5767 );
not ( n5769 , n5585 );
nand ( n5770 , n5467 , n5688 );
nand ( n5771 , n5769 , n5770 );
nand ( n5772 , n5768 , n5575 , n5771 );
and ( n5773 , n1660 , n5772 );
and ( n5774 , n5592 , n5690 );
nor ( n5775 , n5773 , n5774 );
or ( n5776 , n311 , n5775 );
nand ( n5777 , n5466 , n5589 );
nand ( n5778 , n5776 , n5346 , n5777 );
nand ( n5779 , n3899 , n5778 );
nand ( n5780 , n5761 , n5779 );
and ( n5781 , n5221 , n5432 );
not ( n5782 , n5439 );
or ( n5783 , n5445 , n5398 );
nand ( n5784 , n5783 , n5024 );
nand ( n5785 , n5782 , n5784 );
nor ( n5786 , n5781 , n5785 );
or ( n5787 , n2726 , n5786 );
or ( n5788 , n5121 , n5445 );
nand ( n5789 , n5788 , n5152 );
and ( n5790 , n5346 , n5789 );
nand ( n5791 , n2255 , n5398 );
nand ( n5792 , n5787 , n5790 , n5791 );
and ( n5793 , n1135 , n5792 );
not ( n5794 , n358 );
nor ( n5795 , n5793 , n5794 );
not ( n5796 , n5598 );
not ( n5797 , n5796 );
or ( n5798 , n4944 , n5797 );
or ( n5799 , n5103 , n5098 );
not ( n5800 , n5026 );
nand ( n5801 , n5799 , n5800 );
nand ( n5802 , n5798 , n5647 , n5801 );
and ( n5803 , n1218 , n5802 );
or ( n5804 , n5263 , n5637 );
not ( n5805 , n2843 );
not ( n5806 , n5805 );
not ( n5807 , n4941 );
nand ( n5808 , n2763 , n5807 );
nor ( n5809 , n5806 , n5808 );
not ( n5810 , n5545 );
or ( n5811 , n4944 , n5810 );
nand ( n5812 , n5811 , n5041 );
and ( n5813 , n1400 , n5812 );
nor ( n5814 , n5813 , n5563 );
not ( n5815 , n5467 );
nand ( n5816 , n5815 , n5558 );
not ( n5817 , n5568 );
not ( n5818 , n5683 );
not ( n5819 , n5205 );
or ( n5820 , n5818 , n5819 );
nand ( n5821 , n5820 , n5686 );
nand ( n5822 , n5817 , n5821 );
nand ( n5823 , n5814 , n5816 , n5822 );
nor ( n5824 , n5809 , n5823 );
nand ( n5825 , n5804 , n5824 );
nor ( n5826 , n5803 , n5825 );
not ( n5827 , n4976 );
nand ( n5828 , n5221 , n5827 );
or ( n5829 , n4998 , n5019 );
nand ( n5830 , n5829 , n5207 );
nand ( n5831 , n5828 , n5045 , n5830 );
and ( n5832 , n1959 , n5831 );
not ( n5833 , n4924 );
or ( n5834 , n5833 , n4998 );
nand ( n5835 , n5834 , n3755 );
or ( n5836 , n5134 , n5019 );
nand ( n5837 , n5836 , n2251 );
nand ( n5838 , n5835 , n5837 );
nor ( n5839 , n5832 , n5838 );
or ( n5840 , n1136 , n5839 );
or ( n5841 , n5299 , n5090 );
or ( n5842 , n4944 , n5064 );
nand ( n5843 , n5841 , n5842 , n5074 );
nand ( n5844 , n1013 , n5843 );
nand ( n5845 , n5840 , n5844 );
and ( n5846 , n3755 , n5103 );
or ( n5847 , n265 , n5245 );
nand ( n5848 , n5847 , n5111 );
nor ( n5849 , n5846 , n5848 );
nor ( n5850 , n1775 , n5849 );
nor ( n5851 , n5845 , n5850 , n5823 );
nand ( n5852 , n5795 , n5826 , n5307 , n5851 );
or ( n5853 , n5780 , n5852 );
not ( n5854 , n358 );
nand ( n5855 , n3755 , n5470 );
or ( n5856 , n5136 , n5821 );
nand ( n5857 , n5856 , n2251 );
and ( n5858 , n5855 , n5857 );
nor ( n5859 , n5212 , n5210 );
nand ( n5860 , n5544 , n5188 );
not ( n5861 , n5860 );
nand ( n5862 , n5221 , n5861 );
not ( n5863 , n5469 );
or ( n5864 , n5863 , n5821 );
nand ( n5865 , n5864 , n5025 );
nand ( n5866 , n5859 , n5862 , n5865 );
nand ( n5867 , n1660 , n5866 );
and ( n5868 , n5858 , n5867 );
nor ( n5869 , n5868 , n5552 );
not ( n5870 , n5231 );
or ( n5871 , n4944 , n5870 );
and ( n5872 , n5219 , n5074 );
nand ( n5873 , n5097 , n5244 );
nor ( n5874 , n5467 , n5243 );
or ( n5875 , n5873 , n5874 );
nand ( n5876 , n5875 , n5207 );
nand ( n5877 , n5871 , n5872 , n5876 );
nand ( n5878 , n1013 , n5877 );
not ( n5879 , n1524 );
and ( n5880 , n5221 , n5294 );
not ( n5881 , n5174 );
not ( n5882 , n5267 );
nor ( n5883 , n5882 , n4998 );
not ( n5884 , n5883 );
or ( n5885 , n5881 , n5884 );
nand ( n5886 , n5885 , n5024 );
nand ( n5887 , n5278 , n5886 );
nor ( n5888 , n5880 , n5887 );
not ( n5889 , n5888 );
and ( n5890 , n5879 , n5889 );
not ( n5891 , n5256 );
and ( n5892 , n5891 , n5883 );
not ( n5893 , n5118 );
nor ( n5894 , n5892 , n5893 );
nor ( n5895 , n5890 , n5894 );
nand ( n5896 , n5878 , n5895 );
nor ( n5897 , n5869 , n5896 );
and ( n5898 , n5854 , n5897 );
not ( n5899 , n5307 );
or ( n5900 , n5136 , n5873 );
not ( n5901 , n5263 );
nand ( n5902 , n5900 , n5901 );
or ( n5903 , n5256 , n5874 );
nand ( n5904 , n5903 , n4913 );
nand ( n5905 , n5902 , n5904 );
nor ( n5906 , n5899 , n5905 );
or ( n5907 , n1660 , n1204 );
nand ( n5908 , n5907 , n5849 );
and ( n5909 , n2849 , n5908 );
nand ( n5910 , n5453 , n5174 );
and ( n5911 , n5126 , n5910 );
nor ( n5912 , n5909 , n5911 );
or ( n5913 , n4944 , n5369 );
and ( n5914 , n5219 , n5354 );
not ( n5915 , n5336 );
not ( n5916 , n5322 );
or ( n5917 , n5915 , n5916 );
nand ( n5918 , n5917 , n5207 );
nand ( n5919 , n5913 , n5914 , n5918 );
and ( n5920 , n1660 , n5919 );
or ( n5921 , n5134 , n5321 );
nand ( n5922 , n5921 , n2251 );
not ( n5923 , n5922 );
nor ( n5924 , n5920 , n5923 );
or ( n5925 , n311 , n5924 );
or ( n5926 , n2254 , n5336 );
nand ( n5927 , n5925 , n5346 , n5926 );
nand ( n5928 , n948 , n5927 );
nand ( n5929 , n5898 , n5906 , n5912 , n5928 );
nand ( n5930 , n5853 , n5929 );
nand ( n5931 , n5743 , n5930 );
nand ( n5932 , n5681 , n5931 );
nand ( n5933 , n5131 , n4756 , n5932 );
nand ( n5934 , n2436 , n5933 );
not ( n5935 , n5934 );
not ( n5936 , n1076 );
nor ( n5937 , n2596 , n5936 );
not ( n5938 , n5827 );
not ( n5939 , n5938 );
not ( n5940 , n5939 );
and ( n5941 , n5937 , n5940 );
not ( n5942 , n5133 );
nor ( n5943 , n5941 , n5942 );
not ( n5944 , n5839 );
or ( n5945 , n5943 , n5944 );
nand ( n5946 , n5945 , n311 );
buf ( n5947 , n1076 );
buf ( n5948 , n5947 );
and ( n5949 , n5408 , n5420 );
nor ( n5950 , n5949 , n5430 );
nand ( n5951 , n5948 , n5950 );
not ( n5952 , n5951 );
nand ( n5953 , n5952 , n2549 , n5786 );
or ( n5954 , n2596 , n5953 );
nand ( n5955 , n5954 , n5792 );
nand ( n5956 , n5946 , n5955 );
and ( n5957 , n1767 , n5956 );
nand ( n5958 , n1435 , n5850 );
nor ( n5959 , n386 , n5797 );
or ( n5960 , n5959 , n5802 );
nand ( n5961 , n5960 , n2106 );
nand ( n5962 , n5958 , n4756 , n5961 );
nor ( n5963 , n5957 , n5962 , n393 );
nand ( n5964 , n793 , n1961 );
not ( n5965 , n5964 );
not ( n5966 , n5295 );
and ( n5967 , n5965 , n5966 );
nor ( n5968 , n5967 , n1464 );
not ( n5969 , n5520 );
nand ( n5970 , n5948 , n5969 );
not ( n5971 , n5970 );
nand ( n5972 , n5971 , n2550 , n5733 );
or ( n5973 , n2596 , n5972 );
nand ( n5974 , n5973 , n5741 );
and ( n5975 , n5968 , n5974 );
not ( n5976 , n2878 );
nor ( n5977 , n5942 , n5937 );
nand ( n5978 , n5976 , n5977 );
and ( n5979 , n2136 , n5866 );
or ( n5980 , n5552 , n5858 );
not ( n5981 , n358 );
nand ( n5982 , n5980 , n5981 );
nand ( n5983 , n1028 , n5977 );
nor ( n5984 , n386 , n1014 );
and ( n5985 , n5984 , n5231 );
nor ( n5986 , n5985 , n5905 );
nor ( n5987 , n5942 , n5552 );
nand ( n5988 , n5987 , n5861 );
nand ( n5989 , n5983 , n5986 , n5988 , n5878 );
nor ( n5990 , n5979 , n5982 , n5989 );
not ( n5991 , n5936 );
nand ( n5992 , n5991 , n5369 );
not ( n5993 , n5992 );
not ( n5994 , n5919 );
nand ( n5995 , n5922 , n5993 , n281 , n5994 );
or ( n5996 , n2596 , n5995 );
not ( n5997 , n5928 );
nand ( n5998 , n5996 , n5997 );
not ( n5999 , n5690 );
not ( n6000 , n5708 );
nand ( n6001 , n5948 , n6000 );
not ( n6002 , n6001 );
not ( n6003 , n5710 );
nand ( n6004 , n5999 , n6002 , n281 , n6003 );
or ( n6005 , n2596 , n6004 );
not ( n6006 , n3898 );
and ( n6007 , n6006 , n5712 );
nand ( n6008 , n6005 , n6007 );
nand ( n6009 , n5990 , n5998 , n6008 );
nand ( n6010 , n5597 , n1202 );
not ( n6011 , n6010 );
nand ( n6012 , n6011 , n5755 , n281 , n5751 );
and ( n6013 , n6012 , n5759 );
nand ( n6014 , n2665 , n6013 );
not ( n6015 , n5810 );
and ( n6016 , n5987 , n6015 );
nor ( n6017 , n6016 , n5825 );
not ( n6018 , n5064 );
nand ( n6019 , n5984 , n6018 );
nand ( n6020 , n6017 , n5983 , n6019 );
not ( n6021 , n358 );
not ( n6022 , n5844 );
nor ( n6023 , n6020 , n6021 , n6022 );
not ( n6024 , n5948 );
nor ( n6025 , n6024 , n5767 );
not ( n6026 , n5774 );
not ( n6027 , n5772 );
and ( n6028 , n6025 , n6026 , n281 , n6027 );
nor ( n6029 , n5779 , n6028 );
or ( n6030 , n2596 , n6029 );
nand ( n6031 , n6030 , n5780 );
nand ( n6032 , n6014 , n6023 , n6031 );
and ( n6033 , n6009 , n6032 );
nor ( n6034 , n386 , n5286 );
or ( n6035 , n6034 , n5720 );
nand ( n6036 , n6035 , n1218 );
and ( n6037 , n5912 , n6036 );
and ( n6038 , n6037 , n5895 );
nor ( n6039 , n6038 , n358 );
nor ( n6040 , n6033 , n6039 );
nand ( n6041 , n5975 , n5978 , n6040 );
not ( n6042 , n5507 );
not ( n6043 , n5522 );
not ( n6044 , n6043 );
nand ( n6045 , n6044 , n5971 );
not ( n6046 , n6045 );
not ( n6047 , n5525 );
nand ( n6048 , n6042 , n6046 , n281 , n6047 );
not ( n6049 , n6048 );
nand ( n6050 , n6049 , n329 );
and ( n6051 , n6050 , n5529 );
and ( n6052 , n5977 , n2868 , n3771 );
not ( n6053 , n5296 );
and ( n6054 , n5937 , n6053 );
nor ( n6055 , n6054 , n5964 );
nor ( n6056 , n6052 , n6055 );
nand ( n6057 , n1546 , n5046 );
nor ( n6058 , n386 , n4978 );
and ( n6059 , n1546 , n6058 );
or ( n6060 , n2933 , n5066 );
nand ( n6061 , n3388 , n5642 );
nand ( n6062 , n6060 , n6061 );
and ( n6063 , n5133 , n6062 );
nor ( n6064 , n6059 , n6063 , n5650 );
nand ( n6065 , n6056 , n6057 , n5490 , n6064 );
nor ( n6066 , n6051 , n6065 );
nor ( n6067 , n1937 , n5951 );
not ( n6068 , n5450 );
nand ( n6069 , n5457 , n6067 , n281 , n6068 );
or ( n6070 , n2596 , n6069 );
not ( n6071 , n5463 );
nand ( n6072 , n6070 , n6071 );
or ( n6073 , n386 , n5531 );
nand ( n6074 , n6073 , n5538 );
nand ( n6075 , n1947 , n6074 );
and ( n6076 , n5595 , n5634 );
or ( n6077 , n329 , n6076 );
nand ( n6078 , n5948 , n5572 );
not ( n6079 , n6078 );
not ( n6080 , n2548 );
nand ( n6081 , n6079 , n6080 , n5587 );
not ( n6082 , n64 );
and ( n6083 , n6081 , n6082 , n5594 );
and ( n6084 , n2664 , n6083 );
and ( n6085 , n5987 , n5546 );
not ( n6086 , n5128 );
and ( n6087 , n281 , n5093 );
or ( n6088 , n281 , n4942 );
nand ( n6089 , n6088 , n5805 );
nor ( n6090 , n6087 , n6089 );
nor ( n6091 , n6085 , n6086 , n6090 );
not ( n6092 , n5630 );
nor ( n6093 , n6010 , n5371 );
and ( n6094 , n6092 , n6093 , n281 , n5623 );
nor ( n6095 , n5634 , n6094 );
nor ( n6096 , n5569 , n6095 );
nand ( n6097 , n6091 , n358 , n6096 );
nor ( n6098 , n6084 , n6097 );
nand ( n6099 , n6077 , n6098 );
nand ( n6100 , n5669 , n1202 );
not ( n6101 , n6100 );
or ( n6102 , n386 , n6101 );
nand ( n6103 , n6102 , n5675 );
and ( n6104 , n2727 , n6103 );
nor ( n6105 , n6104 , n5665 , n5154 );
not ( n6106 , n6105 );
not ( n6107 , n64 );
nand ( n6108 , n6106 , n6107 , n2664 );
and ( n6109 , n5553 , n5477 );
not ( n6110 , n2914 );
nor ( n6111 , n329 , n6110 );
and ( n6112 , n6111 , n5665 );
and ( n6113 , n2906 , n5977 );
nor ( n6114 , n6109 , n6112 , n6113 );
not ( n6115 , n358 );
nand ( n6116 , n1076 , n5189 );
and ( n6117 , n5987 , n6116 );
nor ( n6118 , n6117 , n5217 );
and ( n6119 , n6108 , n6114 , n6115 , n6118 );
and ( n6120 , n5984 , n5236 );
not ( n6121 , n5305 );
nor ( n6122 , n6120 , n6121 );
or ( n6123 , n5155 , n5676 );
nand ( n6124 , n6123 , n6111 );
not ( n6125 , n5326 );
not ( n6126 , n6024 );
not ( n6127 , n5374 );
nand ( n6128 , n6126 , n6127 );
not ( n6129 , n6128 );
not ( n6130 , n5376 );
nand ( n6131 , n6125 , n6129 , n281 , n6130 );
or ( n6132 , n2596 , n6131 );
not ( n6133 , n5379 );
nand ( n6134 , n6132 , n6133 );
nand ( n6135 , n6119 , n6122 , n6124 , n6134 );
nand ( n6136 , n6099 , n6135 );
nand ( n6137 , n6066 , n6072 , n6075 , n6136 );
nand ( n6138 , n6041 , n6137 );
and ( n6139 , n5963 , n6138 );
not ( n6140 , n715 );
nor ( n6141 , n6139 , n6140 );
nor ( n6142 , n5935 , n6141 );
not ( n6143 , n391 );
not ( n6144 , n5933 );
not ( n6145 , n6144 );
or ( n6146 , n6143 , n6145 );
not ( n6147 , n6029 );
and ( n6148 , n6147 , n6019 , n5851 );
nor ( n6149 , n6148 , n2660 );
and ( n6150 , n6071 , n6069 );
and ( n6151 , n6048 , n5529 );
nor ( n6152 , n6150 , n6151 );
not ( n6153 , n6126 );
nand ( n6154 , n5899 , n2915 , n6153 );
and ( n6155 , n6122 , n6154 , n6118 );
nor ( n6156 , n6155 , n358 );
not ( n6157 , n5491 );
or ( n6158 , n5964 , n6053 );
nand ( n6159 , n6157 , n6158 , n6075 );
not ( n6160 , n3384 );
or ( n6161 , n6160 , n6105 );
nand ( n6162 , n1741 , n5378 , n6131 );
nand ( n6163 , n6161 , n6162 );
nor ( n6164 , n6156 , n6159 , n6163 );
and ( n6165 , n6152 , n6164 );
not ( n6166 , n358 );
and ( n6167 , n6007 , n6004 );
and ( n6168 , n5997 , n5995 );
nor ( n6169 , n6167 , n6168 );
nand ( n6170 , n5947 , n5860 );
and ( n6171 , n5987 , n6170 );
nand ( n6172 , n6154 , n5986 );
nor ( n6173 , n6171 , n6172 );
nand ( n6174 , n6169 , n6173 , n6037 , n5897 );
and ( n6175 , n6166 , n6174 );
and ( n6176 , n5972 , n5741 );
nor ( n6177 , n6175 , n6176 );
and ( n6178 , n5968 , n6177 );
nor ( n6179 , n6165 , n6178 );
nor ( n6180 , n6149 , n6179 );
and ( n6181 , n1767 , n5792 , n5953 );
not ( n6182 , n5130 );
not ( n6183 , n6096 );
or ( n6184 , n6182 , n6183 );
nand ( n6185 , n6184 , n358 );
and ( n6186 , n6064 , n6185 );
nor ( n6187 , n6186 , n372 );
nor ( n6188 , n6181 , n6187 );
nand ( n6189 , n1813 , n6083 );
nand ( n6190 , n1010 , n1768 );
not ( n6191 , n6190 );
or ( n6192 , n265 , n5637 );
nand ( n6193 , n6192 , n5808 );
and ( n6194 , n6191 , n6193 );
not ( n6195 , n5987 );
or ( n6196 , n1075 , n5545 );
nor ( n6197 , n5541 , n6196 );
or ( n6198 , n1760 , n6195 , n6197 );
not ( n6199 , n358 );
or ( n6200 , n6199 , n6154 );
nand ( n6201 , n6198 , n6200 );
nand ( n6202 , n2097 , n6196 );
or ( n6203 , n386 , n6202 );
nand ( n6204 , n6203 , n5961 );
nor ( n6205 , n6194 , n6201 , n6204 );
and ( n6206 , n1769 , n6013 );
nand ( n6207 , n2077 , n1806 );
not ( n6208 , n6207 );
nor ( n6209 , n386 , n5938 );
and ( n6210 , n6208 , n6209 );
nor ( n6211 , n6206 , n6210 );
and ( n6212 , n6188 , n6189 , n6205 , n6211 );
not ( n6213 , n393 );
not ( n6214 , n5934 );
or ( n6215 , n6213 , n6214 );
nand ( n6216 , n6215 , n4756 );
nand ( n6217 , n6180 , n6212 , n6216 );
nand ( n6218 , n6146 , n6217 );
nor ( n6219 , n6142 , n6218 );
and ( n6220 , n2986 , n6219 );
not ( n6221 , n2986 );
and ( n6222 , n6221 , n793 );
nor ( n6223 , n6220 , n6222 );
and ( n6224 , n394 , n396 );
not ( n6225 , n3038 );
not ( n6226 , n408 );
not ( n6227 , n6226 );
and ( n6228 , n6225 , n6227 );
nand ( n6229 , n410 , n411 );
not ( n6230 , n6229 );
nor ( n6231 , n6228 , n6230 );
nand ( n6232 , n736 , n6231 );
and ( n6233 , n416 , n6232 );
not ( n6234 , n6233 );
not ( n6235 , n409 );
not ( n6236 , n755 );
or ( n6237 , n6235 , n6236 );
nand ( n6238 , n6237 , n6231 );
nand ( n6239 , n5704 , n6238 );
not ( n6240 , n6239 );
not ( n6241 , n6240 );
nand ( n6242 , n6234 , n6241 );
buf ( n6243 , n6242 );
nand ( n6244 , n3303 , n6243 );
nand ( n6245 , n956 , n6238 );
not ( n6246 , n6240 );
nand ( n6247 , n6245 , n6246 );
and ( n6248 , n3303 , n6247 );
not ( n6249 , n736 );
nand ( n6250 , n4926 , n6249 );
not ( n6251 , n6250 );
not ( n6252 , n6231 );
or ( n6253 , n6251 , n6252 );
nand ( n6254 , n6253 , n1092 );
not ( n6255 , n6254 );
nand ( n6256 , n402 , n6255 );
not ( n6257 , n6256 );
nor ( n6258 , n6248 , n6257 );
nand ( n6259 , n6244 , n6258 );
not ( n6260 , n6259 );
not ( n6261 , n5289 );
not ( n6262 , n6261 );
not ( n6263 , n6255 );
nand ( n6264 , n3317 , n6240 );
and ( n6265 , n6263 , n6264 );
not ( n6266 , n6265 );
not ( n6267 , n6266 );
or ( n6268 , n6262 , n6267 );
not ( n6269 , n6242 );
nand ( n6270 , n6269 , n6245 );
nand ( n6271 , n3032 , n6270 );
nand ( n6272 , n6268 , n6271 );
not ( n6273 , n6272 );
nand ( n6274 , n6260 , n6273 );
and ( n6275 , n394 , n6274 );
nand ( n6276 , n394 , n769 );
not ( n6277 , n6276 );
not ( n6278 , n6277 );
not ( n6279 , n6265 );
nand ( n6280 , n407 , n6242 );
not ( n6281 , n6280 );
nor ( n6282 , n6279 , n6281 );
nor ( n6283 , n388 , n392 );
nand ( n6284 , n6283 , n2514 );
nor ( n6285 , n6282 , n6284 );
nand ( n6286 , n4948 , n6239 );
not ( n6287 , n6286 );
not ( n6288 , n6287 );
buf ( n6289 , n6288 );
nand ( n6290 , n407 , n6289 );
nor ( n6291 , n6233 , n6286 );
nor ( n6292 , n407 , n6291 );
and ( n6293 , n6292 , n730 );
not ( n6294 , n6255 );
not ( n6295 , n6294 );
nor ( n6296 , n6293 , n6295 );
nand ( n6297 , n6290 , n6296 );
not ( n6298 , n6297 );
not ( n6299 , n6298 );
and ( n6300 , n6285 , n6299 );
not ( n6301 , n6300 );
nand ( n6302 , n6278 , n6301 );
not ( n6303 , n6302 );
not ( n6304 , n6303 );
nor ( n6305 , n6275 , n6304 );
or ( n6306 , n6224 , n6305 );
not ( n6307 , n6224 );
nor ( n6308 , n390 , n6283 );
not ( n6309 , n6308 );
or ( n6310 , n6307 , n6309 );
not ( n6311 , n6298 );
nor ( n6312 , n6281 , n6311 );
not ( n6313 , n6312 );
nand ( n6314 , n6224 , n6313 );
and ( n6315 , n1323 , n6314 );
nand ( n6316 , n6310 , n6315 );
not ( n6317 , n6316 );
nand ( n6318 , n6306 , n6317 );
and ( n6319 , n329 , n2065 , n6318 );
not ( n6320 , n6308 );
and ( n6321 , n6224 , n6320 );
not ( n6322 , n6321 );
not ( n6323 , n3087 );
nor ( n6324 , n3146 , n6291 );
not ( n6325 , n6324 );
or ( n6326 , n6323 , n6325 );
not ( n6327 , n5362 );
nand ( n6328 , n6327 , n6266 );
nand ( n6329 , n6326 , n6328 );
not ( n6330 , n6329 );
not ( n6331 , n6330 );
not ( n6332 , n414 );
not ( n6333 , n6289 );
or ( n6334 , n6332 , n6333 );
not ( n6335 , n1089 );
not ( n6336 , n6287 );
nand ( n6337 , n6335 , n6336 );
not ( n6338 , n6337 );
not ( n6339 , n6338 );
nand ( n6340 , n6334 , n6339 );
not ( n6341 , n3304 );
nand ( n6342 , n6340 , n6341 );
not ( n6343 , n3304 );
and ( n6344 , n6343 , n6338 );
nor ( n6345 , n6344 , n6257 );
and ( n6346 , n6244 , n6345 );
nand ( n6347 , n6342 , n6346 );
nor ( n6348 , n6331 , n6347 );
or ( n6349 , n1847 , n6348 );
buf ( n6350 , n6303 );
nand ( n6351 , n6349 , n6350 );
and ( n6352 , n6322 , n6351 );
not ( n6353 , n6315 );
not ( n6354 , n6353 );
not ( n6355 , n6354 );
nor ( n6356 , n6352 , n6355 );
or ( n6357 , n3562 , n6356 );
not ( n6358 , n810 );
or ( n6359 , n6358 , n6264 );
not ( n6360 , n3028 );
not ( n6361 , n414 );
not ( n6362 , n6289 );
or ( n6363 , n6361 , n6362 );
nand ( n6364 , n6363 , n6245 );
not ( n6365 , n6364 );
nand ( n6366 , n6234 , n6365 );
not ( n6367 , n6366 );
or ( n6368 , n6360 , n6367 );
nand ( n6369 , n6368 , n6294 );
not ( n6370 , n6369 );
nand ( n6371 , n6359 , n6370 );
and ( n6372 , n394 , n6371 );
buf ( n6373 , n6303 );
not ( n6374 , n6373 );
nor ( n6375 , n6372 , n6374 );
or ( n6376 , n6321 , n6375 );
not ( n6377 , n6354 );
not ( n6378 , n6377 );
nand ( n6379 , n6376 , n6378 );
nand ( n6380 , n2606 , n6379 );
nand ( n6381 , n6357 , n6380 );
and ( n6382 , n4084 , n6381 );
nor ( n6383 , n6319 , n6382 );
not ( n6384 , n2072 );
not ( n6385 , n6384 );
nand ( n6386 , n6234 , n6337 );
nand ( n6387 , n3087 , n6386 );
nand ( n6388 , n6387 , n6328 );
not ( n6389 , n6388 );
nand ( n6390 , n6346 , n6389 );
and ( n6391 , n394 , n6390 );
not ( n6392 , n6350 );
nor ( n6393 , n6391 , n6392 );
or ( n6394 , n6321 , n6393 );
not ( n6395 , n6377 );
nand ( n6396 , n6394 , n6395 );
not ( n6397 , n6396 );
or ( n6398 , n6385 , n6397 );
and ( n6399 , n2549 , n6353 );
not ( n6400 , n2254 );
not ( n6401 , n6230 );
or ( n6402 , n6401 , n769 );
nand ( n6403 , n6402 , n6276 );
nand ( n6404 , n2251 , n6403 );
not ( n6405 , n6404 );
or ( n6406 , n6400 , n6405 );
not ( n6407 , n6277 );
not ( n6408 , n6231 );
nand ( n6409 , n6408 , n825 );
and ( n6410 , n6407 , n6409 );
nor ( n6411 , n6410 , n311 );
nand ( n6412 , n6406 , n6411 );
not ( n6413 , n311 );
not ( n6414 , n825 );
not ( n6415 , n6232 );
or ( n6416 , n6414 , n6415 );
nand ( n6417 , n6416 , n6276 );
nand ( n6418 , n3755 , n6417 );
nor ( n6419 , n6413 , n6418 );
nand ( n6420 , n2251 , n5106 );
nor ( n6421 , n410 , n6420 );
nand ( n6422 , n6283 , n6421 );
and ( n6423 , n6422 , n6404 );
not ( n6424 , n311 );
nor ( n6425 , n6423 , n6424 );
nor ( n6426 , n6419 , n6425 );
nand ( n6427 , n6412 , n6426 );
nor ( n6428 , n6399 , n6427 );
not ( n6429 , n6428 );
nand ( n6430 , n6429 , n64 );
not ( n6431 , n6430 );
not ( n6432 , n6224 );
not ( n6433 , n394 );
not ( n6434 , n6259 );
not ( n6435 , n3531 );
not ( n6436 , n6435 );
not ( n6437 , n6436 );
nand ( n6438 , n414 , n6288 );
and ( n6439 , n6438 , n6269 );
not ( n6440 , n6439 );
and ( n6441 , n6437 , n6440 );
nor ( n6442 , n6441 , n6257 );
nand ( n6443 , n6440 , n407 );
not ( n6444 , n860 );
nand ( n6445 , n6444 , n6247 );
nand ( n6446 , n6443 , n6445 );
or ( n6447 , n3471 , n6446 );
nand ( n6448 , n6447 , n6366 , n3484 );
nand ( n6449 , n6442 , n6448 );
not ( n6450 , n6449 );
or ( n6451 , n6434 , n6450 );
nand ( n6452 , n6445 , n6282 );
and ( n6453 , n3129 , n6452 );
and ( n6454 , n892 , n6294 );
and ( n6455 , n6454 , n6439 );
not ( n6456 , n399 );
nor ( n6457 , n6455 , n6456 );
nand ( n6458 , n6457 , n6272 );
not ( n6459 , n6458 );
nor ( n6460 , n6453 , n6459 );
nand ( n6461 , n6451 , n6460 );
not ( n6462 , n6461 );
or ( n6463 , n6433 , n6462 );
nand ( n6464 , n6463 , n6350 );
not ( n6465 , n6464 );
and ( n6466 , n6432 , n6465 );
nor ( n6467 , n6466 , n3019 );
or ( n6468 , n410 , n869 );
nand ( n6469 , n6468 , n6280 );
and ( n6470 , n780 , n6469 );
nor ( n6471 , n6470 , n3129 );
buf ( n6472 , n6266 );
nor ( n6473 , n6472 , n6469 );
or ( n6474 , n6471 , n6473 );
not ( n6475 , n6386 );
or ( n6476 , n3460 , n6475 );
not ( n6477 , n6240 );
not ( n6478 , n6477 );
nand ( n6479 , n3096 , n6478 );
nand ( n6480 , n6454 , n6479 );
and ( n6481 , n6480 , n6388 );
not ( n6482 , n402 );
not ( n6483 , n6280 );
not ( n6484 , n6483 );
nand ( n6485 , n1142 , n6338 );
nand ( n6486 , n6484 , n6485 );
nand ( n6487 , n6482 , n6486 );
and ( n6488 , n3183 , n6487 );
not ( n6489 , n6243 );
buf ( n6490 , n6489 );
nor ( n6491 , n6488 , n6490 );
or ( n6492 , n6481 , n6491 );
nand ( n6493 , n6492 , n399 );
nand ( n6494 , n6474 , n6476 , n6493 );
not ( n6495 , n6437 );
or ( n6496 , n6495 , n6490 );
nand ( n6497 , n6496 , n6256 );
nor ( n6498 , n6494 , n6497 );
or ( n6499 , n1847 , n6498 );
nand ( n6500 , n6499 , n6350 );
and ( n6501 , n1104 , n6500 );
or ( n6502 , n6467 , n6501 );
nand ( n6503 , n6502 , n6322 );
not ( n6504 , n6503 );
or ( n6505 , n6431 , n6504 );
nand ( n6506 , n6505 , n1359 );
nand ( n6507 , n6398 , n6506 );
nand ( n6508 , n1464 , n329 , n6507 );
nand ( n6509 , n6383 , n4684 , n6508 );
not ( n6510 , n2597 );
not ( n6511 , n6301 );
not ( n6512 , n6511 );
and ( n6513 , n6126 , n6312 );
nor ( n6514 , n6513 , n1847 );
not ( n6515 , n6514 );
nand ( n6516 , n6512 , n6515 );
not ( n6517 , n6516 );
or ( n6518 , n6510 , n6517 );
not ( n6519 , n6427 );
nand ( n6520 , n6518 , n6519 );
not ( n6521 , n6520 );
and ( n6522 , n1464 , n6521 );
not ( n6523 , n396 );
not ( n6524 , n402 );
not ( n6525 , n6472 );
not ( n6526 , n6525 );
or ( n6527 , n6526 , n6486 );
nand ( n6528 , n6527 , n3130 );
not ( n6529 , n399 );
not ( n6530 , n3204 );
not ( n6531 , n6489 );
and ( n6532 , n6530 , n6531 );
and ( n6533 , n413 , n6294 );
nand ( n6534 , n6533 , n6479 );
and ( n6535 , n6388 , n6534 );
nor ( n6536 , n6532 , n6535 );
nand ( n6537 , n6487 , n6536 );
nand ( n6538 , n6529 , n6537 );
nand ( n6539 , n6528 , n6538 );
and ( n6540 , n6524 , n6539 );
and ( n6541 , n780 , n6486 );
or ( n6542 , n6436 , n6475 );
not ( n6543 , n3471 );
not ( n6544 , n6242 );
or ( n6545 , n6543 , n6544 );
nand ( n6546 , n6545 , n6256 );
not ( n6547 , n6546 );
nand ( n6548 , n6542 , n6547 );
nor ( n6549 , n6541 , n6548 );
nand ( n6550 , n6549 , n6538 );
nor ( n6551 , n6540 , n6550 );
or ( n6552 , n6551 , n1847 );
not ( n6553 , n6374 );
nand ( n6554 , n6552 , n6553 );
and ( n6555 , n6523 , n6554 );
nor ( n6556 , n6555 , n6316 , n6511 );
or ( n6557 , n1554 , n6556 );
and ( n6558 , n6525 , n6443 );
nor ( n6559 , n1847 , n6558 );
not ( n6560 , n6303 );
nor ( n6561 , n6559 , n6560 );
or ( n6562 , n6321 , n6561 );
nand ( n6563 , n6562 , n6315 );
nand ( n6564 , n1947 , n6563 );
nand ( n6565 , n6557 , n6564 );
not ( n6566 , n6565 );
not ( n6567 , n1070 );
not ( n6568 , n6525 );
nor ( n6569 , n6568 , n6446 );
or ( n6570 , n3130 , n6569 );
not ( n6571 , n6449 );
and ( n6572 , n3032 , n6440 );
nor ( n6573 , n6572 , n6272 );
not ( n6574 , n6573 );
nand ( n6575 , n6457 , n6574 );
nand ( n6576 , n6570 , n6571 , n6575 );
not ( n6577 , n6576 );
or ( n6578 , n6567 , n6577 );
not ( n6579 , n779 );
nand ( n6580 , n6444 , n6340 );
nand ( n6581 , n6443 , n6580 );
not ( n6582 , n6581 );
not ( n6583 , n6582 );
and ( n6584 , n6579 , n6583 );
not ( n6585 , n6525 );
not ( n6586 , n6585 );
nand ( n6587 , n6586 , n6582 );
and ( n6588 , n3129 , n6587 );
nor ( n6589 , n6584 , n6588 );
nand ( n6590 , n6442 , n6589 );
not ( n6591 , n3471 );
not ( n6592 , n6324 );
or ( n6593 , n6591 , n6592 );
not ( n6594 , n402 );
not ( n6595 , n6594 );
not ( n6596 , n6581 );
or ( n6597 , n6595 , n6596 );
and ( n6598 , n6329 , n6480 );
and ( n6599 , n3083 , n6440 );
nor ( n6600 , n6598 , n6599 );
nand ( n6601 , n6597 , n6600 );
nand ( n6602 , n399 , n6601 );
nand ( n6603 , n6593 , n6602 );
or ( n6604 , n6590 , n6603 );
nand ( n6605 , n6604 , n1104 );
nand ( n6606 , n6578 , n6605 );
and ( n6607 , n6606 , n394 );
not ( n6608 , n1069 );
not ( n6609 , n6304 );
or ( n6610 , n6608 , n6609 );
nand ( n6611 , n64 , n6427 );
nand ( n6612 , n6610 , n6611 );
nor ( n6613 , n6607 , n6612 );
or ( n6614 , n6613 , n6321 );
nand ( n6615 , n6614 , n6430 );
nand ( n6616 , n1763 , n6615 );
not ( n6617 , n394 );
not ( n6618 , n6289 );
not ( n6619 , n6618 );
nand ( n6620 , n890 , n6619 );
nand ( n6621 , n6620 , n6256 , n6342 );
nand ( n6622 , n414 , n6621 );
not ( n6623 , n6622 );
not ( n6624 , n402 );
nand ( n6625 , n6485 , n6443 );
nand ( n6626 , n6624 , n6625 );
and ( n6627 , n6534 , n6329 );
not ( n6628 , n3204 );
and ( n6629 , n6628 , n6440 );
nor ( n6630 , n6627 , n6629 );
and ( n6631 , n6626 , n6630 );
nor ( n6632 , n6631 , n399 );
nor ( n6633 , n6623 , n6632 );
not ( n6634 , n402 );
not ( n6635 , n6632 );
or ( n6636 , n6625 , n6568 );
nand ( n6637 , n6636 , n3130 );
nand ( n6638 , n6635 , n6637 );
nand ( n6639 , n6634 , n6638 );
nand ( n6640 , n6633 , n6549 , n6639 );
not ( n6641 , n6640 );
or ( n6642 , n6617 , n6641 );
buf ( n6643 , n6350 );
buf ( n6644 , n6643 );
nand ( n6645 , n6642 , n6644 );
not ( n6646 , n6645 );
or ( n6647 , n6646 , n6321 );
nand ( n6648 , n6647 , n6395 );
nand ( n6649 , n1380 , n6648 );
nand ( n6650 , n1142 , n6247 );
nand ( n6651 , n6443 , n6650 );
not ( n6652 , n6651 );
and ( n6653 , n6652 , n6495 );
nor ( n6654 , n6653 , n3522 );
and ( n6655 , n6270 , n6654 );
nor ( n6656 , n6655 , n6546 );
not ( n6657 , n6533 );
or ( n6658 , n6657 , n6440 );
not ( n6659 , n399 );
nand ( n6660 , n6658 , n6659 );
or ( n6661 , n6573 , n6660 );
and ( n6662 , n6656 , n6661 );
and ( n6663 , n414 , n6449 );
or ( n6664 , n6651 , n6585 );
nand ( n6665 , n6664 , n3130 );
nand ( n6666 , n6665 , n6661 );
not ( n6667 , n6666 );
nor ( n6668 , n402 , n6667 );
nor ( n6669 , n6663 , n6668 );
nand ( n6670 , n6662 , n6669 );
and ( n6671 , n394 , n6670 );
not ( n6672 , n6350 );
nor ( n6673 , n6671 , n6672 );
or ( n6674 , n6321 , n6673 );
nand ( n6675 , n6674 , n6395 );
and ( n6676 , n1961 , n6675 );
not ( n6677 , n1298 );
nand ( n6678 , n6244 , n6282 );
and ( n6679 , n394 , n6678 );
not ( n6680 , n6350 );
nor ( n6681 , n6679 , n6680 );
not ( n6682 , n6681 );
and ( n6683 , n6677 , n6682 );
and ( n6684 , n6650 , n6282 );
nor ( n6685 , n6684 , n3129 );
nor ( n6686 , n6660 , n6273 );
nor ( n6687 , n6685 , n6686 );
or ( n6688 , n402 , n6687 );
not ( n6689 , n6686 );
nand ( n6690 , n6688 , n6689 , n6656 );
nand ( n6691 , n394 , n6690 );
and ( n6692 , n6643 , n6691 );
nor ( n6693 , n6692 , n1547 );
nor ( n6694 , n6683 , n6693 );
nor ( n6695 , n6694 , n6321 );
not ( n6696 , n5705 );
nand ( n6697 , n1210 , n6477 );
not ( n6698 , n6697 );
not ( n6699 , n6698 );
not ( n6700 , n6699 );
nand ( n6701 , n6341 , n6700 );
not ( n6702 , n6701 );
and ( n6703 , n6696 , n6702 );
not ( n6704 , n6558 );
nor ( n6705 , n6703 , n6704 );
or ( n6706 , n1847 , n6705 );
nand ( n6707 , n6706 , n6373 );
nand ( n6708 , n1947 , n6707 );
or ( n6709 , n396 , n6708 );
or ( n6710 , n1538 , n1546 );
nand ( n6711 , n6710 , n6355 );
nand ( n6712 , n6709 , n6711 );
nor ( n6713 , n6676 , n6695 , n6712 );
nand ( n6714 , n6566 , n6616 , n6649 , n6713 );
nand ( n6715 , n329 , n6714 );
and ( n6716 , n6522 , n6715 );
and ( n6717 , n394 , n6638 );
not ( n6718 , n6350 );
nor ( n6719 , n6717 , n6718 );
or ( n6720 , n6321 , n6719 );
nand ( n6721 , n6720 , n6395 );
nand ( n6722 , n3195 , n6721 );
not ( n6723 , n5763 );
not ( n6724 , n6723 );
and ( n6725 , n6724 , n6347 );
not ( n6726 , n6478 );
nor ( n6727 , n5683 , n6726 );
nor ( n6728 , n6725 , n6727 );
and ( n6729 , n6330 , n6728 );
or ( n6730 , n6729 , n1847 );
nand ( n6731 , n6730 , n6373 );
not ( n6732 , n6731 );
or ( n6733 , n6321 , n6732 );
nand ( n6734 , n6733 , n6395 );
and ( n6735 , n2650 , n6734 );
not ( n6736 , n2857 );
or ( n6737 , n1847 , n6687 );
nand ( n6738 , n6737 , n6373 );
and ( n6739 , n6322 , n6738 );
not ( n6740 , n6354 );
nor ( n6741 , n6739 , n6740 );
or ( n6742 , n6736 , n6741 );
not ( n6743 , n394 );
not ( n6744 , n6282 );
not ( n6745 , n6744 );
or ( n6746 , n6743 , n6745 );
nand ( n6747 , n6746 , n6350 );
not ( n6748 , n6747 );
nand ( n6749 , n6748 , n6314 );
nand ( n6750 , n2629 , n6749 );
nand ( n6751 , n6742 , n6750 , n6521 );
nor ( n6752 , n6735 , n6751 , n1464 );
not ( n6753 , n394 );
not ( n6754 , n6539 );
or ( n6755 , n6753 , n6754 );
nand ( n6756 , n6755 , n6553 );
and ( n6757 , n6322 , n6756 );
nor ( n6758 , n6757 , n6355 );
or ( n6759 , n1554 , n6758 );
not ( n6760 , n1359 );
not ( n6761 , n6350 );
not ( n6762 , n6452 );
buf ( n6763 , n3636 );
or ( n6764 , n6762 , n6763 );
nand ( n6765 , n6764 , n6458 );
and ( n6766 , n1010 , n6765 );
not ( n6767 , n6723 );
not ( n6768 , n6767 );
not ( n6769 , n6259 );
or ( n6770 , n6768 , n6769 );
nor ( n6771 , n6727 , n6272 );
nand ( n6772 , n6770 , n6771 );
and ( n6773 , n1252 , n6772 );
nor ( n6774 , n6766 , n6773 );
or ( n6775 , n6728 , n1096 );
nand ( n6776 , n6775 , n6389 );
nand ( n6777 , n1244 , n6776 );
not ( n6778 , n6763 );
not ( n6779 , n6778 );
not ( n6780 , n6473 );
not ( n6781 , n6780 );
or ( n6782 , n6779 , n6781 );
nand ( n6783 , n6782 , n6493 );
nand ( n6784 , n1494 , n6783 );
nand ( n6785 , n6774 , n6777 , n6784 );
nand ( n6786 , n394 , n6785 );
not ( n6787 , n6786 );
or ( n6788 , n6761 , n6787 );
nand ( n6789 , n6788 , n2550 );
not ( n6790 , n6789 );
not ( n6791 , n6790 );
or ( n6792 , n6760 , n6791 );
not ( n6793 , n6612 );
not ( n6794 , n1070 );
not ( n6795 , n6763 );
not ( n6796 , n6795 );
or ( n6797 , n6796 , n6569 );
nand ( n6798 , n6797 , n6575 );
not ( n6799 , n6798 );
or ( n6800 , n6794 , n6799 );
not ( n6801 , n6796 );
nand ( n6802 , n6801 , n6587 );
not ( n6803 , n6802 );
not ( n6804 , n6602 );
or ( n6805 , n6803 , n6804 );
nand ( n6806 , n6805 , n1104 );
nand ( n6807 , n6800 , n6806 );
nand ( n6808 , n394 , n6807 );
nand ( n6809 , n6793 , n6808 );
nand ( n6810 , n1763 , n6809 );
nand ( n6811 , n6792 , n6810 );
nand ( n6812 , n6811 , n6322 );
not ( n6813 , n394 );
not ( n6814 , n6666 );
or ( n6815 , n6813 , n6814 );
nand ( n6816 , n6815 , n6373 );
and ( n6817 , n6432 , n6816 );
nor ( n6818 , n6817 , n6316 );
or ( n6819 , n1962 , n6818 );
nand ( n6820 , n6819 , n6564 );
and ( n6821 , n6724 , n6369 );
not ( n6822 , n6727 );
nand ( n6823 , n6822 , n6573 );
nor ( n6824 , n6821 , n6823 );
or ( n6825 , n6824 , n1847 );
nand ( n6826 , n6825 , n6350 );
and ( n6827 , n6322 , n6826 );
nor ( n6828 , n6827 , n6353 );
or ( n6829 , n2945 , n6828 );
nor ( n6830 , n948 , n1359 );
or ( n6831 , n6830 , n6428 );
nand ( n6832 , n6829 , n6831 );
nor ( n6833 , n6820 , n6832 );
nand ( n6834 , n6759 , n6812 , n6833 );
nand ( n6835 , n329 , n6834 );
and ( n6836 , n6722 , n6752 , n6835 );
nor ( n6837 , n6716 , n6836 );
nor ( n6838 , n6509 , n6837 );
not ( n6839 , n1070 );
not ( n6840 , n6464 );
or ( n6841 , n6839 , n6840 );
nand ( n6842 , n6841 , n6611 );
or ( n6843 , n6842 , n6501 );
nand ( n6844 , n6843 , n1359 );
and ( n6845 , n1380 , n6645 );
and ( n6846 , n1553 , n6554 );
nor ( n6847 , n6845 , n6846 );
or ( n6848 , n2072 , n6393 );
or ( n6849 , n6375 , n2945 );
nand ( n6850 , n6848 , n6849 );
or ( n6851 , n6673 , n1962 );
nand ( n6852 , n6851 , n6708 );
nor ( n6853 , n6850 , n6852 );
nand ( n6854 , n6844 , n6847 , n6694 , n6853 );
nand ( n6855 , n1291 , n6351 );
and ( n6856 , n6613 , n6855 );
nor ( n6857 , n6856 , n1764 );
nor ( n6858 , n6854 , n6857 );
or ( n6859 , n2596 , n6858 );
or ( n6860 , n2837 , n6305 );
nand ( n6861 , n6859 , n6521 , n6860 );
and ( n6862 , n2023 , n6861 );
nand ( n6863 , n403 , n2077 );
not ( n6864 , n6863 );
nor ( n6865 , n329 , n6284 );
not ( n6866 , n6865 );
or ( n6867 , n956 , n6290 );
nand ( n6868 , n6444 , n6697 );
and ( n6869 , n6868 , n6650 );
nand ( n6870 , n6867 , n6869 );
not ( n6871 , n6870 );
not ( n6872 , n6296 );
nand ( n6873 , n3130 , n6872 );
not ( n6874 , n399 );
nand ( n6875 , n417 , n6292 );
nand ( n6876 , n6533 , n6875 );
not ( n6877 , n6876 );
not ( n6878 , n3087 );
not ( n6879 , n6364 );
or ( n6880 , n6878 , n6879 );
and ( n6881 , n746 , n981 );
not ( n6882 , n402 );
nand ( n6883 , n6882 , n6297 );
not ( n6884 , n6883 );
nand ( n6885 , n6881 , n6884 );
nand ( n6886 , n6880 , n6885 );
not ( n6887 , n6886 );
or ( n6888 , n6877 , n6887 );
not ( n6889 , n402 );
and ( n6890 , n6870 , n6889 );
and ( n6891 , n6628 , n6619 );
nor ( n6892 , n6890 , n6891 );
nand ( n6893 , n6888 , n6892 );
nand ( n6894 , n6874 , n6893 );
nand ( n6895 , n6871 , n6873 , n6894 );
nand ( n6896 , n1291 , n6895 );
or ( n6897 , n6866 , n6896 );
not ( n6898 , n64 );
and ( n6899 , n2597 , n6514 );
and ( n6900 , n6898 , n6899 );
nor ( n6901 , n2598 , n6284 );
nand ( n6902 , n64 , n6901 );
not ( n6903 , n6902 );
and ( n6904 , n6903 , n6311 );
nor ( n6905 , n6900 , n6904 );
nand ( n6906 , n6897 , n6905 );
and ( n6907 , n6864 , n6906 );
not ( n6908 , n311 );
nor ( n6909 , n6908 , n6902 );
not ( n6910 , n6872 );
not ( n6911 , n6910 );
nand ( n6912 , n1142 , n6288 );
nand ( n6913 , n6580 , n6912 );
or ( n6914 , n6911 , n6913 );
nand ( n6915 , n6914 , n6795 );
buf ( n6916 , n6915 );
not ( n6917 , n402 );
and ( n6918 , n6917 , n6913 );
and ( n6919 , n892 , n902 , n6619 );
nor ( n6920 , n6918 , n6919 );
not ( n6921 , n6920 );
and ( n6922 , n3032 , n6340 );
not ( n6923 , n3032 );
not ( n6924 , n6883 );
and ( n6925 , n6923 , n6924 );
nor ( n6926 , n6922 , n6925 );
not ( n6927 , n6926 );
or ( n6928 , n6921 , n6927 );
nand ( n6929 , n6928 , n399 );
nand ( n6930 , n6916 , n6929 );
and ( n6931 , n6909 , n6930 );
and ( n6932 , n64 , n6899 );
nor ( n6933 , n6931 , n6932 );
not ( n6934 , n6899 );
nand ( n6935 , n6418 , n6934 );
nand ( n6936 , n1252 , n6935 );
not ( n6937 , n6910 );
and ( n6938 , n6444 , n6364 );
not ( n6939 , n6912 );
nor ( n6940 , n6938 , n6939 );
not ( n6941 , n6940 );
or ( n6942 , n6937 , n6941 );
not ( n6943 , n6763 );
nand ( n6944 , n6942 , n6943 );
nand ( n6945 , n6454 , n6875 );
not ( n6946 , n6945 );
not ( n6947 , n6886 );
or ( n6948 , n6946 , n6947 );
not ( n6949 , n6940 );
not ( n6950 , n402 );
and ( n6951 , n6949 , n6950 );
and ( n6952 , n3083 , n6619 );
nor ( n6953 , n6951 , n6952 );
nand ( n6954 , n6948 , n6953 );
nand ( n6955 , n399 , n6954 );
nand ( n6956 , n6944 , n6955 );
not ( n6957 , n6956 );
not ( n6958 , n6957 );
nor ( n6959 , n311 , n6902 );
nand ( n6960 , n6958 , n6959 );
and ( n6961 , n6933 , n6936 , n6960 );
nor ( n6962 , n2028 , n2660 );
nand ( n6963 , n1027 , n6962 );
nor ( n6964 , n6961 , n6963 );
nor ( n6965 , n6907 , n6964 );
not ( n6966 , n6284 );
and ( n6967 , n396 , n6966 );
nand ( n6968 , n6967 , n6311 );
not ( n6969 , n792 );
or ( n6970 , n396 , n6969 );
not ( n6971 , n6970 );
and ( n6972 , n6971 , n6744 );
nand ( n6973 , n6523 , n6300 );
nand ( n6974 , n6314 , n6278 , n6973 );
not ( n6975 , n6974 );
not ( n6976 , n6975 );
not ( n6977 , n6976 );
not ( n6978 , n6977 );
nor ( n6979 , n6972 , n6978 );
and ( n6980 , n6968 , n6979 );
nor ( n6981 , n6980 , n2338 , n1298 );
and ( n6982 , n329 , n6981 );
nor ( n6983 , n6982 , n4684 );
nor ( n6984 , n6963 , n1565 );
not ( n6985 , n6984 );
not ( n6986 , n6364 );
nor ( n6987 , n6986 , n6881 );
nor ( n6988 , n5683 , n6291 );
not ( n6989 , n6988 );
not ( n6990 , n3087 );
not ( n6991 , n6247 );
or ( n6992 , n6990 , n6991 );
nand ( n6993 , n6992 , n6885 );
not ( n6994 , n6993 );
nand ( n6995 , n6258 , n6994 );
not ( n6996 , n6995 );
nand ( n6997 , n6989 , n6996 );
nor ( n6998 , n6987 , n6997 );
or ( n6999 , n6985 , n6998 );
not ( n7000 , n6926 );
not ( n7001 , n7000 );
and ( n7002 , n1204 , n3133 );
nor ( n7003 , n7002 , n6618 );
nand ( n7004 , n6868 , n6485 );
nor ( n7005 , n7003 , n7004 );
nand ( n7006 , n7001 , n7005 , n6873 );
nand ( n7007 , n1806 , n7006 );
or ( n7008 , n6863 , n7007 );
nand ( n7009 , n6962 , n2136 );
nand ( n7010 , n6256 , n6342 );
nor ( n7011 , n7000 , n7010 );
nand ( n7012 , n6989 , n7011 );
not ( n7013 , n7012 );
or ( n7014 , n7009 , n7013 );
nand ( n7015 , n6999 , n7008 , n7014 );
and ( n7016 , n6865 , n7015 );
nand ( n7017 , n6971 , n6772 );
not ( n7018 , n6978 );
nand ( n7019 , n6967 , n7012 );
and ( n7020 , n7017 , n7018 , n7019 );
nor ( n7021 , n7020 , n2338 , n2837 );
nor ( n7022 , n7016 , n7021 );
nand ( n7023 , n6965 , n6983 , n7022 );
nor ( n7024 , n6862 , n7023 );
and ( n7025 , n2763 , n6411 );
nor ( n7026 , n7025 , n329 , n6427 );
not ( n7027 , n7026 );
nand ( n7028 , n6971 , n1104 );
not ( n7029 , n7028 );
and ( n7030 , n7029 , n6783 );
nor ( n7031 , n6970 , n3019 );
and ( n7032 , n7031 , n6765 );
nor ( n7033 , n7030 , n7032 );
nand ( n7034 , n1069 , n6976 );
and ( n7035 , n6611 , n7034 );
nand ( n7036 , n1070 , n6967 );
not ( n7037 , n7036 );
not ( n7038 , n6930 );
not ( n7039 , n7038 );
and ( n7040 , n7037 , n7039 );
not ( n7041 , n6967 );
nor ( n7042 , n2725 , n7041 );
and ( n7043 , n64 , n7042 );
not ( n7044 , n7043 );
nor ( n7045 , n7044 , n6957 );
nor ( n7046 , n7040 , n7045 );
and ( n7047 , n7033 , n7035 , n7046 );
or ( n7048 , n6963 , n7047 );
not ( n7049 , n64 );
nand ( n7050 , n7049 , n6427 );
nand ( n7051 , n2093 , n6974 );
and ( n7052 , n7050 , n7051 );
not ( n7053 , n7052 );
nor ( n7054 , n6970 , n1565 );
not ( n7055 , n7054 );
not ( n7056 , n6539 );
or ( n7057 , n7055 , n7056 );
nor ( n7058 , n6970 , n1264 );
not ( n7059 , n7058 );
or ( n7060 , n7059 , n6687 );
nand ( n7061 , n7057 , n7060 );
and ( n7062 , n7007 , n6896 );
nor ( n7063 , n7062 , n7041 );
nor ( n7064 , n7053 , n7061 , n7063 );
or ( n7065 , n6863 , n7064 );
nand ( n7066 , n7048 , n7065 );
nand ( n7067 , n7027 , n7066 );
not ( n7068 , n6776 );
or ( n7069 , n6970 , n7068 );
not ( n7070 , n6987 );
nand ( n7071 , n7070 , n6996 );
nand ( n7072 , n6967 , n7071 );
and ( n7073 , n6967 , n6997 );
nor ( n7074 , n7073 , n6978 );
nand ( n7075 , n7069 , n7072 , n7074 );
and ( n7076 , n2894 , n7075 );
or ( n7077 , n6970 , n6729 );
nand ( n7078 , n7077 , n7074 );
and ( n7079 , n2650 , n7078 );
nor ( n7080 , n7076 , n7079 );
not ( n7081 , n6824 );
nand ( n7082 , n7081 , n6971 );
buf ( n7083 , n6339 );
nor ( n7084 , n3031 , n7083 );
not ( n7085 , n7084 );
nand ( n7086 , n3031 , n6924 );
nand ( n7087 , n7085 , n7086 );
not ( n7088 , n7087 );
nand ( n7089 , n6345 , n7088 );
nor ( n7090 , n6988 , n7089 );
not ( n7091 , n7090 );
nand ( n7092 , n7091 , n6967 );
and ( n7093 , n7082 , n7092 , n7018 );
or ( n7094 , n2644 , n7093 );
or ( n7095 , n1764 , n6936 );
or ( n7096 , n6419 , n6899 );
nand ( n7097 , n7096 , n2849 );
nand ( n7098 , n7095 , n7097 );
and ( n7099 , n3770 , n5552 );
nor ( n7100 , n7099 , n2071 );
or ( n7101 , n7100 , n6934 );
not ( n7102 , n6412 );
or ( n7103 , n6425 , n7102 );
nand ( n7104 , n7103 , n1777 );
nand ( n7105 , n7101 , n7104 );
nor ( n7106 , n7098 , n7105 );
nand ( n7107 , n7094 , n7106 );
not ( n7108 , n6901 );
nor ( n7109 , n1378 , n7108 );
not ( n7110 , n7109 );
not ( n7111 , n3130 );
not ( n7112 , n6911 );
nand ( n7113 , n7112 , n6869 );
not ( n7114 , n7113 );
or ( n7115 , n7111 , n7114 );
not ( n7116 , n6700 );
not ( n7117 , n7116 );
or ( n7118 , n7117 , n6892 );
not ( n7119 , n7118 );
nand ( n7120 , n6876 , n6993 );
not ( n7121 , n7120 );
or ( n7122 , n7119 , n7121 );
not ( n7123 , n399 );
nand ( n7124 , n7122 , n7123 );
nand ( n7125 , n7115 , n7124 );
not ( n7126 , n7125 );
or ( n7127 , n7110 , n7126 );
not ( n7128 , n2876 );
nor ( n7129 , n7128 , n6284 );
not ( n7130 , n7129 );
or ( n7131 , n7130 , n7090 );
not ( n7132 , n2939 );
and ( n7133 , n7132 , n6901 , n6997 );
nand ( n7134 , n407 , n6699 );
and ( n7135 , n7134 , n6296 );
nor ( n7136 , n7135 , n2100 , n6902 );
nor ( n7137 , n7133 , n7136 );
nand ( n7138 , n7127 , n7131 , n7137 );
nand ( n7139 , n1763 , n6959 );
nor ( n7140 , n6944 , n7135 );
or ( n7141 , n7117 , n6953 );
not ( n7142 , n7141 );
nand ( n7143 , n6945 , n6993 );
not ( n7144 , n7143 );
or ( n7145 , n7142 , n7144 );
nand ( n7146 , n7145 , n399 );
not ( n7147 , n7146 );
nor ( n7148 , n7140 , n7147 );
or ( n7149 , n7139 , n7148 );
and ( n7150 , n1763 , n6909 );
nor ( n7151 , n7135 , n6915 );
not ( n7152 , n7151 );
not ( n7153 , n6920 );
nand ( n7154 , n7116 , n7153 );
not ( n7155 , n7154 );
not ( n7156 , n6454 );
not ( n7157 , n417 );
nand ( n7158 , n7157 , n6292 );
not ( n7159 , n7158 );
or ( n7160 , n7156 , n7159 );
nand ( n7161 , n7160 , n7087 );
not ( n7162 , n7161 );
or ( n7163 , n7155 , n7162 );
nand ( n7164 , n7163 , n399 );
nand ( n7165 , n7152 , n7164 );
and ( n7166 , n7150 , n7165 );
or ( n7167 , n6970 , n6558 );
or ( n7168 , n7041 , n7135 );
nand ( n7169 , n7167 , n6977 , n7168 );
and ( n7170 , n2814 , n7169 );
nor ( n7171 , n7166 , n7170 );
nor ( n7172 , n2935 , n7108 );
nand ( n7173 , n3130 , n7004 );
not ( n7174 , n7005 );
not ( n7175 , n402 );
nand ( n7176 , n7174 , n7175 , n7116 );
not ( n7177 , n7176 );
not ( n7178 , n6533 );
not ( n7179 , n7158 );
or ( n7180 , n7178 , n7179 );
nand ( n7181 , n7180 , n7087 );
not ( n7182 , n7181 );
or ( n7183 , n7177 , n7182 );
not ( n7184 , n399 );
nand ( n7185 , n7183 , n7184 );
nand ( n7186 , n7173 , n6873 , n7185 );
nand ( n7187 , n7172 , n7186 );
nand ( n7188 , n7149 , n7171 , n7187 );
nor ( n7189 , n7107 , n7138 , n7188 );
not ( n7190 , n7026 );
not ( n7191 , n2685 );
nand ( n7192 , n1959 , n6967 );
nor ( n7193 , n64 , n7192 );
not ( n7194 , n7193 );
not ( n7195 , n7186 );
or ( n7196 , n7194 , n7195 );
not ( n7197 , n64 );
and ( n7198 , n7197 , n7042 );
nand ( n7199 , n7198 , n7125 );
nand ( n7200 , n7196 , n7199 );
not ( n7201 , n7200 );
and ( n7202 , n7054 , n6638 );
and ( n7203 , n7058 , n6666 );
nor ( n7204 , n7202 , n7203 );
nand ( n7205 , n7201 , n7204 , n7052 );
not ( n7206 , n7205 );
or ( n7207 , n7191 , n7206 );
nand ( n7208 , n6971 , n6807 );
not ( n7209 , n7043 );
nor ( n7210 , n7209 , n7148 );
not ( n7211 , n7036 );
and ( n7212 , n7211 , n7165 );
nor ( n7213 , n7210 , n7212 );
nand ( n7214 , n7208 , n7035 , n7213 );
nand ( n7215 , n1763 , n7214 );
nand ( n7216 , n7207 , n7215 );
nand ( n7217 , n7190 , n7216 );
nand ( n7218 , n7080 , n7189 , n7217 );
nand ( n7219 , n1584 , n7218 );
not ( n7220 , n7139 );
not ( n7221 , n402 );
nand ( n7222 , n7221 , n7140 );
nor ( n7223 , n779 , n7134 );
not ( n7224 , n6940 );
and ( n7225 , n7223 , n7224 );
not ( n7226 , n6247 );
or ( n7227 , n3460 , n7226 );
not ( n7228 , n6698 );
and ( n7229 , n6435 , n7228 );
nor ( n7230 , n7229 , n6257 );
nand ( n7231 , n7227 , n7230 );
nor ( n7232 , n7225 , n7231 );
nand ( n7233 , n7222 , n7232 , n7146 );
not ( n7234 , n7233 );
not ( n7235 , n7234 );
and ( n7236 , n7220 , n7235 );
and ( n7237 , n7223 , n6913 );
buf ( n7238 , n7083 );
or ( n7239 , n3460 , n7238 );
nand ( n7240 , n7239 , n7230 );
nor ( n7241 , n7237 , n7240 );
not ( n7242 , n402 );
nand ( n7243 , n7242 , n7151 );
nand ( n7244 , n7164 , n7241 , n7243 );
and ( n7245 , n7150 , n7244 );
nor ( n7246 , n7236 , n7245 );
not ( n7247 , n402 );
not ( n7248 , n7247 );
not ( n7249 , n7006 );
or ( n7250 , n7248 , n7249 );
not ( n7251 , n6621 );
nand ( n7252 , n7250 , n7251 );
and ( n7253 , n6865 , n1546 , n7252 );
or ( n7254 , n2939 , n6996 );
nand ( n7255 , n7254 , n2070 );
buf ( n7256 , n7071 );
and ( n7257 , n7255 , n6901 , n7256 );
nor ( n7258 , n7253 , n7257 );
nand ( n7259 , n6796 , n7113 );
not ( n7260 , n779 );
not ( n7261 , n6869 );
and ( n7262 , n7260 , n7261 );
not ( n7263 , n6437 );
or ( n7264 , n7263 , n7226 );
and ( n7265 , n3471 , n6699 );
nor ( n7266 , n7265 , n6257 );
nand ( n7267 , n7264 , n7266 );
nor ( n7268 , n7262 , n7267 );
nand ( n7269 , n7259 , n7268 , n7124 );
and ( n7270 , n7109 , n7269 );
and ( n7271 , n7129 , n7089 );
and ( n7272 , n6701 , n7136 );
nor ( n7273 , n7271 , n7272 );
not ( n7274 , n6341 );
nor ( n7275 , n7274 , n6619 );
not ( n7276 , n7275 );
nand ( n7277 , n7276 , n3388 , n6311 , n6901 );
not ( n7278 , n358 );
nor ( n7279 , n7278 , n1777 );
nand ( n7280 , n7279 , n6899 );
nand ( n7281 , n7273 , n7277 , n7280 );
nor ( n7282 , n7270 , n7281 );
nand ( n7283 , n7246 , n7106 , n7258 , n7282 );
not ( n7284 , n3732 );
not ( n7285 , n6894 );
nor ( n7286 , n6623 , n7285 );
not ( n7287 , n402 );
nand ( n7288 , n7287 , n6895 );
nand ( n7289 , n7286 , n7268 , n7288 );
and ( n7290 , n7284 , n7289 );
not ( n7291 , n6955 );
nor ( n7292 , n6623 , n7291 );
not ( n7293 , n402 );
nand ( n7294 , n7293 , n6956 );
nand ( n7295 , n7292 , n7232 , n7294 );
not ( n7296 , n7295 );
nor ( n7297 , n1746 , n7296 );
nor ( n7298 , n7290 , n7297 );
or ( n7299 , n7108 , n7298 );
and ( n7300 , n6971 , n6274 );
not ( n7301 , n6977 );
nor ( n7302 , n7041 , n7011 );
nor ( n7303 , n7300 , n7301 , n7302 );
or ( n7304 , n2614 , n7303 );
or ( n7305 , n7108 , n7011 );
not ( n7306 , n6935 );
nand ( n7307 , n7304 , n7305 , n7306 );
nand ( n7308 , n2836 , n7307 );
nand ( n7309 , n7299 , n7308 );
not ( n7310 , n6929 );
nor ( n7311 , n6623 , n7310 );
not ( n7312 , n402 );
and ( n7313 , n7312 , n6930 );
not ( n7314 , n7241 );
nor ( n7315 , n7313 , n7314 );
nand ( n7316 , n7311 , n7315 );
nand ( n7317 , n7316 , n6865 , n1361 );
and ( n7318 , n6971 , n6678 );
nor ( n7319 , n7275 , n6968 );
nor ( n7320 , n7318 , n7319 , n6976 );
or ( n7321 , n1298 , n7320 );
not ( n7322 , n7072 );
and ( n7323 , n6971 , n6390 );
nor ( n7324 , n7323 , n6978 );
not ( n7325 , n7324 );
or ( n7326 , n7322 , n7325 );
nand ( n7327 , n7326 , n6384 );
nand ( n7328 , n7321 , n7327 );
or ( n7329 , n6970 , n6348 );
nand ( n7330 , n6967 , n6995 );
nand ( n7331 , n7329 , n7330 , n6977 );
nand ( n7332 , n1800 , n7331 );
nand ( n7333 , n6967 , n7089 );
and ( n7334 , n6971 , n6371 );
nor ( n7335 , n7334 , n6974 );
nand ( n7336 , n7333 , n7335 );
and ( n7337 , n1807 , n7336 );
or ( n7338 , n6970 , n6705 );
not ( n7339 , n7168 );
nand ( n7340 , n7339 , n6701 );
nand ( n7341 , n7338 , n7340 , n6975 );
and ( n7342 , n7341 , n1947 );
nor ( n7343 , n7337 , n7342 );
nand ( n7344 , n7332 , n7343 );
or ( n7345 , n7328 , n7344 );
nand ( n7346 , n7345 , n329 );
nand ( n7347 , n7317 , n7346 );
nor ( n7348 , n7283 , n7309 , n7347 );
not ( n7349 , n402 );
not ( n7350 , n7349 );
not ( n7351 , n7186 );
or ( n7352 , n7350 , n7351 );
and ( n7353 , n780 , n7004 );
not ( n7354 , n6495 );
not ( n7355 , n7238 );
and ( n7356 , n7354 , n7355 );
nor ( n7357 , n7353 , n7356 );
and ( n7358 , n7357 , n7266 , n7185 );
nand ( n7359 , n7352 , n7358 );
nand ( n7360 , n7172 , n7359 );
not ( n7361 , n7026 );
not ( n7362 , n1763 );
nand ( n7363 , n6971 , n6606 );
and ( n7364 , n7043 , n7233 );
not ( n7365 , n7244 );
nor ( n7366 , n7365 , n7036 );
nor ( n7367 , n7364 , n7366 );
nand ( n7368 , n7035 , n7363 , n7367 );
not ( n7369 , n7368 );
or ( n7370 , n7362 , n7369 );
nand ( n7371 , n7198 , n7289 );
and ( n7372 , n7058 , n6690 );
not ( n7373 , n7054 );
nor ( n7374 , n7373 , n6551 );
nor ( n7375 , n7372 , n7374 );
nand ( n7376 , n7193 , n7252 );
and ( n7377 , n7375 , n7052 , n7376 );
nand ( n7378 , n7371 , n7377 );
nand ( n7379 , n1260 , n7378 );
nand ( n7380 , n7370 , n7379 );
not ( n7381 , n7380 );
and ( n7382 , n7031 , n6461 );
nor ( n7383 , n7028 , n6498 );
nor ( n7384 , n7382 , n7383 );
and ( n7385 , n7043 , n7295 );
not ( n7386 , n7316 );
nor ( n7387 , n7036 , n7386 );
nor ( n7388 , n7385 , n7387 );
nand ( n7389 , n7384 , n7035 , n7388 );
nand ( n7390 , n1359 , n7389 );
not ( n7391 , n7193 );
not ( n7392 , n7359 );
or ( n7393 , n7391 , n7392 );
nand ( n7394 , n7198 , n7269 );
nand ( n7395 , n7393 , n7394 );
not ( n7396 , n7395 );
not ( n7397 , n6670 );
not ( n7398 , n7397 );
not ( n7399 , n7059 );
and ( n7400 , n7398 , n7399 );
and ( n7401 , n7054 , n6640 );
nor ( n7402 , n7400 , n7401 );
nand ( n7403 , n7396 , n7402 , n7052 );
nand ( n7404 , n7403 , n2685 );
nand ( n7405 , n7381 , n7390 , n7404 );
nand ( n7406 , n7361 , n7405 );
nand ( n7407 , n7348 , n7360 , n7406 );
nand ( n7408 , n7407 , n2029 );
and ( n7409 , n7024 , n7067 , n7219 , n7408 );
or ( n7410 , n6838 , n7409 );
not ( n7411 , n6810 );
and ( n7412 , n6789 , n6519 );
nor ( n7413 , n7412 , n1358 );
nor ( n7414 , n7411 , n7413 );
or ( n7415 , n2596 , n7414 );
not ( n7416 , n358 );
and ( n7417 , n2600 , n6731 );
and ( n7418 , n2606 , n6826 );
nor ( n7419 , n7417 , n7418 );
not ( n7420 , n7419 );
and ( n7421 , n7416 , n7420 );
not ( n7422 , n6719 );
and ( n7423 , n3195 , n7422 );
and ( n7424 , n2857 , n6738 );
nor ( n7425 , n7423 , n7424 );
nand ( n7426 , n329 , n1553 , n6756 );
not ( n7427 , n6561 );
and ( n7428 , n2814 , n7427 );
and ( n7429 , n2629 , n6747 );
nor ( n7430 , n7428 , n7429 );
and ( n7431 , n2886 , n6816 );
nor ( n7432 , n7431 , n6520 );
nand ( n7433 , n7425 , n7426 , n7430 , n7432 );
nor ( n7434 , n7421 , n7433 );
nand ( n7435 , n7415 , n7434 );
nand ( n7436 , n372 , n1661 , n2984 , n7435 );
nand ( n7437 , n7410 , n7436 );
nand ( n7438 , n2995 , n7437 );
nand ( n7439 , n6515 , n6973 );
nand ( n7440 , n5510 , n7439 );
and ( n7441 , n6412 , n7440 );
or ( n7442 , n1545 , n7441 );
not ( n7443 , n3900 );
not ( n7444 , n1959 );
not ( n7445 , n7439 );
or ( n7446 , n7444 , n7445 );
nand ( n7447 , n7446 , n6426 );
nand ( n7448 , n7443 , n7447 );
nand ( n7449 , n7442 , n7448 );
or ( n7450 , n1946 , n7168 );
or ( n7451 , n2945 , n7092 );
not ( n7452 , n7447 );
nand ( n7453 , n7441 , n7452 );
and ( n7454 , n1960 , n7453 );
nand ( n7455 , n1069 , n7439 );
and ( n7456 , n6611 , n7455 );
or ( n7457 , n2100 , n7456 );
or ( n7458 , n1740 , n7452 );
nand ( n7459 , n7457 , n7458 );
nor ( n7460 , n7454 , n7459 );
nand ( n7461 , n7450 , n7451 , n7460 );
nor ( n7462 , n7449 , n7461 );
nand ( n7463 , n7198 , n6997 );
nand ( n7464 , n7441 , n7463 , n7213 );
and ( n7465 , n1763 , n7464 );
and ( n7466 , n2685 , n7200 );
nor ( n7467 , n7465 , n7466 );
nand ( n7468 , n7462 , n7467 );
and ( n7469 , n4759 , n7468 );
nor ( n7470 , n4684 , n6863 );
not ( n7471 , n7456 );
and ( n7472 , n7470 , n7471 );
nor ( n7473 , n4684 , n6963 );
not ( n7474 , n7441 );
and ( n7475 , n7473 , n7474 );
nor ( n7476 , n7472 , n7475 );
not ( n7477 , n6968 );
nand ( n7478 , n7477 , n4759 , n1538 );
not ( n7479 , n6516 );
or ( n7480 , n2551 , n7479 );
nand ( n7481 , n7480 , n6519 );
and ( n7482 , n4756 , n7481 );
not ( n7483 , n64 );
nand ( n7484 , n7483 , n7470 );
nand ( n7485 , n64 , n7473 );
and ( n7486 , n7484 , n7485 );
nor ( n7487 , n7486 , n7452 );
nor ( n7488 , n7482 , n7487 );
nand ( n7489 , n7476 , n7478 , n7488 );
not ( n7490 , n7485 );
not ( n7491 , n7038 );
and ( n7492 , n7490 , n7491 );
not ( n7493 , n7484 );
and ( n7494 , n7493 , n7006 );
nor ( n7495 , n7492 , n7494 );
or ( n7496 , n7192 , n7495 );
not ( n7497 , n2096 );
not ( n7498 , n7019 );
and ( n7499 , n7497 , n7498 );
not ( n7500 , n7042 );
nor ( n7501 , n7500 , n2070 );
not ( n7502 , n6998 );
and ( n7503 , n7501 , n7502 );
nor ( n7504 , n7499 , n7503 );
or ( n7505 , n4758 , n7504 );
nand ( n7506 , n7496 , n7505 );
nor ( n7507 , n7469 , n7489 , n7506 );
not ( n7508 , n6895 );
or ( n7509 , n7484 , n7508 );
or ( n7510 , n7485 , n6957 );
nand ( n7511 , n7509 , n7510 );
nand ( n7512 , n7042 , n7511 );
and ( n7513 , n2691 , n7453 );
and ( n7514 , n7501 , n7256 );
not ( n7515 , n1538 );
not ( n7516 , n7319 );
or ( n7517 , n7515 , n7516 );
or ( n7518 , n1946 , n7340 );
nand ( n7519 , n7517 , n7518 );
nor ( n7520 , n7513 , n7514 , n7519 );
not ( n7521 , n3393 );
and ( n7522 , n7521 , n7474 );
and ( n7523 , n7497 , n7302 );
nor ( n7524 , n7522 , n7523 );
not ( n7525 , n7367 );
nand ( n7526 , n1763 , n7525 );
nand ( n7527 , n2685 , n7395 );
nand ( n7528 , n7520 , n7524 , n7526 , n7527 );
not ( n7529 , n7388 );
and ( n7530 , n1359 , n7529 );
nand ( n7531 , n7448 , n7460 );
nor ( n7532 , n7530 , n7531 );
not ( n7533 , n7333 );
nand ( n7534 , n1807 , n7533 );
or ( n7535 , n2166 , n7330 );
and ( n7536 , n7452 , n7376 );
nand ( n7537 , n7536 , n7456 , n7371 );
nand ( n7538 , n1260 , n7537 );
nand ( n7539 , n7532 , n7534 , n7535 , n7538 );
or ( n7540 , n7528 , n7539 );
nand ( n7541 , n7540 , n4685 );
nand ( n7542 , n7507 , n7512 , n7541 );
and ( n7543 , n2987 , n7542 );
and ( n7544 , n4242 , n6734 );
and ( n7545 , n2106 , n6749 );
nor ( n7546 , n7544 , n7545 );
or ( n7547 , n2166 , n6356 );
and ( n7548 , n1807 , n6379 );
not ( n7549 , n7497 );
not ( n7550 , n6318 );
or ( n7551 , n7549 , n7550 );
nand ( n7552 , n1778 , n1740 , n6427 );
nand ( n7553 , n7551 , n7552 );
nor ( n7554 , n7548 , n7553 );
nand ( n7555 , n7547 , n7554 , n1464 );
nor ( n7556 , n7555 , n6507 );
not ( n7557 , n7556 );
not ( n7558 , n6714 );
not ( n7559 , n7558 );
or ( n7560 , n7557 , n7559 );
and ( n7561 , n1380 , n6721 );
and ( n7562 , n6830 , n6427 );
nor ( n7563 , n7561 , n7562 );
nand ( n7564 , n372 , n6833 , n7563 , n6812 );
nand ( n7565 , n7560 , n7564 );
and ( n7566 , n7546 , n7565 );
nand ( n7567 , n393 , n395 );
not ( n7568 , n7567 );
xor ( n7569 , n1734 , n7568 );
nand ( n7570 , n714 , n7569 );
nor ( n7571 , n3001 , n7570 );
nand ( n7572 , n4684 , n7571 );
nor ( n7573 , n7566 , n7572 );
nor ( n7574 , n7543 , n7573 );
or ( n7575 , n2945 , n7093 );
not ( n7576 , n7216 );
nand ( n7577 , n7575 , n7576 );
nand ( n7578 , n1584 , n7577 );
not ( n7579 , n7344 );
nor ( n7580 , n358 , n2926 );
nand ( n7581 , n7580 , n6427 );
not ( n7582 , n7405 );
nand ( n7583 , n7579 , n7581 , n7582 );
nand ( n7584 , n2029 , n7583 );
not ( n7585 , n2096 );
not ( n7586 , n7303 );
and ( n7587 , n7585 , n7586 );
nor ( n7588 , n7587 , n7328 );
or ( n7589 , n7588 , n372 );
nand ( n7590 , n4242 , n7078 );
nand ( n7591 , n7589 , n7590 , n403 );
nand ( n7592 , n372 , n1947 );
or ( n7593 , n7592 , n6561 );
and ( n7594 , n6208 , n6738 );
and ( n7595 , n2106 , n6747 );
nor ( n7596 , n7594 , n7595 , n403 );
and ( n7597 , n311 , n6826 );
not ( n7598 , n311 );
and ( n7599 , n7598 , n6731 );
nor ( n7600 , n7597 , n7599 );
or ( n7601 , n7600 , n358 , n720 );
or ( n7602 , n1379 , n6719 );
nand ( n7603 , n7601 , n7602 );
and ( n7604 , n372 , n7603 );
nor ( n7605 , n2660 , n2282 );
and ( n7606 , n7605 , n6756 );
nor ( n7607 , n7604 , n7606 );
nand ( n7608 , n7593 , n7596 , n7607 );
and ( n7609 , n7591 , n7608 );
nor ( n7610 , n7609 , n7066 );
and ( n7611 , n6984 , n7075 );
or ( n7612 , n7414 , n2408 );
and ( n7613 , n7169 , n1584 , n1947 );
and ( n7614 , n24 , n2407 );
not ( n7615 , n6963 );
nor ( n7616 , n7614 , n7615 );
or ( n7617 , n64 , n7616 );
not ( n7618 , n7580 );
nand ( n7619 , n7618 , n3389 );
and ( n7620 , n372 , n7619 );
and ( n7621 , n2029 , n7279 );
nor ( n7622 , n7620 , n7621 );
nand ( n7623 , n7617 , n7622 );
and ( n7624 , n7623 , n6427 );
nor ( n7625 , n7613 , n7624 );
and ( n7626 , n2407 , n1961 , n6816 );
nor ( n7627 , n7626 , n6981 );
nand ( n7628 , n7612 , n7625 , n7627 );
nor ( n7629 , n7009 , n7020 );
nor ( n7630 , n7611 , n7628 , n7629 );
not ( n7631 , n6305 );
nand ( n7632 , n7631 , n7497 );
nand ( n7633 , n6858 , n7632 , n7552 );
nand ( n7634 , n2023 , n7633 );
and ( n7635 , n7610 , n7630 , n7634 );
nand ( n7636 , n7578 , n7584 , n7635 );
not ( n7637 , n4684 );
nand ( n7638 , n7636 , n7637 , n7571 );
and ( n7639 , n394 , n2977 );
nor ( n7640 , n6207 , n7572 , n6741 );
not ( n7641 , n7605 );
nor ( n7642 , n7641 , n7572 , n6758 );
nor ( n7643 , n7639 , n7640 , n7642 );
nand ( n7644 , n7438 , n7574 , n7638 , n7643 );
not ( n7645 , n396 );
not ( n7646 , n6320 );
or ( n7647 , n7645 , n7646 );
nand ( n7648 , n7647 , n793 );
not ( n7649 , n6126 );
nor ( n7650 , n5222 , n5234 );
not ( n7651 , n7650 );
or ( n7652 , n7649 , n7651 );
nand ( n7653 , n7652 , n6523 );
not ( n7654 , n7653 );
or ( n7655 , n7648 , n7654 );
nand ( n7656 , n396 , n5236 );
or ( n7657 , n386 , n7656 );
and ( n7658 , n396 , n793 );
nand ( n7659 , n390 , n7658 );
nand ( n7660 , n7655 , n7657 , n7659 );
and ( n7661 , n1925 , n7660 );
nand ( n7662 , n396 , n5296 );
or ( n7663 , n386 , n7662 );
not ( n7664 , n7648 );
buf ( n7665 , n1206 );
nand ( n7666 , n7665 , n5293 );
or ( n7667 , n5282 , n7666 );
nand ( n7668 , n7667 , n6523 );
nand ( n7669 , n7664 , n7668 );
nand ( n7670 , n7663 , n7659 , n7669 );
and ( n7671 , n1961 , n7670 );
nor ( n7672 , n7661 , n7671 );
or ( n7673 , n793 , n1855 );
nor ( n7674 , n1412 , n7673 );
nand ( n7675 , n6523 , n6128 );
nand ( n7676 , n7674 , n7675 );
and ( n7677 , n281 , n3068 );
not ( n7678 , n7677 );
or ( n7679 , n7678 , n5374 );
nand ( n7680 , n265 , n396 );
not ( n7681 , n7680 );
nand ( n7682 , n7679 , n7681 );
nand ( n7683 , n396 , n6129 );
nand ( n7684 , n7683 , n5133 , n7675 );
nand ( n7685 , n7676 , n7682 , n7684 );
and ( n7686 , n3730 , n7685 );
nor ( n7687 , n6523 , n5671 );
and ( n7688 , n7132 , n7687 );
nor ( n7689 , n7686 , n7688 );
and ( n7690 , n7677 , n5433 );
nor ( n7691 , n7690 , n7680 );
not ( n7692 , n7674 );
nand ( n7693 , n396 , n5952 );
or ( n7694 , n1937 , n7693 );
nand ( n7695 , n7694 , n5133 );
and ( n7696 , n7692 , n7695 );
nor ( n7697 , n396 , n6067 );
nor ( n7698 , n7696 , n7697 );
nor ( n7699 , n7691 , n7698 );
not ( n7700 , n7699 );
nand ( n7701 , n7700 , n7284 );
or ( n7702 , n7678 , n5523 );
nand ( n7703 , n7702 , n7681 );
not ( n7704 , n7692 );
nand ( n7705 , n396 , n5971 );
or ( n7706 , n6043 , n7705 );
nand ( n7707 , n7706 , n5133 );
not ( n7708 , n7707 );
or ( n7709 , n7704 , n7708 );
nand ( n7710 , n6523 , n6045 );
nand ( n7711 , n7709 , n7710 );
nand ( n7712 , n7703 , n7711 );
and ( n7713 , n3731 , n7712 );
and ( n7714 , n5948 , n5066 );
nor ( n7715 , n7714 , n396 );
or ( n7716 , n7648 , n7715 );
or ( n7717 , n390 , n5065 );
nand ( n7718 , n7717 , n7658 );
nand ( n7719 , n7716 , n7718 );
and ( n7720 , n1361 , n7719 );
nand ( n7721 , n6523 , n6116 );
not ( n7722 , n7721 );
or ( n7723 , n7648 , n7722 );
nor ( n7724 , n6523 , n5189 );
not ( n7725 , n7724 );
or ( n7726 , n386 , n7725 );
nand ( n7727 , n7723 , n7726 , n7659 );
and ( n7728 , n1807 , n7727 );
nor ( n7729 , n7720 , n7728 );
or ( n7730 , n396 , n6197 );
not ( n7731 , n7730 );
or ( n7732 , n7648 , n7731 );
nand ( n7733 , n396 , n5546 );
or ( n7734 , n386 , n7733 );
nand ( n7735 , n7732 , n7734 , n7659 );
and ( n7736 , n7497 , n7735 );
and ( n7737 , n6523 , n6100 );
or ( n7738 , n7648 , n7737 );
nand ( n7739 , n793 , n7687 );
nand ( n7740 , n7738 , n7659 , n7739 );
and ( n7741 , n1800 , n7740 );
nor ( n7742 , n7736 , n7741 );
not ( n7743 , n5948 );
or ( n7744 , n7743 , n4977 );
nand ( n7745 , n7744 , n6523 );
not ( n7746 , n7745 );
or ( n7747 , n7648 , n7746 );
nand ( n7748 , n396 , n6058 );
nand ( n7749 , n7747 , n7659 , n7748 );
and ( n7750 , n1546 , n7749 );
and ( n7751 , n6523 , n6078 );
or ( n7752 , n7648 , n7751 );
nand ( n7753 , n396 , n5573 );
or ( n7754 , n386 , n7753 );
nand ( n7755 , n7752 , n7754 , n7659 );
and ( n7756 , n6384 , n7755 );
nor ( n7757 , n7750 , n7756 );
and ( n7758 , n7729 , n7742 , n7757 );
not ( n7759 , n1746 );
not ( n7760 , n5600 );
or ( n7761 , n7678 , n7760 );
nand ( n7762 , n7761 , n7681 );
nand ( n7763 , n396 , n6011 );
not ( n7764 , n7763 );
and ( n7765 , n7764 , n5372 );
nor ( n7766 , n7765 , n5942 );
or ( n7767 , n7674 , n7766 );
not ( n7768 , n6093 );
nand ( n7769 , n7768 , n6523 );
nand ( n7770 , n7767 , n7769 );
nand ( n7771 , n7762 , n7770 );
and ( n7772 , n7759 , n7771 );
nand ( n7773 , n2690 , n1741 );
or ( n7774 , n7773 , n7650 );
nor ( n7775 , n6523 , n265 );
or ( n7776 , n7775 , n2935 );
or ( n7777 , n7776 , n6053 );
not ( n7778 , n6061 );
not ( n7779 , n2938 );
not ( n7780 , n2844 );
and ( n7781 , n7779 , n7780 );
nor ( n7782 , n7781 , n7677 );
nor ( n7783 , n7778 , n7782 );
not ( n7784 , n358 );
nor ( n7785 , n7784 , n7775 );
nand ( n7786 , n2906 , n7785 , n5065 );
and ( n7787 , n7783 , n265 , n7786 );
nand ( n7788 , n7774 , n7777 , n7787 );
nand ( n7789 , n396 , n7788 );
not ( n7790 , n2070 );
not ( n7791 , n7753 );
and ( n7792 , n7790 , n7791 );
nand ( n7793 , n7785 , n1137 );
not ( n7794 , n7793 );
nor ( n7795 , n6523 , n4978 );
and ( n7796 , n7794 , n7795 );
nor ( n7797 , n7792 , n7796 );
nor ( n7798 , n1946 , n7648 );
nand ( n7799 , n6523 , n1212 );
nand ( n7800 , n7798 , n7799 );
not ( n7801 , n2836 );
nor ( n7802 , n7680 , n7801 );
and ( n7803 , n7802 , n5546 );
or ( n7804 , n6523 , n1945 , n5531 );
and ( n7805 , n3388 , n7674 );
nor ( n7806 , n1298 , n7648 );
nor ( n7807 , n7805 , n7806 );
not ( n7808 , n5642 );
nand ( n7809 , n5991 , n7808 );
and ( n7810 , n6523 , n7809 );
or ( n7811 , n7807 , n7810 );
nand ( n7812 , n7804 , n7811 );
nand ( n7813 , n265 , n3729 );
nor ( n7814 , n7813 , n7725 );
nor ( n7815 , n7803 , n7812 , n7814 );
nand ( n7816 , n7789 , n7797 , n7800 , n7815 );
not ( n7817 , n2070 );
not ( n7818 , n7751 );
and ( n7819 , n7817 , n7818 );
and ( n7820 , n2836 , n7730 );
nor ( n7821 , n7819 , n7820 );
nand ( n7822 , n3729 , n7721 );
and ( n7823 , n5480 , n7799 );
nor ( n7824 , n2939 , n7737 );
nor ( n7825 , n7823 , n7824 );
nand ( n7826 , n7822 , n7825 );
not ( n7827 , n7826 );
and ( n7828 , n7821 , n7827 );
nor ( n7829 , n7828 , n7692 );
nor ( n7830 , n7772 , n7816 , n7829 );
nand ( n7831 , n7758 , n7830 );
nor ( n7832 , n1924 , n7654 );
not ( n7833 , n7832 );
nand ( n7834 , n1546 , n7745 );
nor ( n7835 , n1362 , n7715 );
not ( n7836 , n7835 );
nand ( n7837 , n1961 , n7668 );
and ( n7838 , n7834 , n7836 , n7837 );
and ( n7839 , n7833 , n7838 );
nor ( n7840 , n7839 , n7673 );
nor ( n7841 , n7713 , n7831 , n7840 );
nand ( n7842 , n7672 , n7689 , n7701 , n7841 );
and ( n7843 , n7842 , n4685 , n3004 );
nand ( n7844 , n6523 , n6196 );
and ( n7845 , n2836 , n7844 );
nor ( n7846 , n396 , n6025 );
or ( n7847 , n2070 , n7846 );
and ( n7848 , n6523 , n7666 );
or ( n7849 , n2935 , n7848 );
nand ( n7850 , n7847 , n7849 );
nor ( n7851 , n7845 , n7850 );
or ( n7852 , n396 , n7665 );
nand ( n7853 , n5480 , n7852 );
not ( n7854 , n358 );
not ( n7855 , n5553 );
nand ( n7856 , n6523 , n6170 );
not ( n7857 , n7856 );
or ( n7858 , n7855 , n7857 );
nand ( n7859 , n6523 , n6001 );
nand ( n7860 , n2938 , n7859 );
nand ( n7861 , n7858 , n7860 );
nand ( n7862 , n7854 , n7861 );
nand ( n7863 , n7851 , n7853 , n7862 );
and ( n7864 , n2550 , n7863 );
and ( n7865 , n5991 , n5064 );
nor ( n7866 , n7865 , n396 );
or ( n7867 , n1362 , n7866 );
nand ( n7868 , n5947 , n4976 );
nand ( n7869 , n6523 , n7868 );
nand ( n7870 , n1546 , n7869 );
nand ( n7871 , n7867 , n7870 );
not ( n7872 , n7871 );
and ( n7873 , n5948 , n5870 );
nor ( n7874 , n7873 , n396 );
or ( n7875 , n1924 , n7874 );
nand ( n7876 , n7872 , n7875 );
nor ( n7877 , n7864 , n7876 );
or ( n7878 , n7673 , n7877 );
nor ( n7879 , n396 , n5952 );
not ( n7880 , n7879 );
nand ( n7881 , n7880 , n7674 );
or ( n7882 , n7678 , n5432 );
nand ( n7883 , n7882 , n7681 );
not ( n7884 , n7879 );
nand ( n7885 , n7884 , n7693 , n5133 );
and ( n7886 , n7881 , n7883 , n7885 );
or ( n7887 , n3732 , n7886 );
nand ( n7888 , n7878 , n7887 );
and ( n7889 , n6523 , n5970 );
or ( n7890 , n7692 , n7889 );
or ( n7891 , n7678 , n5520 );
nand ( n7892 , n7891 , n7681 );
not ( n7893 , n7889 );
nand ( n7894 , n7893 , n7705 , n5133 );
nand ( n7895 , n7890 , n7892 , n7894 );
and ( n7896 , n3731 , n7895 );
not ( n7897 , n358 );
not ( n7898 , n7897 );
not ( n7899 , n1013 );
or ( n7900 , n7648 , n7874 );
nand ( n7901 , n396 , n5231 );
or ( n7902 , n386 , n7901 );
nand ( n7903 , n7900 , n7902 , n7659 );
not ( n7904 , n7903 );
or ( n7905 , n7899 , n7904 );
not ( n7906 , n7664 );
not ( n7907 , n7856 );
or ( n7908 , n7906 , n7907 );
or ( n7909 , n390 , n5861 );
nand ( n7910 , n7909 , n7658 );
nand ( n7911 , n7908 , n7910 );
nand ( n7912 , n2136 , n7911 );
nand ( n7913 , n7905 , n7912 );
not ( n7914 , n7913 );
or ( n7915 , n7898 , n7914 );
nand ( n7916 , n6523 , n5992 );
nand ( n7917 , n7674 , n7916 );
not ( n7918 , n7677 );
not ( n7919 , n5369 );
or ( n7920 , n7918 , n7919 );
nand ( n7921 , n7920 , n7681 );
nor ( n7922 , n6523 , n5992 );
not ( n7923 , n7922 );
nand ( n7924 , n7923 , n5133 , n7916 );
nand ( n7925 , n7917 , n7921 , n7924 );
and ( n7926 , n3730 , n7925 );
nand ( n7927 , n396 , n5708 );
nor ( n7928 , n2939 , n7927 );
nor ( n7929 , n7926 , n7928 );
nand ( n7930 , n7915 , n7929 );
nor ( n7931 , n7896 , n7930 );
and ( n7932 , n7664 , n7871 );
not ( n7933 , n396 );
not ( n7934 , n6209 );
or ( n7935 , n7933 , n7934 );
nand ( n7936 , n7935 , n7659 );
and ( n7937 , n1546 , n7936 );
nor ( n7938 , n7932 , n7937 );
or ( n7939 , n7648 , n7846 );
nand ( n7940 , n396 , n5767 );
or ( n7941 , n386 , n7940 );
nand ( n7942 , n7939 , n7941 , n7659 );
and ( n7943 , n6384 , n7942 );
nor ( n7944 , n6523 , n5064 );
nand ( n7945 , n793 , n7944 );
and ( n7946 , n7659 , n7945 );
nor ( n7947 , n7946 , n1362 );
nor ( n7948 , n7943 , n7947 );
nand ( n7949 , n7938 , n7948 );
not ( n7950 , n7759 );
nand ( n7951 , n6523 , n6010 );
nand ( n7952 , n7674 , n7951 );
or ( n7953 , n7678 , n5599 );
nand ( n7954 , n7953 , n7681 );
nand ( n7955 , n7763 , n5133 , n7951 );
nand ( n7956 , n7952 , n7954 , n7955 );
not ( n7957 , n7956 );
or ( n7958 , n7950 , n7957 );
not ( n7959 , n6523 );
not ( n7960 , n358 );
nand ( n7961 , n414 , n7960 );
or ( n7962 , n746 , n7961 );
nand ( n7963 , n7962 , n5797 );
and ( n7964 , n2849 , n7963 );
or ( n7965 , n7793 , n5938 );
or ( n7966 , n7776 , n5295 );
nand ( n7967 , n7965 , n7966 , n5262 );
nor ( n7968 , n7964 , n7967 , n7782 );
not ( n7969 , n7968 );
and ( n7970 , n7959 , n7969 );
not ( n7971 , n358 );
not ( n7972 , n386 );
not ( n7973 , n7927 );
and ( n7974 , n7972 , n7973 );
and ( n7975 , n7664 , n7859 );
nor ( n7976 , n7974 , n7975 );
and ( n7977 , n7659 , n7976 );
nor ( n7978 , n7977 , n1345 );
and ( n7979 , n7971 , n7978 );
nor ( n7980 , n7970 , n7979 );
nand ( n7981 , n7958 , n7980 );
or ( n7982 , n7648 , n7848 );
or ( n7983 , n390 , n5294 );
nand ( n7984 , n7983 , n7658 );
nand ( n7985 , n7982 , n7984 );
nand ( n7986 , n1961 , n7985 );
and ( n7987 , n2692 , n7944 );
or ( n7988 , n7773 , n7901 );
or ( n7989 , n2070 , n7940 );
nand ( n7990 , n7988 , n7989 );
nor ( n7991 , n7987 , n7990 );
and ( n7992 , n7798 , n7852 );
or ( n7993 , n1068 , n7659 );
not ( n7994 , n7775 );
nand ( n7995 , n7993 , n7994 );
and ( n7996 , n2685 , n7995 );
nor ( n7997 , n7992 , n7996 );
not ( n7998 , n6196 );
and ( n7999 , n396 , n7998 );
nor ( n8000 , n7999 , n5942 );
and ( n8001 , n8000 , n7845 );
and ( n8002 , n7802 , n6015 );
nand ( n8003 , n5544 , n7724 );
or ( n8004 , n7813 , n8003 );
not ( n8005 , n7995 );
or ( n8006 , n1297 , n8005 );
and ( n8007 , n6523 , n1203 );
or ( n8008 , n8007 , n7807 );
nand ( n8009 , n8004 , n8006 , n8008 );
nor ( n8010 , n8001 , n8002 , n8009 );
nand ( n8011 , n7986 , n7991 , n7997 , n8010 );
nor ( n8012 , n7949 , n7981 , n8011 );
nand ( n8013 , n7931 , n8012 );
nor ( n8014 , n7888 , n8013 );
or ( n8015 , n8014 , n4758 , n3003 );
or ( n8016 , n6523 , n2986 );
nand ( n8017 , n8015 , n8016 );
nor ( n8018 , n7843 , n8017 );
not ( n8019 , n724 );
not ( n8020 , n8019 );
not ( n8021 , n8020 );
nand ( n8022 , n8021 , n5971 );
and ( n8023 , n8022 , n2226 , n1246 );
and ( n8024 , n8019 , n1074 );
not ( n8025 , n5599 );
and ( n8026 , n8024 , n8025 );
nor ( n8027 , n8026 , n1105 );
and ( n8028 , n7473 , n8027 );
and ( n8029 , n8021 , n1202 );
nor ( n8030 , n8029 , n2105 );
nor ( n8031 , n8028 , n8030 );
or ( n8032 , n2226 , n1770 );
not ( n8033 , n2549 );
nand ( n8034 , n8032 , n8033 );
nand ( n8035 , n8031 , n4757 , n8034 );
nor ( n8036 , n8023 , n8035 );
or ( n8037 , n6523 , n8036 );
not ( n8038 , n2548 );
not ( n8039 , n2109 );
or ( n8040 , n6523 , n8024 );
not ( n8041 , n8040 );
nor ( n8042 , n8041 , n7795 );
or ( n8043 , n1251 , n8039 , n8042 );
nor ( n8044 , n8041 , n7944 );
or ( n8045 , n6190 , n8044 );
nand ( n8046 , n8043 , n8045 );
and ( n8047 , n8038 , n8046 );
not ( n8048 , n8024 );
not ( n8049 , n5523 );
not ( n8050 , n8049 );
or ( n8051 , n8048 , n8050 );
nand ( n8052 , n8051 , n396 );
or ( n8053 , n2120 , n2282 , n8052 );
nand ( n8054 , n8040 , n7733 );
nand ( n8055 , n2065 , n8054 );
nand ( n8056 , n8053 , n8055 );
and ( n8057 , n8040 , n7725 );
not ( n8058 , n2228 );
nor ( n8059 , n8057 , n8058 );
nor ( n8060 , n8047 , n8056 , n8059 );
nand ( n8061 , n8040 , n7753 );
and ( n8062 , n2073 , n8061 );
nor ( n8063 , n6523 , n1021 );
and ( n8064 , n8063 , n2101 );
nor ( n8065 , n8062 , n8064 );
not ( n8066 , n8021 );
or ( n8067 , n8066 , n7868 );
nand ( n8068 , n8067 , n396 );
or ( n8069 , n6207 , n8068 );
nand ( n8070 , n8024 , n5295 );
nand ( n8071 , n396 , n2226 , n1138 , n8070 );
nand ( n8072 , n8060 , n8065 , n8069 , n8071 );
and ( n8073 , n8021 , n6129 );
nor ( n8074 , n8073 , n6523 );
and ( n8075 , n2174 , n8074 );
nand ( n8076 , n8024 , n5950 );
and ( n8077 , n396 , n8076 );
and ( n8078 , n7605 , n8077 );
nor ( n8079 , n8075 , n8078 );
not ( n8080 , n766 );
not ( n8081 , n721 );
or ( n8082 , n8080 , n8081 );
nand ( n8083 , n8082 , n396 );
and ( n8084 , n6320 , n8083 );
nand ( n8085 , n8084 , n7650 );
and ( n8086 , n1464 , n8085 , n7832 );
nand ( n8087 , n8084 , n5066 );
and ( n8088 , n1464 , n8087 , n7835 );
nor ( n8089 , n8086 , n8088 );
nand ( n8090 , n8079 , n8089 );
not ( n8091 , n1212 );
and ( n8092 , n8021 , n8091 );
nor ( n8093 , n8092 , n6523 );
nand ( n8094 , n1464 , n1947 , n8093 );
nand ( n8095 , n8040 , n8003 );
and ( n8096 , n1807 , n8095 );
or ( n8097 , n6308 , n6015 );
nand ( n8098 , n8097 , n396 );
nand ( n8099 , n8083 , n8098 );
and ( n8100 , n7497 , n8099 );
nor ( n8101 , n8096 , n8100 );
not ( n8102 , n8101 );
not ( n8103 , n8021 );
not ( n8104 , n5993 );
or ( n8105 , n8103 , n8104 );
nand ( n8106 , n8105 , n1743 );
and ( n8107 , n2166 , n8106 );
nand ( n8108 , n1743 , n5992 );
and ( n8109 , n8021 , n8108 , n6002 );
nor ( n8110 , n8107 , n8109 );
and ( n8111 , n396 , n8110 );
nor ( n8112 , n8111 , n1464 );
not ( n8113 , n8112 );
or ( n8114 , n8102 , n8113 );
and ( n8115 , n8084 , n6053 );
or ( n8116 , n8115 , n7837 );
or ( n8117 , n1937 , n8076 );
nand ( n8118 , n8117 , n396 );
or ( n8119 , n1554 , n8118 );
nand ( n8120 , n8116 , n8119 , n1464 );
nand ( n8121 , n8114 , n8120 );
and ( n8122 , n8024 , n7808 );
nand ( n8123 , n396 , n1759 );
nor ( n8124 , n8122 , n8123 , n1217 );
not ( n8125 , n7852 );
and ( n8126 , n8084 , n5286 );
nor ( n8127 , n7592 , n8125 , n8126 );
nor ( n8128 , n8124 , n8127 );
not ( n8129 , n2224 );
nor ( n8130 , n8041 , n7687 );
not ( n8131 , n8130 );
and ( n8132 , n8129 , n8131 );
and ( n8133 , n8021 , n6093 );
nor ( n8134 , n8133 , n8123 , n952 );
nor ( n8135 , n8132 , n8134 );
nand ( n8136 , n8094 , n8121 , n8128 , n8135 );
nor ( n8137 , n8072 , n8090 , n8136 );
or ( n8138 , n4756 , n8137 );
nand ( n8139 , n8040 , n7901 );
and ( n8140 , n2143 , n8139 );
nand ( n8141 , n8040 , n7940 );
and ( n8142 , n2132 , n8141 );
nor ( n8143 , n8140 , n8142 );
or ( n8144 , n401 , n8143 );
nand ( n8145 , n8037 , n8138 , n8144 );
nand ( n8146 , n2987 , n8145 );
or ( n8147 , n1464 , n1378 , n7894 );
or ( n8148 , n2250 , n7924 );
not ( n8149 , n7978 );
nand ( n8150 , n1427 , n792 );
not ( n8151 , n8150 );
not ( n8152 , n2250 );
not ( n8153 , n8152 );
not ( n8154 , n7916 );
or ( n8155 , n8153 , n8154 );
not ( n8156 , n7861 );
nand ( n8157 , n8155 , n8156 );
nand ( n8158 , n8151 , n8157 );
nor ( n8159 , n6969 , n7874 );
or ( n8160 , n8159 , n7903 );
nand ( n8161 , n8160 , n1013 );
and ( n8162 , n8148 , n8149 , n8158 , n8161 );
and ( n8163 , n1218 , n792 , n7852 );
and ( n8164 , n2251 , n1135 );
nor ( n8165 , n8164 , n6523 );
nor ( n8166 , n8163 , n8165 );
and ( n8167 , n8162 , n8166 , n7912 );
nor ( n8168 , n8167 , n358 );
and ( n8169 , n1748 , n7951 );
nor ( n8170 , n8169 , n7871 );
not ( n8171 , n7879 );
nand ( n8172 , n8171 , n1553 );
not ( n8173 , n7889 );
nand ( n8174 , n8173 , n3731 );
not ( n8175 , n8174 );
not ( n8176 , n7850 );
not ( n8177 , n8176 );
or ( n8178 , n8175 , n8177 );
not ( n8179 , n8033 );
nand ( n8180 , n8178 , n8179 );
and ( n8181 , n8170 , n8172 , n8180 );
nor ( n8182 , n8181 , n6969 );
nor ( n8183 , n1746 , n7955 );
nor ( n8184 , n3732 , n7885 );
nor ( n8185 , n8183 , n8184 , n7949 );
not ( n8186 , n3389 );
not ( n8187 , n8150 );
and ( n8188 , n8186 , n8187 );
nor ( n8189 , n8188 , n7806 );
or ( n8190 , n8189 , n8007 );
and ( n8191 , n1218 , n6034 );
nor ( n8192 , n8191 , n358 );
or ( n8193 , n6523 , n8192 );
nand ( n8194 , n8190 , n8193 , n7997 );
not ( n8195 , n7845 );
not ( n8196 , n8150 );
nor ( n8197 , n8196 , n8000 );
nor ( n8198 , n8195 , n8197 );
nor ( n8199 , n8194 , n1464 , n8198 );
nand ( n8200 , n8185 , n7986 , n8199 );
nor ( n8201 , n8168 , n8182 , n8200 );
nand ( n8202 , n3731 , n7710 );
or ( n8203 , n7707 , n8202 );
not ( n8204 , n7695 );
nor ( n8205 , n3732 , n7697 );
nand ( n8206 , n8204 , n8205 );
nand ( n8207 , n8203 , n8150 , n8206 );
not ( n8208 , n8205 );
nand ( n8209 , n3730 , n7675 );
not ( n8210 , n2696 );
nand ( n8211 , n8210 , n7653 );
nand ( n8212 , n8209 , n8211 );
not ( n8213 , n8212 );
nand ( n8214 , n8208 , n7821 , n8213 , n8202 );
and ( n8215 , n8207 , n8214 );
not ( n8216 , n7684 );
and ( n8217 , n3730 , n8216 );
not ( n8218 , n7766 );
and ( n8219 , n7759 , n7769 );
not ( n8220 , n8219 );
or ( n8221 , n8218 , n8220 );
or ( n8222 , n8189 , n7809 );
nand ( n8223 , n8221 , n8222 );
or ( n8224 , n8219 , n7826 );
nand ( n8225 , n8224 , n1695 );
and ( n8226 , n8225 , n7838 );
nor ( n8227 , n8226 , n6969 );
nor ( n8228 , n8217 , n8223 , n8227 );
nor ( n8229 , n372 , n396 );
nand ( n8230 , n7758 , n8228 , n8229 , n7800 );
not ( n8231 , n7672 );
nor ( n8232 , n8215 , n8230 , n8231 );
or ( n8233 , n8201 , n8232 );
nand ( n8234 , n8147 , n8233 );
nand ( n8235 , n8234 , n4756 , n3004 );
or ( n8236 , n3562 , n7846 );
not ( n8237 , n7866 );
and ( n8238 , n2615 , n8237 );
and ( n8239 , n2606 , n7844 );
nor ( n8240 , n8238 , n8239 );
nand ( n8241 , n8236 , n8240 );
and ( n8242 , n358 , n8241 );
and ( n8243 , n3165 , n7916 );
nor ( n8244 , n8242 , n8243 );
and ( n8245 , n2888 , n7951 );
or ( n8246 , n2630 , n8007 );
and ( n8247 , n2814 , n7852 );
nor ( n8248 , n6523 , n2613 );
nor ( n8249 , n8247 , n8248 );
nand ( n8250 , n8246 , n8249 );
nor ( n8251 , n8245 , n8250 , n1464 );
nand ( n8252 , n8174 , n7849 , n7862 );
nand ( n8253 , n2550 , n8252 );
nand ( n8254 , n7870 , n7875 , n8172 , n8253 );
nand ( n8255 , n329 , n8254 );
and ( n8256 , n8244 , n8251 , n8255 );
not ( n8257 , n7821 );
not ( n8258 , n8219 );
nand ( n8259 , n8258 , n7825 );
nor ( n8260 , n8257 , n8259 , n8205 , n8212 );
or ( n8261 , n2551 , n8260 );
nand ( n8262 , n8261 , n7838 );
and ( n8263 , n329 , n8262 );
not ( n8264 , n8248 );
or ( n8265 , n2630 , n7810 );
not ( n8266 , n7822 );
not ( n8267 , n8202 );
or ( n8268 , n8266 , n8267 );
nand ( n8269 , n8268 , n2613 );
nand ( n8270 , n8264 , n8265 , n1464 , n8269 );
nor ( n8271 , n8263 , n8270 );
nor ( n8272 , n8256 , n8271 );
or ( n8273 , n4757 , n8272 );
not ( n8274 , n7929 );
and ( n8275 , n329 , n8274 );
and ( n8276 , n396 , n2596 );
and ( n8277 , n8276 , n8110 );
not ( n8278 , n6523 );
nand ( n8279 , n396 , n2603 );
not ( n8280 , n8279 );
nor ( n8281 , n8280 , n2604 );
nand ( n8282 , n24 , n8281 );
or ( n8283 , n8282 , n5295 );
nand ( n8284 , n2596 , n1138 );
nand ( n8285 , n8283 , n8284 );
and ( n8286 , n8070 , n8285 );
nor ( n8287 , n329 , n1565 );
nand ( n8288 , n24 , n8287 );
not ( n8289 , n8288 );
and ( n8290 , n8289 , n8022 );
nor ( n8291 , n8286 , n8290 );
not ( n8292 , n8291 );
and ( n8293 , n8278 , n8292 );
nor ( n8294 , n2786 , n2868 );
and ( n8295 , n8294 , n7895 );
nor ( n8296 , n8293 , n8295 );
and ( n8297 , n6523 , n2613 );
and ( n8298 , n1244 , n8297 );
nand ( n8299 , n24 , n8298 , n5971 );
not ( n8300 , n2768 );
or ( n8301 , n8300 , n8126 );
nand ( n8302 , n2849 , n8297 );
not ( n8303 , n8276 );
nand ( n8304 , n8303 , n2849 );
not ( n8305 , n8304 );
nand ( n8306 , n8305 , n6308 );
and ( n8307 , n8302 , n8306 );
nand ( n8308 , n8301 , n8307 );
and ( n8309 , n7852 , n8308 );
not ( n8310 , n2603 );
nand ( n8311 , n6523 , n8310 );
and ( n8312 , n8311 , n6320 );
and ( n8313 , n8312 , n8003 );
not ( n8314 , n7856 );
nor ( n8315 , n8313 , n8314 );
and ( n8316 , n8281 , n8315 );
and ( n8317 , n2874 , n8095 );
nor ( n8318 , n8316 , n8317 );
or ( n8319 , n24 , n8318 );
or ( n8320 , n6523 , n8304 );
or ( n8321 , n8320 , n5286 );
nor ( n8322 , n8280 , n8312 );
not ( n8323 , n8322 );
nor ( n8324 , n2604 , n8323 );
nand ( n8325 , n24 , n8324 );
or ( n8326 , n8325 , n7848 );
nand ( n8327 , n8319 , n8321 , n8326 );
not ( n8328 , n8063 );
or ( n8329 , n2596 , n8083 );
and ( n8330 , n8328 , n8329 );
not ( n8331 , n64 );
nor ( n8332 , n8330 , n8331 );
not ( n8333 , n64 );
and ( n8334 , n8333 , n8063 );
nor ( n8335 , n1264 , n8329 );
nor ( n8336 , n8334 , n8335 );
not ( n8337 , n8336 );
or ( n8338 , n8332 , n8337 );
nand ( n8339 , n8338 , n24 );
not ( n8340 , n8339 );
nor ( n8341 , n8309 , n8327 , n8340 );
and ( n8342 , n8296 , n8299 , n8341 );
nor ( n8343 , n8342 , n358 );
nor ( n8344 , n8275 , n8277 , n8343 );
not ( n8345 , n358 );
nor ( n8346 , n8276 , n2868 , n6320 );
not ( n8347 , n8346 );
not ( n8348 , n8297 );
nand ( n8349 , n8347 , n8348 );
not ( n8350 , n7860 );
nand ( n8351 , n8345 , n8349 , n8350 );
not ( n8352 , n2764 );
nor ( n8353 , n8352 , n7773 );
not ( n8354 , n8353 );
not ( n8355 , n8139 );
or ( n8356 , n8354 , n8355 );
and ( n8357 , n8297 , n3730 , n5993 );
not ( n8358 , n8329 );
and ( n8359 , n1244 , n8358 );
nor ( n8360 , n8359 , n8063 );
or ( n8361 , n1764 , n8360 );
not ( n8362 , n7773 );
not ( n8363 , n7813 );
or ( n8364 , n8362 , n8363 );
nor ( n8365 , n2603 , n8083 );
nand ( n8366 , n8364 , n8365 );
nand ( n8367 , n8361 , n8366 );
nor ( n8368 , n8357 , n8367 );
nand ( n8369 , n8356 , n8368 );
and ( n8370 , n8312 , n7901 );
not ( n8371 , n7773 );
nand ( n8372 , n8279 , n8371 );
nor ( n8373 , n8370 , n8372 , n7874 );
nor ( n8374 , n8369 , n1464 , n8373 );
nand ( n8375 , n8344 , n8351 , n8374 );
not ( n8376 , n8375 );
not ( n8377 , n8209 );
not ( n8378 , n8074 );
or ( n8379 , n2598 , n8378 );
nand ( n8380 , n8379 , n8348 );
and ( n8381 , n8377 , n8380 );
not ( n8382 , n2598 );
not ( n8383 , n8130 );
and ( n8384 , n8382 , n8383 );
not ( n8385 , n8349 );
nor ( n8386 , n8385 , n7737 );
nor ( n8387 , n8384 , n8386 );
or ( n8388 , n2939 , n8387 );
nand ( n8389 , n8388 , n1464 );
and ( n8390 , n8322 , n7721 );
or ( n8391 , n329 , n8040 );
nand ( n8392 , n8391 , n7725 );
and ( n8393 , n281 , n8392 );
nor ( n8394 , n8390 , n8393 );
or ( n8395 , n7813 , n8394 );
and ( n8396 , n8353 , n8085 );
and ( n8397 , n8312 , n7656 );
nor ( n8398 , n8397 , n8372 );
nor ( n8399 , n8396 , n8398 );
or ( n8400 , n7654 , n8399 );
not ( n8401 , n8367 );
nand ( n8402 , n8395 , n8400 , n8401 );
nor ( n8403 , n8381 , n8389 , n8402 );
not ( n8404 , n2596 );
not ( n8405 , n7689 );
and ( n8406 , n8404 , n8405 );
not ( n8407 , n6043 );
not ( n8408 , n8299 );
and ( n8409 , n8407 , n8408 );
or ( n8410 , n8288 , n8052 );
not ( n8411 , n2768 );
not ( n8412 , n8093 );
or ( n8413 , n8411 , n8412 );
nand ( n8414 , n8413 , n8339 );
or ( n8415 , n8282 , n7662 );
or ( n8416 , n8320 , n5531 );
not ( n8417 , n7799 );
or ( n8418 , n8307 , n8417 );
nand ( n8419 , n8415 , n8416 , n8418 );
nor ( n8420 , n8414 , n8419 );
nand ( n8421 , n8410 , n8420 );
nor ( n8422 , n8409 , n8421 );
and ( n8423 , n8294 , n7712 );
or ( n8424 , n8284 , n8115 );
nand ( n8425 , n8424 , n8325 );
and ( n8426 , n7668 , n8425 );
nor ( n8427 , n8423 , n8426 );
and ( n8428 , n8422 , n8427 );
nor ( n8429 , n8428 , n358 );
nor ( n8430 , n8406 , n8429 );
nand ( n8431 , n8403 , n8430 );
not ( n8432 , n8431 );
or ( n8433 , n8376 , n8432 );
nand ( n8434 , n329 , n1244 );
or ( n8435 , n8434 , n7699 );
not ( n8436 , n8118 );
and ( n8437 , n8287 , n8436 );
and ( n8438 , n8298 , n6067 );
nor ( n8439 , n8437 , n8438 );
not ( n8440 , n8042 );
and ( n8441 , n2874 , n8440 );
and ( n8442 , n2605 , n7795 );
not ( n8443 , n8324 );
or ( n8444 , n8443 , n7746 );
nand ( n8445 , n8444 , n8336 );
nor ( n8446 , n8441 , n8442 , n8445 );
nand ( n8447 , n8435 , n8439 , n8446 );
and ( n8448 , n2109 , n8447 );
and ( n8449 , n2605 , n5939 );
nor ( n8450 , n8449 , n2874 );
or ( n8451 , n8068 , n8450 );
nand ( n8452 , n8451 , n8443 );
and ( n8453 , n7869 , n8452 );
nor ( n8454 , n8453 , n8337 );
and ( n8455 , n8287 , n8077 );
and ( n8456 , n8298 , n5952 );
nor ( n8457 , n8455 , n8456 );
nand ( n8458 , n8454 , n8457 );
nor ( n8459 , n8434 , n7886 );
nor ( n8460 , n8458 , n8459 );
or ( n8461 , n1766 , n8460 );
and ( n8462 , n2764 , n8087 );
nor ( n8463 , n2603 , n5066 );
nor ( n8464 , n8462 , n8322 , n8463 );
or ( n8465 , n7715 , n8464 );
not ( n8466 , n8365 );
nand ( n8467 , n8465 , n8466 );
and ( n8468 , n5805 , n8467 );
nor ( n8469 , n8298 , n8346 );
not ( n8470 , n8469 );
not ( n8471 , n7751 );
and ( n8472 , n8470 , n8471 );
and ( n8473 , n8287 , n8061 );
nor ( n8474 , n8472 , n8473 );
not ( n8475 , n8434 );
not ( n8476 , n7753 );
and ( n8477 , n8475 , n8476 );
and ( n8478 , n2874 , n8054 );
nor ( n8479 , n8477 , n8478 );
and ( n8480 , n8324 , n7730 );
not ( n8481 , n7733 );
and ( n8482 , n2605 , n8481 );
nor ( n8483 , n8480 , n8482 );
and ( n8484 , n8474 , n8479 , n8483 );
nor ( n8485 , n8484 , n24 );
nor ( n8486 , n6308 , n5796 );
and ( n8487 , n4949 , n8486 );
nor ( n8488 , n8487 , n8320 );
nor ( n8489 , n8468 , n8485 , n8488 );
or ( n8490 , n1760 , n8489 );
nand ( n8491 , n8297 , n2129 , n6011 );
not ( n8492 , n8007 );
or ( n8493 , n8486 , n2660 , n8304 );
or ( n8494 , n1766 , n8302 );
nand ( n8495 , n8493 , n8494 );
and ( n8496 , n8492 , n8495 );
and ( n8497 , n1260 , n8332 );
nor ( n8498 , n8496 , n8497 );
not ( n8499 , n8360 );
or ( n8500 , n8335 , n8499 );
nand ( n8501 , n8500 , n1359 );
nand ( n8502 , n8491 , n8498 , n4757 , n8501 );
and ( n8503 , n396 , n8030 );
nor ( n8504 , n8503 , n8124 , n8134 );
or ( n8505 , n329 , n8504 );
nand ( n8506 , n2759 , n1769 , n7944 );
nand ( n8507 , n8505 , n8506 );
nor ( n8508 , n8502 , n8507 );
not ( n8509 , n1494 );
nor ( n8510 , n2596 , n8509 );
and ( n8511 , n8510 , n1813 , n7771 );
or ( n8512 , n8352 , n8044 );
or ( n8513 , n8323 , n7866 );
nand ( n8514 , n8512 , n8513 , n8466 );
and ( n8515 , n1769 , n2690 , n8514 );
nor ( n8516 , n8511 , n8515 );
not ( n8517 , n1695 );
not ( n8518 , n8219 );
or ( n8519 , n8517 , n8518 );
nand ( n8520 , n8519 , n8265 );
nand ( n8521 , n8520 , n329 , n8229 );
and ( n8522 , n8276 , n8027 );
and ( n8523 , n2874 , n8099 );
nor ( n8524 , n8522 , n8523 );
and ( n8525 , n8287 , n8141 );
or ( n8526 , n8311 , n6196 );
nand ( n8527 , n8526 , n8098 );
and ( n8528 , n8281 , n8527 );
nor ( n8529 , n8525 , n8528 );
nand ( n8530 , n8524 , n8529 );
or ( n8531 , n8469 , n7846 );
or ( n8532 , n8434 , n7940 );
nand ( n8533 , n8510 , n7956 );
nand ( n8534 , n8531 , n8532 , n8533 );
or ( n8535 , n8530 , n8534 );
nand ( n8536 , n8535 , n1768 );
and ( n8537 , n8508 , n8516 , n8521 , n8536 );
nand ( n8538 , n8461 , n8490 , n8537 );
nor ( n8539 , n8448 , n8538 );
nand ( n8540 , n8433 , n8539 );
nand ( n8541 , n8273 , n8540 , n2995 );
nand ( n8542 , n8018 , n8146 , n8235 , n8541 );
not ( n8543 , n385 );
and ( n8544 , n405 , n8543 );
not ( n8545 , n400 );
and ( n8546 , n388 , n8545 );
and ( n8547 , n5268 , n5006 );
and ( n8548 , n387 , n8546 , n8547 );
nor ( n8549 , n8548 , n766 );
or ( n8550 , n385 , n8549 );
nand ( n8551 , n385 , n390 );
nand ( n8552 , n8550 , n8551 );
nand ( n8553 , n397 , n8552 );
not ( n8554 , n4755 );
not ( n8555 , n1677 );
or ( n8556 , n8554 , n8555 );
not ( n8557 , n401 );
and ( n8558 , n8557 , n1661 );
and ( n8559 , n8558 , n1671 );
nand ( n8560 , n403 , n406 );
and ( n8561 , n8560 , n2984 );
nor ( n8562 , n8559 , n8561 );
nand ( n8563 , n8556 , n8562 );
not ( n8564 , n8563 );
not ( n8565 , n401 );
and ( n8566 , n403 , n1423 );
nor ( n8567 , n8565 , n8566 );
nor ( n8568 , n406 , n8567 );
not ( n8569 , n8568 );
not ( n8570 , n1656 );
or ( n8571 , n8569 , n8570 );
nand ( n8572 , n8571 , n1843 );
nand ( n8573 , n1634 , n1649 );
and ( n8574 , n8564 , n8572 , n8573 );
nor ( n8575 , n8574 , n7570 );
not ( n8576 , n8575 );
not ( n8577 , n1705 );
and ( n8578 , n344 , n8577 );
not ( n8579 , n1707 );
nor ( n8580 , n8578 , n8579 );
or ( n8581 , n1633 , n8580 );
or ( n8582 , n390 , n1686 );
nand ( n8583 , n8582 , n4798 );
nand ( n8584 , n2534 , n4709 );
nand ( n8585 , n8581 , n8583 , n8584 );
and ( n8586 , n1041 , n8585 );
nand ( n8587 , n8561 , n1327 );
not ( n8588 , n8587 );
nor ( n8589 , n8586 , n8588 );
nor ( n8590 , n1424 , n401 );
not ( n8591 , n8590 );
nor ( n8592 , n8591 , n4747 );
or ( n8593 , n2570 , n8592 );
or ( n8594 , n8579 , n1408 );
nand ( n8595 , n8593 , n8594 );
nor ( n8596 , n1633 , n2553 );
not ( n8597 , n8596 );
not ( n8598 , n8597 );
not ( n8599 , n8564 );
or ( n8600 , n8598 , n8599 );
nand ( n8601 , n8600 , n1042 );
and ( n8602 , n8589 , n8595 , n8601 );
not ( n8603 , n4619 );
nor ( n8604 , n8602 , n8603 );
not ( n8605 , n2578 );
not ( n8606 , n8585 );
not ( n8607 , n8606 );
and ( n8608 , n8605 , n8607 );
not ( n8609 , n2510 );
not ( n8610 , n8561 );
nand ( n8611 , n8609 , n406 , n8610 );
not ( n8612 , n2535 );
nand ( n8613 , n8612 , n1677 );
not ( n8614 , n1019 );
not ( n8615 , n2985 );
not ( n8616 , n8568 );
or ( n8617 , n8615 , n8616 );
nand ( n8618 , n1707 , n8587 );
nand ( n8619 , n8617 , n8618 );
not ( n8620 , n8619 );
or ( n8621 , n8614 , n8620 );
not ( n8622 , n8562 );
nand ( n8623 , n8621 , n8622 );
nand ( n8624 , n8611 , n8613 , n8623 );
and ( n8625 , n2576 , n8624 );
nor ( n8626 , n8608 , n8625 );
nor ( n8627 , n1626 , n2448 );
or ( n8628 , n8588 , n8627 );
and ( n8629 , n389 , n2495 );
nand ( n8630 , n8628 , n8629 );
not ( n8631 , n2510 );
nand ( n8632 , n8631 , n2576 , n8567 );
not ( n8633 , n2577 );
not ( n8634 , n8573 );
and ( n8635 , n8633 , n8634 );
and ( n8636 , n2444 , n8629 );
and ( n8637 , n8636 , n8563 );
nor ( n8638 , n8635 , n8637 );
nand ( n8639 , n8632 , n8638 );
and ( n8640 , n8636 , n8596 );
not ( n8641 , n8592 );
nor ( n8642 , n8641 , n2448 );
and ( n8643 , n8629 , n8642 );
nor ( n8644 , n8640 , n8643 );
not ( n8645 , n8644 );
and ( n8646 , n8639 , n8645 );
not ( n8647 , n8639 );
and ( n8648 , n8647 , n8644 );
nor ( n8649 , n8646 , n8648 );
and ( n8650 , n8626 , n8630 , n8649 );
nor ( n8651 , n8650 , n391 );
nor ( n8652 , n8604 , n8651 );
not ( n8653 , n8619 );
or ( n8654 , n8653 , n8585 );
and ( n8655 , n1734 , n7568 );
or ( n8656 , n8655 , n4860 );
nand ( n8657 , n8654 , n8656 );
nand ( n8658 , n8576 , n8652 , n8657 );
or ( n8659 , n385 , n8658 );
not ( n8660 , n7570 );
not ( n8661 , n8618 );
not ( n8662 , n8661 );
or ( n8663 , n8660 , n8662 );
not ( n8664 , n1843 );
not ( n8665 , n7570 );
and ( n8666 , n8664 , n8610 , n8665 );
nor ( n8667 , n8666 , n8543 );
nand ( n8668 , n8663 , n8667 );
not ( n8669 , n8668 );
nor ( n8670 , n8669 , n397 );
nand ( n8671 , n8659 , n8670 );
and ( n8672 , n8553 , n8671 );
nor ( n8673 , n8672 , n405 );
nor ( n8674 , n8544 , n8673 );
not ( n8675 , n400 );
not ( n8676 , n405 );
or ( n8677 , n8675 , n8676 );
and ( n8678 , n8545 , n8658 );
nand ( n8679 , n385 , n387 );
not ( n8680 , n3763 );
nand ( n8681 , n1418 , n8680 );
not ( n8682 , n1736 );
nand ( n8683 , n8682 , n401 );
not ( n8684 , n1042 );
not ( n8685 , n2971 );
and ( n8686 , n8684 , n8685 );
nor ( n8687 , n373 , n2499 );
nor ( n8688 , n8686 , n8687 );
or ( n8689 , n8683 , n8688 );
nand ( n8690 , n8689 , n2585 );
and ( n8691 , n8681 , n8690 );
not ( n8692 , n4722 );
not ( n8693 , n2565 );
or ( n8694 , n8692 , n8693 );
not ( n8695 , n1734 );
not ( n8696 , n2972 );
and ( n8697 , n8695 , n8696 );
nor ( n8698 , n8697 , n4619 );
or ( n8699 , n1626 , n8698 );
nand ( n8700 , n8694 , n8699 );
and ( n8701 , n1327 , n8700 );
nor ( n8702 , n8691 , n8701 );
and ( n8703 , n1041 , n2499 );
and ( n8704 , n1019 , n2971 );
nor ( n8705 , n8703 , n8704 );
not ( n8706 , n4709 );
or ( n8707 , n4803 , n1736 , n8706 );
or ( n8708 , n344 , n8683 , n1365 );
nand ( n8709 , n8707 , n8708 );
and ( n8710 , n8705 , n8709 );
nand ( n8711 , n1042 , n716 );
nor ( n8712 , n714 , n8711 );
and ( n8713 , n4805 , n4709 );
nor ( n8714 , n8713 , n1710 );
not ( n8715 , n8714 );
and ( n8716 , n8712 , n8715 );
nor ( n8717 , n8710 , n8716 );
and ( n8718 , n4718 , n2566 , n4709 );
not ( n8719 , n2031 );
not ( n8720 , n8681 );
or ( n8721 , n8719 , n8720 );
not ( n8722 , n1670 );
nand ( n8723 , n44 , n403 );
nand ( n8724 , n2028 , n1666 );
and ( n8725 , n8723 , n8724 );
nor ( n8726 , n8725 , n2024 );
not ( n8727 , n8726 );
or ( n8728 , n8722 , n8727 );
not ( n8729 , n401 );
nand ( n8730 , n8728 , n8729 );
nand ( n8731 , n8721 , n8730 );
and ( n8732 , n8698 , n8731 );
nor ( n8733 , n8718 , n8732 );
or ( n8734 , n1019 , n8603 );
nand ( n8735 , n8734 , n2496 );
or ( n8736 , n2444 , n8730 );
or ( n8737 , n2453 , n8714 );
not ( n8738 , n401 );
and ( n8739 , n344 , n2028 );
nor ( n8740 , n8739 , n2024 );
nor ( n8741 , n8740 , n1365 );
nand ( n8742 , n8738 , n8741 );
nand ( n8743 , n8736 , n8737 , n8742 );
and ( n8744 , n8735 , n8743 );
or ( n8745 , n2444 , n8741 );
nand ( n8746 , n8745 , n4619 );
and ( n8747 , n4796 , n8746 );
and ( n8748 , n373 , n8715 );
or ( n8749 , n373 , n8730 );
nand ( n8750 , n8749 , n8742 );
nor ( n8751 , n8748 , n8750 );
nor ( n8752 , n8747 , n8751 );
nor ( n8753 , n8744 , n8752 );
nand ( n8754 , n8702 , n8717 , n8733 , n8753 );
and ( n8755 , n8679 , n8754 );
and ( n8756 , n400 , n8668 );
nor ( n8757 , n8756 , n8679 );
nor ( n8758 , n8755 , n8757 );
nor ( n8759 , n8678 , n8758 );
or ( n8760 , n397 , n8759 );
and ( n8761 , n397 , n766 );
nor ( n8762 , n8761 , n8679 );
or ( n8763 , n400 , n8679 );
not ( n8764 , n2980 );
nand ( n8765 , n8763 , n397 , n8764 );
not ( n8766 , n8765 );
and ( n8767 , n8762 , n8766 );
nor ( n8768 , n8543 , n1638 , n8547 );
nand ( n8769 , n400 , n8768 );
not ( n8770 , n8769 );
nand ( n8771 , n8770 , n397 );
nand ( n8772 , n2976 , n8771 );
nor ( n8773 , n400 , n8762 );
nor ( n8774 , n8767 , n8772 , n8773 );
nand ( n8775 , n8760 , n8774 );
nand ( n8776 , n8677 , n8775 );
not ( n8777 , n8658 );
or ( n8778 , n397 , n8777 );
nand ( n8779 , n8778 , n2976 );
and ( n8780 , n2978 , n8779 );
nand ( n8781 , n8543 , n8754 );
and ( n8782 , n8781 , n387 , n8670 );
nand ( n8783 , n387 , n8551 );
not ( n8784 , n397 );
or ( n8785 , n388 , n400 );
and ( n8786 , n390 , n2978 );
nand ( n8787 , n8785 , n8786 );
not ( n8788 , n8787 );
or ( n8789 , n8784 , n8788 );
nand ( n8790 , n8789 , n385 );
and ( n8791 , n8783 , n8790 );
nor ( n8792 , n8782 , n8791 );
nand ( n8793 , n397 , n2536 , n8547 );
not ( n8794 , n8793 );
nand ( n8795 , n8794 , n2979 );
and ( n8796 , n8792 , n8771 , n8795 );
nor ( n8797 , n8796 , n405 );
nor ( n8798 , n8780 , n8797 );
nand ( n8799 , n7568 , n2435 );
nor ( n8800 , n2977 , n8799 );
nand ( n8801 , n2980 , n8800 );
not ( n8802 , n4740 );
or ( n8803 , n1019 , n8802 );
and ( n8804 , n8566 , n8590 );
nand ( n8805 , n8803 , n8804 );
not ( n8806 , n4741 );
and ( n8807 , n8805 , n414 , n8806 );
or ( n8808 , n2509 , n4740 );
and ( n8809 , n1019 , n3242 );
and ( n8810 , n44 , n373 );
nor ( n8811 , n8809 , n8810 , n6320 );
or ( n8812 , n414 , n8811 );
and ( n8813 , n8811 , n4710 );
not ( n8814 , n8804 );
nor ( n8815 , n8813 , n8814 );
nand ( n8816 , n8812 , n8815 );
nand ( n8817 , n8808 , n8816 );
nor ( n8818 , n8807 , n8817 );
or ( n8819 , n8801 , n8818 );
nand ( n8820 , n8810 , n1707 );
nor ( n8821 , n8814 , n8801 );
nand ( n8822 , n392 , n8821 );
or ( n8823 , n8820 , n8822 );
not ( n8824 , n8799 );
nand ( n8825 , n394 , n8802 );
nor ( n8826 , n8825 , n8814 );
or ( n8827 , n8824 , n8826 );
and ( n8828 , n2986 , n2980 );
nand ( n8829 , n8827 , n8828 );
and ( n8830 , n414 , n8829 );
nand ( n8831 , n44 , n8828 );
nand ( n8832 , n8799 , n8826 );
nor ( n8833 , n8831 , n8832 );
nor ( n8834 , n8830 , n8833 );
nand ( n8835 , n8819 , n8823 , n8834 );
nor ( n8836 , n401 , n2977 );
not ( n8837 , n8836 );
nor ( n8838 , n8837 , n8726 );
nor ( n8839 , n1323 , n8765 );
and ( n8840 , n385 , n8546 );
and ( n8841 , n394 , n2978 , n8768 );
nor ( n8842 , n8841 , n8545 );
nor ( n8843 , n8840 , n8842 , n8553 );
and ( n8844 , n8839 , n8843 );
nand ( n8845 , n8566 , n1830 );
and ( n8846 , n401 , n8845 );
not ( n8847 , n8560 );
nor ( n8848 , n8846 , n397 , n8847 );
nor ( n8849 , n8844 , n8848 );
nor ( n8850 , n405 , n8838 , n8849 );
nor ( n8851 , n397 , n8712 , n2579 );
not ( n8852 , n1842 );
or ( n8853 , n8783 , n8852 , n8793 );
nand ( n8854 , n1323 , n8786 );
or ( n8855 , n388 , n8543 , n8854 );
nand ( n8856 , n8853 , n8855 );
and ( n8857 , n8545 , n8856 );
or ( n8858 , n8854 , n8769 );
nand ( n8859 , n8858 , n397 );
nor ( n8860 , n8857 , n8859 );
nor ( n8861 , n405 , n8851 , n8860 );
or ( n8862 , n413 , n4741 , n8826 );
or ( n8863 , n359 , n8806 );
nand ( n8864 , n8862 , n8863 );
nand ( n8865 , n1644 , n8826 );
not ( n8866 , n8801 );
nand ( n8867 , n8865 , n8866 );
or ( n8868 , n8864 , n8867 );
and ( n8869 , n1040 , n4740 , n8821 );
not ( n8870 , n8828 );
nor ( n8871 , n8869 , n8870 );
or ( n8872 , n892 , n8871 );
buf ( n8873 , n8800 );
buf ( n8874 , n8873 );
not ( n8875 , n8874 );
not ( n8876 , n8875 );
not ( n8877 , n1842 );
nor ( n8878 , n1644 , n8814 );
not ( n8879 , n8878 );
nor ( n8880 , n8877 , n8879 );
and ( n8881 , n3243 , n8828 , n8880 );
and ( n8882 , n413 , n8865 );
nor ( n8883 , n8881 , n8882 );
or ( n8884 , n8876 , n8883 );
nand ( n8885 , n8868 , n8872 , n8884 );
not ( n8886 , n6283 );
not ( n8887 , n5003 );
not ( n8888 , n727 );
nor ( n8889 , n8887 , n8888 );
and ( n8890 , n871 , n1025 , n8889 );
nor ( n8891 , n8890 , n2977 );
not ( n8892 , n8891 );
or ( n8893 , n8886 , n8892 );
nand ( n8894 , n8893 , n766 );
not ( n8895 , n402 );
nand ( n8896 , n1707 , n792 );
or ( n8897 , n8896 , n8814 );
and ( n8898 , n8799 , n8897 );
nand ( n8899 , n8828 , n8822 );
nor ( n8900 , n8898 , n8899 );
or ( n8901 , n8895 , n8900 );
nand ( n8902 , n5035 , n2514 );
and ( n8903 , n402 , n8814 , n8902 );
not ( n8904 , n8820 );
and ( n8905 , n791 , n8904 );
and ( n8906 , n402 , n6320 );
nor ( n8907 , n8905 , n8906 );
or ( n8908 , n8814 , n8907 );
or ( n8909 , n3261 , n2515 );
nand ( n8910 , n8908 , n8909 );
nor ( n8911 , n8903 , n8910 );
or ( n8912 , n8801 , n8911 );
or ( n8913 , n1019 , n8799 );
not ( n8914 , n8897 );
nand ( n8915 , n8913 , n8914 );
or ( n8916 , n8831 , n8915 );
nand ( n8917 , n8901 , n8912 , n8916 );
not ( n8918 , n311 );
or ( n8919 , n8918 , n913 );
not ( n8920 , n311 );
and ( n8921 , n8920 , n981 );
not ( n8922 , n64 );
nor ( n8923 , n8922 , n399 );
nor ( n8924 , n8921 , n8923 );
nand ( n8925 , n8919 , n8924 );
nor ( n8926 , n402 , n24 , n8925 );
not ( n8927 , n3130 );
not ( n8928 , n8925 );
and ( n8929 , n8927 , n8928 );
and ( n8930 , n791 , n2536 );
nor ( n8931 , n8929 , n8930 );
and ( n8932 , n8931 , n372 , n407 );
not ( n8933 , n399 );
and ( n8934 , n8933 , n8924 );
not ( n8935 , n402 );
nor ( n8936 , n8935 , n372 );
and ( n8937 , n730 , n8936 );
nand ( n8938 , n407 , n3261 );
nor ( n8939 , n8934 , n8937 , n8938 );
nor ( n8940 , n8932 , n8939 );
or ( n8941 , n8926 , n8940 );
and ( n8942 , n8923 , n3544 );
nor ( n8943 , n8942 , n8938 );
and ( n8944 , n8943 , n1464 , n8925 );
nor ( n8945 , n390 , n3261 );
nor ( n8946 , n8944 , n8945 );
nand ( n8947 , n8941 , n8946 );
not ( n8948 , n399 );
and ( n8949 , n8948 , n8902 , n8897 );
nor ( n8950 , n359 , n8902 );
nor ( n8951 , n8949 , n8950 );
nand ( n8952 , n359 , n8878 );
not ( n8953 , n8897 );
nand ( n8954 , n8953 , n1644 );
and ( n8955 , n8951 , n8952 , n8954 );
not ( n8956 , n399 );
not ( n8957 , n8945 );
and ( n8958 , n8956 , n8957 );
nor ( n8959 , n8958 , n8952 );
nor ( n8960 , n8955 , n8959 );
or ( n8961 , n8801 , n8960 );
not ( n8962 , n399 );
and ( n8963 , n8799 , n8954 );
nor ( n8964 , n8963 , n8870 );
or ( n8965 , n8962 , n8964 );
nand ( n8966 , n792 , n8799 , n8828 , n8880 );
nand ( n8967 , n8961 , n8965 , n8966 );
or ( n8968 , n2028 , n2986 );
nor ( n8969 , n8847 , n4747 );
or ( n8970 , n8723 , n1655 );
nand ( n8971 , n723 , n2984 );
and ( n8972 , n8591 , n8971 );
nor ( n8973 , n1424 , n403 );
nor ( n8974 , n8972 , n8973 );
nor ( n8975 , n8558 , n8974 );
nand ( n8976 , n8970 , n8975 );
and ( n8977 , n8969 , n8838 , n8976 );
and ( n8978 , n8975 , n2028 , n2986 );
nor ( n8979 , n8977 , n8978 );
nand ( n8980 , n8968 , n8979 );
nand ( n8981 , n714 , n1848 );
not ( n8982 , n716 );
or ( n8983 , n8981 , n8982 );
nand ( n8984 , n329 , n2995 );
not ( n8985 , n8984 );
not ( n8986 , n2987 );
nor ( n8987 , n8986 , n2579 );
or ( n8988 , n393 , n8985 , n8987 );
nand ( n8989 , n8988 , n3001 );
nand ( n8990 , n8983 , n8989 );
nor ( n8991 , n1425 , n2977 );
not ( n8992 , n8991 );
nor ( n8993 , n8992 , n8845 );
not ( n8994 , n401 );
not ( n8995 , n8847 );
nor ( n8996 , n8995 , n2977 );
and ( n8997 , n398 , n8996 );
nor ( n8998 , n8993 , n8994 , n8997 );
and ( n8999 , n8991 , n8998 );
nor ( n9000 , n8999 , n8836 , n8973 );
or ( n9001 , n8976 , n9000 );
or ( n9002 , n1424 , n2986 );
nand ( n9003 , n9001 , n9002 );
and ( n9004 , n311 , n409 );
not ( n9005 , n311 );
and ( n9006 , n9005 , n757 );
nor ( n9007 , n9004 , n9006 );
not ( n9008 , n64 );
and ( n9009 , n9008 , n892 );
and ( n9010 , n413 , n1027 );
nor ( n9011 , n9009 , n9010 );
or ( n9012 , n9007 , n9011 );
or ( n9013 , n409 , n2070 );
nand ( n9014 , n9012 , n9013 );
and ( n9015 , n956 , n9014 );
not ( n9016 , n7961 );
nor ( n9017 , n9015 , n9016 );
or ( n9018 , n415 , n9017 );
nand ( n9019 , n9018 , n416 , n3242 );
nand ( n9020 , n4740 , n9019 );
not ( n9021 , n8987 );
or ( n9022 , n7569 , n9021 );
or ( n9023 , n1734 , n2986 );
nand ( n9024 , n9022 , n9023 );
and ( n9025 , n311 , n7157 );
or ( n9026 , n7157 , n746 , n311 );
nand ( n9027 , n9026 , n3023 );
nand ( n9028 , n2 , n1027 );
nor ( n9029 , n9025 , n9027 , n9028 );
or ( n9030 , n8936 , n9029 );
nor ( n9031 , n404 , n8938 );
nand ( n9032 , n9030 , n9031 );
not ( n9033 , n759 );
and ( n9034 , n409 , n7157 );
and ( n9035 , n417 , n757 );
nor ( n9036 , n9034 , n9035 );
or ( n9037 , n730 , n388 );
not ( n9038 , n8945 );
nand ( n9039 , n9037 , n9038 );
and ( n9040 , n9033 , n9036 , n9039 );
not ( n9041 , n9036 );
or ( n9042 , n790 , n9041 );
nand ( n9043 , n9042 , n407 );
and ( n9044 , n9043 , n404 , n3261 );
nor ( n9045 , n9040 , n9044 );
nand ( n9046 , n9032 , n9045 );
not ( n9047 , n401 );
not ( n9048 , n9047 );
not ( n9049 , n8997 );
or ( n9050 , n9048 , n9049 );
not ( n9051 , n8998 );
nand ( n9052 , n9050 , n9051 );
nand ( n9053 , n416 , n750 );
nor ( n9054 , n3243 , n9053 );
not ( n9055 , n9054 );
or ( n9056 , n7961 , n9055 );
not ( n9057 , n727 );
or ( n9058 , n388 , n9057 , n5763 );
and ( n9059 , n416 , n9041 );
nor ( n9060 , n9059 , n750 , n3243 );
not ( n9061 , n5762 );
nand ( n9062 , n1707 , n9036 );
and ( n9063 , n9061 , n9062 );
and ( n9064 , n388 , n4930 );
nor ( n9065 , n9063 , n9064 );
or ( n9066 , n9060 , n9065 );
nand ( n9067 , n9058 , n9066 );
and ( n9068 , n9053 , n727 );
not ( n9069 , n9028 );
nor ( n9070 , n9068 , n9069 , n7961 );
not ( n9071 , n5492 );
nor ( n9072 , n9071 , n9028 , n9053 , n9007 );
or ( n9073 , n9070 , n9072 );
or ( n9074 , n3242 , n9065 );
nand ( n9075 , n9073 , n9074 );
nand ( n9076 , n9056 , n9067 , n9075 );
not ( n9077 , n395 );
not ( n9078 , n3001 );
or ( n9079 , n9077 , n9078 );
not ( n9080 , n8981 );
nor ( n9081 , n9080 , n8705 );
or ( n9082 , n8687 , n9081 );
nand ( n9083 , n9082 , n3002 );
nand ( n9084 , n9079 , n9083 );
not ( n9085 , n389 );
not ( n9086 , n7571 );
or ( n9087 , n9085 , n9086 );
and ( n9088 , n4858 , n8711 );
nor ( n9089 , n9088 , n3001 );
or ( n9090 , n714 , n9089 );
nand ( n9091 , n9087 , n9090 );
nand ( n9092 , n359 , n373 );
not ( n9093 , n8873 );
nor ( n9094 , n2444 , n9093 );
and ( n9095 , n9092 , n9094 );
or ( n9096 , n4144 , n3003 );
nand ( n9097 , n9096 , n8984 );
nor ( n9098 , n9092 , n8875 );
and ( n9099 , n8836 , n8726 );
nor ( n9100 , n398 , n8996 );
nor ( n9101 , n9099 , n8997 , n9100 );
not ( n9102 , n411 );
not ( n9103 , n6421 );
not ( n9104 , n9103 );
or ( n9105 , n9102 , n9104 );
not ( n9106 , n311 );
or ( n9107 , n9106 , n9103 );
nand ( n9108 , n9105 , n9107 );
not ( n9109 , n408 );
nand ( n9110 , n862 , n5342 );
not ( n9111 , n9110 );
or ( n9112 , n9109 , n9111 );
not ( n9113 , n311 );
or ( n9114 , n9113 , n9110 );
nand ( n9115 , n9112 , n9114 );
nor ( n9116 , n373 , n8875 );
and ( n9117 , n374 , n8874 );
and ( n9118 , n152 , n8874 );
buf ( n9119 , n8873 );
and ( n9120 , n282 , n9119 );
and ( n9121 , n345 , n8874 );
and ( n9122 , n296 , n8874 );
and ( n9123 , n360 , n9119 );
and ( n9124 , n330 , n9119 );
and ( n9125 , n266 , n9119 );
not ( n9126 , n5341 );
nor ( n9127 , n2975 , n405 );
and ( n9128 , n2978 , n8545 , n385 , n9127 );
and ( n9129 , n9126 , n9128 );
not ( n9130 , n5342 );
and ( n9131 , n862 , n9130 );
nor ( n9132 , n9129 , n9131 );
and ( n9133 , n106 , n9119 );
and ( n9134 , n313 , n8874 );
and ( n9135 , n267 , n9119 );
and ( n9136 , n85 , n9119 );
and ( n9137 , n361 , n9119 );
and ( n9138 , n283 , n8874 );
and ( n9139 , n86 , n9119 );
and ( n9140 , n331 , n8874 );
and ( n9141 , n129 , n9119 );
and ( n9142 , n128 , n9119 );
and ( n9143 , n346 , n9119 );
and ( n9144 , n297 , n8874 );
and ( n9145 , n375 , n9119 );
and ( n9146 , n312 , n9119 );
and ( n9147 , n332 , n9119 );
and ( n9148 , n151 , n9119 );
and ( n9149 , n2986 , n8804 );
not ( n9150 , n9149 );
nor ( n9151 , n1889 , n9150 );
nor ( n9152 , n44 , n9150 );
nor ( n9153 , n1830 , n9150 );
nor ( n9154 , n1642 , n9150 );
and ( n9155 , n164 , n9149 );
and ( n9156 , n199 , n9149 );
and ( n9157 , n33 , n9149 );
and ( n9158 , n181 , n9149 );
and ( n9159 , n52 , n9149 );
and ( n9160 , n95 , n9149 );
and ( n9161 , n190 , n9149 );
and ( n9162 , n162 , n9149 );
and ( n9163 , n141 , n9149 );
and ( n9164 , n32 , n9149 );
and ( n9165 , n206 , n9149 );
and ( n9166 , n74 , n9149 );
and ( n9167 , n139 , n9149 );
and ( n9168 , n116 , n9149 );
not ( n9169 , n409 );
not ( n9170 , n4740 );
or ( n9171 , n9169 , n9170 );
nand ( n9172 , n9171 , n8825 );
and ( n9173 , n118 , n9149 );
and ( n9174 , n94 , n9149 );
and ( n9175 , n140 , n9149 );
not ( n9176 , n5106 );
and ( n9177 , n9176 , n9128 );
not ( n9178 , n410 );
and ( n9179 , n9178 , n6420 );
nor ( n9180 , n9177 , n9179 );
and ( n9181 , n96 , n9149 );
and ( n9182 , n117 , n9149 );
and ( n9183 , n53 , n9149 );
and ( n9184 , n10 , n9149 );
and ( n9185 , n11 , n9149 );
and ( n9186 , n163 , n9149 );
and ( n9187 , n73 , n9149 );
not ( n9188 , n8991 );
nor ( n9189 , n9188 , n8971 );
or ( n9190 , n7157 , n8945 );
nand ( n9191 , n9190 , n8896 );
endmodule

