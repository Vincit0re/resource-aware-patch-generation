module top ( g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 , g98 , g99 , g100 , g101 , g102 , g103 , g104 , g105 , g106 , g107 , g108 , g109 , g110 , g111 , g112 , g113 , g114 , g115 , g116 , g117 , g118 , g119 , g120 , g121 , g122 , g123 , g124 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g136 , g137 , g138 , g139 , g140 , g141 , g142 , g143 , g144 , g145 , g146 , g147 , g148 , g149 , g150 , g151 , g152 , g153 , g154 , g155 , g156 , g157 , g158 , g159 , g160 , g161 , g162 , g163 , g164 , g165 , g166 , g167 , g168 , g169 , g170 , g171 , g172 , g173 , g174 , g175 , g176 , g177 , g178 , g179 , g180 , g181 , g182 , g183 , g184 , g185 , g186 , g187 , g188 , g189 , g190 , g191 , g192 , g193 , g194 , g195 , g196 , g197 , g198 , g199 , g200 , g201 , g202 , g203 , g204 , g205 , g206 , g207 , g208 , g209 , g210 , g211 , g212 , g213 , g214 , g215 , g216 , g217 , g218 , g219 , g220 , g221 , g222 , g223 , g224 , g225 , g226 );
input g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 , g98 ;
output g99 , g100 , g101 , g102 , g103 , g104 , g105 , g106 , g107 , g108 , g109 , g110 , g111 , g112 , g113 , g114 , g115 , g116 , g117 , g118 , g119 , g120 , g121 , g122 , g123 , g124 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g136 , g137 , g138 , g139 , g140 , g141 , g142 , g143 , g144 , g145 , g146 , g147 , g148 , g149 , g150 , g151 , g152 , g153 , g154 , g155 , g156 , g157 , g158 , g159 , g160 , g161 , g162 , g163 , g164 , g165 , g166 , g167 , g168 , g169 , g170 , g171 , g172 , g173 , g174 , g175 , g176 , g177 , g178 , g179 , g180 , g181 , g182 , g183 , g184 , g185 , g186 , g187 , g188 , g189 , g190 , g191 , g192 , g193 , g194 , g195 , g196 , g197 , g198 , g199 , g200 , g201 , g202 , g203 , g204 , g205 , g206 , g207 , g208 , g209 , g210 , g211 , g212 , g213 , g214 , g215 , g216 , g217 , g218 , g219 , g220 , g221 , g222 , g223 , g224 , g225 , g226 ;

wire n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , 
     n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , 
     n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , 
     n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , 
     n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , 
     n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , 
     n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , 
     n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , 
     n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , 
     n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , 
     n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , 
     n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , 
     n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , 
     n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , 
     n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , 
     n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , 
     n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , 
     n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , 
     n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , 
     n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , 
     n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , 
     n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , 
     n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , 
     n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , 
     n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , 
     n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , 
     n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , 
     n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , 
     n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , 
     n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , 
     n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , 
     n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , 
     n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , 
     n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , 
     n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , 
     n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , 
     n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , 
     n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , 
     n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , 
     n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , 
     n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , 
     n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , 
     n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , 
     n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , 
     n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , 
     n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , 
     n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , 
     n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , 
     n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , 
     n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , 
     n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , 
     n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , 
     n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , 
     n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , 
     n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , 
     n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , 
     n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , 
     n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , 
     n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , 
     n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , 
     n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , 
     n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , 
     n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , 
     n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , 
     n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , 
     n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , 
     n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , 
     n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , 
     n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , 
     n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , 
     n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , 
     n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , 
     n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , 
     n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , 
     n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , 
     n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , 
     n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , 
     n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , 
     n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , 
     n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , 
     n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , 
     n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , 
     n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , 
     n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , 
     n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , 
     n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , 
     n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , 
     n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , 
     n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , 
     n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , 
     n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , 
     n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , 
     n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , 
     n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , 
     n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , 
     n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , 
     n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , 
     n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , 
     n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , 
     n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , 
     n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , 
     n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , 
     n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , 
     n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , 
     n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , 
     n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , 
     n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , 
     n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , 
     n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , 
     n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , 
     n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , 
     n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , 
     n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , 
     n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , 
     n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , 
     n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , 
     n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , 
     n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , 
     n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , 
     n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , 
     n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , 
     n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , 
     n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , 
     n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , 
     n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , 
     n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , 
     n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , 
     n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , 
     n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , 
     n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , 
     n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , 
     n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , 
     n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , 
     n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , 
     n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , 
     n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , 
     n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , 
     n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , 
     n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , 
     n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , 
     n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , 
     n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , 
     n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , 
     n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , 
     n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , 
     n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , 
     n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , 
     n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , 
     n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , 
     n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , 
     n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , 
     n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , 
     n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , 
     n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , 
     n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , 
     n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , 
     n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , 
     n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , 
     n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , 
     n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , 
     n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , 
     n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , 
     n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , 
     n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , 
     n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , 
     n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , 
     n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , 
     n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , 
     n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , 
     n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , 
     n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , 
     n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , 
     n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , 
     n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , 
     n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , 
     n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , 
     n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , 
     n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , 
     n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , 
     n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , 
     n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , 
     n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , 
     n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , 
     n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , 
     n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , 
     n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , 
     n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , 
     n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , 
     n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , 
     n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , 
     n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , 
     n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , 
     n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , 
     n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , 
     n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , 
     n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , 
     n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , 
     n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , 
     n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , 
     n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , 
     n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , 
     n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , 
     n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , 
     n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , 
     n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , 
     n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , 
     n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , 
     n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , 
     n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , 
     n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , 
     n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , 
     n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , 
     n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , 
     n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , 
     n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , 
     n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , 
     n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , 
     n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , 
     n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , 
     n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , 
     n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , 
     n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , 
     n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , 
     n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , 
     n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , 
     n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , 
     n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , 
     n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , 
     n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , 
     n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , 
     n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , 
     n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , 
     n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , 
     n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , 
     n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , 
     n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , 
     n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , 
     n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , 
     n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , 
     n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , 
     n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , 
     n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , 
     n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , 
     n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , 
     n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , 
     n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , 
     n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , 
     n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , 
     n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , 
     n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , 
     n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , 
     n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , 
     n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , 
     n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , 
     n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , 
     n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , 
     n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , 
     n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , 
     n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , 
     n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , 
     n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , 
     n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , 
     n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , 
     n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , 
     n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , 
     n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , 
     n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , 
     n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , 
     n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , 
     n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , 
     n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , 
     n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , 
     n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , 
     n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , 
     n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , 
     n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , 
     n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , 
     n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , 
     n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , 
     n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , 
     n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , 
     n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , 
     n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , 
     n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , 
     n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , 
     n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , 
     n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , 
     n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , 
     n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , 
     n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , 
     n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , 
     n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , 
     n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , 
     n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , 
     n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , 
     n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , 
     n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , 
     n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , 
     n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , 
     n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , 
     n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , 
     n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , 
     n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , 
     n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , 
     n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , 
     n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , 
     n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , 
     n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , 
     n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , 
     n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , 
     n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , 
     n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , 
     n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , 
     n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , 
     n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , 
     n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , 
     n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , 
     n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , 
     n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , 
     n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , 
     n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , 
     n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , 
     n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , 
     n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , 
     n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , 
     n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , 
     n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , 
     n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , 
     n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , 
     n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , 
     n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , 
     n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , 
     n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , 
     n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , 
     n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , 
     n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , 
     n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , 
     n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , 
     n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , 
     n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , 
     n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , 
     n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , 
     n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , 
     n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , 
     n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , 
     n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , 
     n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , 
     n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , 
     n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , 
     n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , 
     n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , 
     n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , 
     n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , 
     n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , 
     n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , 
     n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , 
     n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , 
     n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , 
     n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , 
     n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , 
     n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , 
     n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , 
     n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , 
     n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , 
     n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , 
     n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , 
     n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , 
     n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , 
     n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , 
     n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , 
     n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , 
     n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , 
     n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , 
     n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , 
     n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , 
     n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , 
     n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , 
     n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , 
     n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , 
     n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , 
     n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , 
     n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , 
     n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , 
     n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , 
     n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , 
     n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , 
     n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , 
     n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , 
     n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , 
     n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , 
     n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , 
     n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , 
     n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , 
     n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , 
     n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , 
     n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , 
     n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , 
     n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , 
     n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , 
     n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , 
     n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , 
     n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , 
     n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , 
     n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , 
     n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , 
     n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , 
     n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , 
     n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , 
     n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , 
     n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , 
     n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , 
     n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , 
     n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , 
     n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , 
     n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , 
     n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , 
     n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , 
     n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , 
     n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , 
     n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , 
     n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , 
     n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , 
     n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , 
     n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , 
     n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , 
     n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , 
     n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , 
     n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , 
     n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , 
     n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , 
     n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , 
     n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , 
     n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , 
     n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , 
     n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , 
     n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , 
     n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , 
     n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , 
     n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , 
     n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , 
     n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , 
     n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , 
     n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , 
     n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , 
     n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , 
     n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , 
     n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , 
     n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , 
     n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , 
     n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , 
     n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , 
     n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , 
     n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , 
     n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , 
     n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , 
     n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , 
     n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , 
     n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , 
     n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , 
     n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , 
     n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , 
     n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , 
     n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , 
     n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , 
     n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , 
     n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , 
     n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , 
     n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , 
     n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , 
     n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , 
     n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , 
     n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , 
     n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , 
     n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , 
     n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , 
     n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , 
     n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , 
     n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , 
     n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , 
     n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , 
     n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , 
     n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , 
     n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , 
     n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , 
     n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , 
     n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , 
     n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , 
     n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , 
     n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , 
     n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , 
     n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , 
     n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , 
     n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , 
     n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , 
     n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , 
     n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , 
     n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , 
     n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , 
     n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , 
     n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , 
     n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , 
     n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , 
     n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , 
     n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , 
     n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , 
     n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , 
     n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , 
     n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , 
     n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , 
     n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , 
     n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , 
     n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , 
     n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , 
     n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , 
     n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , 
     n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , 
     n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , 
     n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , 
     n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , 
     n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , 
     n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , 
     n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , 
     n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , 
     n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , 
     n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , 
     n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , 
     n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , 
     n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , 
     n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , 
     n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , 
     n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , 
     n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , 
     n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , 
     n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , 
     n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , 
     n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , 
     n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , 
     n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , 
     n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , 
     n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , 
     n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , 
     n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , 
     n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , 
     n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , 
     n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , 
     n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , 
     n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , 
     n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , 
     n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , 
     n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , 
     n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , 
     n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , 
     n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , 
     n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , 
     n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , 
     n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , 
     n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , 
     n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , 
     n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , 
     n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , 
     n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , 
     n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , 
     n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , 
     n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , 
     n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , 
     n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , 
     n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , 
     n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , 
     n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , 
     n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , 
     n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , 
     n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , 
     n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , 
     n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , 
     n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , 
     n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , 
     n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , 
     n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , 
     n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , 
     n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , 
     n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , 
     n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , 
     n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , 
     n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , 
     n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , 
     n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , 
     n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , 
     n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , 
     n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , 
     n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , 
     n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , 
     n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , 
     n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , 
     n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , 
     n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , 
     n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , 
     n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , 
     n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , 
     n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , 
     n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , 
     n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , 
     n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , 
     n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , 
     n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , 
     n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , 
     n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , 
     n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , 
     n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , 
     n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , 
     n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , 
     n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , 
     n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , 
     n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , 
     n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , 
     n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , 
     n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , 
     n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , 
     n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , 
     n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , 
     n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , 
     n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , 
     n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , 
     n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , 
     n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , 
     n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , 
     n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , 
     n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , 
     n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , 
     n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , 
     n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , 
     n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , 
     n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , 
     n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , 
     n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , 
     n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , 
     n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , 
     n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , 
     n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , 
     n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , 
     n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , 
     n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , 
     n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , 
     n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , 
     n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , 
     n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , 
     n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , 
     n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , 
     n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , 
     n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , 
     n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , 
     n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , 
     n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , 
     n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , 
     n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , 
     n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , 
     n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , 
     n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , 
     n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , 
     n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , 
     n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , 
     n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , 
     n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , 
     n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , 
     n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , 
     n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , 
     n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , 
     n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , 
     n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , 
     n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , 
     n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , 
     n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , 
     n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , 
     n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , 
     n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , 
     n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , 
     n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , 
     n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , 
     n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , 
     n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , 
     n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , 
     n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , 
     n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , 
     n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , 
     n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , 
     n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , 
     n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , 
     n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , 
     n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , 
     n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , 
     n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , 
     n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , 
     n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , 
     n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , 
     n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , 
     n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , 
     n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , 
     n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , 
     n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , 
     n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , 
     n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , 
     n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , 
     n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , 
     n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , 
     n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , 
     n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , 
     n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , 
     n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , 
     n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , 
     n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , 
     n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , 
     n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , 
     n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , 
     n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , 
     n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , 
     n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , 
     n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , 
     n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , 
     n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , 
     n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , 
     n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , 
     n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , 
     n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , 
     n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , 
     n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , 
     n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , 
     n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , 
     n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , 
     n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , 
     n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , 
     n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , 
     n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , 
     n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , 
     n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , 
     n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , 
     n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , 
     n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , 
     n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , 
     n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , 
     n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , 
     n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , 
     n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , 
     n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , 
     n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , 
     n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , 
     n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , 
     n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , 
     n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , 
     n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , 
     n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , 
     n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , 
     n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , 
     n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , 
     n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , 
     n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , 
     n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , 
     n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , 
     n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , 
     n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , 
     n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , 
     n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , 
     n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , 
     n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , 
     n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , 
     n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , 
     n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , 
     n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , 
     n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , 
     n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , 
     n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , 
     n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , 
     n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , 
     n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , 
     n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , 
     n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , 
     n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , 
     n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , 
     n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , 
     n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , 
     n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , 
     n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , 
     n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , 
     n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , 
     n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , 
     n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , 
     n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , 
     n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , 
     n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , 
     n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , 
     n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , 
     n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , 
     n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , 
     n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , 
     n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , 
     n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , 
     n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , 
     n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , 
     n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , 
     n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , 
     n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , 
     n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , 
     n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , 
     n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , 
     n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , 
     n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , 
     n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , 
     n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , 
     n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , 
     n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , 
     n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , 
     n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , 
     n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , 
     n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , 
     n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , 
     n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , 
     n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , 
     n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , 
     n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , 
     n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , 
     n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , 
     n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , 
     n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , 
     n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , 
     n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , 
     n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , 
     n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , 
     n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , 
     n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , 
     n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , 
     n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , 
     n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , 
     n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , 
     n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , 
     n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , 
     n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , 
     n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , 
     n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , 
     n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , 
     n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , 
     n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , 
     n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , 
     n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , 
     n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , 
     n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , 
     n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , 
     n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , 
     n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , 
     n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , 
     n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , 
     n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , 
     n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , 
     n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , 
     n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , 
     n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , 
     n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , 
     n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , 
     n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , 
     n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , 
     n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , 
     n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , 
     n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , 
     n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , 
     n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , 
     n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , 
     n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , 
     n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , 
     n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , 
     n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , 
     n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , 
     n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , 
     n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , 
     n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , 
     n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , 
     n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , 
     n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , 
     n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , 
     n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , 
     n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , 
     n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , 
     n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , 
     n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , 
     n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , 
     n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , 
     n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , 
     n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , 
     n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , 
     n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , 
     n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , 
     n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , 
     n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , 
     n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , 
     n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , 
     n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , 
     n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , 
     n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , 
     n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , 
     n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , 
     n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , 
     n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , 
     n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , 
     n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , 
     n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , 
     n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , 
     n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , 
     n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , 
     n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , 
     n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , 
     n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , 
     n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , 
     n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , 
     n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , 
     n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , 
     n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , 
     n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , 
     n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , 
     n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , 
     n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , 
     n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , 
     n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , 
     n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , 
     n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , 
     n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , 
     n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , 
     n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , 
     n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , 
     n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , 
     n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , 
     n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , 
     n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , 
     n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , 
     n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , 
     n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , 
     n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , 
     n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , 
     n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , 
     n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , 
     n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , 
     n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , 
     n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , 
     n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , 
     n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , 
     n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , 
     n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , 
     n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , 
     n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , 
     n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , 
     n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , 
     n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , 
     n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , 
     n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , 
     n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , 
     n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , 
     n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , 
     n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , 
     n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , 
     n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , 
     n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , 
     n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , 
     n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , 
     n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , 
     n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , 
     n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , 
     n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , 
     n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , 
     n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , 
     n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , 
     n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , 
     n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , 
     n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , 
     n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , 
     n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , 
     n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , 
     n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , 
     n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , 
     n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , 
     n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , 
     n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , 
     n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , 
     n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , 
     n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , 
     n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , 
     n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , 
     n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , 
     n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , 
     n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , 
     n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , 
     n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , 
     n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , 
     n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , 
     n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , 
     n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , 
     n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , 
     n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , 
     n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , 
     n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , 
     n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , 
     n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , 
     n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , 
     n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , 
     n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , 
     n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , 
     n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , 
     n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , 
     n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , 
     n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , 
     n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , 
     n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , 
     n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , 
     n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , 
     n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , 
     n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , 
     n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , 
     n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , 
     n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , 
     n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , 
     n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , 
     n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , 
     n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , 
     n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , 
     n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , 
     n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , 
     n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , 
     n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , 
     n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , 
     n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , 
     n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , 
     n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , 
     n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , 
     n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , 
     n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , 
     n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , 
     n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , 
     n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , 
     n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , 
     n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , 
     n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , 
     n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , 
     n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , 
     n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , 
     n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , 
     n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , 
     n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , 
     n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , 
     n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , 
     n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , 
     n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , 
     n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , 
     n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , 
     n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , 
     n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , 
     n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , 
     n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , 
     n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , 
     n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , 
     n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , 
     n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , 
     n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , 
     n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , 
     n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , 
     n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , 
     n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , 
     n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , 
     n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , 
     n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , 
     n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , 
     n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , 
     n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , 
     n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , 
     n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , 
     n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , 
     n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , 
     n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , 
     n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , 
     n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , 
     n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , 
     n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , 
     n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , 
     n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , 
     n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , 
     n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , 
     n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , 
     n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , 
     n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , 
     n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , 
     n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , 
     n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , 
     n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , 
     n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , 
     n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , 
     n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , 
     n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , 
     n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , 
     n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , 
     n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , 
     n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , 
     n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , 
     n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , 
     n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , 
     n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , 
     n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , 
     n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , 
     n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , 
     n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , 
     n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , 
     n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , 
     n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , 
     n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , 
     n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , 
     n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , 
     n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , 
     n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , 
     n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , 
     n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , 
     n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , 
     n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , 
     n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , 
     n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , 
     n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , 
     n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , 
     n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , 
     n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , 
     n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , 
     n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , 
     n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , 
     n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , 
     n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , 
     n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , 
     n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , 
     n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , 
     n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , 
     n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , 
     n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , 
     n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , 
     n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , 
     n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , 
     n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , 
     n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , 
     n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , 
     n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , 
     n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , 
     n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , 
     n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , 
     n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , 
     n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , 
     n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , 
     n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , 
     n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , 
     n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , 
     n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , 
     n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , 
     n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , 
     n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , 
     n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , 
     n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , 
     n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , 
     n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , 
     n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , 
     n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , 
     n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , 
     n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , 
     n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , 
     n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , 
     n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , 
     n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , 
     n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , 
     n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , 
     n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , 
     n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , 
     n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , 
     n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , 
     n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , 
     n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , 
     n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , 
     n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , 
     n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , 
     n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , 
     n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , 
     n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , 
     n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , 
     n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , 
     n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , 
     n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , 
     n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , 
     n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , 
     n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , 
     n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , 
     n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , 
     n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , 
     n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , 
     n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , 
     n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , 
     n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , 
     n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , 
     n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , 
     n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , 
     n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , 
     n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , 
     n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , 
     n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , 
     n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , 
     n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , 
     n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , 
     n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , 
     n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , 
     n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , 
     n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , 
     n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , 
     n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , 
     n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , 
     n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , 
     n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , 
     n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , 
     n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , 
     n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , 
     n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , 
     n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , 
     n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , 
     n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , 
     n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , 
     n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , 
     n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , 
     n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , 
     n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , 
     n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , 
     n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , 
     n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , 
     n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , 
     n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , 
     n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , 
     n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , 
     n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , 
     n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , 
     n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , 
     n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , 
     n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , 
     n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , 
     n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , 
     n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , 
     n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , 
     n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , 
     n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , 
     n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , 
     n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , 
     n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , 
     n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , 
     n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , 
     n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , 
     n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , 
     n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , 
     n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , 
     n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , 
     n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , 
     n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , 
     n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , 
     n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , 
     n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , 
     n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , 
     n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , 
     n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , 
     n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , 
     n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , 
     n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , 
     n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , 
     n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , 
     n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , 
     n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , 
     n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , 
     n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , 
     n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , 
     n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , 
     n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , 
     n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , 
     n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , 
     n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , 
     n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , 
     n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , 
     n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , 
     n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , 
     n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , 
     n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , 
     n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , 
     n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , 
     n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , 
     n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , 
     n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , 
     n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , 
     n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , 
     n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , 
     n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , 
     n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , 
     n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , 
     n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , 
     n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , 
     n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , 
     n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , 
     n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , 
     n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , 
     n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , 
     n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , 
     n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , 
     n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , 
     n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , 
     n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , 
     n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , 
     n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , 
     n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , 
     n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , 
     n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , 
     n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , 
     n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , 
     n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , 
     n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , 
     n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , 
     n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , 
     n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , 
     n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , 
     n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , 
     n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , 
     n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , 
     n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , 
     n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , 
     n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , 
     n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , 
     n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , 
     n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , 
     n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , 
     n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , 
     n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , 
     n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , 
     n13280 , n13281 , n13282 , n13283 ;
wire t_0 , t_1 , t_2 , t_3 ;
buf ( n1 , g0 );
buf ( n2 , g1 );
buf ( n3 , g2 );
buf ( n4 , g3 );
buf ( n5 , g4 );
buf ( n6 , g5 );
buf ( n7 , g6 );
buf ( n8 , g7 );
buf ( n9 , g8 );
buf ( n10 , g9 );
buf ( n11 , g10 );
buf ( n12 , g11 );
buf ( n13 , g12 );
buf ( n14 , g13 );
buf ( n15 , g14 );
buf ( n16 , g15 );
buf ( n17 , g16 );
buf ( n18 , g17 );
buf ( n19 , g18 );
buf ( n20 , g19 );
buf ( n21 , g20 );
buf ( n22 , g21 );
buf ( n23 , g22 );
buf ( n24 , g23 );
buf ( n25 , g24 );
buf ( n26 , g25 );
buf ( n27 , g26 );
buf ( n28 , g27 );
buf ( n29 , g28 );
buf ( n30 , g29 );
buf ( n31 , g30 );
buf ( n32 , g31 );
buf ( n33 , g32 );
buf ( n34 , g33 );
buf ( n35 , g34 );
buf ( n36 , g35 );
buf ( n37 , g36 );
buf ( n38 , g37 );
buf ( n39 , g38 );
buf ( n40 , g39 );
buf ( n41 , g40 );
buf ( n42 , g41 );
buf ( n43 , g42 );
buf ( n44 , g43 );
buf ( n45 , g44 );
buf ( n46 , g45 );
buf ( n47 , g46 );
buf ( n48 , g47 );
buf ( n49 , g48 );
buf ( n50 , g49 );
buf ( n51 , g50 );
buf ( n52 , g51 );
buf ( n53 , g52 );
buf ( n54 , g53 );
buf ( n55 , g54 );
buf ( n56 , g55 );
buf ( n57 , g56 );
buf ( n58 , g57 );
buf ( n59 , g58 );
buf ( n60 , g59 );
buf ( n61 , g60 );
buf ( n62 , g61 );
buf ( n63 , g62 );
buf ( n64 , g63 );
buf ( n65 , g64 );
buf ( n66 , g65 );
buf ( n67 , g66 );
buf ( n68 , g67 );
buf ( n69 , g68 );
buf ( n70 , g69 );
buf ( n71 , g70 );
buf ( n72 , g71 );
buf ( n73 , g72 );
buf ( n74 , g73 );
buf ( n75 , g74 );
buf ( n76 , g75 );
buf ( n77 , g76 );
buf ( n78 , g77 );
buf ( n79 , g78 );
buf ( n80 , g79 );
buf ( n81 , g80 );
buf ( n82 , g81 );
buf ( n83 , g82 );
buf ( n84 , g83 );
buf ( n85 , g84 );
buf ( n86 , g85 );
buf ( n87 , g86 );
buf ( n88 , g87 );
buf ( n89 , g88 );
buf ( n90 , g89 );
buf ( n91 , g90 );
buf ( n92 , g91 );
buf ( n93 , g92 );
buf ( n94 , g93 );
buf ( n95 , g94 );
buf ( n96 , g95 );
buf ( n97 , g96 );
buf ( n98 , g97 );
buf ( n99 , g98 );
buf ( g99 , n100 );
buf ( g100 , n101 );
buf ( g101 , n102 );
buf ( g102 , n103 );
buf ( g103 , n104 );
buf ( g104 , n105 );
buf ( g105 , n106 );
buf ( g106 , n107 );
buf ( g107 , n108 );
buf ( g108 , n109 );
buf ( g109 , n110 );
buf ( g110 , n111 );
buf ( g111 , n112 );
buf ( g112 , n113 );
buf ( g113 , n114 );
buf ( g114 , n115 );
buf ( g115 , n116 );
buf ( g116 , n117 );
buf ( g117 , n118 );
buf ( g118 , n119 );
buf ( g119 , n120 );
buf ( g120 , n121 );
buf ( g121 , n122 );
buf ( g122 , n123 );
buf ( g123 , n124 );
buf ( g124 , n125 );
buf ( g125 , n126 );
buf ( g126 , n127 );
buf ( g127 , n128 );
buf ( g128 , n129 );
buf ( g129 , n130 );
buf ( g130 , n131 );
buf ( g131 , n132 );
buf ( g132 , n133 );
buf ( g133 , n134 );
buf ( g134 , n135 );
buf ( g135 , n136 );
buf ( g136 , n137 );
buf ( g137 , n138 );
buf ( g138 , n139 );
buf ( g139 , n140 );
buf ( g140 , n141 );
buf ( g141 , n142 );
buf ( g142 , n143 );
buf ( g143 , n144 );
buf ( g144 , n145 );
buf ( g145 , n146 );
buf ( g146 , n147 );
buf ( g147 , n148 );
buf ( g148 , n149 );
buf ( g149 , n150 );
buf ( g150 , n151 );
buf ( g151 , n152 );
buf ( g152 , n153 );
buf ( g153 , n154 );
buf ( g154 , n155 );
buf ( g155 , n156 );
buf ( g156 , n157 );
buf ( g157 , n158 );
buf ( g158 , n159 );
buf ( g159 , n160 );
buf ( g160 , n161 );
buf ( g161 , n162 );
buf ( g162 , n163 );
buf ( g163 , n164 );
buf ( g164 , n165 );
buf ( g165 , n166 );
buf ( g166 , n167 );
buf ( g167 , n168 );
buf ( g168 , n169 );
buf ( g169 , n170 );
buf ( g170 , n171 );
buf ( g171 , n172 );
buf ( g172 , n173 );
buf ( g173 , n174 );
buf ( g174 , n175 );
buf ( g175 , n176 );
buf ( g176 , n177 );
buf ( g177 , n178 );
buf ( g178 , n179 );
buf ( g179 , n180 );
buf ( g180 , n181 );
buf ( g181 , n182 );
buf ( g182 , n183 );
buf ( g183 , n184 );
buf ( g184 , n185 );
buf ( g185 , n186 );
buf ( g186 , n187 );
buf ( g187 , n188 );
buf ( g188 , n189 );
buf ( g189 , n190 );
buf ( g190 , n191 );
buf ( g191 , n192 );
buf ( g192 , n193 );
buf ( g193 , n194 );
buf ( g194 , n195 );
buf ( g195 , n196 );
buf ( g196 , n197 );
buf ( g197 , n198 );
buf ( g198 , n199 );
buf ( g199 , n200 );
buf ( g200 , n201 );
buf ( g201 , n202 );
buf ( g202 , n203 );
buf ( g203 , n204 );
buf ( g204 , n205 );
buf ( g205 , n206 );
buf ( g206 , n207 );
buf ( g207 , n208 );
buf ( g208 , n209 );
buf ( g209 , n210 );
buf ( g210 , n211 );
buf ( g211 , n212 );
buf ( g212 , n213 );
buf ( g213 , n214 );
buf ( g214 , n215 );
buf ( g215 , n216 );
buf ( g216 , n217 );
buf ( g217 , n218 );
buf ( g218 , n219 );
buf ( g219 , n220 );
buf ( g220 , n221 );
buf ( g221 , n222 );
buf ( g222 , n223 );
buf ( g223 , n224 );
buf ( g224 , n225 );
buf ( g225 , n226 );
buf ( g226 , n227 );
buf ( n100 , 1'b0 );
buf ( n101 , 1'b0 );
buf ( n102 , 1'b0 );
buf ( n103 , 1'b0 );
buf ( n104 , 1'b0 );
buf ( n105 , 1'b0 );
buf ( n106 , 1'b0 );
buf ( n107 , 1'b0 );
buf ( n108 , 1'b0 );
buf ( n109 , 1'b0 );
buf ( n110 , 1'b0 );
buf ( n111 , 1'b0 );
buf ( n112 , 1'b0 );
buf ( n113 , 1'b0 );
buf ( n114 , 1'b0 );
buf ( n115 , 1'b0 );
buf ( n116 , 1'b0 );
buf ( n117 , 1'b0 );
buf ( n118 , 1'b0 );
buf ( n119 , 1'b0 );
buf ( n120 , 1'b0 );
buf ( n121 , 1'b0 );
buf ( n122 , 1'b0 );
buf ( n123 , 1'b0 );
buf ( n124 , 1'b0 );
buf ( n125 , 1'b0 );
buf ( n126 , 1'b0 );
buf ( n127 , 1'b0 );
buf ( n128 , 1'b0 );
buf ( n129 , 1'b0 );
buf ( n130 , 1'b0 );
buf ( n131 , n10553 );
buf ( n132 , n10084 );
buf ( n133 , n12778 );
buf ( n134 , n10129 );
buf ( n135 , n12852 );
buf ( n136 , n13282 );
buf ( n137 , n12908 );
buf ( n138 , n13283 );
buf ( n139 , n12888 );
buf ( n140 , n12891 );
buf ( n141 , n12953 );
buf ( n142 , n12955 );
buf ( n143 , n13020 );
buf ( n144 , n10233 );
buf ( n145 , n10453 );
buf ( n146 , n10254 );
buf ( n147 , n10262 );
buf ( n148 , n10402 );
buf ( n149 , n13008 );
buf ( n150 , n10421 );
buf ( n151 , n10276 );
buf ( n152 , n10293 );
buf ( n153 , n10367 );
buf ( n154 , n10377 );
buf ( n155 , n10357 );
buf ( n156 , n10352 );
buf ( n157 , n10331 );
buf ( n158 , n10315 );
buf ( n159 , n13249 );
buf ( n160 , n13262 );
buf ( n161 , n13268 );
buf ( n162 , n13275 );
buf ( n163 , n13281 );
buf ( n164 , 1'b0 );
buf ( n165 , 1'b0 );
buf ( n166 , 1'b0 );
buf ( n167 , 1'b0 );
buf ( n168 , 1'b0 );
buf ( n169 , 1'b0 );
buf ( n170 , 1'b0 );
buf ( n171 , 1'b0 );
buf ( n172 , 1'b0 );
buf ( n173 , 1'b0 );
buf ( n174 , 1'b0 );
buf ( n175 , 1'b0 );
buf ( n176 , 1'b0 );
buf ( n177 , 1'b0 );
buf ( n178 , 1'b0 );
buf ( n179 , 1'b0 );
buf ( n180 , 1'b0 );
buf ( n181 , 1'b0 );
buf ( n182 , 1'b0 );
buf ( n183 , 1'b0 );
buf ( n184 , 1'b0 );
buf ( n185 , 1'b0 );
buf ( n186 , 1'b0 );
buf ( n187 , 1'b0 );
buf ( n188 , 1'b0 );
buf ( n189 , 1'b0 );
buf ( n190 , 1'b0 );
buf ( n191 , 1'b0 );
buf ( n192 , 1'b0 );
buf ( n193 , 1'b0 );
buf ( n194 , 1'b0 );
buf ( n195 , 1'b0 );
buf ( n196 , 1'b0 );
buf ( n197 , 1'b0 );
buf ( n198 , n13119 );
buf ( n199 , n12829 );
buf ( n200 , n12740 );
buf ( n201 , n12768 );
buf ( n202 , n12790 );
buf ( n203 , n12847 );
buf ( n204 , n12876 );
buf ( n205 , n12887 );
buf ( n206 , n12928 );
buf ( n207 , n12940 );
buf ( n208 , n12907 );
buf ( n209 , n12952 );
buf ( n210 , n12967 );
buf ( n211 , n12992 );
buf ( n212 , n13033 );
buf ( n213 , n13019 );
buf ( n214 , n13051 );
buf ( n215 , n13070 );
buf ( n216 , n13080 );
buf ( n217 , n13136 );
buf ( n218 , n13148 );
buf ( n219 , n13156 );
buf ( n220 , n13168 );
buf ( n221 , n13181 );
buf ( n222 , n13192 );
buf ( n223 , n13205 );
buf ( n224 , n13216 );
buf ( n225 , n13231 );
buf ( n226 , n13238 );
buf ( n227 , n13243 );
or ( n295 , n68 , n84 );
not ( n296 , n68 );
not ( n297 , n84 );
nor ( n298 , n296 , n297 );
not ( n299 , n298 );
nand ( n300 , n295 , n299 );
not ( n301 , n300 );
xor ( n302 , n85 , n86 );
not ( n303 , n302 );
xor ( n304 , n84 , n85 );
nand ( n305 , n303 , n304 );
not ( n306 , n305 );
not ( n307 , n306 );
not ( n308 , n307 );
not ( n309 , n308 );
not ( n310 , n309 );
not ( n311 , n310 );
not ( n312 , n311 );
and ( n313 , n301 , n312 );
and ( n314 , n84 , n302 );
nor ( n315 , n313 , n314 );
nand ( n316 , n69 , n84 );
and ( n317 , n315 , n316 );
not ( n318 , n315 );
not ( n319 , n316 );
and ( n320 , n318 , n319 );
nor ( n321 , n317 , n320 );
xor ( n322 , n87 , n88 );
not ( n323 , n322 );
not ( n324 , n323 );
buf ( n325 , n324 );
not ( n326 , n325 );
not ( n327 , n326 );
not ( n328 , n327 );
not ( n329 , n328 );
not ( n330 , n322 );
xor ( n331 , n86 , n87 );
nand ( n332 , n330 , n331 );
not ( n333 , n332 );
buf ( n334 , n333 );
buf ( n335 , n334 );
buf ( n336 , n335 );
buf ( n337 , n336 );
buf ( n338 , n337 );
buf ( n339 , n338 );
buf ( n340 , n339 );
or ( n341 , n329 , n340 );
nand ( n342 , n341 , n86 );
or ( n343 , n69 , n84 );
nand ( n344 , n343 , n316 );
or ( n345 , n344 , n311 );
not ( n346 , n302 );
or ( n347 , n346 , n300 );
nand ( n348 , n345 , n347 );
and ( n349 , n70 , n84 );
xor ( n350 , n348 , n349 );
and ( n351 , n342 , n350 );
and ( n352 , n349 , n348 );
nor ( n353 , n351 , n352 );
or ( n354 , n321 , n353 );
and ( n355 , n321 , n353 );
nor ( n356 , n355 , n1 );
nand ( n357 , n354 , n356 );
not ( n358 , n86 );
and ( n359 , n296 , n358 );
and ( n360 , n68 , n86 );
nor ( n361 , n359 , n360 );
and ( n362 , n361 , n340 );
and ( n363 , n86 , n329 );
nor ( n364 , n362 , n363 );
or ( n365 , n70 , n84 );
not ( n366 , n349 );
nand ( n367 , n365 , n366 );
or ( n368 , n367 , n311 );
or ( n369 , n346 , n344 );
nand ( n370 , n368 , n369 );
and ( n371 , n71 , n84 );
xor ( n372 , n370 , n371 );
and ( n373 , n364 , n372 );
and ( n374 , n371 , n370 );
nor ( n375 , n373 , n374 );
nor ( n376 , n364 , n375 );
xnor ( n377 , n342 , n350 );
xnor ( n378 , n375 , n364 );
nor ( n379 , n377 , n378 );
or ( n380 , n376 , n379 );
not ( n381 , n1 );
nand ( n382 , n380 , n381 );
nor ( n383 , n357 , n382 );
not ( n384 , n383 );
and ( n385 , n357 , n382 );
not ( n386 , n385 );
and ( n387 , n377 , n378 );
nor ( n388 , n387 , n1 , n379 );
not ( n389 , n69 );
and ( n390 , n389 , n358 );
and ( n391 , n69 , n86 );
nor ( n392 , n390 , n391 );
and ( n393 , n392 , n340 );
and ( n394 , n329 , n361 );
nor ( n395 , n393 , n394 );
nand ( n396 , n72 , n84 );
not ( n397 , n89 );
nand ( n398 , n397 , n90 );
not ( n399 , n90 );
nand ( n400 , n89 , n399 );
nand ( n401 , n398 , n400 );
not ( n402 , n401 );
not ( n403 , n402 );
not ( n404 , n403 );
not ( n405 , n404 );
not ( n406 , n405 );
not ( n407 , n88 );
not ( n408 , n89 );
and ( n409 , n407 , n408 );
and ( n410 , n88 , n89 );
nor ( n411 , n409 , n410 );
and ( n412 , n411 , n398 , n400 );
not ( n413 , n412 );
not ( n414 , n413 );
not ( n415 , n414 );
not ( n416 , n415 );
not ( n417 , n416 );
and ( n418 , n406 , n417 );
not ( n419 , n88 );
nor ( n420 , n418 , n419 );
xnor ( n421 , n396 , n420 );
or ( n422 , n395 , n421 );
or ( n423 , n396 , n420 );
nand ( n424 , n422 , n423 );
xor ( n425 , n372 , n364 );
and ( n426 , n424 , n425 );
and ( n427 , n296 , n419 );
and ( n428 , n68 , n88 );
nor ( n429 , n427 , n428 );
and ( n430 , n429 , n416 );
and ( n431 , n88 , n405 );
nor ( n432 , n430 , n431 );
or ( n433 , n71 , n84 );
not ( n434 , n371 );
nand ( n435 , n433 , n434 );
or ( n436 , n435 , n309 );
or ( n437 , n346 , n367 );
nand ( n438 , n436 , n437 );
and ( n439 , n432 , n438 );
not ( n440 , n432 );
not ( n441 , n438 );
and ( n442 , n440 , n441 );
nor ( n443 , n439 , n442 );
not ( n444 , n70 );
and ( n445 , n444 , n358 );
and ( n446 , n70 , n86 );
nor ( n447 , n445 , n446 );
and ( n448 , n447 , n339 );
and ( n449 , n329 , n392 );
nor ( n450 , n448 , n449 );
not ( n451 , n450 );
or ( n452 , n72 , n84 );
nand ( n453 , n452 , n396 );
or ( n454 , n453 , n309 );
or ( n455 , n346 , n435 );
nand ( n456 , n454 , n455 );
nand ( n457 , n73 , n84 );
not ( n458 , n457 );
xnor ( n459 , n456 , n458 );
not ( n460 , n459 );
and ( n461 , n451 , n460 );
and ( n462 , n458 , n456 );
nor ( n463 , n461 , n462 );
or ( n464 , n443 , n463 );
or ( n465 , n432 , n441 );
nand ( n466 , n464 , n465 );
xor ( n467 , n425 , n424 );
and ( n468 , n466 , n467 );
nor ( n469 , n426 , n468 );
nor ( n470 , n1 , n469 );
nor ( n471 , n388 , n470 );
not ( n472 , n471 );
not ( n473 , n472 );
not ( n474 , n1 );
not ( n475 , n2 );
xor ( n476 , n37 , n38 );
buf ( n477 , n476 );
buf ( n478 , n477 );
not ( n479 , n478 );
not ( n480 , n479 );
buf ( n481 , n480 );
not ( n482 , n481 );
not ( n483 , n482 );
not ( n484 , n483 );
nand ( n485 , n36 , n37 );
nor ( n486 , n36 , n37 );
not ( n487 , n486 );
not ( n488 , n476 );
and ( n489 , n485 , n487 , n488 );
buf ( n490 , n489 );
not ( n491 , n490 );
not ( n492 , n491 );
not ( n493 , n492 );
not ( n494 , n493 );
not ( n495 , n494 );
and ( n496 , n484 , n495 );
not ( n497 , n36 );
nor ( n498 , n496 , n497 );
not ( n499 , n498 );
and ( n500 , n3 , n4 );
not ( n501 , n3 );
and ( n502 , n501 , n20 );
nor ( n503 , n500 , n502 );
not ( n504 , n503 );
buf ( n505 , n504 );
buf ( n506 , n505 );
and ( n507 , n36 , n506 );
not ( n508 , n507 );
and ( n509 , n3 , n5 );
not ( n510 , n3 );
and ( n511 , n510 , n21 );
nor ( n512 , n509 , n511 );
not ( n513 , n512 );
not ( n514 , n513 );
not ( n515 , n514 );
not ( n516 , n515 );
not ( n517 , n516 );
not ( n518 , n517 );
buf ( n519 , n518 );
not ( n520 , n519 );
and ( n521 , n36 , n520 );
not ( n522 , n521 );
not ( n523 , n522 );
and ( n524 , n508 , n523 );
not ( n525 , n508 );
and ( n526 , n525 , n522 );
nor ( n527 , n524 , n526 );
not ( n528 , n527 );
and ( n529 , n499 , n528 );
and ( n530 , n498 , n527 );
nor ( n531 , n529 , n530 );
buf ( n532 , n505 );
not ( n533 , n532 );
and ( n534 , n497 , n533 );
nor ( n535 , n534 , n507 );
not ( n536 , n535 );
or ( n537 , n495 , n536 );
nand ( n538 , n36 , n483 );
nand ( n539 , n537 , n538 );
or ( n540 , n523 , n539 );
nand ( n541 , n523 , n539 );
nand ( n542 , n540 , n541 );
not ( n543 , n520 );
and ( n544 , n497 , n543 );
nor ( n545 , n544 , n521 );
and ( n546 , n494 , n545 );
and ( n547 , n483 , n535 );
nor ( n548 , n546 , n547 );
and ( n549 , n3 , n6 );
not ( n550 , n3 );
and ( n551 , n550 , n22 );
nor ( n552 , n549 , n551 );
not ( n553 , n552 );
buf ( n554 , n553 );
not ( n555 , n554 );
buf ( n556 , n555 );
not ( n557 , n556 );
nand ( n558 , n36 , n557 );
xor ( n559 , n39 , n40 );
buf ( n560 , n559 );
not ( n561 , n560 );
not ( n562 , n561 );
buf ( n563 , n562 );
not ( n564 , n563 );
not ( n565 , n38 );
not ( n566 , n39 );
or ( n567 , n565 , n566 );
xor ( n568 , n39 , n40 );
nor ( n569 , n38 , n39 );
nor ( n570 , n568 , n569 );
nand ( n571 , n567 , n570 );
not ( n572 , n571 );
buf ( n573 , n572 );
not ( n574 , n573 );
not ( n575 , n574 );
not ( n576 , n575 );
nand ( n577 , n564 , n576 );
and ( n578 , n38 , n577 );
xnor ( n579 , n558 , n578 );
or ( n580 , n548 , n579 );
or ( n581 , n558 , n578 );
nand ( n582 , n580 , n581 );
and ( n583 , n542 , n582 );
and ( n584 , n522 , n539 );
nor ( n585 , n583 , n584 );
xor ( n586 , n531 , n585 );
not ( n587 , n586 );
xor ( n588 , n582 , n542 );
not ( n589 , n588 );
and ( n590 , n497 , n557 );
not ( n591 , n556 );
not ( n592 , n591 );
and ( n593 , n36 , n592 );
nor ( n594 , n590 , n593 );
not ( n595 , n594 );
and ( n596 , n494 , n595 );
and ( n597 , n483 , n545 );
nor ( n598 , n596 , n597 );
and ( n599 , n3 , n7 );
not ( n600 , n3 );
and ( n601 , n600 , n23 );
nor ( n602 , n599 , n601 );
not ( n603 , n602 );
not ( n604 , n603 );
not ( n605 , n604 );
nand ( n606 , n36 , n605 );
not ( n607 , n574 );
not ( n608 , n607 );
not ( n609 , n38 );
buf ( n610 , n506 );
and ( n611 , n609 , n610 );
and ( n612 , n38 , n533 );
nor ( n613 , n611 , n612 );
or ( n614 , n608 , n613 );
not ( n615 , n563 );
or ( n616 , n615 , n609 );
nand ( n617 , n614 , n616 );
not ( n618 , n617 );
and ( n619 , n606 , n618 );
not ( n620 , n606 );
and ( n621 , n620 , n617 );
nor ( n622 , n619 , n621 );
or ( n623 , n598 , n622 );
or ( n624 , n606 , n617 );
nand ( n625 , n623 , n624 );
xor ( n626 , n548 , n579 );
and ( n627 , n626 , n617 );
not ( n628 , n626 );
and ( n629 , n628 , n618 );
nor ( n630 , n627 , n629 );
and ( n631 , n625 , n630 );
and ( n632 , n617 , n626 );
nor ( n633 , n631 , n632 );
nand ( n634 , n589 , n633 );
not ( n635 , n634 );
xor ( n636 , n41 , n42 );
buf ( n637 , n636 );
buf ( n638 , n637 );
buf ( n639 , n638 );
not ( n640 , n639 );
and ( n641 , n3 , n10 );
not ( n642 , n3 );
and ( n643 , n642 , n26 );
nor ( n644 , n641 , n643 );
buf ( n645 , n644 );
not ( n646 , n645 );
not ( n647 , n40 );
nand ( n648 , n646 , n647 );
nand ( n649 , n3 , n10 );
not ( n650 , n3 );
nand ( n651 , n650 , n26 );
nand ( n652 , n40 , n649 , n651 );
and ( n653 , n648 , n652 );
or ( n654 , n640 , n653 );
and ( n655 , n3 , n11 );
not ( n656 , n3 );
and ( n657 , n656 , n27 );
nor ( n658 , n655 , n657 );
not ( n659 , n658 );
not ( n660 , n659 );
not ( n661 , n660 );
not ( n662 , n661 );
not ( n663 , n40 );
and ( n664 , n662 , n663 );
not ( n665 , n660 );
and ( n666 , n665 , n40 );
nor ( n667 , n664 , n666 );
nand ( n668 , n40 , n41 );
not ( n669 , n41 );
nand ( n670 , n42 , n669 );
nor ( n671 , n40 , n42 );
not ( n672 , n671 );
nand ( n673 , n668 , n670 , n672 );
not ( n674 , n673 );
nand ( n675 , n667 , n674 );
nand ( n676 , n654 , n675 );
buf ( n677 , n44 );
not ( n678 , n677 );
not ( n679 , n45 );
or ( n680 , n678 , n679 );
buf ( n681 , n44 );
nor ( n682 , n681 , n45 );
xor ( n683 , n45 , n46 );
nor ( n684 , n682 , n683 );
nand ( n685 , n680 , n684 );
not ( n686 , n685 );
not ( n687 , n686 );
buf ( n688 , n44 );
not ( n689 , n688 );
not ( n690 , n689 );
and ( n691 , n3 , n7 );
not ( n692 , n3 );
and ( n693 , n692 , n23 );
nor ( n694 , n691 , n693 );
not ( n695 , n694 );
not ( n696 , n695 );
or ( n697 , n690 , n696 );
buf ( n698 , n44 );
not ( n699 , n698 );
or ( n700 , n699 , n695 );
nand ( n701 , n697 , n700 );
not ( n702 , n701 );
or ( n703 , n687 , n702 );
buf ( n704 , n683 );
buf ( n705 , n704 );
not ( n706 , n699 );
buf ( n707 , n553 );
not ( n708 , n707 );
or ( n709 , n706 , n708 );
buf ( n710 , n698 );
not ( n711 , n710 );
or ( n712 , n711 , n554 );
nand ( n713 , n709 , n712 );
nand ( n714 , n705 , n713 );
nand ( n715 , n703 , n714 );
not ( n716 , n715 );
and ( n717 , n3 , n16 );
not ( n718 , n3 );
and ( n719 , n718 , n32 );
nor ( n720 , n717 , n719 );
buf ( n721 , n720 );
not ( n722 , n721 );
not ( n723 , n722 );
or ( n724 , n497 , n723 );
nand ( n725 , n716 , n724 );
and ( n726 , n676 , n725 );
not ( n727 , n715 );
nor ( n728 , n727 , n724 );
nor ( n729 , n726 , n728 );
xor ( n730 , n47 , n48 );
xnor ( n731 , n46 , n47 );
nor ( n732 , n730 , n731 );
buf ( n733 , n732 );
buf ( n734 , n733 );
not ( n735 , n734 );
not ( n736 , n46 );
not ( n737 , n503 );
not ( n738 , n737 );
not ( n739 , n738 );
or ( n740 , n736 , n739 );
or ( n741 , n46 , n738 );
nand ( n742 , n740 , n741 );
not ( n743 , n742 );
or ( n744 , n735 , n743 );
buf ( n745 , n730 );
not ( n746 , n745 );
not ( n747 , n746 );
nand ( n748 , n46 , n747 );
nand ( n749 , n744 , n748 );
and ( n750 , n729 , n749 );
not ( n751 , n729 );
not ( n752 , n749 );
and ( n753 , n751 , n752 );
nor ( n754 , n750 , n753 );
buf ( n755 , n730 );
not ( n756 , n755 );
not ( n757 , n756 );
not ( n758 , n757 );
not ( n759 , n742 );
or ( n760 , n758 , n759 );
not ( n761 , n733 );
not ( n762 , n761 );
not ( n763 , n46 );
not ( n764 , n763 );
not ( n765 , n514 );
not ( n766 , n765 );
or ( n767 , n764 , n766 );
or ( n768 , n763 , n515 );
nand ( n769 , n767 , n768 );
nand ( n770 , n762 , n769 );
nand ( n771 , n760 , n770 );
not ( n772 , n771 );
xnor ( n773 , n43 , n44 );
xor ( n774 , n42 , n43 );
nand ( n775 , n773 , n774 );
buf ( n776 , n775 );
not ( n777 , n776 );
not ( n778 , n777 );
and ( n779 , n3 , n9 );
not ( n780 , n3 );
and ( n781 , n780 , n25 );
nor ( n782 , n779 , n781 );
not ( n783 , n782 );
xor ( n784 , n783 , n42 );
not ( n785 , n784 );
or ( n786 , n778 , n785 );
xor ( n787 , n43 , n44 );
buf ( n788 , n787 );
not ( n789 , n788 );
not ( n790 , n789 );
and ( n791 , n3 , n8 );
not ( n792 , n3 );
and ( n793 , n792 , n24 );
nor ( n794 , n791 , n793 );
not ( n795 , n794 );
xor ( n796 , n42 , n795 );
nand ( n797 , n790 , n796 );
nand ( n798 , n786 , n797 );
xor ( n799 , n49 , n50 );
buf ( n800 , n799 );
not ( n801 , n800 );
not ( n802 , n801 );
xor ( n803 , n49 , n50 );
not ( n804 , n803 );
xor ( n805 , n48 , n49 );
nand ( n806 , n804 , n805 );
buf ( n807 , n806 );
not ( n808 , n807 );
or ( n809 , n802 , n808 );
nand ( n810 , n809 , n48 );
xor ( n811 , n798 , n810 );
not ( n812 , n811 );
or ( n813 , n772 , n812 );
buf ( n814 , n798 );
nand ( n815 , n810 , n814 );
nand ( n816 , n813 , n815 );
not ( n817 , n816 );
and ( n818 , n754 , n817 );
not ( n819 , n754 );
and ( n820 , n819 , n816 );
nor ( n821 , n818 , n820 );
xor ( n822 , n810 , n814 );
xor ( n823 , n822 , n771 );
not ( n824 , n823 );
not ( n825 , n733 );
not ( n826 , n46 );
not ( n827 , n554 );
not ( n828 , n827 );
or ( n829 , n826 , n828 );
and ( n830 , n3 , n6 );
not ( n831 , n3 );
and ( n832 , n831 , n22 );
or ( n833 , n830 , n832 );
nand ( n834 , n833 , n763 );
nand ( n835 , n829 , n834 );
not ( n836 , n835 );
or ( n837 , n825 , n836 );
nand ( n838 , n747 , n769 );
nand ( n839 , n837 , n838 );
not ( n840 , n839 );
and ( n841 , n3 , n17 );
not ( n842 , n3 );
and ( n843 , n842 , n33 );
nor ( n844 , n841 , n843 );
buf ( n845 , n844 );
not ( n846 , n845 );
nand ( n847 , n36 , n846 );
not ( n848 , n847 );
not ( n849 , n848 );
and ( n850 , n3 , n10 );
not ( n851 , n3 );
and ( n852 , n851 , n26 );
or ( n853 , n850 , n852 );
xor ( n854 , n853 , n42 );
nand ( n855 , n777 , n854 );
buf ( n856 , n788 );
nand ( n857 , n856 , n784 );
nand ( n858 , n849 , n855 , n857 );
not ( n859 , n858 );
or ( n860 , n840 , n859 );
not ( n861 , n847 );
buf ( n862 , n788 );
not ( n863 , n862 );
not ( n864 , n784 );
or ( n865 , n863 , n864 );
nand ( n866 , n865 , n855 );
nand ( n867 , n861 , n866 );
nand ( n868 , n860 , n867 );
not ( n869 , n868 );
not ( n870 , n673 );
buf ( n871 , n870 );
not ( n872 , n871 );
not ( n873 , n40 );
and ( n874 , n3 , n12 );
not ( n875 , n3 );
and ( n876 , n875 , n28 );
nor ( n877 , n874 , n876 );
buf ( n878 , n877 );
not ( n879 , n878 );
or ( n880 , n873 , n879 );
or ( n881 , n40 , n878 );
nand ( n882 , n880 , n881 );
not ( n883 , n882 );
or ( n884 , n872 , n883 );
not ( n885 , n637 );
buf ( n886 , n885 );
not ( n887 , n886 );
nand ( n888 , n887 , n667 );
nand ( n889 , n884 , n888 );
not ( n890 , n889 );
not ( n891 , n559 );
not ( n892 , n609 );
and ( n893 , n3 , n13 );
not ( n894 , n3 );
and ( n895 , n894 , n29 );
nor ( n896 , n893 , n895 );
not ( n897 , n896 );
not ( n898 , n897 );
or ( n899 , n892 , n898 );
and ( n900 , n3 , n13 );
not ( n901 , n3 );
and ( n902 , n901 , n29 );
nor ( n903 , n900 , n902 );
not ( n904 , n903 );
or ( n905 , n609 , n904 );
nand ( n906 , n899 , n905 );
not ( n907 , n906 );
or ( n908 , n891 , n907 );
not ( n909 , n571 );
not ( n910 , n38 );
not ( n911 , n14 );
and ( n912 , n3 , n911 );
not ( n913 , n3 );
not ( n914 , n30 );
and ( n915 , n913 , n914 );
nor ( n916 , n912 , n915 );
not ( n917 , n916 );
not ( n918 , n917 );
or ( n919 , n910 , n918 );
and ( n920 , n3 , n14 );
not ( n921 , n3 );
and ( n922 , n921 , n30 );
or ( n923 , n920 , n922 );
nand ( n924 , n609 , n923 );
nand ( n925 , n919 , n924 );
nand ( n926 , n909 , n925 );
nand ( n927 , n908 , n926 );
not ( n928 , n704 );
not ( n929 , n701 );
or ( n930 , n928 , n929 );
not ( n931 , n685 );
not ( n932 , n688 );
and ( n933 , n3 , n8 );
not ( n934 , n3 );
and ( n935 , n934 , n24 );
nor ( n936 , n933 , n935 );
not ( n937 , n936 );
or ( n938 , n932 , n937 );
not ( n939 , n698 );
not ( n940 , n936 );
nand ( n941 , n939 , n940 );
nand ( n942 , n938 , n941 );
nand ( n943 , n931 , n942 );
nand ( n944 , n930 , n943 );
and ( n945 , n927 , n944 );
not ( n946 , n927 );
not ( n947 , n944 );
and ( n948 , n946 , n947 );
nor ( n949 , n945 , n948 );
not ( n950 , n949 );
or ( n951 , n890 , n950 );
not ( n952 , n947 );
nand ( n953 , n952 , n927 );
nand ( n954 , n951 , n953 );
not ( n955 , n954 );
and ( n956 , n869 , n955 );
not ( n957 , n869 );
not ( n958 , n955 );
and ( n959 , n957 , n958 );
nor ( n960 , n956 , n959 );
not ( n961 , n960 );
or ( n962 , n824 , n961 );
not ( n963 , n869 );
nand ( n964 , n963 , n958 );
nand ( n965 , n962 , n964 );
xor ( n966 , n821 , n965 );
not ( n967 , n480 );
not ( n968 , n497 );
buf ( n969 , n917 );
not ( n970 , n969 );
not ( n971 , n970 );
or ( n972 , n968 , n971 );
buf ( n973 , n969 );
nand ( n974 , n36 , n973 );
nand ( n975 , n972 , n974 );
not ( n976 , n975 );
or ( n977 , n967 , n976 );
not ( n978 , n36 );
and ( n979 , n3 , n15 );
not ( n980 , n3 );
and ( n981 , n980 , n31 );
nor ( n982 , n979 , n981 );
not ( n983 , n982 );
not ( n984 , n983 );
not ( n985 , n984 );
or ( n986 , n978 , n985 );
buf ( n987 , n982 );
or ( n988 , n36 , n987 );
nand ( n989 , n986 , n988 );
nand ( n990 , n490 , n989 );
nand ( n991 , n977 , n990 );
nand ( n992 , n49 , n50 );
not ( n993 , n992 );
nor ( n994 , n49 , n50 );
not ( n995 , n994 );
not ( n996 , n995 );
or ( n997 , n993 , n996 );
nand ( n998 , n997 , n805 );
not ( n999 , n998 );
not ( n1000 , n999 );
not ( n1001 , n48 );
and ( n1002 , n3 , n4 );
not ( n1003 , n3 );
and ( n1004 , n1003 , n20 );
nor ( n1005 , n1002 , n1004 );
not ( n1006 , n1005 );
or ( n1007 , n1001 , n1006 );
not ( n1008 , n48 );
and ( n1009 , n3 , n4 );
not ( n1010 , n3 );
and ( n1011 , n1010 , n20 );
or ( n1012 , n1009 , n1011 );
nand ( n1013 , n1008 , n1012 );
nand ( n1014 , n1007 , n1013 );
not ( n1015 , n1014 );
or ( n1016 , n1000 , n1015 );
buf ( n1017 , n799 );
buf ( n1018 , n1017 );
nand ( n1019 , n1018 , n48 );
nand ( n1020 , n1016 , n1019 );
buf ( n1021 , n559 );
buf ( n1022 , n1021 );
not ( n1023 , n1022 );
not ( n1024 , n38 );
not ( n1025 , n878 );
or ( n1026 , n1024 , n1025 );
buf ( n1027 , n877 );
not ( n1028 , n1027 );
nand ( n1029 , n609 , n1028 );
nand ( n1030 , n1026 , n1029 );
not ( n1031 , n1030 );
or ( n1032 , n1023 , n1031 );
nand ( n1033 , n573 , n906 );
nand ( n1034 , n1032 , n1033 );
xor ( n1035 , n1020 , n1034 );
and ( n1036 , n991 , n1035 );
and ( n1037 , n1020 , n1034 );
nor ( n1038 , n1036 , n1037 );
not ( n1039 , n987 );
nand ( n1040 , n1039 , n36 );
not ( n1041 , n862 );
not ( n1042 , n42 );
not ( n1043 , n602 );
not ( n1044 , n1043 );
not ( n1045 , n1044 );
or ( n1046 , n1042 , n1045 );
or ( n1047 , n42 , n1044 );
nand ( n1048 , n1046 , n1047 );
not ( n1049 , n1048 );
or ( n1050 , n1041 , n1049 );
not ( n1051 , n776 );
nand ( n1052 , n1051 , n796 );
nand ( n1053 , n1050 , n1052 );
not ( n1054 , n1053 );
xor ( n1055 , n1040 , n1054 );
not ( n1056 , n490 );
not ( n1057 , n975 );
or ( n1058 , n1056 , n1057 );
not ( n1059 , n479 );
not ( n1060 , n36 );
buf ( n1061 , n903 );
not ( n1062 , n1061 );
or ( n1063 , n1060 , n1062 );
or ( n1064 , n36 , n1061 );
nand ( n1065 , n1063 , n1064 );
nand ( n1066 , n1059 , n1065 );
nand ( n1067 , n1058 , n1066 );
xnor ( n1068 , n1055 , n1067 );
xor ( n1069 , n1038 , n1068 );
not ( n1070 , n871 );
not ( n1071 , n653 );
not ( n1072 , n1071 );
or ( n1073 , n1070 , n1072 );
not ( n1074 , n886 );
not ( n1075 , n40 );
and ( n1076 , n3 , n9 );
not ( n1077 , n3 );
and ( n1078 , n1077 , n25 );
nor ( n1079 , n1076 , n1078 );
buf ( n1080 , n1079 );
not ( n1081 , n1080 );
or ( n1082 , n1075 , n1081 );
or ( n1083 , n40 , n1080 );
nand ( n1084 , n1082 , n1083 );
nand ( n1085 , n1074 , n1084 );
nand ( n1086 , n1073 , n1085 );
not ( n1087 , n572 );
not ( n1088 , n1087 );
and ( n1089 , n1088 , n1030 );
xnor ( n1090 , n609 , n660 );
nor ( n1091 , n561 , n1090 );
nor ( n1092 , n1089 , n1091 );
not ( n1093 , n1092 );
xor ( n1094 , n1086 , n1093 );
buf ( n1095 , n931 );
not ( n1096 , n1095 );
not ( n1097 , n713 );
or ( n1098 , n1096 , n1097 );
buf ( n1099 , n704 );
buf ( n1100 , n1099 );
not ( n1101 , n765 );
buf ( n1102 , n698 );
not ( n1103 , n1102 );
and ( n1104 , n1101 , n1103 );
not ( n1105 , n1101 );
buf ( n1106 , n681 );
buf ( n1107 , n1106 );
and ( n1108 , n1105 , n1107 );
nor ( n1109 , n1104 , n1108 );
nand ( n1110 , n1100 , n1109 );
nand ( n1111 , n1098 , n1110 );
not ( n1112 , n1111 );
not ( n1113 , n1112 );
and ( n1114 , n1094 , n1113 );
not ( n1115 , n1094 );
not ( n1116 , n1113 );
and ( n1117 , n1115 , n1116 );
nor ( n1118 , n1114 , n1117 );
and ( n1119 , n1069 , n1118 );
not ( n1120 , n1069 );
not ( n1121 , n1118 );
and ( n1122 , n1120 , n1121 );
nor ( n1123 , n1119 , n1122 );
xnor ( n1124 , n966 , n1123 );
not ( n1125 , n1124 );
not ( n1126 , n705 );
not ( n1127 , n1126 );
not ( n1128 , n1127 );
buf ( n1129 , n681 );
buf ( n1130 , n1129 );
not ( n1131 , n1130 );
not ( n1132 , n1080 );
or ( n1133 , n1131 , n1132 );
not ( n1134 , n1103 );
or ( n1135 , n1134 , n1080 );
nand ( n1136 , n1133 , n1135 );
not ( n1137 , n1136 );
or ( n1138 , n1128 , n1137 );
buf ( n1139 , n686 );
not ( n1140 , n644 );
and ( n1141 , n1140 , n688 );
not ( n1142 , n1140 );
and ( n1143 , n1142 , n689 );
nor ( n1144 , n1141 , n1143 );
nand ( n1145 , n1139 , n1144 );
nand ( n1146 , n1138 , n1145 );
not ( n1147 , n1146 );
not ( n1148 , n776 );
and ( n1149 , n3 , n12 );
not ( n1150 , n3 );
and ( n1151 , n1150 , n28 );
nor ( n1152 , n1149 , n1151 );
xnor ( n1153 , n1152 , n42 );
and ( n1154 , n1148 , n1153 );
buf ( n1155 , n787 );
not ( n1156 , n42 );
not ( n1157 , n658 );
or ( n1158 , n1156 , n1157 );
nand ( n1159 , n3 , n11 );
not ( n1160 , n1159 );
not ( n1161 , n27 );
nor ( n1162 , n1161 , n3 );
or ( n1163 , n1160 , n1162 );
not ( n1164 , n42 );
nand ( n1165 , n1163 , n1164 );
nand ( n1166 , n1158 , n1165 );
nand ( n1167 , n1155 , n1166 );
not ( n1168 , n1167 );
nor ( n1169 , n1154 , n1168 );
not ( n1170 , n1169 );
not ( n1171 , n477 );
and ( n1172 , n3 , n17 );
not ( n1173 , n3 );
and ( n1174 , n1173 , n33 );
nor ( n1175 , n1172 , n1174 );
xor ( n1176 , n497 , n1175 );
not ( n1177 , n1176 );
or ( n1178 , n1171 , n1177 );
not ( n1179 , n476 );
and ( n1180 , n485 , n487 , n1179 );
and ( n1181 , n3 , n18 );
not ( n1182 , n3 );
and ( n1183 , n1182 , n34 );
nor ( n1184 , n1181 , n1183 );
and ( n1185 , n36 , n1184 );
not ( n1186 , n36 );
not ( n1187 , n18 );
and ( n1188 , n3 , n1187 );
not ( n1189 , n3 );
not ( n1190 , n34 );
and ( n1191 , n1189 , n1190 );
nor ( n1192 , n1188 , n1191 );
and ( n1193 , n1186 , n1192 );
or ( n1194 , n1185 , n1193 );
nand ( n1195 , n1180 , n1194 );
nand ( n1196 , n1178 , n1195 );
not ( n1197 , n1196 );
or ( n1198 , n1170 , n1197 );
not ( n1199 , n776 );
and ( n1200 , n1199 , n1153 );
nor ( n1201 , n1200 , n1168 );
or ( n1202 , n1201 , n1196 );
nand ( n1203 , n1198 , n1202 );
not ( n1204 , n1203 );
or ( n1205 , n1147 , n1204 );
not ( n1206 , n1201 );
nand ( n1207 , n1206 , n1196 );
nand ( n1208 , n1205 , n1207 );
not ( n1209 , n1208 );
not ( n1210 , n50 );
nor ( n1211 , n503 , n51 );
nor ( n1212 , n1210 , n1211 );
not ( n1213 , n1212 );
not ( n1214 , n19 );
and ( n1215 , n3 , n1214 );
not ( n1216 , n3 );
not ( n1217 , n35 );
and ( n1218 , n1216 , n1217 );
nor ( n1219 , n1215 , n1218 );
not ( n1220 , n1219 );
not ( n1221 , n1220 );
nand ( n1222 , n36 , n1221 );
not ( n1223 , n1222 );
and ( n1224 , n1213 , n1223 );
not ( n1225 , n1213 );
and ( n1226 , n1225 , n1222 );
nor ( n1227 , n1224 , n1226 );
not ( n1228 , n1227 );
not ( n1229 , n999 );
not ( n1230 , n552 );
not ( n1231 , n1230 );
not ( n1232 , n48 );
not ( n1233 , n1232 );
and ( n1234 , n1231 , n1233 );
not ( n1235 , n48 );
and ( n1236 , n1235 , n1230 );
nor ( n1237 , n1234 , n1236 );
or ( n1238 , n1229 , n1237 );
xor ( n1239 , n513 , n48 );
nand ( n1240 , n800 , n1239 );
nand ( n1241 , n1238 , n1240 );
and ( n1242 , n1228 , n1241 );
not ( n1243 , n1223 );
nor ( n1244 , n1243 , n1213 );
nor ( n1245 , n1242 , n1244 );
not ( n1246 , n1245 );
xnor ( n1247 , n897 , n40 );
not ( n1248 , n1247 );
not ( n1249 , n637 );
not ( n1250 , n1249 );
and ( n1251 , n1248 , n1250 );
nand ( n1252 , n668 , n670 , n672 );
not ( n1253 , n1252 );
not ( n1254 , n647 );
not ( n1255 , n923 );
or ( n1256 , n1254 , n1255 );
or ( n1257 , n647 , n916 );
nand ( n1258 , n1256 , n1257 );
and ( n1259 , n1253 , n1258 );
nor ( n1260 , n1251 , n1259 );
not ( n1261 , n1260 );
not ( n1262 , n1261 );
and ( n1263 , n3 , n15 );
not ( n1264 , n3 );
and ( n1265 , n1264 , n31 );
nor ( n1266 , n1263 , n1265 );
xnor ( n1267 , n609 , n1266 );
not ( n1268 , n1267 );
not ( n1269 , n559 );
not ( n1270 , n1269 );
and ( n1271 , n1268 , n1270 );
not ( n1272 , n571 );
and ( n1273 , n3 , n16 );
not ( n1274 , n3 );
and ( n1275 , n1274 , n32 );
nor ( n1276 , n1273 , n1275 );
and ( n1277 , n609 , n1276 );
not ( n1278 , n609 );
not ( n1279 , n1276 );
and ( n1280 , n1278 , n1279 );
nor ( n1281 , n1277 , n1280 );
and ( n1282 , n1272 , n1281 );
nor ( n1283 , n1271 , n1282 );
not ( n1284 , n1283 );
not ( n1285 , n1284 );
or ( n1286 , n1262 , n1285 );
not ( n1287 , n1260 );
not ( n1288 , n1283 );
or ( n1289 , n1287 , n1288 );
not ( n1290 , n755 );
not ( n1291 , n763 );
not ( n1292 , n695 );
or ( n1293 , n1291 , n1292 );
or ( n1294 , n763 , n603 );
nand ( n1295 , n1293 , n1294 );
not ( n1296 , n1295 );
or ( n1297 , n1290 , n1296 );
not ( n1298 , n936 );
and ( n1299 , n763 , n1298 );
not ( n1300 , n763 );
and ( n1301 , n1300 , n794 );
or ( n1302 , n1299 , n1301 );
nand ( n1303 , n1302 , n733 );
nand ( n1304 , n1297 , n1303 );
nand ( n1305 , n1289 , n1304 );
nand ( n1306 , n1286 , n1305 );
not ( n1307 , n1306 );
or ( n1308 , n1246 , n1307 );
or ( n1309 , n1245 , n1306 );
nand ( n1310 , n1308 , n1309 );
not ( n1311 , n1310 );
or ( n1312 , n1209 , n1311 );
not ( n1313 , n1245 );
nand ( n1314 , n1313 , n1306 );
nand ( n1315 , n1312 , n1314 );
not ( n1316 , n1315 );
xor ( n1317 , n861 , n839 );
not ( n1318 , n866 );
xnor ( n1319 , n1317 , n1318 );
not ( n1320 , n1319 );
not ( n1321 , n1320 );
not ( n1322 , n1139 );
not ( n1323 , n1136 );
or ( n1324 , n1322 , n1323 );
not ( n1325 , n1126 );
nand ( n1326 , n1325 , n942 );
nand ( n1327 , n1324 , n1326 );
not ( n1328 , n1327 );
not ( n1329 , n478 );
not ( n1330 , n989 );
or ( n1331 , n1329 , n1330 );
and ( n1332 , n721 , n497 );
not ( n1333 , n721 );
and ( n1334 , n1333 , n36 );
nor ( n1335 , n1332 , n1334 );
nand ( n1336 , n490 , n1335 );
nand ( n1337 , n1331 , n1336 );
not ( n1338 , n1337 );
not ( n1339 , n1020 );
or ( n1340 , n1338 , n1339 );
or ( n1341 , n1020 , n1337 );
nand ( n1342 , n1340 , n1341 );
xor ( n1343 , n1328 , n1342 );
not ( n1344 , n1343 );
not ( n1345 , n1344 );
or ( n1346 , n1321 , n1345 );
nand ( n1347 , n1319 , n1343 );
nand ( n1348 , n1346 , n1347 );
not ( n1349 , n1348 );
or ( n1350 , n1316 , n1349 );
nand ( n1351 , n1319 , n1344 );
nand ( n1352 , n1350 , n1351 );
not ( n1353 , n1352 );
and ( n1354 , n949 , n889 );
not ( n1355 , n949 );
not ( n1356 , n889 );
and ( n1357 , n1355 , n1356 );
nor ( n1358 , n1354 , n1357 );
not ( n1359 , n1358 );
not ( n1360 , n755 );
not ( n1361 , n835 );
or ( n1362 , n1360 , n1361 );
nand ( n1363 , n733 , n1295 );
nand ( n1364 , n1362 , n1363 );
not ( n1365 , n1364 );
and ( n1366 , n788 , n854 );
not ( n1367 , n775 );
nand ( n1368 , n1367 , n1166 );
not ( n1369 , n1368 );
nor ( n1370 , n1366 , n1369 );
not ( n1371 , n1370 );
not ( n1372 , n799 );
not ( n1373 , n1014 );
or ( n1374 , n1372 , n1373 );
not ( n1375 , n998 );
nand ( n1376 , n1239 , n1375 );
nand ( n1377 , n1374 , n1376 );
not ( n1378 , n1377 );
or ( n1379 , n1371 , n1378 );
and ( n1380 , n788 , n854 );
nor ( n1381 , n1380 , n1369 );
or ( n1382 , n1381 , n1377 );
nand ( n1383 , n1379 , n1382 );
not ( n1384 , n1383 );
or ( n1385 , n1365 , n1384 );
not ( n1386 , n1381 );
nand ( n1387 , n1386 , n1377 );
nand ( n1388 , n1385 , n1387 );
not ( n1389 , n1388 );
and ( n1390 , n3 , n18 );
not ( n1391 , n3 );
and ( n1392 , n1391 , n34 );
nor ( n1393 , n1390 , n1392 );
buf ( n1394 , n1393 );
not ( n1395 , n1394 );
nand ( n1396 , n36 , n1395 );
nand ( n1397 , n50 , n1396 );
not ( n1398 , n1397 );
not ( n1399 , n489 );
not ( n1400 , n1176 );
or ( n1401 , n1399 , n1400 );
nand ( n1402 , n477 , n1335 );
nand ( n1403 , n1401 , n1402 );
not ( n1404 , n1403 );
or ( n1405 , n1398 , n1404 );
not ( n1406 , n50 );
not ( n1407 , n1396 );
nand ( n1408 , n1406 , n1407 );
nand ( n1409 , n1405 , n1408 );
not ( n1410 , n1409 );
not ( n1411 , n1410 );
and ( n1412 , n1389 , n1411 );
not ( n1413 , n1409 );
and ( n1414 , n1413 , n1388 );
nor ( n1415 , n1412 , n1414 );
not ( n1416 , n1415 );
not ( n1417 , n1416 );
or ( n1418 , n1359 , n1417 );
not ( n1419 , n1413 );
nand ( n1420 , n1419 , n1388 );
nand ( n1421 , n1418 , n1420 );
not ( n1422 , n1421 );
not ( n1423 , n1422 );
not ( n1424 , n868 );
xor ( n1425 , n1424 , n955 );
xnor ( n1426 , n1425 , n823 );
not ( n1427 , n1426 );
not ( n1428 , n1427 );
or ( n1429 , n1423 , n1428 );
nand ( n1430 , n1421 , n1426 );
nand ( n1431 , n1429 , n1430 );
not ( n1432 , n1431 );
or ( n1433 , n1353 , n1432 );
nand ( n1434 , n1421 , n1427 );
nand ( n1435 , n1433 , n1434 );
xor ( n1436 , n727 , n724 );
xor ( n1437 , n1436 , n676 );
not ( n1438 , n1437 );
not ( n1439 , n1327 );
not ( n1440 , n1342 );
or ( n1441 , n1439 , n1440 );
not ( n1442 , n1020 );
nand ( n1443 , n1442 , n1337 );
nand ( n1444 , n1441 , n1443 );
not ( n1445 , n1444 );
not ( n1446 , n991 );
and ( n1447 , n1035 , n1446 );
not ( n1448 , n1035 );
and ( n1449 , n1448 , n991 );
nor ( n1450 , n1447 , n1449 );
not ( n1451 , n1450 );
and ( n1452 , n1445 , n1451 );
and ( n1453 , n1444 , n1450 );
nor ( n1454 , n1452 , n1453 );
not ( n1455 , n1454 );
not ( n1456 , n1455 );
or ( n1457 , n1438 , n1456 );
not ( n1458 , n1444 );
or ( n1459 , n1458 , n1450 );
nand ( n1460 , n1457 , n1459 );
not ( n1461 , n1460 );
not ( n1462 , n1461 );
and ( n1463 , n1435 , n1462 );
not ( n1464 , n1435 );
and ( n1465 , n1464 , n1461 );
nor ( n1466 , n1463 , n1465 );
not ( n1467 , n1466 );
or ( n1468 , n1125 , n1467 );
nand ( n1469 , n1462 , n1435 );
nand ( n1470 , n1468 , n1469 );
not ( n1471 , n477 );
not ( n1472 , n1471 );
not ( n1473 , n1472 );
not ( n1474 , n36 );
not ( n1475 , n878 );
or ( n1476 , n1474 , n1475 );
or ( n1477 , n36 , n878 );
nand ( n1478 , n1476 , n1477 );
not ( n1479 , n1478 );
or ( n1480 , n1473 , n1479 );
nand ( n1481 , n490 , n1065 );
nand ( n1482 , n1480 , n1481 );
not ( n1483 , n856 );
not ( n1484 , n554 );
nor ( n1485 , n42 , n1484 );
not ( n1486 , n1485 );
nand ( n1487 , n42 , n555 );
nand ( n1488 , n1486 , n1487 );
not ( n1489 , n1488 );
or ( n1490 , n1483 , n1489 );
buf ( n1491 , n776 );
not ( n1492 , n1491 );
nand ( n1493 , n1492 , n1048 );
nand ( n1494 , n1490 , n1493 );
xor ( n1495 , n1482 , n1494 );
not ( n1496 , n562 );
not ( n1497 , n38 );
buf ( n1498 , n644 );
buf ( n1499 , n1498 );
not ( n1500 , n1499 );
or ( n1501 , n1497 , n1500 );
or ( n1502 , n38 , n1499 );
nand ( n1503 , n1501 , n1502 );
not ( n1504 , n1503 );
or ( n1505 , n1496 , n1504 );
not ( n1506 , n1087 );
buf ( n1507 , n1506 );
not ( n1508 , n1090 );
nand ( n1509 , n1507 , n1508 );
nand ( n1510 , n1505 , n1509 );
xor ( n1511 , n1495 , n1510 );
not ( n1512 , n1511 );
not ( n1513 , n1512 );
not ( n1514 , n871 );
not ( n1515 , n1514 );
not ( n1516 , n1515 );
not ( n1517 , n1084 );
or ( n1518 , n1516 , n1517 );
not ( n1519 , n640 );
not ( n1520 , n795 );
xnor ( n1521 , n40 , n1520 );
nand ( n1522 , n1519 , n1521 );
nand ( n1523 , n1518 , n1522 );
not ( n1524 , n1100 );
not ( n1525 , n1107 );
not ( n1526 , n738 );
or ( n1527 , n1525 , n1526 );
not ( n1528 , n710 );
nand ( n1529 , n1528 , n504 );
nand ( n1530 , n1527 , n1529 );
not ( n1531 , n1530 );
or ( n1532 , n1524 , n1531 );
nand ( n1533 , n1095 , n1109 );
nand ( n1534 , n1532 , n1533 );
not ( n1535 , n756 );
not ( n1536 , n761 );
or ( n1537 , n1535 , n1536 );
nand ( n1538 , n1537 , n46 );
and ( n1539 , n1534 , n1538 );
not ( n1540 , n1534 );
not ( n1541 , n1538 );
and ( n1542 , n1540 , n1541 );
nor ( n1543 , n1539 , n1542 );
xor ( n1544 , n1523 , n1543 );
not ( n1545 , n1067 );
not ( n1546 , n1054 );
not ( n1547 , n1040 );
and ( n1548 , n1546 , n1547 );
not ( n1549 , n1546 );
and ( n1550 , n1549 , n1040 );
nor ( n1551 , n1548 , n1550 );
not ( n1552 , n1551 );
or ( n1553 , n1545 , n1552 );
nand ( n1554 , n1547 , n1546 );
nand ( n1555 , n1553 , n1554 );
and ( n1556 , n1544 , n1555 );
not ( n1557 , n1544 );
not ( n1558 , n1555 );
and ( n1559 , n1557 , n1558 );
nor ( n1560 , n1556 , n1559 );
not ( n1561 , n1560 );
or ( n1562 , n1513 , n1561 );
not ( n1563 , n1560 );
nand ( n1564 , n1511 , n1563 );
nand ( n1565 , n1562 , n1564 );
not ( n1566 , n1118 );
not ( n1567 , n1069 );
or ( n1568 , n1566 , n1567 );
not ( n1569 , n1038 );
not ( n1570 , n1068 );
nand ( n1571 , n1569 , n1570 );
nand ( n1572 , n1568 , n1571 );
not ( n1573 , n1572 );
not ( n1574 , n1573 );
buf ( n1575 , n973 );
not ( n1576 , n1575 );
nand ( n1577 , n36 , n1576 );
not ( n1578 , n1577 );
not ( n1579 , n749 );
or ( n1580 , n1578 , n1579 );
or ( n1581 , n1577 , n749 );
nand ( n1582 , n1580 , n1581 );
not ( n1583 , n1093 );
not ( n1584 , n1113 );
or ( n1585 , n1583 , n1584 );
not ( n1586 , n1092 );
not ( n1587 , n1112 );
or ( n1588 , n1586 , n1587 );
nand ( n1589 , n1588 , n1086 );
nand ( n1590 , n1585 , n1589 );
not ( n1591 , n1590 );
and ( n1592 , n1582 , n1591 );
not ( n1593 , n1582 );
and ( n1594 , n1593 , n1590 );
nor ( n1595 , n1592 , n1594 );
not ( n1596 , n1595 );
not ( n1597 , n816 );
not ( n1598 , n754 );
or ( n1599 , n1597 , n1598 );
not ( n1600 , n729 );
nand ( n1601 , n752 , n1600 );
nand ( n1602 , n1599 , n1601 );
not ( n1603 , n1602 );
or ( n1604 , n1596 , n1603 );
or ( n1605 , n1595 , n1602 );
nand ( n1606 , n1604 , n1605 );
not ( n1607 , n1606 );
or ( n1608 , n1574 , n1607 );
not ( n1609 , n1606 );
nand ( n1610 , n1609 , n1572 );
nand ( n1611 , n1608 , n1610 );
not ( n1612 , n1611 );
xor ( n1613 , n1565 , n1612 );
not ( n1614 , n1123 );
not ( n1615 , n821 );
and ( n1616 , n965 , n1615 );
not ( n1617 , n965 );
and ( n1618 , n1617 , n821 );
nor ( n1619 , n1616 , n1618 );
not ( n1620 , n1619 );
or ( n1621 , n1614 , n1620 );
nand ( n1622 , n1615 , n965 );
nand ( n1623 , n1621 , n1622 );
xnor ( n1624 , n1613 , n1623 );
nand ( n1625 , n1470 , n1624 );
xor ( n1626 , n1565 , n1611 );
and ( n1627 , n1623 , n1626 );
and ( n1628 , n1565 , n1611 );
nor ( n1629 , n1627 , n1628 );
not ( n1630 , n1510 );
not ( n1631 , n1495 );
or ( n1632 , n1630 , n1631 );
nand ( n1633 , n1482 , n1494 );
nand ( n1634 , n1632 , n1633 );
not ( n1635 , n1523 );
not ( n1636 , n1543 );
or ( n1637 , n1635 , n1636 );
not ( n1638 , n1541 );
nand ( n1639 , n1638 , n1534 );
nand ( n1640 , n1637 , n1639 );
not ( n1641 , n1640 );
and ( n1642 , n1634 , n1641 );
not ( n1643 , n1634 );
and ( n1644 , n1643 , n1640 );
nor ( n1645 , n1642 , n1644 );
not ( n1646 , n1139 );
not ( n1647 , n1530 );
or ( n1648 , n1646 , n1647 );
not ( n1649 , n1130 );
not ( n1650 , n1649 );
nand ( n1651 , n1650 , n1100 );
nand ( n1652 , n1648 , n1651 );
not ( n1653 , n38 );
not ( n1654 , n1080 );
or ( n1655 , n1653 , n1654 );
or ( n1656 , n38 , n1080 );
nand ( n1657 , n1655 , n1656 );
nand ( n1658 , n1022 , n1657 );
nand ( n1659 , n1088 , n1503 );
nand ( n1660 , n1658 , n1659 );
xor ( n1661 , n1652 , n1660 );
not ( n1662 , n490 );
not ( n1663 , n1478 );
or ( n1664 , n1662 , n1663 );
not ( n1665 , n665 );
and ( n1666 , n1665 , n497 );
not ( n1667 , n1665 );
and ( n1668 , n1667 , n36 );
nor ( n1669 , n1666 , n1668 );
nand ( n1670 , n478 , n1669 );
nand ( n1671 , n1664 , n1670 );
xor ( n1672 , n1661 , n1671 );
and ( n1673 , n1645 , n1672 );
not ( n1674 , n1645 );
not ( n1675 , n1672 );
and ( n1676 , n1674 , n1675 );
nor ( n1677 , n1673 , n1676 );
not ( n1678 , n1572 );
not ( n1679 , n1606 );
or ( n1680 , n1678 , n1679 );
not ( n1681 , n1595 );
nand ( n1682 , n1681 , n1602 );
nand ( n1683 , n1680 , n1682 );
not ( n1684 , n1683 );
xor ( n1685 , n1677 , n1684 );
not ( n1686 , n1061 );
not ( n1687 , n1686 );
not ( n1688 , n1687 );
and ( n1689 , n1688 , n36 );
buf ( n1690 , n1199 );
not ( n1691 , n1690 );
not ( n1692 , n1488 );
or ( n1693 , n1691 , n1692 );
buf ( n1694 , n862 );
not ( n1695 , n42 );
not ( n1696 , n516 );
or ( n1697 , n1695 , n1696 );
or ( n1698 , n42 , n516 );
nand ( n1699 , n1697 , n1698 );
nand ( n1700 , n1694 , n1699 );
nand ( n1701 , n1693 , n1700 );
not ( n1702 , n1701 );
xor ( n1703 , n1689 , n1702 );
not ( n1704 , n1515 );
not ( n1705 , n1521 );
or ( n1706 , n1704 , n1705 );
buf ( n1707 , n640 );
not ( n1708 , n1707 );
not ( n1709 , n40 );
not ( n1710 , n1044 );
or ( n1711 , n1709 , n1710 );
or ( n1712 , n40 , n604 );
nand ( n1713 , n1711 , n1712 );
nand ( n1714 , n1708 , n1713 );
nand ( n1715 , n1706 , n1714 );
xnor ( n1716 , n1703 , n1715 );
not ( n1717 , n1716 );
not ( n1718 , n1582 );
not ( n1719 , n1591 );
not ( n1720 , n1719 );
or ( n1721 , n1718 , n1720 );
not ( n1722 , n1577 );
not ( n1723 , n752 );
nand ( n1724 , n1722 , n1723 );
nand ( n1725 , n1721 , n1724 );
not ( n1726 , n1725 );
or ( n1727 , n1717 , n1726 );
or ( n1728 , n1716 , n1725 );
nand ( n1729 , n1727 , n1728 );
not ( n1730 , n1511 );
not ( n1731 , n1560 );
or ( n1732 , n1730 , n1731 );
not ( n1733 , n1558 );
nand ( n1734 , n1733 , n1544 );
nand ( n1735 , n1732 , n1734 );
xor ( n1736 , n1729 , n1735 );
xnor ( n1737 , n1685 , n1736 );
nor ( n1738 , n1629 , n1737 );
not ( n1739 , n1736 );
not ( n1740 , n1677 );
and ( n1741 , n1683 , n1740 );
not ( n1742 , n1683 );
and ( n1743 , n1742 , n1677 );
nor ( n1744 , n1741 , n1743 );
not ( n1745 , n1744 );
or ( n1746 , n1739 , n1745 );
not ( n1747 , n1684 );
nand ( n1748 , n1740 , n1747 );
nand ( n1749 , n1746 , n1748 );
not ( n1750 , n1749 );
not ( n1751 , n479 );
buf ( n1752 , n1499 );
xnor ( n1753 , n36 , n1752 );
and ( n1754 , n1751 , n1753 );
not ( n1755 , n1669 );
nor ( n1756 , n491 , n1755 );
nor ( n1757 , n1754 , n1756 );
not ( n1758 , n1757 );
not ( n1759 , n878 );
not ( n1760 , n1759 );
not ( n1761 , n1760 );
nand ( n1762 , n1761 , n36 );
not ( n1763 , n1762 );
not ( n1764 , n1763 );
not ( n1765 , n639 );
not ( n1766 , n40 );
not ( n1767 , n555 );
or ( n1768 , n1766 , n1767 );
or ( n1769 , n40 , n555 );
nand ( n1770 , n1768 , n1769 );
not ( n1771 , n1770 );
or ( n1772 , n1765 , n1771 );
nand ( n1773 , n871 , n1713 );
nand ( n1774 , n1772 , n1773 );
not ( n1775 , n1774 );
not ( n1776 , n1775 );
or ( n1777 , n1764 , n1776 );
not ( n1778 , n1762 );
or ( n1779 , n1778 , n1775 );
nand ( n1780 , n1777 , n1779 );
not ( n1781 , n1780 );
and ( n1782 , n1758 , n1781 );
and ( n1783 , n1757 , n1780 );
nor ( n1784 , n1782 , n1783 );
not ( n1785 , n1702 );
not ( n1786 , n1652 );
not ( n1787 , n1660 );
or ( n1788 , n1786 , n1787 );
or ( n1789 , n1652 , n1660 );
nand ( n1790 , n1789 , n1671 );
nand ( n1791 , n1788 , n1790 );
xor ( n1792 , n1785 , n1791 );
xor ( n1793 , n1784 , n1792 );
not ( n1794 , n1793 );
and ( n1795 , n1715 , n1703 );
and ( n1796 , n1689 , n1702 );
nor ( n1797 , n1795 , n1796 );
not ( n1798 , n1797 );
not ( n1799 , n1126 );
not ( n1800 , n1139 );
not ( n1801 , n1800 );
or ( n1802 , n1799 , n1801 );
nand ( n1803 , n1802 , n1650 );
not ( n1804 , n1694 );
not ( n1805 , n42 );
not ( n1806 , n504 );
not ( n1807 , n1806 );
or ( n1808 , n1805 , n1807 );
or ( n1809 , n42 , n1806 );
nand ( n1810 , n1808 , n1809 );
not ( n1811 , n1810 );
or ( n1812 , n1804 , n1811 );
nand ( n1813 , n1690 , n1699 );
nand ( n1814 , n1812 , n1813 );
xor ( n1815 , n1803 , n1814 );
not ( n1816 , n1507 );
not ( n1817 , n1657 );
or ( n1818 , n1816 , n1817 );
buf ( n1819 , n1022 );
buf ( n1820 , n1520 );
and ( n1821 , n1820 , n609 );
not ( n1822 , n1820 );
and ( n1823 , n1822 , n38 );
nor ( n1824 , n1821 , n1823 );
nand ( n1825 , n1819 , n1824 );
nand ( n1826 , n1818 , n1825 );
and ( n1827 , n1815 , n1826 );
not ( n1828 , n1815 );
not ( n1829 , n1826 );
and ( n1830 , n1828 , n1829 );
nor ( n1831 , n1827 , n1830 );
not ( n1832 , n1831 );
or ( n1833 , n1798 , n1832 );
or ( n1834 , n1797 , n1831 );
nand ( n1835 , n1833 , n1834 );
not ( n1836 , n1835 );
or ( n1837 , n1794 , n1836 );
or ( n1838 , n1835 , n1793 );
nand ( n1839 , n1837 , n1838 );
not ( n1840 , n1672 );
not ( n1841 , n1645 );
not ( n1842 , n1841 );
or ( n1843 , n1840 , n1842 );
not ( n1844 , n1641 );
nand ( n1845 , n1844 , n1634 );
nand ( n1846 , n1843 , n1845 );
and ( n1847 , n1839 , n1846 );
not ( n1848 , n1839 );
not ( n1849 , n1846 );
and ( n1850 , n1848 , n1849 );
nor ( n1851 , n1847 , n1850 );
not ( n1852 , n1851 );
not ( n1853 , n1729 );
not ( n1854 , n1735 );
or ( n1855 , n1853 , n1854 );
not ( n1856 , n1716 );
nand ( n1857 , n1856 , n1725 );
nand ( n1858 , n1855 , n1857 );
not ( n1859 , n1858 );
not ( n1860 , n1859 );
and ( n1861 , n1852 , n1860 );
and ( n1862 , n1859 , n1851 );
nor ( n1863 , n1861 , n1862 );
nor ( n1864 , n1750 , n1863 );
nor ( n1865 , n1738 , n1864 );
nand ( n1866 , n1625 , n1865 );
not ( n1867 , n1866 );
and ( n1868 , n1454 , n1437 );
not ( n1869 , n1454 );
not ( n1870 , n1437 );
and ( n1871 , n1869 , n1870 );
nor ( n1872 , n1868 , n1871 );
not ( n1873 , n762 );
xor ( n1874 , n763 , n1079 );
not ( n1875 , n1874 );
or ( n1876 , n1873 , n1875 );
buf ( n1877 , n1302 );
nand ( n1878 , n757 , n1877 );
nand ( n1879 , n1876 , n1878 );
not ( n1880 , n1879 );
not ( n1881 , n870 );
and ( n1882 , n40 , n983 );
not ( n1883 , n40 );
and ( n1884 , n3 , n15 );
not ( n1885 , n3 );
and ( n1886 , n1885 , n31 );
nor ( n1887 , n1884 , n1886 );
and ( n1888 , n1883 , n1887 );
nor ( n1889 , n1882 , n1888 );
not ( n1890 , n1889 );
or ( n1891 , n1881 , n1890 );
not ( n1892 , n885 );
nand ( n1893 , n1892 , n1258 );
nand ( n1894 , n1891 , n1893 );
not ( n1895 , n776 );
not ( n1896 , n1895 );
and ( n1897 , n42 , n903 );
not ( n1898 , n42 );
and ( n1899 , n1898 , n904 );
or ( n1900 , n1897 , n1899 );
not ( n1901 , n1900 );
or ( n1902 , n1896 , n1901 );
buf ( n1903 , n1155 );
nand ( n1904 , n1903 , n1153 );
nand ( n1905 , n1902 , n1904 );
and ( n1906 , n1894 , n1905 );
not ( n1907 , n1894 );
not ( n1908 , n1905 );
and ( n1909 , n1907 , n1908 );
nor ( n1910 , n1906 , n1909 );
not ( n1911 , n1910 );
or ( n1912 , n1880 , n1911 );
not ( n1913 , n1908 );
nand ( n1914 , n1894 , n1913 );
nand ( n1915 , n1912 , n1914 );
not ( n1916 , n1915 );
buf ( n1917 , n1221 );
nand ( n1918 , n37 , n38 );
not ( n1919 , n1918 );
or ( n1920 , n1917 , n1919 );
nor ( n1921 , n37 , n38 );
not ( n1922 , n1921 );
nand ( n1923 , n1920 , n1922 );
nand ( n1924 , n1923 , n36 );
not ( n1925 , n1924 );
not ( n1926 , n51 );
not ( n1927 , n1406 );
not ( n1928 , n737 );
or ( n1929 , n1927 , n1928 );
or ( n1930 , n1406 , n504 );
nand ( n1931 , n1929 , n1930 );
not ( n1932 , n1931 );
or ( n1933 , n1926 , n1932 );
not ( n1934 , n51 );
nand ( n1935 , n1934 , n50 );
buf ( n1936 , n1935 );
not ( n1937 , n1936 );
and ( n1938 , n1406 , n514 );
not ( n1939 , n1406 );
and ( n1940 , n1939 , n765 );
nor ( n1941 , n1938 , n1940 );
nand ( n1942 , n1937 , n1941 );
nand ( n1943 , n1933 , n1942 );
not ( n1944 , n1943 );
not ( n1945 , n1944 );
nand ( n1946 , n1925 , n1945 );
not ( n1947 , n1946 );
not ( n1948 , n1947 );
not ( n1949 , n1144 );
not ( n1950 , n1099 );
or ( n1951 , n1949 , n1950 );
not ( n1952 , n689 );
not ( n1953 , n659 );
or ( n1954 , n1952 , n1953 );
or ( n1955 , n699 , n659 );
nand ( n1956 , n1954 , n1955 );
nand ( n1957 , n686 , n1956 );
nand ( n1958 , n1951 , n1957 );
not ( n1959 , n1237 );
not ( n1960 , n1017 );
not ( n1961 , n1960 );
and ( n1962 , n1959 , n1961 );
not ( n1963 , n48 );
not ( n1964 , n1963 );
not ( n1965 , n695 );
or ( n1966 , n1964 , n1965 );
not ( n1967 , n48 );
or ( n1968 , n1967 , n603 );
nand ( n1969 , n1966 , n1968 );
and ( n1970 , n999 , n1969 );
nor ( n1971 , n1962 , n1970 );
not ( n1972 , n1971 );
nand ( n1973 , n1958 , n1972 );
not ( n1974 , n1958 );
not ( n1975 , n1974 );
not ( n1976 , n1971 );
or ( n1977 , n1975 , n1976 );
not ( n1978 , n1180 );
not ( n1979 , n497 );
not ( n1980 , n19 );
and ( n1981 , n3 , n1980 );
not ( n1982 , n3 );
not ( n1983 , n35 );
and ( n1984 , n1982 , n1983 );
nor ( n1985 , n1981 , n1984 );
not ( n1986 , n1985 );
or ( n1987 , n1979 , n1986 );
or ( n1988 , n497 , n1985 );
nand ( n1989 , n1987 , n1988 );
not ( n1990 , n1989 );
or ( n1991 , n1978 , n1990 );
nand ( n1992 , n477 , n1194 );
nand ( n1993 , n1991 , n1992 );
nand ( n1994 , n1977 , n1993 );
nand ( n1995 , n1973 , n1994 );
not ( n1996 , n1995 );
not ( n1997 , n1996 );
or ( n1998 , n1948 , n1997 );
not ( n1999 , n1973 );
not ( n2000 , n1994 );
or ( n2001 , n1999 , n2000 );
nand ( n2002 , n2001 , n1946 );
nand ( n2003 , n1998 , n2002 );
not ( n2004 , n2003 );
or ( n2005 , n1916 , n2004 );
nand ( n2006 , n1947 , n1995 );
nand ( n2007 , n2005 , n2006 );
not ( n2008 , n2007 );
not ( n2009 , n50 );
not ( n2010 , n1396 );
or ( n2011 , n2009 , n2010 );
nand ( n2012 , n1406 , n1407 );
nand ( n2013 , n2011 , n2012 );
not ( n2014 , n1403 );
and ( n2015 , n2013 , n2014 );
not ( n2016 , n2013 );
and ( n2017 , n2016 , n1403 );
nor ( n2018 , n2015 , n2017 );
not ( n2019 , n2018 );
not ( n2020 , n1364 );
and ( n2021 , n1383 , n2020 );
not ( n2022 , n1383 );
and ( n2023 , n2022 , n1364 );
nor ( n2024 , n2021 , n2023 );
not ( n2025 , n2024 );
or ( n2026 , n2019 , n2025 );
or ( n2027 , n2018 , n2024 );
nand ( n2028 , n2026 , n2027 );
not ( n2029 , n2028 );
or ( n2030 , n2008 , n2029 );
not ( n2031 , n2024 );
nand ( n2032 , n2018 , n2031 );
nand ( n2033 , n2030 , n2032 );
not ( n2034 , n2033 );
xor ( n2035 , n1358 , n1416 );
not ( n2036 , n1328 );
not ( n2037 , n639 );
not ( n2038 , n882 );
or ( n2039 , n2037 , n2038 );
not ( n2040 , n1247 );
nand ( n2041 , n674 , n2040 );
nand ( n2042 , n2039 , n2041 );
not ( n2043 , n573 );
not ( n2044 , n1267 );
not ( n2045 , n2044 );
or ( n2046 , n2043 , n2045 );
nand ( n2047 , n1022 , n925 );
nand ( n2048 , n2046 , n2047 );
xor ( n2049 , n2042 , n2048 );
not ( n2050 , n2049 );
or ( n2051 , n2036 , n2050 );
nand ( n2052 , n2042 , n2048 );
nand ( n2053 , n2051 , n2052 );
not ( n2054 , n2053 );
xnor ( n2055 , n2035 , n2054 );
not ( n2056 , n2055 );
or ( n2057 , n2034 , n2056 );
not ( n2058 , n2054 );
xor ( n2059 , n1416 , n1358 );
nand ( n2060 , n2058 , n2059 );
nand ( n2061 , n2057 , n2060 );
not ( n2062 , n2061 );
xor ( n2063 , n1872 , n2062 );
and ( n2064 , n1431 , n1352 );
not ( n2065 , n1431 );
not ( n2066 , n1352 );
and ( n2067 , n2065 , n2066 );
nor ( n2068 , n2064 , n2067 );
xnor ( n2069 , n2063 , n2068 );
xor ( n2070 , n2055 , n2033 );
and ( n2071 , n1348 , n1315 );
not ( n2072 , n1348 );
not ( n2073 , n1315 );
and ( n2074 , n2072 , n2073 );
nor ( n2075 , n2071 , n2074 );
xor ( n2076 , n1304 , n1261 );
xor ( n2077 , n2076 , n1284 );
not ( n2078 , n1227 );
not ( n2079 , n2078 );
not ( n2080 , n1241 );
not ( n2081 , n2080 );
or ( n2082 , n2079 , n2081 );
or ( n2083 , n2080 , n2078 );
nand ( n2084 , n2082 , n2083 );
xor ( n2085 , n1146 , n1203 );
xor ( n2086 , n2084 , n2085 );
and ( n2087 , n2077 , n2086 );
and ( n2088 , n2084 , n2085 );
nor ( n2089 , n2087 , n2088 );
not ( n2090 , n2089 );
not ( n2091 , n2090 );
not ( n2092 , n1327 );
not ( n2093 , n2049 );
or ( n2094 , n2092 , n2093 );
or ( n2095 , n1327 , n2049 );
nand ( n2096 , n2094 , n2095 );
not ( n2097 , n2096 );
not ( n2098 , n1208 );
not ( n2099 , n1310 );
not ( n2100 , n2099 );
or ( n2101 , n2098 , n2100 );
not ( n2102 , n1208 );
nand ( n2103 , n2102 , n1310 );
nand ( n2104 , n2101 , n2103 );
not ( n2105 , n2104 );
not ( n2106 , n2105 );
or ( n2107 , n2097 , n2106 );
not ( n2108 , n2104 );
or ( n2109 , n2096 , n2108 );
nand ( n2110 , n2107 , n2109 );
not ( n2111 , n2110 );
or ( n2112 , n2091 , n2111 );
not ( n2113 , n2108 );
nand ( n2114 , n2096 , n2113 );
nand ( n2115 , n2112 , n2114 );
xor ( n2116 , n2075 , n2115 );
and ( n2117 , n2070 , n2116 );
and ( n2118 , n2075 , n2115 );
nor ( n2119 , n2117 , n2118 );
and ( n2120 , n2069 , n2119 );
and ( n2121 , n2007 , n2028 );
not ( n2122 , n2007 );
not ( n2123 , n2028 );
and ( n2124 , n2122 , n2123 );
nor ( n2125 , n2121 , n2124 );
not ( n2126 , n2110 );
not ( n2127 , n2089 );
and ( n2128 , n2126 , n2127 );
and ( n2129 , n2089 , n2110 );
nor ( n2130 , n2128 , n2129 );
not ( n2131 , n2130 );
xor ( n2132 , n2125 , n2131 );
and ( n2133 , n1910 , n1879 );
not ( n2134 , n1910 );
not ( n2135 , n1879 );
and ( n2136 , n2134 , n2135 );
nor ( n2137 , n2133 , n2136 );
not ( n2138 , n2137 );
xor ( n2139 , n1993 , n1958 );
xor ( n2140 , n2139 , n1972 );
not ( n2141 , n2140 );
not ( n2142 , n733 );
not ( n2143 , n46 );
not ( n2144 , n645 );
or ( n2145 , n2143 , n2144 );
or ( n2146 , n46 , n1498 );
nand ( n2147 , n2145 , n2146 );
not ( n2148 , n2147 );
or ( n2149 , n2142 , n2148 );
not ( n2150 , n745 );
not ( n2151 , n2150 );
nand ( n2152 , n2151 , n1874 );
nand ( n2153 , n2149 , n2152 );
not ( n2154 , n2153 );
not ( n2155 , n2154 );
not ( n2156 , n2155 );
not ( n2157 , n1199 );
not ( n2158 , n42 );
not ( n2159 , n969 );
or ( n2160 , n2158 , n2159 );
or ( n2161 , n42 , n969 );
nand ( n2162 , n2160 , n2161 );
not ( n2163 , n2162 );
or ( n2164 , n2157 , n2163 );
buf ( n2165 , n788 );
nand ( n2166 , n2165 , n1900 );
nand ( n2167 , n2164 , n2166 );
not ( n2168 , n2167 );
or ( n2169 , n2156 , n2168 );
not ( n2170 , n2154 );
not ( n2171 , n2167 );
not ( n2172 , n2171 );
or ( n2173 , n2170 , n2172 );
not ( n2174 , n1139 );
not ( n2175 , n1102 );
not ( n2176 , n1027 );
or ( n2177 , n2175 , n2176 );
or ( n2178 , n710 , n1027 );
nand ( n2179 , n2177 , n2178 );
not ( n2180 , n2179 );
or ( n2181 , n2174 , n2180 );
not ( n2182 , n1126 );
nand ( n2183 , n2182 , n1956 );
nand ( n2184 , n2181 , n2183 );
nand ( n2185 , n2173 , n2184 );
nand ( n2186 , n2169 , n2185 );
not ( n2187 , n2186 );
not ( n2188 , n2187 );
or ( n2189 , n2141 , n2188 );
not ( n2190 , n2186 );
or ( n2191 , n2190 , n2140 );
nand ( n2192 , n2189 , n2191 );
not ( n2193 , n2192 );
or ( n2194 , n2138 , n2193 );
not ( n2195 , n2190 );
nand ( n2196 , n2195 , n2140 );
nand ( n2197 , n2194 , n2196 );
not ( n2198 , n2197 );
xor ( n2199 , n1915 , n2003 );
not ( n2200 , n800 );
not ( n2201 , n1969 );
or ( n2202 , n2200 , n2201 );
and ( n2203 , n48 , n794 );
not ( n2204 , n48 );
and ( n2205 , n2204 , n1298 );
or ( n2206 , n2203 , n2205 );
nand ( n2207 , n804 , n805 );
not ( n2208 , n2207 );
nand ( n2209 , n2206 , n2208 );
nand ( n2210 , n2202 , n2209 );
not ( n2211 , n1937 );
not ( n2212 , n1406 );
not ( n2213 , n707 );
or ( n2214 , n2212 , n2213 );
or ( n2215 , n1406 , n707 );
nand ( n2216 , n2214 , n2215 );
not ( n2217 , n2216 );
or ( n2218 , n2211 , n2217 );
nand ( n2219 , n51 , n1941 );
nand ( n2220 , n2218 , n2219 );
xor ( n2221 , n2210 , n2220 );
not ( n2222 , n1220 );
not ( n2223 , n2222 );
not ( n2224 , n2223 );
and ( n2225 , n1472 , n2224 );
and ( n2226 , n2221 , n2225 );
and ( n2227 , n2210 , n2220 );
or ( n2228 , n2226 , n2227 );
not ( n2229 , n2228 );
not ( n2230 , n1506 );
not ( n2231 , n38 );
not ( n2232 , n845 );
or ( n2233 , n2231 , n2232 );
or ( n2234 , n38 , n845 );
nand ( n2235 , n2233 , n2234 );
not ( n2236 , n2235 );
or ( n2237 , n2230 , n2236 );
nand ( n2238 , n1022 , n1281 );
nand ( n2239 , n2237 , n2238 );
not ( n2240 , n2239 );
and ( n2241 , n1944 , n1925 );
not ( n2242 , n1944 );
and ( n2243 , n2242 , n1924 );
nor ( n2244 , n2241 , n2243 );
not ( n2245 , n2244 );
and ( n2246 , n2240 , n2245 );
not ( n2247 , n2240 );
and ( n2248 , n2247 , n2244 );
nor ( n2249 , n2246 , n2248 );
not ( n2250 , n2249 );
not ( n2251 , n2250 );
or ( n2252 , n2229 , n2251 );
not ( n2253 , n2240 );
nand ( n2254 , n2253 , n2245 );
nand ( n2255 , n2252 , n2254 );
not ( n2256 , n2255 );
and ( n2257 , n2199 , n2256 );
not ( n2258 , n2199 );
and ( n2259 , n2258 , n2255 );
nor ( n2260 , n2257 , n2259 );
not ( n2261 , n2260 );
not ( n2262 , n2261 );
or ( n2263 , n2198 , n2262 );
not ( n2264 , n2256 );
nand ( n2265 , n2264 , n2199 );
nand ( n2266 , n2263 , n2265 );
xnor ( n2267 , n2132 , n2266 );
not ( n2268 , n2077 );
and ( n2269 , n2086 , n2268 );
not ( n2270 , n2086 );
and ( n2271 , n2270 , n2077 );
nor ( n2272 , n2269 , n2271 );
not ( n2273 , n800 );
not ( n2274 , n2206 );
or ( n2275 , n2273 , n2274 );
not ( n2276 , n2207 );
not ( n2277 , n782 );
and ( n2278 , n48 , n2277 );
not ( n2279 , n48 );
and ( n2280 , n2279 , n782 );
nor ( n2281 , n2278 , n2280 );
nand ( n2282 , n2276 , n2281 );
nand ( n2283 , n2275 , n2282 );
not ( n2284 , n2283 );
not ( n2285 , n2284 );
not ( n2286 , n856 );
not ( n2287 , n2162 );
or ( n2288 , n2286 , n2287 );
not ( n2289 , n1491 );
and ( n2290 , n982 , n42 );
not ( n2291 , n982 );
not ( n2292 , n42 );
and ( n2293 , n2291 , n2292 );
nor ( n2294 , n2290 , n2293 );
not ( n2295 , n2294 );
nand ( n2296 , n2289 , n2295 );
nand ( n2297 , n2288 , n2296 );
not ( n2298 , n2297 );
not ( n2299 , n2298 );
or ( n2300 , n2285 , n2299 );
not ( n2301 , n2283 );
not ( n2302 , n2297 );
or ( n2303 , n2301 , n2302 );
buf ( n2304 , n704 );
not ( n2305 , n2304 );
not ( n2306 , n2179 );
or ( n2307 , n2305 , n2306 );
not ( n2308 , n710 );
not ( n2309 , n904 );
not ( n2310 , n2309 );
or ( n2311 , n2308 , n2310 );
not ( n2312 , n1129 );
not ( n2313 , n2312 );
or ( n2314 , n2313 , n2309 );
nand ( n2315 , n2311 , n2314 );
nand ( n2316 , n1095 , n2315 );
nand ( n2317 , n2307 , n2316 );
not ( n2318 , n2317 );
nand ( n2319 , n2303 , n2318 );
nand ( n2320 , n2300 , n2319 );
not ( n2321 , n2320 );
not ( n2322 , n2321 );
xor ( n2323 , n2210 , n2220 );
xor ( n2324 , n2323 , n2225 );
not ( n2325 , n2324 );
not ( n2326 , n2325 );
not ( n2327 , n2326 );
or ( n2328 , n2322 , n2327 );
not ( n2329 , n2320 );
not ( n2330 , n2325 );
or ( n2331 , n2329 , n2330 );
not ( n2332 , n746 );
not ( n2333 , n2332 );
not ( n2334 , n2147 );
or ( n2335 , n2333 , n2334 );
not ( n2336 , n46 );
buf ( n2337 , n660 );
not ( n2338 , n2337 );
or ( n2339 , n2336 , n2338 );
or ( n2340 , n46 , n2337 );
nand ( n2341 , n2339 , n2340 );
nand ( n2342 , n734 , n2341 );
nand ( n2343 , n2335 , n2342 );
not ( n2344 , n2343 );
not ( n2345 , n638 );
and ( n2346 , n40 , n1279 );
not ( n2347 , n40 );
and ( n2348 , n2347 , n721 );
nor ( n2349 , n2346 , n2348 );
not ( n2350 , n2349 );
or ( n2351 , n2345 , n2350 );
and ( n2352 , n40 , n1175 );
not ( n2353 , n40 );
and ( n2354 , n3 , n17 );
not ( n2355 , n3 );
and ( n2356 , n2355 , n33 );
or ( n2357 , n2354 , n2356 );
and ( n2358 , n2353 , n2357 );
or ( n2359 , n2352 , n2358 );
nand ( n2360 , n1253 , n2359 );
nand ( n2361 , n2351 , n2360 );
not ( n2362 , n2361 );
not ( n2363 , n1021 );
not ( n2364 , n38 );
not ( n2365 , n1184 );
or ( n2366 , n2364 , n2365 );
or ( n2367 , n1184 , n38 );
nand ( n2368 , n2366 , n2367 );
not ( n2369 , n2368 );
or ( n2370 , n2363 , n2369 );
not ( n2371 , n609 );
not ( n2372 , n1985 );
or ( n2373 , n2371 , n2372 );
or ( n2374 , n609 , n1221 );
nand ( n2375 , n2373 , n2374 );
nand ( n2376 , n572 , n2375 );
nand ( n2377 , n2370 , n2376 );
not ( n2378 , n2377 );
and ( n2379 , n2362 , n2378 );
not ( n2380 , n2362 );
and ( n2381 , n2380 , n2377 );
nor ( n2382 , n2379 , n2381 );
not ( n2383 , n2382 );
or ( n2384 , n2344 , n2383 );
not ( n2385 , n2362 );
nand ( n2386 , n2385 , n2377 );
nand ( n2387 , n2384 , n2386 );
nand ( n2388 , n2331 , n2387 );
nand ( n2389 , n2328 , n2388 );
not ( n2390 , n2389 );
xor ( n2391 , n2228 , n2250 );
not ( n2392 , n51 );
not ( n2393 , n2216 );
or ( n2394 , n2392 , n2393 );
not ( n2395 , n1935 );
not ( n2396 , n50 );
not ( n2397 , n1043 );
not ( n2398 , n2397 );
or ( n2399 , n2396 , n2398 );
not ( n2400 , n50 );
not ( n2401 , n7 );
nand ( n2402 , n3 , n2401 );
not ( n2403 , n3 );
not ( n2404 , n23 );
nand ( n2405 , n2403 , n2404 );
nand ( n2406 , n2400 , n2402 , n2405 );
nand ( n2407 , n2399 , n2406 );
nand ( n2408 , n2395 , n2407 );
nand ( n2409 , n2394 , n2408 );
nor ( n2410 , n39 , n40 );
not ( n2411 , n2410 );
not ( n2412 , n2411 );
buf ( n2413 , n1220 );
not ( n2414 , n2413 );
not ( n2415 , n2414 );
or ( n2416 , n2412 , n2415 );
nand ( n2417 , n39 , n40 );
and ( n2418 , n38 , n2417 );
nand ( n2419 , n2416 , n2418 );
not ( n2420 , n2419 );
nand ( n2421 , n2409 , n2420 );
not ( n2422 , n2421 );
not ( n2423 , n2422 );
not ( n2424 , n870 );
not ( n2425 , n2349 );
or ( n2426 , n2424 , n2425 );
nand ( n2427 , n638 , n1889 );
nand ( n2428 , n2426 , n2427 );
not ( n2429 , n2428 );
not ( n2430 , n1021 );
not ( n2431 , n2235 );
or ( n2432 , n2430 , n2431 );
not ( n2433 , n571 );
nand ( n2434 , n2433 , n2368 );
nand ( n2435 , n2432 , n2434 );
not ( n2436 , n2435 );
not ( n2437 , n2436 );
or ( n2438 , n2429 , n2437 );
not ( n2439 , n2435 );
or ( n2440 , n2428 , n2439 );
nand ( n2441 , n2438 , n2440 );
not ( n2442 , n2441 );
or ( n2443 , n2423 , n2442 );
not ( n2444 , n2439 );
nand ( n2445 , n2428 , n2444 );
nand ( n2446 , n2443 , n2445 );
not ( n2447 , n2446 );
xnor ( n2448 , n2391 , n2447 );
not ( n2449 , n2448 );
or ( n2450 , n2390 , n2449 );
not ( n2451 , n2228 );
nand ( n2452 , n2451 , n2250 );
not ( n2453 , n2452 );
nand ( n2454 , n2228 , n2249 );
not ( n2455 , n2454 );
or ( n2456 , n2453 , n2455 );
not ( n2457 , n2447 );
nand ( n2458 , n2456 , n2457 );
nand ( n2459 , n2450 , n2458 );
not ( n2460 , n2459 );
nand ( n2461 , n2272 , n2460 );
not ( n2462 , n2197 );
not ( n2463 , n2462 );
not ( n2464 , n2261 );
or ( n2465 , n2463 , n2464 );
nand ( n2466 , n2197 , n2260 );
nand ( n2467 , n2465 , n2466 );
and ( n2468 , n2461 , n2467 );
nor ( n2469 , n2272 , n2460 );
nor ( n2470 , n2468 , n2469 );
nand ( n2471 , n2267 , n2470 );
not ( n2472 , n2471 );
nor ( n2473 , n2120 , n2472 );
nor ( n2474 , n2267 , n2470 );
not ( n2475 , n2474 );
not ( n2476 , n2459 );
xor ( n2477 , n2272 , n2476 );
xnor ( n2478 , n2477 , n2467 );
not ( n2479 , n2389 );
xor ( n2480 , n2448 , n2479 );
not ( n2481 , n2480 );
not ( n2482 , n2481 );
xnor ( n2483 , n2192 , n2137 );
not ( n2484 , n2483 );
not ( n2485 , n1139 );
not ( n2486 , n1649 );
not ( n2487 , n970 );
or ( n2488 , n2486 , n2487 );
nand ( n2489 , n1134 , n973 );
nand ( n2490 , n2488 , n2489 );
not ( n2491 , n2490 );
or ( n2492 , n2485 , n2491 );
nand ( n2493 , n1325 , n2315 );
nand ( n2494 , n2492 , n2493 );
not ( n2495 , n2494 );
nand ( n2496 , n1022 , n2224 );
not ( n2497 , n2496 );
not ( n2498 , n806 );
not ( n2499 , n2498 );
not ( n2500 , n48 );
not ( n2501 , n1498 );
or ( n2502 , n2500 , n2501 );
or ( n2503 , n48 , n1498 );
nand ( n2504 , n2502 , n2503 );
not ( n2505 , n2504 );
or ( n2506 , n2499 , n2505 );
buf ( n2507 , n1017 );
nand ( n2508 , n2507 , n2281 );
nand ( n2509 , n2506 , n2508 );
not ( n2510 , n2509 );
or ( n2511 , n2497 , n2510 );
or ( n2512 , n2496 , n2509 );
nand ( n2513 , n2511 , n2512 );
not ( n2514 , n2513 );
or ( n2515 , n2495 , n2514 );
not ( n2516 , n2496 );
nand ( n2517 , n2516 , n2509 );
nand ( n2518 , n2515 , n2517 );
not ( n2519 , n2518 );
not ( n2520 , n2419 );
not ( n2521 , n2409 );
or ( n2522 , n2520 , n2521 );
or ( n2523 , n2419 , n2409 );
nand ( n2524 , n2522 , n2523 );
not ( n2525 , n2524 );
and ( n2526 , n51 , n2407 );
xor ( n2527 , n50 , n794 );
nor ( n2528 , n1936 , n2527 );
nor ( n2529 , n2526 , n2528 );
not ( n2530 , n2529 );
not ( n2531 , n2530 );
not ( n2532 , n776 );
not ( n2533 , n42 );
not ( n2534 , n2533 );
not ( n2535 , n722 );
or ( n2536 , n2534 , n2535 );
not ( n2537 , n721 );
not ( n2538 , n42 );
or ( n2539 , n2537 , n2538 );
nand ( n2540 , n2536 , n2539 );
and ( n2541 , n2532 , n2540 );
not ( n2542 , n1155 );
nor ( n2543 , n2542 , n2294 );
nor ( n2544 , n2541 , n2543 );
not ( n2545 , n2544 );
not ( n2546 , n2545 );
or ( n2547 , n2531 , n2546 );
not ( n2548 , n2529 );
not ( n2549 , n2544 );
or ( n2550 , n2548 , n2549 );
not ( n2551 , n1892 );
not ( n2552 , n2359 );
or ( n2553 , n2551 , n2552 );
not ( n2554 , n40 );
not ( n2555 , n1394 );
or ( n2556 , n2554 , n2555 );
or ( n2557 , n40 , n1394 );
nand ( n2558 , n2556 , n2557 );
nand ( n2559 , n674 , n2558 );
nand ( n2560 , n2553 , n2559 );
nand ( n2561 , n2550 , n2560 );
nand ( n2562 , n2547 , n2561 );
not ( n2563 , n2562 );
not ( n2564 , n2563 );
or ( n2565 , n2525 , n2564 );
not ( n2566 , n2562 );
or ( n2567 , n2524 , n2566 );
nand ( n2568 , n2565 , n2567 );
not ( n2569 , n2568 );
or ( n2570 , n2519 , n2569 );
not ( n2571 , n2566 );
nand ( n2572 , n2524 , n2571 );
nand ( n2573 , n2570 , n2572 );
not ( n2574 , n2573 );
not ( n2575 , n2441 );
not ( n2576 , n2421 );
and ( n2577 , n2575 , n2576 );
and ( n2578 , n2421 , n2441 );
nor ( n2579 , n2577 , n2578 );
and ( n2580 , n2167 , n2153 );
not ( n2581 , n2167 );
and ( n2582 , n2581 , n2154 );
nor ( n2583 , n2580 , n2582 );
and ( n2584 , n2583 , n2184 );
not ( n2585 , n2583 );
not ( n2586 , n2184 );
and ( n2587 , n2585 , n2586 );
nor ( n2588 , n2584 , n2587 );
xnor ( n2589 , n2579 , n2588 );
not ( n2590 , n2589 );
or ( n2591 , n2574 , n2590 );
not ( n2592 , n2579 );
nand ( n2593 , n2592 , n2588 );
nand ( n2594 , n2591 , n2593 );
not ( n2595 , n2594 );
or ( n2596 , n2484 , n2595 );
or ( n2597 , n2483 , n2594 );
nand ( n2598 , n2596 , n2597 );
not ( n2599 , n2598 );
or ( n2600 , n2482 , n2599 );
not ( n2601 , n2483 );
nand ( n2602 , n2601 , n2594 );
nand ( n2603 , n2600 , n2602 );
not ( n2604 , n2603 );
nor ( n2605 , n2478 , n2604 );
not ( n2606 , n2605 );
and ( n2607 , n2475 , n2606 );
not ( n2608 , n2266 );
not ( n2609 , n2125 );
not ( n2610 , n2609 );
not ( n2611 , n2130 );
not ( n2612 , n2611 );
or ( n2613 , n2610 , n2612 );
or ( n2614 , n2609 , n2611 );
nand ( n2615 , n2613 , n2614 );
not ( n2616 , n2615 );
or ( n2617 , n2608 , n2616 );
not ( n2618 , n2609 );
nand ( n2619 , n2618 , n2611 );
nand ( n2620 , n2617 , n2619 );
not ( n2621 , n2070 );
not ( n2622 , n2621 );
not ( n2623 , n2116 );
or ( n2624 , n2622 , n2623 );
not ( n2625 , n2070 );
or ( n2626 , n2625 , n2116 );
nand ( n2627 , n2624 , n2626 );
nor ( n2628 , n2620 , n2627 );
nor ( n2629 , n2607 , n2628 );
nand ( n2630 , n2473 , n2629 );
not ( n2631 , n2069 );
not ( n2632 , n2119 );
nand ( n2633 , n2631 , n2632 );
nand ( n2634 , n1867 , n2630 , n2633 );
not ( n2635 , n1470 );
not ( n2636 , n1624 );
nand ( n2637 , n2635 , n2636 );
not ( n2638 , n2637 );
not ( n2639 , n1435 );
xor ( n2640 , n1461 , n2639 );
xnor ( n2641 , n2640 , n1124 );
not ( n2642 , n2068 );
not ( n2643 , n1872 );
and ( n2644 , n2643 , n2061 );
not ( n2645 , n2643 );
and ( n2646 , n2645 , n2062 );
nor ( n2647 , n2644 , n2646 );
not ( n2648 , n2647 );
or ( n2649 , n2642 , n2648 );
nand ( n2650 , n2643 , n2061 );
nand ( n2651 , n2649 , n2650 );
not ( n2652 , n2651 );
nor ( n2653 , n2641 , n2652 );
not ( n2654 , n2653 );
or ( n2655 , n2638 , n2654 );
not ( n2656 , n2120 );
and ( n2657 , n2620 , n2627 );
nand ( n2658 , n2656 , n2657 );
nand ( n2659 , n2655 , n2658 );
or ( n2660 , n2634 , n2659 );
nand ( n2661 , n1629 , n1737 );
not ( n2662 , n2661 );
buf ( n2663 , n2662 );
not ( n2664 , n1865 );
not ( n2665 , n2664 );
nand ( n2666 , n2663 , n2665 );
nand ( n2667 , n2660 , n2666 );
not ( n2668 , n1625 );
nor ( n2669 , n2668 , n2664 );
not ( n2670 , n2669 );
nand ( n2671 , n2641 , n2652 );
not ( n2672 , n1470 );
not ( n2673 , n1624 );
nand ( n2674 , n2672 , n2673 );
nand ( n2675 , n2671 , n2674 );
not ( n2676 , n2675 );
or ( n2677 , n2670 , n2676 );
not ( n2678 , n1750 );
not ( n2679 , n1863 );
nor ( n2680 , n2678 , n2679 );
not ( n2681 , n2680 );
nand ( n2682 , n2677 , n2681 );
or ( n2683 , n2667 , n2682 );
not ( n2684 , n2471 );
not ( n2685 , n2478 );
not ( n2686 , n2604 );
nor ( n2687 , n2685 , n2686 );
nor ( n2688 , n2684 , n2687 );
not ( n2689 , n2628 );
nand ( n2690 , n2688 , n2689 , n2656 );
not ( n2691 , n2690 );
or ( n2692 , n41 , n42 );
not ( n2693 , n2692 );
not ( n2694 , n2413 );
not ( n2695 , n2694 );
or ( n2696 , n2693 , n2695 );
nand ( n2697 , n41 , n42 );
not ( n2698 , n2697 );
nor ( n2699 , n647 , n2698 );
nand ( n2700 , n2696 , n2699 );
not ( n2701 , n2700 );
not ( n2702 , n801 );
not ( n2703 , n2702 );
not ( n2704 , n2504 );
or ( n2705 , n2703 , n2704 );
and ( n2706 , n659 , n48 );
not ( n2707 , n659 );
not ( n2708 , n48 );
and ( n2709 , n2707 , n2708 );
nor ( n2710 , n2706 , n2709 );
nand ( n2711 , n2498 , n2710 );
nand ( n2712 , n2705 , n2711 );
not ( n2713 , n2712 );
or ( n2714 , n2701 , n2713 );
or ( n2715 , n2700 , n2712 );
nand ( n2716 , n2714 , n2715 );
not ( n2717 , n2716 );
not ( n2718 , n755 );
not ( n2719 , n2718 );
not ( n2720 , n763 );
not ( n2721 , n1027 );
not ( n2722 , n2721 );
or ( n2723 , n2720 , n2722 );
or ( n2724 , n1759 , n763 );
nand ( n2725 , n2723 , n2724 );
and ( n2726 , n2719 , n2725 );
and ( n2727 , n1061 , n46 );
not ( n2728 , n1061 );
and ( n2729 , n2728 , n763 );
nor ( n2730 , n2727 , n2729 );
nor ( n2731 , n761 , n2730 );
nor ( n2732 , n2726 , n2731 );
not ( n2733 , n2732 );
not ( n2734 , n871 );
not ( n2735 , n2413 );
and ( n2736 , n2735 , n40 );
not ( n2737 , n2735 );
and ( n2738 , n2737 , n647 );
nor ( n2739 , n2736 , n2738 );
not ( n2740 , n2739 );
or ( n2741 , n2734 , n2740 );
not ( n2742 , n886 );
nand ( n2743 , n2742 , n2558 );
nand ( n2744 , n2741 , n2743 );
and ( n2745 , n2733 , n2744 );
not ( n2746 , n2733 );
not ( n2747 , n2744 );
and ( n2748 , n2746 , n2747 );
nor ( n2749 , n2745 , n2748 );
not ( n2750 , n2749 );
not ( n2751 , n2750 );
or ( n2752 , n2717 , n2751 );
not ( n2753 , n2716 );
nand ( n2754 , n2753 , n2749 );
nand ( n2755 , n2752 , n2754 );
not ( n2756 , n51 );
not ( n2757 , n646 );
not ( n2758 , n2757 );
not ( n2759 , n1406 );
and ( n2760 , n2758 , n2759 );
not ( n2761 , n646 );
and ( n2762 , n2761 , n1406 );
nor ( n2763 , n2760 , n2762 );
not ( n2764 , n2763 );
or ( n2765 , n2756 , n2764 );
not ( n2766 , n1936 );
buf ( n2767 , n2766 );
not ( n2768 , n50 );
not ( n2769 , n2337 );
not ( n2770 , n2769 );
not ( n2771 , n2770 );
or ( n2772 , n2768 , n2771 );
or ( n2773 , n50 , n2770 );
nand ( n2774 , n2772 , n2773 );
nand ( n2775 , n2767 , n2774 );
nand ( n2776 , n2765 , n2775 );
not ( n2777 , n2776 );
not ( n2778 , n2182 );
not ( n2779 , n1107 );
not ( n2780 , n723 );
or ( n2781 , n2779 , n2780 );
nand ( n2782 , n1528 , n2537 );
nand ( n2783 , n2781 , n2782 );
not ( n2784 , n2783 );
or ( n2785 , n2778 , n2784 );
not ( n2786 , n1107 );
not ( n2787 , n845 );
or ( n2788 , n2786 , n2787 );
not ( n2789 , n845 );
not ( n2790 , n2789 );
or ( n2791 , n1130 , n2790 );
nand ( n2792 , n2788 , n2791 );
nand ( n2793 , n1139 , n2792 );
nand ( n2794 , n2785 , n2793 );
buf ( n2795 , n1903 );
not ( n2796 , n2795 );
and ( n2797 , n42 , n1394 );
not ( n2798 , n42 );
and ( n2799 , n2798 , n1395 );
nor ( n2800 , n2797 , n2799 );
not ( n2801 , n2800 );
not ( n2802 , n2801 );
or ( n2803 , n2796 , n2802 );
not ( n2804 , n42 );
not ( n2805 , n2223 );
or ( n2806 , n2804 , n2805 );
or ( n2807 , n42 , n2223 );
nand ( n2808 , n2806 , n2807 );
nand ( n2809 , n2289 , n2808 );
nand ( n2810 , n2803 , n2809 );
and ( n2811 , n2794 , n2810 );
not ( n2812 , n2794 );
not ( n2813 , n2810 );
and ( n2814 , n2812 , n2813 );
nor ( n2815 , n2811 , n2814 );
not ( n2816 , n2815 );
or ( n2817 , n2777 , n2816 );
not ( n2818 , n2813 );
nand ( n2819 , n2818 , n2794 );
nand ( n2820 , n2817 , n2819 );
not ( n2821 , n2820 );
nor ( n2822 , n43 , n677 );
not ( n2823 , n2822 );
not ( n2824 , n2823 );
not ( n2825 , n2224 );
or ( n2826 , n2824 , n2825 );
nand ( n2827 , n43 , n1129 );
and ( n2828 , n42 , n2827 );
nand ( n2829 , n2826 , n2828 );
not ( n2830 , n2829 );
not ( n2831 , n2830 );
not ( n2832 , n2702 );
xnor ( n2833 , n48 , n1152 );
not ( n2834 , n2833 );
or ( n2835 , n2832 , n2834 );
not ( n2836 , n807 );
not ( n2837 , n48 );
not ( n2838 , n1061 );
or ( n2839 , n2837 , n2838 );
or ( n2840 , n48 , n1061 );
nand ( n2841 , n2839 , n2840 );
nand ( n2842 , n2836 , n2841 );
nand ( n2843 , n2835 , n2842 );
not ( n2844 , n2843 );
nor ( n2845 , n2831 , n2844 );
not ( n2846 , n2845 );
and ( n2847 , n637 , n2222 );
not ( n2848 , n999 );
not ( n2849 , n2833 );
or ( n2850 , n2848 , n2849 );
nand ( n2851 , n800 , n2710 );
nand ( n2852 , n2850 , n2851 );
not ( n2853 , n2852 );
xor ( n2854 , n2847 , n2853 );
not ( n2855 , n1139 );
not ( n2856 , n2783 );
or ( n2857 , n2855 , n2856 );
not ( n2858 , n1107 );
not ( n2859 , n984 );
or ( n2860 , n2858 , n2859 );
or ( n2861 , n1130 , n984 );
nand ( n2862 , n2860 , n2861 );
nand ( n2863 , n1100 , n2862 );
nand ( n2864 , n2857 , n2863 );
xnor ( n2865 , n2854 , n2864 );
not ( n2866 , n2865 );
not ( n2867 , n2866 );
or ( n2868 , n2846 , n2867 );
not ( n2869 , n2845 );
nand ( n2870 , n2869 , n2865 );
nand ( n2871 , n2868 , n2870 );
not ( n2872 , n2871 );
or ( n2873 , n2821 , n2872 );
nand ( n2874 , n2845 , n2865 );
nand ( n2875 , n2873 , n2874 );
not ( n2876 , n2875 );
xor ( n2877 , n2755 , n2876 );
not ( n2878 , n1903 );
not ( n2879 , n42 );
not ( n2880 , n845 );
or ( n2881 , n2879 , n2880 );
or ( n2882 , n845 , n42 );
nand ( n2883 , n2881 , n2882 );
not ( n2884 , n2883 );
nor ( n2885 , n2878 , n2884 );
nor ( n2886 , n1491 , n2800 );
nor ( n2887 , n2885 , n2886 );
not ( n2888 , n2887 );
not ( n2889 , n2888 );
and ( n2890 , n46 , n969 );
not ( n2891 , n46 );
not ( n2892 , n969 );
and ( n2893 , n2891 , n2892 );
nor ( n2894 , n2890 , n2893 );
nor ( n2895 , n761 , n2894 );
nor ( n2896 , n2730 , n756 );
nor ( n2897 , n2895 , n2896 );
not ( n2898 , n2897 );
not ( n2899 , n2898 );
or ( n2900 , n2889 , n2899 );
not ( n2901 , n2887 );
not ( n2902 , n2897 );
or ( n2903 , n2901 , n2902 );
not ( n2904 , n1937 );
not ( n2905 , n2904 );
not ( n2906 , n2905 );
not ( n2907 , n2763 );
or ( n2908 , n2906 , n2907 );
not ( n2909 , n50 );
not ( n2910 , n1079 );
or ( n2911 , n2909 , n2910 );
not ( n2912 , n50 );
and ( n2913 , n3 , n9 );
not ( n2914 , n3 );
and ( n2915 , n2914 , n25 );
or ( n2916 , n2913 , n2915 );
nand ( n2917 , n2912 , n2916 );
nand ( n2918 , n2911 , n2917 );
nand ( n2919 , n51 , n2918 );
nand ( n2920 , n2908 , n2919 );
nand ( n2921 , n2903 , n2920 );
nand ( n2922 , n2900 , n2921 );
not ( n2923 , n2922 );
not ( n2924 , n2864 );
not ( n2925 , n2853 );
and ( n2926 , n2847 , n2925 );
not ( n2927 , n2847 );
and ( n2928 , n2927 , n2853 );
nor ( n2929 , n2926 , n2928 );
not ( n2930 , n2929 );
or ( n2931 , n2924 , n2930 );
not ( n2932 , n2853 );
nand ( n2933 , n2847 , n2932 );
nand ( n2934 , n2931 , n2933 );
not ( n2935 , n2934 );
xor ( n2936 , n2923 , n2935 );
not ( n2937 , n1937 );
not ( n2938 , n2918 );
or ( n2939 , n2937 , n2938 );
not ( n2940 , n2527 );
nand ( n2941 , n51 , n2940 );
nand ( n2942 , n2939 , n2941 );
not ( n2943 , n2942 );
not ( n2944 , n2943 );
not ( n2945 , n856 );
not ( n2946 , n2540 );
or ( n2947 , n2945 , n2946 );
nand ( n2948 , n1051 , n2883 );
nand ( n2949 , n2947 , n2948 );
not ( n2950 , n2949 );
or ( n2951 , n2944 , n2950 );
not ( n2952 , n2942 );
or ( n2953 , n2952 , n2949 );
nand ( n2954 , n2951 , n2953 );
not ( n2955 , n1325 );
not ( n2956 , n2490 );
or ( n2957 , n2955 , n2956 );
nand ( n2958 , n1139 , n2862 );
nand ( n2959 , n2957 , n2958 );
and ( n2960 , n2954 , n2959 );
not ( n2961 , n2954 );
not ( n2962 , n2959 );
and ( n2963 , n2961 , n2962 );
nor ( n2964 , n2960 , n2963 );
xnor ( n2965 , n2936 , n2964 );
xnor ( n2966 , n2877 , n2965 );
not ( n2967 , n2820 );
and ( n2968 , n2871 , n2967 );
not ( n2969 , n2871 );
and ( n2970 , n2969 , n2820 );
nor ( n2971 , n2968 , n2970 );
not ( n2972 , n2971 );
xor ( n2973 , n2920 , n2888 );
xor ( n2974 , n2973 , n2898 );
not ( n2975 , n2767 );
not ( n2976 , n1406 );
not ( n2977 , n1759 );
or ( n2978 , n2976 , n2977 );
nand ( n2979 , n3 , n12 );
not ( n2980 , n3 );
nand ( n2981 , n2980 , n28 );
nand ( n2982 , n50 , n2979 , n2981 );
nand ( n2983 , n2978 , n2982 );
not ( n2984 , n2983 );
or ( n2985 , n2975 , n2984 );
nand ( n2986 , n51 , n2774 );
nand ( n2987 , n2985 , n2986 );
not ( n2988 , n2987 );
and ( n2989 , n2795 , n2224 );
not ( n2990 , n2989 );
not ( n2991 , n1100 );
not ( n2992 , n2792 );
or ( n2993 , n2991 , n2992 );
not ( n2994 , n2313 );
not ( n2995 , n1394 );
or ( n2996 , n2994 , n2995 );
or ( n2997 , n1107 , n1394 );
nand ( n2998 , n2996 , n2997 );
nand ( n2999 , n1139 , n2998 );
nand ( n3000 , n2993 , n2999 );
not ( n3001 , n3000 );
not ( n3002 , n3001 );
or ( n3003 , n2990 , n3002 );
not ( n3004 , n2694 );
nor ( n3005 , n2878 , n3004 );
not ( n3006 , n3005 );
nand ( n3007 , n3006 , n3000 );
nand ( n3008 , n3003 , n3007 );
not ( n3009 , n3008 );
or ( n3010 , n2988 , n3009 );
nand ( n3011 , n2989 , n3000 );
nand ( n3012 , n3010 , n3011 );
not ( n3013 , n3012 );
not ( n3014 , n2718 );
buf ( n3015 , n3014 );
not ( n3016 , n3015 );
not ( n3017 , n2894 );
not ( n3018 , n3017 );
or ( n3019 , n3016 , n3018 );
not ( n3020 , n46 );
not ( n3021 , n987 );
or ( n3022 , n3020 , n3021 );
or ( n3023 , n46 , n987 );
nand ( n3024 , n3022 , n3023 );
nand ( n3025 , n762 , n3024 );
nand ( n3026 , n3019 , n3025 );
not ( n3027 , n3026 );
not ( n3028 , n3027 );
not ( n3029 , n2830 );
not ( n3030 , n2843 );
not ( n3031 , n3030 );
and ( n3032 , n3029 , n3031 );
and ( n3033 , n2830 , n2844 );
nor ( n3034 , n3032 , n3033 );
not ( n3035 , n3034 );
not ( n3036 , n3035 );
or ( n3037 , n3028 , n3036 );
nand ( n3038 , n3026 , n3034 );
nand ( n3039 , n3037 , n3038 );
not ( n3040 , n3039 );
or ( n3041 , n3013 , n3040 );
nand ( n3042 , n3026 , n3035 );
nand ( n3043 , n3041 , n3042 );
xor ( n3044 , n2974 , n3043 );
and ( n3045 , n2972 , n3044 );
and ( n3046 , n2974 , n3043 );
nor ( n3047 , n3045 , n3046 );
nand ( n3048 , n2966 , n3047 );
not ( n3049 , n3047 );
not ( n3050 , n3049 );
not ( n3051 , n2966 );
not ( n3052 , n3051 );
or ( n3053 , n3050 , n3052 );
not ( n3054 , n3012 );
and ( n3055 , n3039 , n3054 );
not ( n3056 , n3039 );
and ( n3057 , n3056 , n3012 );
nor ( n3058 , n3055 , n3057 );
not ( n3059 , n3058 );
not ( n3060 , n3059 );
nand ( n3061 , n45 , n46 );
not ( n3062 , n3061 );
not ( n3063 , n2222 );
not ( n3064 , n3063 );
or ( n3065 , n3062 , n3064 );
nor ( n3066 , n45 , n46 );
not ( n3067 , n3066 );
nand ( n3068 , n3065 , n3067 );
and ( n3069 , n1650 , n3068 );
not ( n3070 , n51 );
not ( n3071 , n2983 );
or ( n3072 , n3070 , n3071 );
not ( n3073 , n50 );
not ( n3074 , n2309 );
or ( n3075 , n3073 , n3074 );
or ( n3076 , n50 , n903 );
nand ( n3077 , n3075 , n3076 );
nand ( n3078 , n2767 , n3077 );
nand ( n3079 , n3072 , n3078 );
and ( n3080 , n3069 , n3079 );
not ( n3081 , n3080 );
not ( n3082 , n807 );
not ( n3083 , n3082 );
not ( n3084 , n48 );
not ( n3085 , n969 );
or ( n3086 , n3084 , n3085 );
not ( n3087 , n48 );
not ( n3088 , n969 );
nand ( n3089 , n3087 , n3088 );
nand ( n3090 , n3086 , n3089 );
not ( n3091 , n3090 );
or ( n3092 , n3083 , n3091 );
not ( n3093 , n800 );
not ( n3094 , n3093 );
nand ( n3095 , n3094 , n2841 );
nand ( n3096 , n3092 , n3095 );
not ( n3097 , n3096 );
not ( n3098 , n734 );
not ( n3099 , n46 );
buf ( n3100 , n721 );
not ( n3101 , n3100 );
or ( n3102 , n3099 , n3101 );
nand ( n3103 , n763 , n2537 );
nand ( n3104 , n3102 , n3103 );
not ( n3105 , n3104 );
or ( n3106 , n3098 , n3105 );
nand ( n3107 , n3014 , n3024 );
nand ( n3108 , n3106 , n3107 );
not ( n3109 , n3108 );
not ( n3110 , n3109 );
or ( n3111 , n3097 , n3110 );
not ( n3112 , n3108 );
or ( n3113 , n3096 , n3112 );
nand ( n3114 , n3111 , n3113 );
not ( n3115 , n3114 );
or ( n3116 , n3081 , n3115 );
not ( n3117 , n3112 );
nand ( n3118 , n3096 , n3117 );
nand ( n3119 , n3116 , n3118 );
not ( n3120 , n3119 );
not ( n3121 , n3120 );
not ( n3122 , n2776 );
and ( n3123 , n2815 , n3122 );
not ( n3124 , n2815 );
and ( n3125 , n3124 , n2776 );
nor ( n3126 , n3123 , n3125 );
not ( n3127 , n3126 );
not ( n3128 , n3127 );
or ( n3129 , n3121 , n3128 );
nand ( n3130 , n3119 , n3126 );
nand ( n3131 , n3129 , n3130 );
not ( n3132 , n3131 );
or ( n3133 , n3060 , n3132 );
not ( n3134 , n3120 );
not ( n3135 , n3126 );
nand ( n3136 , n3134 , n3135 );
nand ( n3137 , n3133 , n3136 );
not ( n3138 , n2971 );
not ( n3139 , n3044 );
or ( n3140 , n3138 , n3139 );
or ( n3141 , n2971 , n3044 );
nand ( n3142 , n3140 , n3141 );
nand ( n3143 , n3137 , n3142 );
nand ( n3144 , n3053 , n3143 );
nand ( n3145 , n3048 , n3144 );
not ( n3146 , n3063 );
nand ( n3147 , n3146 , n2304 );
not ( n3148 , n3147 );
not ( n3149 , n51 );
not ( n3150 , n3077 );
or ( n3151 , n3149 , n3150 );
not ( n3152 , n50 );
not ( n3153 , n969 );
or ( n3154 , n3152 , n3153 );
or ( n3155 , n50 , n969 );
nand ( n3156 , n3154 , n3155 );
nand ( n3157 , n2766 , n3156 );
nand ( n3158 , n3151 , n3157 );
nor ( n3159 , n3148 , n3158 );
not ( n3160 , n801 );
not ( n3161 , n3160 );
not ( n3162 , n48 );
not ( n3163 , n987 );
or ( n3164 , n3162 , n3163 );
or ( n3165 , n48 , n987 );
nand ( n3166 , n3164 , n3165 );
not ( n3167 , n3166 );
or ( n3168 , n3161 , n3167 );
not ( n3169 , n48 );
and ( n3170 , n723 , n3169 );
not ( n3171 , n723 );
and ( n3172 , n3171 , n48 );
nor ( n3173 , n3170 , n3172 );
nand ( n3174 , n3082 , n3173 );
nand ( n3175 , n3168 , n3174 );
not ( n3176 , n3175 );
or ( n3177 , n3159 , n3176 );
not ( n3178 , n3147 );
nand ( n3179 , n3178 , n3158 );
nand ( n3180 , n3177 , n3179 );
not ( n3181 , n3180 );
xor ( n3182 , n3069 , n3079 );
and ( n3183 , n3181 , n3182 );
not ( n3184 , n3181 );
not ( n3185 , n3182 );
and ( n3186 , n3184 , n3185 );
nor ( n3187 , n3183 , n3186 );
not ( n3188 , n3187 );
buf ( n3189 , n705 );
not ( n3190 , n3189 );
not ( n3191 , n2998 );
or ( n3192 , n3190 , n3191 );
not ( n3193 , n1528 );
not ( n3194 , n1917 );
or ( n3195 , n3193 , n3194 );
not ( n3196 , n2413 );
or ( n3197 , n1649 , n3196 );
nand ( n3198 , n3195 , n3197 );
nand ( n3199 , n1095 , n3198 );
nand ( n3200 , n3192 , n3199 );
not ( n3201 , n747 );
not ( n3202 , n3104 );
or ( n3203 , n3201 , n3202 );
xnor ( n3204 , n46 , n845 );
nand ( n3205 , n734 , n3204 );
nand ( n3206 , n3203 , n3205 );
and ( n3207 , n3200 , n3206 );
not ( n3208 , n3200 );
not ( n3209 , n3206 );
and ( n3210 , n3208 , n3209 );
nor ( n3211 , n3207 , n3210 );
not ( n3212 , n3094 );
not ( n3213 , n3090 );
or ( n3214 , n3212 , n3213 );
not ( n3215 , n806 );
not ( n3216 , n3215 );
not ( n3217 , n3216 );
nand ( n3218 , n3217 , n3166 );
nand ( n3219 , n3214 , n3218 );
and ( n3220 , n3211 , n3219 );
not ( n3221 , n3211 );
not ( n3222 , n3219 );
and ( n3223 , n3221 , n3222 );
nor ( n3224 , n3220 , n3223 );
and ( n3225 , n3188 , n3224 );
nor ( n3226 , n3185 , n3181 );
nor ( n3227 , n3225 , n3226 );
not ( n3228 , n3227 );
xor ( n3229 , n3114 , n3080 );
not ( n3230 , n3229 );
not ( n3231 , n3219 );
not ( n3232 , n3211 );
or ( n3233 , n3231 , n3232 );
not ( n3234 , n3209 );
nand ( n3235 , n3234 , n3200 );
nand ( n3236 , n3233 , n3235 );
not ( n3237 , n3236 );
and ( n3238 , n3008 , n2987 );
not ( n3239 , n3008 );
not ( n3240 , n2987 );
and ( n3241 , n3239 , n3240 );
nor ( n3242 , n3238 , n3241 );
and ( n3243 , n3237 , n3242 );
not ( n3244 , n3237 );
not ( n3245 , n3242 );
and ( n3246 , n3244 , n3245 );
nor ( n3247 , n3243 , n3246 );
not ( n3248 , n3247 );
or ( n3249 , n3230 , n3248 );
or ( n3250 , n3229 , n3247 );
nand ( n3251 , n3249 , n3250 );
nand ( n3252 , n3228 , n3251 );
not ( n3253 , n3252 );
not ( n3254 , n3229 );
not ( n3255 , n3247 );
not ( n3256 , n3255 );
or ( n3257 , n3254 , n3256 );
nand ( n3258 , n3242 , n3236 );
nand ( n3259 , n3257 , n3258 );
not ( n3260 , n3058 );
not ( n3261 , n3131 );
or ( n3262 , n3260 , n3261 );
or ( n3263 , n3058 , n3131 );
nand ( n3264 , n3262 , n3263 );
nand ( n3265 , n3259 , n3264 );
not ( n3266 , n3265 );
or ( n3267 , n3253 , n3266 );
not ( n3268 , n3264 );
not ( n3269 , n3259 );
nand ( n3270 , n3268 , n3269 );
nand ( n3271 , n3267 , n3270 );
not ( n3272 , n3271 );
nor ( n3273 , n3137 , n3142 );
not ( n3274 , n3273 );
nand ( n3275 , n3272 , n3274 , n3048 );
nand ( n3276 , n47 , n48 );
and ( n3277 , n3276 , n3063 );
nor ( n3278 , n47 , n48 );
not ( n3279 , n3278 );
not ( n3280 , n3279 );
nor ( n3281 , n3277 , n3280 );
nor ( n3282 , n763 , n3281 );
not ( n3283 , n2766 );
not ( n3284 , n50 );
not ( n3285 , n987 );
or ( n3286 , n3284 , n3285 );
or ( n3287 , n50 , n987 );
nand ( n3288 , n3286 , n3287 );
not ( n3289 , n3288 );
or ( n3290 , n3283 , n3289 );
nand ( n3291 , n51 , n3156 );
nand ( n3292 , n3290 , n3291 );
xnor ( n3293 , n3282 , n3292 );
not ( n3294 , n3293 );
not ( n3295 , n3294 );
not ( n3296 , n3093 );
not ( n3297 , n3296 );
not ( n3298 , n3173 );
or ( n3299 , n3297 , n3298 );
not ( n3300 , n3216 );
not ( n3301 , n48 );
not ( n3302 , n3301 );
not ( n3303 , n2789 );
or ( n3304 , n3302 , n3303 );
not ( n3305 , n48 );
or ( n3306 , n3305 , n2789 );
nand ( n3307 , n3304 , n3306 );
nand ( n3308 , n3300 , n3307 );
nand ( n3309 , n3299 , n3308 );
not ( n3310 , n3309 );
not ( n3311 , n3310 );
not ( n3312 , n2718 );
not ( n3313 , n763 );
not ( n3314 , n1394 );
not ( n3315 , n3314 );
or ( n3316 , n3313 , n3315 );
not ( n3317 , n1394 );
or ( n3318 , n763 , n3317 );
nand ( n3319 , n3316 , n3318 );
and ( n3320 , n3312 , n3319 );
not ( n3321 , n763 );
not ( n3322 , n1917 );
and ( n3323 , n3321 , n3322 );
and ( n3324 , n763 , n2694 );
nor ( n3325 , n3323 , n3324 );
nor ( n3326 , n761 , n3325 );
nor ( n3327 , n3320 , n3326 );
not ( n3328 , n3327 );
not ( n3329 , n3328 );
or ( n3330 , n3311 , n3329 );
nand ( n3331 , n3309 , n3327 );
nand ( n3332 , n3330 , n3331 );
not ( n3333 , n3332 );
or ( n3334 , n3295 , n3333 );
nand ( n3335 , n3309 , n3328 );
nand ( n3336 , n3334 , n3335 );
xor ( n3337 , n3147 , n3158 );
xnor ( n3338 , n3337 , n3175 );
and ( n3339 , n3282 , n3292 );
not ( n3340 , n762 );
not ( n3341 , n3319 );
or ( n3342 , n3340 , n3341 );
nand ( n3343 , n757 , n3204 );
nand ( n3344 , n3342 , n3343 );
not ( n3345 , n3344 );
and ( n3346 , n3339 , n3345 );
not ( n3347 , n3339 );
and ( n3348 , n3347 , n3344 );
nor ( n3349 , n3346 , n3348 );
not ( n3350 , n3349 );
and ( n3351 , n3338 , n3350 );
not ( n3352 , n3338 );
and ( n3353 , n3352 , n3349 );
nor ( n3354 , n3351 , n3353 );
nor ( n3355 , n3336 , n3354 );
not ( n3356 , n3187 );
not ( n3357 , n3356 );
not ( n3358 , n3224 );
not ( n3359 , n3358 );
or ( n3360 , n3357 , n3359 );
nand ( n3361 , n3187 , n3224 );
nand ( n3362 , n3360 , n3361 );
not ( n3363 , n3350 );
not ( n3364 , n3338 );
or ( n3365 , n3363 , n3364 );
nand ( n3366 , n3339 , n3344 );
nand ( n3367 , n3365 , n3366 );
nor ( n3368 , n3362 , n3367 );
nor ( n3369 , n3355 , n3368 );
not ( n3370 , n3369 );
and ( n3371 , n51 , n3288 );
not ( n3372 , n2905 );
not ( n3373 , n1406 );
not ( n3374 , n3100 );
not ( n3375 , n3374 );
or ( n3376 , n3373 , n3375 );
not ( n3377 , n3100 );
or ( n3378 , n1406 , n3377 );
nand ( n3379 , n3376 , n3378 );
not ( n3380 , n3379 );
nor ( n3381 , n3372 , n3380 );
nor ( n3382 , n3371 , n3381 );
not ( n3383 , n3382 );
not ( n3384 , n3004 );
nand ( n3385 , n2719 , n3384 );
not ( n3386 , n3385 );
not ( n3387 , n2702 );
not ( n3388 , n3307 );
or ( n3389 , n3387 , n3388 );
not ( n3390 , n807 );
not ( n3391 , n48 );
not ( n3392 , n3391 );
not ( n3393 , n1394 );
not ( n3394 , n3393 );
or ( n3395 , n3392 , n3394 );
not ( n3396 , n48 );
or ( n3397 , n3396 , n1395 );
nand ( n3398 , n3395 , n3397 );
nand ( n3399 , n3390 , n3398 );
nand ( n3400 , n3389 , n3399 );
not ( n3401 , n3400 );
and ( n3402 , n3386 , n3401 );
and ( n3403 , n3385 , n3400 );
nor ( n3404 , n3402 , n3403 );
not ( n3405 , n3404 );
and ( n3406 , n3383 , n3405 );
not ( n3407 , n3400 );
nor ( n3408 , n3385 , n3407 );
nor ( n3409 , n3406 , n3408 );
not ( n3410 , n3409 );
not ( n3411 , n3293 );
not ( n3412 , n3332 );
or ( n3413 , n3411 , n3412 );
or ( n3414 , n3293 , n3332 );
nand ( n3415 , n3413 , n3414 );
nand ( n3416 , n3410 , n3415 );
not ( n3417 , n3336 );
not ( n3418 , n3417 );
nand ( n3419 , n3418 , n3354 );
not ( n3420 , n3415 );
nand ( n3421 , n3420 , n3409 );
not ( n3422 , n50 );
not ( n3423 , n3317 );
not ( n3424 , n3423 );
or ( n3425 , n3422 , n3424 );
not ( n3426 , n3004 );
not ( n3427 , n3426 );
nand ( n3428 , n3425 , n3427 );
not ( n3429 , n3094 );
nand ( n3430 , n3429 , n3426 );
not ( n3431 , n51 );
not ( n3432 , n1406 );
not ( n3433 , n846 );
or ( n3434 , n3432 , n3433 );
or ( n3435 , n1406 , n846 );
nand ( n3436 , n3434 , n3435 );
not ( n3437 , n3436 );
or ( n3438 , n3431 , n3437 );
nand ( n3439 , n2767 , n3423 );
nand ( n3440 , n3438 , n3439 );
and ( n3441 , n3428 , n3430 , n3440 );
not ( n3442 , n3217 );
and ( n3443 , n48 , n3004 );
not ( n3444 , n48 );
and ( n3445 , n3444 , n3426 );
nor ( n3446 , n3443 , n3445 );
or ( n3447 , n3442 , n3446 );
not ( n3448 , n3398 );
or ( n3449 , n3429 , n3448 );
nand ( n3450 , n3447 , n3449 );
not ( n3451 , n3450 );
not ( n3452 , n51 );
not ( n3453 , n3379 );
or ( n3454 , n3452 , n3453 );
not ( n3455 , n2904 );
nand ( n3456 , n3455 , n3436 );
nand ( n3457 , n3454 , n3456 );
not ( n3458 , n3457 );
nand ( n3459 , n49 , n50 );
not ( n3460 , n3459 );
not ( n3461 , n3063 );
or ( n3462 , n3460 , n3461 );
not ( n3463 , n994 );
nand ( n3464 , n3462 , n3463 );
nand ( n3465 , n48 , n3464 );
not ( n3466 , n3465 );
and ( n3467 , n3458 , n3466 );
and ( n3468 , n3465 , n3457 );
nor ( n3469 , n3467 , n3468 );
nand ( n3470 , n3451 , n3469 );
and ( n3471 , n3441 , n3470 );
not ( n3472 , n3450 );
nor ( n3473 , n3472 , n3469 );
nor ( n3474 , n3471 , n3473 );
not ( n3475 , n3465 );
and ( n3476 , n3475 , n3457 );
not ( n3477 , n3382 );
not ( n3478 , n3404 );
not ( n3479 , n3478 );
or ( n3480 , n3477 , n3479 );
not ( n3481 , n3382 );
nand ( n3482 , n3481 , n3404 );
nand ( n3483 , n3480 , n3482 );
nor ( n3484 , n3476 , n3483 );
or ( n3485 , n3474 , n3484 );
nand ( n3486 , n3476 , n3483 );
nand ( n3487 , n3485 , n3486 );
nand ( n3488 , n3421 , n3487 );
nand ( n3489 , n3416 , n3419 , n3488 );
not ( n3490 , n3489 );
or ( n3491 , n3370 , n3490 );
not ( n3492 , n3367 );
not ( n3493 , n3492 );
nand ( n3494 , n3493 , n3362 );
nand ( n3495 , n3491 , n3494 );
not ( n3496 , n3495 );
not ( n3497 , n3268 );
not ( n3498 , n3269 );
or ( n3499 , n3497 , n3498 );
not ( n3500 , n3251 );
nand ( n3501 , n3500 , n3227 );
nand ( n3502 , n3499 , n3501 );
nor ( n3503 , n3496 , n3502 );
nand ( n3504 , n3503 , n3274 , n3048 );
nand ( n3505 , n3145 , n3275 , n3504 );
not ( n3506 , n3505 );
not ( n3507 , n762 );
not ( n3508 , n2725 );
or ( n3509 , n3507 , n3508 );
nand ( n3510 , n3015 , n2341 );
nand ( n3511 , n3509 , n3510 );
not ( n3512 , n3511 );
not ( n3513 , n3512 );
not ( n3514 , n3513 );
not ( n3515 , n2700 );
and ( n3516 , n3515 , n2712 );
not ( n3517 , n3516 );
or ( n3518 , n3514 , n3517 );
and ( n3519 , n3516 , n3511 );
not ( n3520 , n3516 );
and ( n3521 , n3520 , n3512 );
nor ( n3522 , n3519 , n3521 );
not ( n3523 , n2959 );
not ( n3524 , n2954 );
or ( n3525 , n3523 , n3524 );
not ( n3526 , n2952 );
nand ( n3527 , n3526 , n2949 );
nand ( n3528 , n3525 , n3527 );
nand ( n3529 , n3522 , n3528 );
nand ( n3530 , n3518 , n3529 );
xor ( n3531 , n2343 , n2382 );
xor ( n3532 , n2283 , n2317 );
xor ( n3533 , n3532 , n2298 );
xnor ( n3534 , n3531 , n3533 );
xor ( n3535 , n3530 , n3534 );
not ( n3536 , n3535 );
xor ( n3537 , n2545 , n2560 );
not ( n3538 , n2530 );
xnor ( n3539 , n3537 , n3538 );
not ( n3540 , n3539 );
nand ( n3541 , n2747 , n2732 );
and ( n3542 , n3541 , n2716 );
nor ( n3543 , n2747 , n2732 );
nor ( n3544 , n3542 , n3543 );
not ( n3545 , n3544 );
not ( n3546 , n3545 );
not ( n3547 , n2494 );
not ( n3548 , n3547 );
not ( n3549 , n2513 );
or ( n3550 , n3548 , n3549 );
or ( n3551 , n3547 , n2513 );
nand ( n3552 , n3550 , n3551 );
not ( n3553 , n3552 );
not ( n3554 , n3553 );
or ( n3555 , n3546 , n3554 );
nand ( n3556 , n3544 , n3552 );
nand ( n3557 , n3555 , n3556 );
not ( n3558 , n3557 );
or ( n3559 , n3540 , n3558 );
nand ( n3560 , n3545 , n3552 );
nand ( n3561 , n3559 , n3560 );
xor ( n3562 , n2518 , n2568 );
and ( n3563 , n3561 , n3562 );
not ( n3564 , n3561 );
not ( n3565 , n3562 );
and ( n3566 , n3564 , n3565 );
nor ( n3567 , n3563 , n3566 );
not ( n3568 , n3567 );
or ( n3569 , n3536 , n3568 );
not ( n3570 , n3565 );
not ( n3571 , n3561 );
not ( n3572 , n3571 );
nand ( n3573 , n3570 , n3572 );
nand ( n3574 , n3569 , n3573 );
not ( n3575 , n3574 );
not ( n3576 , n2387 );
not ( n3577 , n2324 );
or ( n3578 , n3576 , n3577 );
or ( n3579 , n2324 , n2387 );
nand ( n3580 , n3578 , n3579 );
and ( n3581 , n3580 , n2320 );
not ( n3582 , n3580 );
and ( n3583 , n3582 , n2321 );
nor ( n3584 , n3581 , n3583 );
not ( n3585 , n3584 );
not ( n3586 , n3585 );
not ( n3587 , n3530 );
not ( n3588 , n3534 );
or ( n3589 , n3587 , n3588 );
not ( n3590 , n3533 );
nand ( n3591 , n3531 , n3590 );
nand ( n3592 , n3589 , n3591 );
not ( n3593 , n3592 );
or ( n3594 , n3586 , n3593 );
not ( n3595 , n3584 );
or ( n3596 , n3595 , n3592 );
nand ( n3597 , n3594 , n3596 );
not ( n3598 , n3597 );
xor ( n3599 , n2589 , n2573 );
not ( n3600 , n3599 );
not ( n3601 , n3600 );
and ( n3602 , n3598 , n3601 );
not ( n3603 , n3599 );
and ( n3604 , n3603 , n3597 );
nor ( n3605 , n3602 , n3604 );
nand ( n3606 , n3575 , n3605 );
not ( n3607 , n3599 );
not ( n3608 , n3597 );
or ( n3609 , n3607 , n3608 );
not ( n3610 , n3595 );
nand ( n3611 , n3610 , n3592 );
nand ( n3612 , n3609 , n3611 );
not ( n3613 , n3612 );
not ( n3614 , n2598 );
not ( n3615 , n2480 );
and ( n3616 , n3614 , n3615 );
and ( n3617 , n2480 , n2598 );
nor ( n3618 , n3616 , n3617 );
nand ( n3619 , n3613 , n3618 );
nand ( n3620 , n3606 , n3619 );
not ( n3621 , n2964 );
and ( n3622 , n2934 , n2922 );
not ( n3623 , n2934 );
and ( n3624 , n3623 , n2923 );
nor ( n3625 , n3622 , n3624 );
not ( n3626 , n3625 );
or ( n3627 , n3621 , n3626 );
nand ( n3628 , n2922 , n2934 );
nand ( n3629 , n3627 , n3628 );
not ( n3630 , n3528 );
and ( n3631 , n3522 , n3630 );
not ( n3632 , n3522 );
and ( n3633 , n3632 , n3528 );
nor ( n3634 , n3631 , n3633 );
not ( n3635 , n3539 );
and ( n3636 , n3557 , n3635 );
not ( n3637 , n3557 );
and ( n3638 , n3637 , n3539 );
nor ( n3639 , n3636 , n3638 );
nand ( n3640 , n3634 , n3639 );
and ( n3641 , n3629 , n3640 );
nor ( n3642 , n3634 , n3639 );
nor ( n3643 , n3641 , n3642 );
not ( n3644 , n3643 );
not ( n3645 , n3644 );
not ( n3646 , n3645 );
xor ( n3647 , n3562 , n3571 );
xnor ( n3648 , n3647 , n3535 );
not ( n3649 , n3648 );
not ( n3650 , n3649 );
or ( n3651 , n3646 , n3650 );
not ( n3652 , n3639 );
not ( n3653 , n3629 );
not ( n3654 , n3634 );
or ( n3655 , n3653 , n3654 );
or ( n3656 , n3634 , n3629 );
nand ( n3657 , n3655 , n3656 );
nor ( n3658 , n3652 , n3657 );
not ( n3659 , n3658 );
nand ( n3660 , n3652 , n3657 );
nand ( n3661 , n3659 , n3660 );
not ( n3662 , n2965 );
not ( n3663 , n3662 );
not ( n3664 , n2876 );
and ( n3665 , n2755 , n3664 );
not ( n3666 , n2755 );
not ( n3667 , n3664 );
and ( n3668 , n3666 , n3667 );
nor ( n3669 , n3665 , n3668 );
not ( n3670 , n3669 );
or ( n3671 , n3663 , n3670 );
not ( n3672 , n3667 );
nand ( n3673 , n2755 , n3672 );
nand ( n3674 , n3671 , n3673 );
not ( n3675 , n3674 );
nand ( n3676 , n3661 , n3675 );
nand ( n3677 , n3651 , n3676 );
nor ( n3678 , n3620 , n3677 );
not ( n3679 , n3678 );
or ( n3680 , n3506 , n3679 );
not ( n3681 , n3620 );
not ( n3682 , n3658 );
nand ( n3683 , n3660 , n3682 , n3674 );
nand ( n3684 , n3644 , n3648 );
and ( n3685 , n3683 , n3684 );
not ( n3686 , n3643 );
nor ( n3687 , n3686 , n3648 );
nor ( n3688 , n3685 , n3687 );
and ( n3689 , n3681 , n3688 );
not ( n3690 , n3619 );
not ( n3691 , n3605 );
not ( n3692 , n3575 );
nand ( n3693 , n3691 , n3692 );
or ( n3694 , n3690 , n3693 );
not ( n3695 , n3613 );
not ( n3696 , n3618 );
nand ( n3697 , n3695 , n3696 );
nand ( n3698 , n3694 , n3697 );
nor ( n3699 , n3689 , n3698 );
nand ( n3700 , n3680 , n3699 );
nor ( n3701 , n2662 , n2680 );
not ( n3702 , n2675 );
nand ( n3703 , n2691 , n3700 , n3701 , n3702 );
nand ( n3704 , n2683 , n3703 );
buf ( n3705 , n3704 );
and ( n3706 , n497 , n605 );
not ( n3707 , n497 );
not ( n3708 , n604 );
not ( n3709 , n3708 );
and ( n3710 , n3707 , n3709 );
nor ( n3711 , n3706 , n3710 );
or ( n3712 , n493 , n3711 );
not ( n3713 , n481 );
or ( n3714 , n594 , n3713 );
nand ( n3715 , n3712 , n3714 );
xor ( n3716 , n40 , n505 );
not ( n3717 , n3716 );
not ( n3718 , n1515 );
or ( n3719 , n3717 , n3718 );
or ( n3720 , n647 , n1707 );
nand ( n3721 , n3719 , n3720 );
and ( n3722 , n3715 , n3721 );
not ( n3723 , n3715 );
not ( n3724 , n3721 );
and ( n3725 , n3723 , n3724 );
nor ( n3726 , n3722 , n3725 );
not ( n3727 , n607 );
not ( n3728 , n38 );
not ( n3729 , n556 );
or ( n3730 , n3728 , n3729 );
not ( n3731 , n556 );
nand ( n3732 , n609 , n3731 );
nand ( n3733 , n3730 , n3732 );
not ( n3734 , n3733 );
or ( n3735 , n3727 , n3734 );
and ( n3736 , n38 , n519 );
not ( n3737 , n516 );
not ( n3738 , n3737 );
not ( n3739 , n3738 );
and ( n3740 , n609 , n3739 );
nor ( n3741 , n3736 , n3740 );
or ( n3742 , n3741 , n564 );
nand ( n3743 , n3735 , n3742 );
not ( n3744 , n481 );
not ( n3745 , n3711 );
not ( n3746 , n3745 );
or ( n3747 , n3744 , n3746 );
xor ( n3748 , n36 , n795 );
nand ( n3749 , n492 , n3748 );
nand ( n3750 , n3747 , n3749 );
not ( n3751 , n1080 );
not ( n3752 , n3751 );
not ( n3753 , n3752 );
and ( n3754 , n36 , n3753 );
and ( n3755 , n3750 , n3754 );
not ( n3756 , n3750 );
not ( n3757 , n3754 );
and ( n3758 , n3756 , n3757 );
nor ( n3759 , n3755 , n3758 );
and ( n3760 , n3743 , n3759 );
and ( n3761 , n3754 , n3750 );
nor ( n3762 , n3760 , n3761 );
not ( n3763 , n3762 );
and ( n3764 , n3726 , n3763 );
and ( n3765 , n3721 , n3715 );
nor ( n3766 , n3764 , n3765 );
or ( n3767 , n608 , n3741 );
or ( n3768 , n615 , n613 );
nand ( n3769 , n3767 , n3768 );
not ( n3770 , n1707 );
not ( n3771 , n1514 );
or ( n3772 , n3770 , n3771 );
nand ( n3773 , n3772 , n40 );
not ( n3774 , n1820 );
and ( n3775 , n36 , n3774 );
xor ( n3776 , n3773 , n3775 );
and ( n3777 , n3769 , n3776 );
and ( n3778 , n3775 , n3773 );
nor ( n3779 , n3777 , n3778 );
xor ( n3780 , n3766 , n3779 );
xnor ( n3781 , n598 , n622 );
xor ( n3782 , n3780 , n3781 );
and ( n3783 , n3726 , n3762 );
not ( n3784 , n3726 );
and ( n3785 , n3784 , n3763 );
nor ( n3786 , n3783 , n3785 );
buf ( n3787 , n3786 );
not ( n3788 , n3787 );
xnor ( n3789 , n3776 , n3769 );
and ( n3790 , n3759 , n3743 );
not ( n3791 , n3759 );
not ( n3792 , n3743 );
and ( n3793 , n3791 , n3792 );
nor ( n3794 , n3790 , n3793 );
not ( n3795 , n3794 );
and ( n3796 , n1708 , n3716 );
not ( n3797 , n517 );
not ( n3798 , n647 );
and ( n3799 , n3797 , n3798 );
and ( n3800 , n647 , n3737 );
nor ( n3801 , n3799 , n3800 );
nor ( n3802 , n1514 , n3801 );
nor ( n3803 , n3796 , n3802 );
not ( n3804 , n3803 );
not ( n3805 , n3804 );
not ( n3806 , n2878 );
not ( n3807 , n1491 );
or ( n3808 , n3806 , n3807 );
nand ( n3809 , n3808 , n42 );
not ( n3810 , n490 );
not ( n3811 , n36 );
not ( n3812 , n1080 );
or ( n3813 , n3811 , n3812 );
or ( n3814 , n36 , n1080 );
nand ( n3815 , n3813 , n3814 );
not ( n3816 , n3815 );
or ( n3817 , n3810 , n3816 );
nand ( n3818 , n478 , n3748 );
nand ( n3819 , n3817 , n3818 );
xor ( n3820 , n3809 , n3819 );
not ( n3821 , n3820 );
or ( n3822 , n3805 , n3821 );
not ( n3823 , n3809 );
not ( n3824 , n3823 );
nand ( n3825 , n3824 , n3819 );
nand ( n3826 , n3822 , n3825 );
and ( n3827 , n3826 , n3721 );
not ( n3828 , n3826 );
and ( n3829 , n3828 , n3724 );
or ( n3830 , n3827 , n3829 );
not ( n3831 , n3830 );
or ( n3832 , n3795 , n3831 );
nand ( n3833 , n3724 , n3826 );
nand ( n3834 , n3832 , n3833 );
xnor ( n3835 , n3789 , n3834 );
and ( n3836 , n3788 , n3835 );
not ( n3837 , n3789 );
and ( n3838 , n3837 , n3834 );
nor ( n3839 , n3836 , n3838 );
nand ( n3840 , n3782 , n3839 );
xor ( n3841 , n3766 , n3779 );
and ( n3842 , n3841 , n3781 );
and ( n3843 , n3766 , n3779 );
or ( n3844 , n3842 , n3843 );
xnor ( n3845 , n630 , n625 );
nand ( n3846 , n3844 , n3845 );
not ( n3847 , n492 );
not ( n3848 , n1753 );
or ( n3849 , n3847 , n3848 );
nand ( n3850 , n481 , n3815 );
nand ( n3851 , n3849 , n3850 );
not ( n3852 , n3851 );
not ( n3853 , n1665 );
nand ( n3854 , n36 , n3853 );
not ( n3855 , n3854 );
not ( n3856 , n1690 );
not ( n3857 , n1810 );
or ( n3858 , n3856 , n3857 );
nand ( n3859 , n1694 , n42 );
nand ( n3860 , n3858 , n3859 );
not ( n3861 , n3860 );
or ( n3862 , n3855 , n3861 );
or ( n3863 , n3854 , n3860 );
nand ( n3864 , n3862 , n3863 );
not ( n3865 , n3864 );
or ( n3866 , n3852 , n3865 );
not ( n3867 , n3854 );
nand ( n3868 , n3867 , n3860 );
nand ( n3869 , n3866 , n3868 );
not ( n3870 , n3869 );
not ( n3871 , n3870 );
not ( n3872 , n3820 );
not ( n3873 , n3803 );
and ( n3874 , n3872 , n3873 );
and ( n3875 , n3803 , n3820 );
nor ( n3876 , n3874 , n3875 );
not ( n3877 , n3876 );
and ( n3878 , n3871 , n3877 );
not ( n3879 , n3869 );
not ( n3880 , n3876 );
nand ( n3881 , n3879 , n3880 );
not ( n3882 , n3881 );
not ( n3883 , n3876 );
nor ( n3884 , n3883 , n3870 );
nor ( n3885 , n3882 , n3884 );
not ( n3886 , n3885 );
not ( n3887 , n38 );
not ( n3888 , n3709 );
or ( n3889 , n3887 , n3888 );
or ( n3890 , n38 , n3709 );
nand ( n3891 , n3889 , n3890 );
not ( n3892 , n3891 );
or ( n3893 , n608 , n3892 );
not ( n3894 , n3733 );
or ( n3895 , n615 , n3894 );
nand ( n3896 , n3893 , n3895 );
not ( n3897 , n3896 );
buf ( n3898 , n1499 );
not ( n3899 , n3898 );
nand ( n3900 , n3899 , n36 );
not ( n3901 , n1515 );
not ( n3902 , n1770 );
or ( n3903 , n3901 , n3902 );
not ( n3904 , n3801 );
nand ( n3905 , n1519 , n3904 );
nand ( n3906 , n3903 , n3905 );
nand ( n3907 , n3900 , n3906 );
not ( n3908 , n3907 );
not ( n3909 , n3900 );
not ( n3910 , n3906 );
and ( n3911 , n3909 , n3910 );
nor ( n3912 , n3908 , n3911 );
not ( n3913 , n3912 );
or ( n3914 , n3897 , n3913 );
or ( n3915 , n3896 , n3912 );
nand ( n3916 , n3914 , n3915 );
and ( n3917 , n3886 , n3916 );
nor ( n3918 , n3878 , n3917 );
not ( n3919 , n3900 );
not ( n3920 , n3910 );
not ( n3921 , n3920 );
not ( n3922 , n3921 );
and ( n3923 , n3919 , n3922 );
not ( n3924 , n3912 );
and ( n3925 , n3896 , n3924 );
nor ( n3926 , n3923 , n3925 );
not ( n3927 , n3794 );
and ( n3928 , n3830 , n3927 );
not ( n3929 , n3830 );
and ( n3930 , n3929 , n3794 );
nor ( n3931 , n3928 , n3930 );
not ( n3932 , n3931 );
and ( n3933 , n3926 , n3932 );
not ( n3934 , n3926 );
and ( n3935 , n3934 , n3931 );
nor ( n3936 , n3933 , n3935 );
xnor ( n3937 , n3918 , n3936 );
not ( n3938 , n1829 );
and ( n3939 , n3938 , n1815 );
and ( n3940 , n1803 , n1814 );
nor ( n3941 , n3939 , n3940 );
not ( n3942 , n3941 );
xor ( n3943 , n3851 , n3864 );
not ( n3944 , n3943 );
and ( n3945 , n3942 , n3944 );
and ( n3946 , n3941 , n3943 );
nor ( n3947 , n3945 , n3946 );
not ( n3948 , n3947 );
not ( n3949 , n3948 );
not ( n3950 , n563 );
not ( n3951 , n3891 );
or ( n3952 , n3950 , n3951 );
nand ( n3953 , n575 , n1824 );
nand ( n3954 , n3952 , n3953 );
and ( n3955 , n3954 , n3920 );
not ( n3956 , n3954 );
and ( n3957 , n3956 , n3910 );
or ( n3958 , n3955 , n3957 );
not ( n3959 , n1757 );
not ( n3960 , n3959 );
not ( n3961 , n1780 );
or ( n3962 , n3960 , n3961 );
nand ( n3963 , n1778 , n1774 );
nand ( n3964 , n3962 , n3963 );
xor ( n3965 , n3958 , n3964 );
not ( n3966 , n3965 );
or ( n3967 , n3949 , n3966 );
not ( n3968 , n3941 );
nand ( n3969 , n3968 , n3943 );
nand ( n3970 , n3967 , n3969 );
not ( n3971 , n3970 );
not ( n3972 , n3916 );
not ( n3973 , n3885 );
or ( n3974 , n3972 , n3973 );
or ( n3975 , n3916 , n3885 );
nand ( n3976 , n3974 , n3975 );
not ( n3977 , n3976 );
and ( n3978 , n3921 , n3954 );
and ( n3979 , n3958 , n3964 );
nor ( n3980 , n3978 , n3979 );
not ( n3981 , n3980 );
and ( n3982 , n3977 , n3981 );
and ( n3983 , n3980 , n3976 );
nor ( n3984 , n3982 , n3983 );
not ( n3985 , n3984 );
not ( n3986 , n3985 );
or ( n3987 , n3971 , n3986 );
not ( n3988 , n3980 );
nand ( n3989 , n3988 , n3976 );
nand ( n3990 , n3987 , n3989 );
not ( n3991 , n3990 );
nand ( n3992 , n3937 , n3991 );
not ( n3993 , n3786 );
not ( n3994 , n3835 );
or ( n3995 , n3993 , n3994 );
or ( n3996 , n3787 , n3835 );
nand ( n3997 , n3995 , n3996 );
not ( n3998 , n3997 );
or ( n3999 , n3918 , n3936 );
or ( n4000 , n3926 , n3931 );
nand ( n4001 , n3999 , n4000 );
not ( n4002 , n4001 );
nand ( n4003 , n3998 , n4002 );
not ( n4004 , n3970 );
not ( n4005 , n3984 );
or ( n4006 , n4004 , n4005 );
or ( n4007 , n3970 , n3984 );
nand ( n4008 , n4006 , n4007 );
not ( n4009 , n1835 );
not ( n4010 , n1793 );
not ( n4011 , n4010 );
or ( n4012 , n4009 , n4011 );
not ( n4013 , n1797 );
nand ( n4014 , n4013 , n1831 );
nand ( n4015 , n4012 , n4014 );
not ( n4016 , n4015 );
not ( n4017 , n1784 );
and ( n4018 , n4017 , n1792 );
and ( n4019 , n1785 , n1791 );
nor ( n4020 , n4018 , n4019 );
not ( n4021 , n4020 );
not ( n4022 , n3965 );
not ( n4023 , n3947 );
or ( n4024 , n4022 , n4023 );
or ( n4025 , n3965 , n3947 );
nand ( n4026 , n4024 , n4025 );
not ( n4027 , n4026 );
or ( n4028 , n4021 , n4027 );
or ( n4029 , n4020 , n4026 );
nand ( n4030 , n4028 , n4029 );
not ( n4031 , n4030 );
or ( n4032 , n4016 , n4031 );
not ( n4033 , n4020 );
nand ( n4034 , n4033 , n4026 );
nand ( n4035 , n4032 , n4034 );
nor ( n4036 , n4008 , n4035 );
xor ( n4037 , n4015 , n4030 );
not ( n4038 , n1858 );
not ( n4039 , n1851 );
or ( n4040 , n4038 , n4039 );
not ( n4041 , n1849 );
nand ( n4042 , n4041 , n1839 );
nand ( n4043 , n4040 , n4042 );
nor ( n4044 , n4037 , n4043 );
nor ( n4045 , n4036 , n4044 );
nand ( n4046 , n3992 , n4003 , n4045 );
or ( n4047 , n3782 , n3839 );
nand ( n4048 , n4001 , n3997 );
not ( n4049 , n3992 );
nand ( n4050 , n4037 , n4043 );
or ( n4051 , n4050 , n4036 );
nand ( n4052 , n4035 , n4008 );
nand ( n4053 , n4051 , n4052 );
not ( n4054 , n4053 );
or ( n4055 , n4049 , n4054 );
not ( n4056 , n3937 );
nand ( n4057 , n4056 , n3990 );
nand ( n4058 , n4055 , n4057 );
nand ( n4059 , n4058 , n4003 );
nor ( n4060 , n3844 , n3845 );
not ( n4061 , t_0 );
or ( n4062 , n635 , n4061 );
not ( n4063 , n633 );
nand ( n4064 , n588 , n4063 );
nand ( n4065 , n4062 , n4064 );
not ( n4066 , n4065 );
or ( n4067 , n587 , n4066 );
or ( n4068 , n586 , n4065 );
nand ( n4069 , n4067 , n4068 );
not ( n4070 , n4069 );
or ( n4071 , n475 , n4070 );
nand ( n4072 , n36 , n53 );
not ( n4073 , n4072 );
nand ( n4074 , n36 , n52 );
not ( n4075 , n4074 );
not ( n4076 , n476 );
nand ( n4077 , n36 , n37 );
buf ( n4078 , n4077 );
nor ( n4079 , n36 , n37 );
not ( n4080 , n4079 );
nand ( n4081 , n4076 , n4078 , n4080 );
not ( n4082 , n4081 );
not ( n4083 , n4082 );
not ( n4084 , n4083 );
buf ( n4085 , n4084 );
not ( n4086 , n4085 );
not ( n4087 , n4086 );
or ( n4088 , n483 , n4087 );
nand ( n4089 , n4088 , n36 );
not ( n4090 , n4089 );
or ( n4091 , n4075 , n4090 );
or ( n4092 , n4074 , n4089 );
nand ( n4093 , n4091 , n4092 );
not ( n4094 , n4093 );
and ( n4095 , n4073 , n4094 );
and ( n4096 , n4072 , n4093 );
nor ( n4097 , n4095 , n4096 );
not ( n4098 , n4097 );
or ( n4099 , n36 , n52 );
nand ( n4100 , n4099 , n4074 );
or ( n4101 , n4100 , n4086 );
nand ( n4102 , n4101 , n538 );
xor ( n4103 , n4102 , n4072 );
nand ( n4104 , n38 , n577 );
not ( n4105 , n53 );
and ( n4106 , n36 , n4105 );
and ( n4107 , n53 , n497 );
nor ( n4108 , n4106 , n4107 );
or ( n4109 , n4108 , n4086 );
or ( n4110 , n482 , n4100 );
nand ( n4111 , n4109 , n4110 );
nand ( n4112 , n36 , n54 );
not ( n4113 , n4112 );
xor ( n4114 , n4111 , n4113 );
and ( n4115 , n4104 , n4114 );
and ( n4116 , n4113 , n4111 );
nor ( n4117 , n4115 , n4116 );
not ( n4118 , n4117 );
and ( n4119 , n4103 , n4118 );
and ( n4120 , n4072 , n4102 );
nor ( n4121 , n4119 , n4120 );
not ( n4122 , n4121 );
or ( n4123 , n4098 , n4122 );
or ( n4124 , n4097 , n4121 );
nand ( n4125 , n4123 , n4124 );
not ( n4126 , n4125 );
not ( n4127 , n4126 );
nand ( n4128 , n36 , n55 );
nor ( n4129 , n36 , n55 );
not ( n4130 , n4129 );
nand ( n4131 , n4128 , n4130 );
not ( n4132 , n4085 );
or ( n4133 , n4131 , n4132 );
not ( n4134 , n480 );
or ( n4135 , n36 , n54 );
nand ( n4136 , n4135 , n4112 );
or ( n4137 , n4134 , n4136 );
nand ( n4138 , n4133 , n4137 );
not ( n4139 , n4138 );
not ( n4140 , n40 );
not ( n4141 , n52 );
and ( n4142 , n4140 , n4141 );
and ( n4143 , n40 , n52 );
nor ( n4144 , n4142 , n4143 );
not ( n4145 , n4144 );
not ( n4146 , n40 );
not ( n4147 , n41 );
or ( n4148 , n4146 , n4147 );
nor ( n4149 , n40 , n41 );
nor ( n4150 , n4149 , n636 );
nand ( n4151 , n4148 , n4150 );
not ( n4152 , n4151 );
buf ( n4153 , n4152 );
not ( n4154 , n4153 );
not ( n4155 , n4154 );
not ( n4156 , n4155 );
or ( n4157 , n4145 , n4156 );
nand ( n4158 , n40 , n1519 );
nand ( n4159 , n4157 , n4158 );
not ( n4160 , n4159 );
nand ( n4161 , n4139 , n4160 );
not ( n4162 , n38 );
not ( n4163 , n54 );
and ( n4164 , n4162 , n4163 );
and ( n4165 , n38 , n54 );
nor ( n4166 , n4164 , n4165 );
and ( n4167 , n4166 , n575 );
not ( n4168 , n38 );
not ( n4169 , n53 );
and ( n4170 , n4168 , n4169 );
and ( n4171 , n38 , n53 );
nor ( n4172 , n4170 , n4171 );
and ( n4173 , n1819 , n4172 );
nor ( n4174 , n4167 , n4173 );
not ( n4175 , n4174 );
not ( n4176 , n4175 );
nand ( n4177 , n36 , n57 );
not ( n4178 , n4177 );
and ( n4179 , n36 , n56 );
not ( n4180 , n36 );
not ( n4181 , n56 );
and ( n4182 , n4180 , n4181 );
nor ( n4183 , n4179 , n4182 );
not ( n4184 , n4183 );
not ( n4185 , n4084 );
or ( n4186 , n4184 , n4185 );
not ( n4187 , n4131 );
nand ( n4188 , n4187 , n1472 );
nand ( n4189 , n4186 , n4188 );
not ( n4190 , n4189 );
or ( n4191 , n4178 , n4190 );
or ( n4192 , n4177 , n4189 );
nand ( n4193 , n4191 , n4192 );
not ( n4194 , n4193 );
or ( n4195 , n4176 , n4194 );
not ( n4196 , n4177 );
nand ( n4197 , n4196 , n4189 );
nand ( n4198 , n4195 , n4197 );
and ( n4199 , n4161 , n4198 );
and ( n4200 , n4159 , n4138 );
nor ( n4201 , n4199 , n4200 );
not ( n4202 , n1708 );
not ( n4203 , n4155 );
and ( n4204 , n4202 , n4203 );
nor ( n4205 , n4204 , n647 );
nand ( n4206 , n36 , n56 );
xor ( n4207 , n4205 , n4206 );
and ( n4208 , n4172 , n607 );
not ( n4209 , n52 );
and ( n4210 , n609 , n4209 );
and ( n4211 , n38 , n52 );
nor ( n4212 , n4210 , n4211 );
and ( n4213 , n563 , n4212 );
nor ( n4214 , n4208 , n4213 );
and ( n4215 , n4207 , n4214 );
and ( n4216 , n4205 , n4206 );
or ( n4217 , n4215 , n4216 );
xor ( n4218 , n4201 , n4217 );
or ( n4219 , n4136 , n4086 );
or ( n4220 , n482 , n4108 );
nand ( n4221 , n4219 , n4220 );
and ( n4222 , n4221 , n4128 );
not ( n4223 , n4221 );
not ( n4224 , n4128 );
and ( n4225 , n4223 , n4224 );
nor ( n4226 , n4222 , n4225 );
and ( n4227 , n607 , n4212 );
and ( n4228 , n38 , n1819 );
nor ( n4229 , n4227 , n4228 );
and ( n4230 , n4226 , n4229 );
not ( n4231 , n4226 );
not ( n4232 , n4229 );
and ( n4233 , n4231 , n4232 );
nor ( n4234 , n4230 , n4233 );
and ( n4235 , n4218 , n4234 );
and ( n4236 , n4201 , n4217 );
or ( n4237 , n4235 , n4236 );
or ( n4238 , n4128 , n4232 );
or ( n4239 , n4224 , n4229 );
nand ( n4240 , n4239 , n4221 );
nand ( n4241 , n4238 , n4240 );
and ( n4242 , n4241 , n4232 );
not ( n4243 , n4241 );
and ( n4244 , n4243 , n4229 );
nor ( n4245 , n4242 , n4244 );
xor ( n4246 , n4114 , n4104 );
xnor ( n4247 , n4245 , n4246 );
nor ( n4248 , n4237 , n4247 );
not ( n4249 , n4248 );
or ( n4250 , n67 , n2698 );
nand ( n4251 , n4250 , n2692 );
and ( n4252 , n40 , n4251 );
xor ( n4253 , n48 , n59 );
not ( n4254 , n4253 );
not ( n4255 , n3217 );
or ( n4256 , n4254 , n4255 );
xor ( n4257 , n48 , n58 );
nand ( n4258 , n3094 , n4257 );
nand ( n4259 , n4256 , n4258 );
nand ( n4260 , n4252 , n4259 );
not ( n4261 , n4260 );
xnor ( n4262 , n46 , n60 );
not ( n4263 , n46 );
nand ( n4264 , n4263 , n48 , n47 );
not ( n4265 , n48 );
not ( n4266 , n47 );
nand ( n4267 , n4265 , n4266 , n46 );
nand ( n4268 , n4264 , n4267 );
buf ( n4269 , n4268 );
not ( n4270 , n4269 );
not ( n4271 , n4270 );
not ( n4272 , n4271 );
or ( n4273 , n4262 , n4272 );
not ( n4274 , n3015 );
xnor ( n4275 , n46 , n59 );
or ( n4276 , n4274 , n4275 );
nand ( n4277 , n4273 , n4276 );
nand ( n4278 , n4261 , n4277 );
not ( n4279 , n4277 );
buf ( n4280 , n4260 );
nand ( n4281 , n4279 , n4280 );
not ( n4282 , n51 );
xor ( n4283 , n50 , n56 );
not ( n4284 , n4283 );
or ( n4285 , n4282 , n4284 );
not ( n4286 , n51 );
nand ( n4287 , n50 , n4286 );
not ( n4288 , n4287 );
xor ( n4289 , n50 , n57 );
nand ( n4290 , n4288 , n4289 );
nand ( n4291 , n4285 , n4290 );
not ( n4292 , n677 );
nand ( n4293 , n4292 , n63 );
not ( n4294 , n63 );
nand ( n4295 , n4294 , n698 );
nand ( n4296 , n4293 , n4295 );
not ( n4297 , n44 );
nand ( n4298 , n4297 , n46 , n45 );
not ( n4299 , n46 );
not ( n4300 , n45 );
nand ( n4301 , n4299 , n44 , n4300 );
nand ( n4302 , n4298 , n4301 );
buf ( n4303 , n4302 );
buf ( n4304 , n4303 );
and ( n4305 , n4296 , n4304 );
xor ( n4306 , n62 , n1107 );
and ( n4307 , n1100 , n4306 );
nor ( n4308 , n4305 , n4307 );
not ( n4309 , n4308 );
nand ( n4310 , n4291 , n4309 );
xnor ( n4311 , n42 , n65 );
not ( n4312 , n4311 );
not ( n4313 , n4312 );
not ( n4314 , n1491 );
not ( n4315 , n4314 );
or ( n4316 , n4313 , n4315 );
not ( n4317 , n2878 );
xor ( n4318 , n42 , n64 );
nand ( n4319 , n4317 , n4318 );
nand ( n4320 , n4316 , n4319 );
not ( n4321 , n4291 );
nand ( n4322 , n4321 , n4308 );
nand ( n4323 , n4320 , n4322 );
nand ( n4324 , n4310 , n4323 );
nand ( n4325 , n4281 , n4324 );
nand ( n4326 , n4278 , n4325 );
not ( n4327 , n4326 );
xor ( n4328 , n42 , n63 );
not ( n4329 , n4328 );
not ( n4330 , n4314 );
or ( n4331 , n4329 , n4330 );
xor ( n4332 , n42 , n62 );
nand ( n4333 , n1694 , n4332 );
nand ( n4334 , n4331 , n4333 );
not ( n4335 , n4334 );
not ( n4336 , n4335 );
and ( n4337 , n61 , n2312 );
not ( n4338 , n61 );
and ( n4339 , n4338 , n1107 );
or ( n4340 , n4337 , n4339 );
not ( n4341 , n4340 );
buf ( n4342 , n4303 );
not ( n4343 , n4342 );
or ( n4344 , n4341 , n4343 );
xor ( n4345 , n1129 , n60 );
nand ( n4346 , n1100 , n4345 );
nand ( n4347 , n4344 , n4346 );
not ( n4348 , n4347 );
not ( n4349 , n4348 );
xor ( n4350 , n48 , n57 );
not ( n4351 , n4350 );
not ( n4352 , n3082 );
or ( n4353 , n4351 , n4352 );
xor ( n4354 , n48 , n56 );
nand ( n4355 , n3160 , n4354 );
nand ( n4356 , n4353 , n4355 );
not ( n4357 , n4356 );
or ( n4358 , n4349 , n4357 );
or ( n4359 , n4348 , n4356 );
nand ( n4360 , n4358 , n4359 );
not ( n4361 , n4360 );
or ( n4362 , n4336 , n4361 );
or ( n4363 , n4335 , n4360 );
nand ( n4364 , n4362 , n4363 );
xor ( n4365 , n38 , n66 );
not ( n4366 , n4365 );
or ( n4367 , n561 , n4366 );
nand ( n4368 , n38 , n67 );
or ( n4369 , n38 , n67 );
nand ( n4370 , n4368 , n4369 , n1506 );
nand ( n4371 , n4367 , n4370 );
not ( n4372 , n4371 );
not ( n4373 , n4372 );
not ( n4374 , n4275 );
not ( n4375 , n4374 );
not ( n4376 , n4271 );
or ( n4377 , n4375 , n4376 );
xor ( n4378 , n46 , n58 );
not ( n4379 , n4378 );
not ( n4380 , n4379 );
nand ( n4381 , n4380 , n2332 );
nand ( n4382 , n4377 , n4381 );
xor ( n4383 , n40 , n65 );
not ( n4384 , n4383 );
not ( n4385 , n4153 );
or ( n4386 , n4384 , n4385 );
xor ( n4387 , n40 , n64 );
nand ( n4388 , n1074 , n4387 );
nand ( n4389 , n4386 , n4388 );
xor ( n4390 , n4382 , n4389 );
not ( n4391 , n4390 );
or ( n4392 , n4373 , n4391 );
or ( n4393 , n4372 , n4390 );
nand ( n4394 , n4392 , n4393 );
xor ( n4395 , n4364 , n4394 );
not ( n4396 , n4395 );
or ( n4397 , n4327 , n4396 );
nand ( n4398 , n4364 , n4394 );
nand ( n4399 , n4397 , n4398 );
not ( n4400 , n4399 );
not ( n4401 , n67 );
nand ( n4402 , n4401 , n2417 );
nand ( n4403 , n2411 , n4402 );
nand ( n4404 , n38 , n4403 );
not ( n4405 , n4404 );
not ( n4406 , n4405 );
not ( n4407 , n51 );
xor ( n4408 , n50 , n54 );
not ( n4409 , n4408 );
or ( n4410 , n4407 , n4409 );
not ( n4411 , n51 );
xor ( n4412 , n50 , n55 );
nand ( n4413 , n4411 , n50 , n4412 );
nand ( n4414 , n4410 , n4413 );
not ( n4415 , n4414 );
not ( n4416 , n4415 );
or ( n4417 , n4406 , n4416 );
nand ( n4418 , n4404 , n4414 );
nand ( n4419 , n4417 , n4418 );
not ( n4420 , n4306 );
not ( n4421 , n4342 );
or ( n4422 , n4420 , n4421 );
nand ( n4423 , n3189 , n4340 );
nand ( n4424 , n4422 , n4423 );
not ( n4425 , n4424 );
nand ( n4426 , n67 , n1021 );
not ( n4427 , n4257 );
not ( n4428 , n2207 );
not ( n4429 , n4428 );
or ( n4430 , n4427 , n4429 );
nand ( n4431 , n1017 , n4350 );
nand ( n4432 , n4430 , n4431 );
xnor ( n4433 , n4426 , n4432 );
not ( n4434 , n4433 );
or ( n4435 , n4425 , n4434 );
not ( n4436 , n4426 );
nand ( n4437 , n4436 , n4432 );
nand ( n4438 , n4435 , n4437 );
xor ( n4439 , n4419 , n4438 );
and ( n4440 , n40 , n66 );
not ( n4441 , n40 );
not ( n4442 , n66 );
and ( n4443 , n4441 , n4442 );
nor ( n4444 , n4440 , n4443 );
not ( n4445 , n4444 );
not ( n4446 , n4153 );
or ( n4447 , n4445 , n4446 );
nand ( n4448 , n2742 , n4383 );
nand ( n4449 , n4447 , n4448 );
not ( n4450 , n4449 );
not ( n4451 , n51 );
not ( n4452 , n4412 );
or ( n4453 , n4451 , n4452 );
nand ( n4454 , n4288 , n4283 );
nand ( n4455 , n4453 , n4454 );
not ( n4456 , n4455 );
not ( n4457 , n4318 );
not ( n4458 , n777 );
or ( n4459 , n4457 , n4458 );
nand ( n4460 , n862 , n4328 );
nand ( n4461 , n4459 , n4460 );
not ( n4462 , n4461 );
not ( n4463 , n4462 );
or ( n4464 , n4456 , n4463 );
not ( n4465 , n4455 );
nand ( n4466 , n4465 , n4461 );
nand ( n4467 , n4464 , n4466 );
not ( n4468 , n4467 );
or ( n4469 , n4450 , n4468 );
nand ( n4470 , n4455 , n4461 );
nand ( n4471 , n4469 , n4470 );
and ( n4472 , n4439 , n4471 );
and ( n4473 , n4419 , n4438 );
nor ( n4474 , n4472 , n4473 );
not ( n4475 , n4474 );
not ( n4476 , n4475 );
nand ( n4477 , n4414 , n4405 );
not ( n4478 , n4477 );
not ( n4479 , n4365 );
not ( n4480 , n2433 );
or ( n4481 , n4479 , n4480 );
xor ( n4482 , n38 , n65 );
nand ( n4483 , n560 , n4482 );
nand ( n4484 , n4481 , n4483 );
not ( n4485 , n4387 );
not ( n4486 , n4152 );
or ( n4487 , n4485 , n4486 );
xor ( n4488 , n40 , n63 );
nand ( n4489 , n1892 , n4488 );
nand ( n4490 , n4487 , n4489 );
xor ( n4491 , n4484 , n4490 );
not ( n4492 , n4491 );
or ( n4493 , n4478 , n4492 );
or ( n4494 , n4477 , n4491 );
nand ( n4495 , n4493 , n4494 );
not ( n4496 , n4495 );
not ( n4497 , n4332 );
not ( n4498 , n1690 );
or ( n4499 , n4497 , n4498 );
not ( n4500 , n42 );
not ( n4501 , n61 );
and ( n4502 , n4500 , n4501 );
and ( n4503 , n42 , n61 );
nor ( n4504 , n4502 , n4503 );
nand ( n4505 , n2795 , n4504 );
nand ( n4506 , n4499 , n4505 );
not ( n4507 , n4269 );
or ( n4508 , n4379 , n4507 );
xor ( n4509 , n46 , n57 );
nand ( n4510 , n755 , n4509 );
nand ( n4511 , n4508 , n4510 );
not ( n4512 , n4511 );
not ( n4513 , n4303 );
not ( n4514 , n4345 );
or ( n4515 , n4513 , n4514 );
xor ( n4516 , n1106 , n59 );
nand ( n4517 , n1099 , n4516 );
nand ( n4518 , n4515 , n4517 );
not ( n4519 , n4518 );
not ( n4520 , n4519 );
or ( n4521 , n4512 , n4520 );
not ( n4522 , n4518 );
or ( n4523 , n4522 , n4511 );
nand ( n4524 , n4521 , n4523 );
xnor ( n4525 , n4506 , n4524 );
not ( n4526 , n4525 );
or ( n4527 , n4496 , n4526 );
or ( n4528 , n4525 , n4495 );
nand ( n4529 , n4527 , n4528 );
not ( n4530 , n4529 );
not ( n4531 , n4530 );
or ( n4532 , n4476 , n4531 );
nand ( n4533 , n4474 , n4529 );
nand ( n4534 , n4532 , n4533 );
not ( n4535 , n4347 );
not ( n4536 , n4356 );
or ( n4537 , n4535 , n4536 );
not ( n4538 , n4348 );
not ( n4539 , n4356 );
not ( n4540 , n4539 );
or ( n4541 , n4538 , n4540 );
nand ( n4542 , n4541 , n4334 );
nand ( n4543 , n4537 , n4542 );
not ( n4544 , n4543 );
not ( n4545 , n4354 );
not ( n4546 , n3300 );
or ( n4547 , n4545 , n4546 );
xor ( n4548 , n48 , n55 );
nand ( n4549 , n3296 , n4548 );
nand ( n4550 , n4547 , n4549 );
not ( n4551 , n1471 );
nand ( n4552 , n67 , n4551 );
not ( n4553 , n4552 );
not ( n4554 , n4553 );
not ( n4555 , n4288 );
not ( n4556 , n4408 );
or ( n4557 , n4555 , n4556 );
xor ( n4558 , n50 , n53 );
nand ( n4559 , n51 , n4558 );
nand ( n4560 , n4557 , n4559 );
not ( n4561 , n4560 );
not ( n4562 , n4561 );
or ( n4563 , n4554 , n4562 );
nand ( n4564 , n4552 , n4560 );
nand ( n4565 , n4563 , n4564 );
xnor ( n4566 , n4550 , n4565 );
not ( n4567 , n4566 );
and ( n4568 , n4544 , n4567 );
and ( n4569 , n4543 , n4566 );
nor ( n4570 , n4568 , n4569 );
not ( n4571 , n4371 );
not ( n4572 , n4390 );
or ( n4573 , n4571 , n4572 );
nand ( n4574 , n4382 , n4389 );
nand ( n4575 , n4573 , n4574 );
not ( n4576 , n4575 );
and ( n4577 , n4570 , n4576 );
not ( n4578 , n4570 );
and ( n4579 , n4578 , n4575 );
nor ( n4580 , n4577 , n4579 );
not ( n4581 , n4580 );
and ( n4582 , n4534 , n4581 );
not ( n4583 , n4534 );
and ( n4584 , n4583 , n4580 );
nor ( n4585 , n4582 , n4584 );
not ( n4586 , n4585 );
and ( n4587 , n4400 , n4586 );
not ( n4588 , n4400 );
and ( n4589 , n4588 , n4585 );
nor ( n4590 , n4587 , n4589 );
not ( n4591 , n4326 );
not ( n4592 , n4591 );
not ( n4593 , n4395 );
and ( n4594 , n4592 , n4593 );
and ( n4595 , n4591 , n4395 );
nor ( n4596 , n4594 , n4595 );
not ( n4597 , n4596 );
and ( n4598 , n4439 , n4471 );
not ( n4599 , n4439 );
not ( n4600 , n4471 );
and ( n4601 , n4599 , n4600 );
nor ( n4602 , n4598 , n4601 );
not ( n4603 , n4252 );
not ( n4604 , n4259 );
not ( n4605 , n4604 );
or ( n4606 , n4603 , n4605 );
not ( n4607 , n4252 );
nand ( n4608 , n4607 , n4259 );
nand ( n4609 , n4606 , n4608 );
not ( n4610 , n4609 );
not ( n4611 , n640 );
not ( n4612 , n4611 );
not ( n4613 , n4444 );
or ( n4614 , n4612 , n4613 );
nand ( n4615 , n40 , n67 );
or ( n4616 , n40 , n67 );
nand ( n4617 , n4615 , n4616 , n4153 );
nand ( n4618 , n4614 , n4617 );
xor ( n4619 , n46 , n61 );
not ( n4620 , n4619 );
not ( n4621 , n4271 );
or ( n4622 , n4620 , n4621 );
not ( n4623 , n4262 );
nand ( n4624 , n4623 , n3312 );
nand ( n4625 , n4622 , n4624 );
and ( n4626 , n4618 , n4625 );
not ( n4627 , n4618 );
not ( n4628 , n4625 );
and ( n4629 , n4627 , n4628 );
nor ( n4630 , n4626 , n4629 );
not ( n4631 , n4630 );
or ( n4632 , n4610 , n4631 );
not ( n4633 , n4628 );
nand ( n4634 , n4633 , n4618 );
nand ( n4635 , n4632 , n4634 );
not ( n4636 , n4635 );
xor ( n4637 , n4424 , n4433 );
not ( n4638 , n4637 );
not ( n4639 , n4449 );
not ( n4640 , n4639 );
not ( n4641 , n4467 );
or ( n4642 , n4640 , n4641 );
or ( n4643 , n4639 , n4467 );
nand ( n4644 , n4642 , n4643 );
not ( n4645 , n4644 );
not ( n4646 , n4645 );
or ( n4647 , n4638 , n4646 );
not ( n4648 , n4637 );
nand ( n4649 , n4648 , n4644 );
nand ( n4650 , n4647 , n4649 );
not ( n4651 , n4650 );
or ( n4652 , n4636 , n4651 );
nand ( n4653 , n4637 , n4644 );
nand ( n4654 , n4652 , n4653 );
xor ( n4655 , n4602 , n4654 );
and ( n4656 , n4597 , n4655 );
and ( n4657 , n4602 , n4654 );
nor ( n4658 , n4656 , n4657 );
nand ( n4659 , n4590 , n4658 );
not ( n4660 , n4399 );
not ( n4661 , n4585 );
not ( n4662 , n4661 );
or ( n4663 , n4660 , n4662 );
not ( n4664 , n4581 );
nand ( n4665 , n4664 , n4534 );
nand ( n4666 , n4663 , n4665 );
not ( n4667 , n4666 );
not ( n4668 , n4506 );
not ( n4669 , n4524 );
or ( n4670 , n4668 , n4669 );
not ( n4671 , n4522 );
nand ( n4672 , n4671 , n4511 );
nand ( n4673 , n4670 , n4672 );
not ( n4674 , n4673 );
not ( n4675 , n4674 );
not ( n4676 , n774 );
not ( n4677 , n4676 );
nand ( n4678 , n4677 , n4504 );
or ( n4679 , n2795 , n4678 );
xor ( n4680 , n42 , n60 );
nand ( n4681 , n862 , n4680 );
nand ( n4682 , n4679 , n4681 );
not ( n4683 , n4682 );
not ( n4684 , n755 );
xor ( n4685 , n46 , n56 );
not ( n4686 , n4685 );
or ( n4687 , n4684 , n4686 );
not ( n4688 , n731 );
nand ( n4689 , n4509 , n4688 );
not ( n4690 , n4689 );
nand ( n4691 , n746 , n4690 );
nand ( n4692 , n4687 , n4691 );
not ( n4693 , n4488 );
not ( n4694 , n4152 );
or ( n4695 , n4693 , n4694 );
xor ( n4696 , n40 , n62 );
nand ( n4697 , n1892 , n4696 );
nand ( n4698 , n4695 , n4697 );
xor ( n4699 , n4692 , n4698 );
xor ( n4700 , n4683 , n4699 );
not ( n4701 , n4516 );
not ( n4702 , n4302 );
or ( n4703 , n4701 , n4702 );
xor ( n4704 , n58 , n698 );
nand ( n4705 , n704 , n4704 );
nand ( n4706 , n4703 , n4705 );
not ( n4707 , n477 );
xor ( n4708 , n36 , n66 );
not ( n4709 , n4708 );
or ( n4710 , n4707 , n4709 );
not ( n4711 , n476 );
nand ( n4712 , n4711 , n4078 , n4080 );
not ( n4713 , n4712 );
nor ( n4714 , n36 , n67 );
not ( n4715 , n4714 );
nand ( n4716 , n36 , n67 );
nand ( n4717 , n4713 , n4715 , n4716 );
nand ( n4718 , n4710 , n4717 );
not ( n4719 , n4718 );
xor ( n4720 , n4706 , n4719 );
not ( n4721 , n4548 );
not ( n4722 , n2276 );
or ( n4723 , n4721 , n4722 );
xor ( n4724 , n48 , n54 );
nand ( n4725 , n1017 , n4724 );
nand ( n4726 , n4723 , n4725 );
not ( n4727 , n4726 );
not ( n4728 , n4727 );
xnor ( n4729 , n4720 , n4728 );
xnor ( n4730 , n4700 , n4729 );
buf ( n4731 , n4730 );
not ( n4732 , n4731 );
or ( n4733 , n4675 , n4732 );
or ( n4734 , n4731 , n4674 );
nand ( n4735 , n4733 , n4734 );
not ( n4736 , n4475 );
not ( n4737 , n4529 );
or ( n4738 , n4736 , n4737 );
not ( n4739 , n4525 );
nand ( n4740 , n4739 , n4495 );
nand ( n4741 , n4738 , n4740 );
not ( n4742 , n4741 );
and ( n4743 , n4735 , n4742 );
not ( n4744 , n4735 );
and ( n4745 , n4744 , n4741 );
nor ( n4746 , n4743 , n4745 );
not ( n4747 , n4746 );
not ( n4748 , n4477 );
and ( n4749 , n4748 , n4491 );
and ( n4750 , n4484 , n4490 );
nor ( n4751 , n4749 , n4750 );
not ( n4752 , n4751 );
not ( n4753 , n4550 );
not ( n4754 , n4565 );
or ( n4755 , n4753 , n4754 );
nand ( n4756 , n4553 , n4560 );
nand ( n4757 , n4755 , n4756 );
not ( n4758 , n4482 );
not ( n4759 , n1088 );
or ( n4760 , n4758 , n4759 );
xor ( n4761 , n38 , n64 );
nand ( n4762 , n1022 , n4761 );
nand ( n4763 , n4760 , n4762 );
not ( n4764 , n4763 );
not ( n4765 , n1922 );
not ( n4766 , n67 );
nand ( n4767 , n4766 , n1918 );
not ( n4768 , n4767 );
or ( n4769 , n4765 , n4768 );
nand ( n4770 , n4769 , n36 );
not ( n4771 , n4770 );
not ( n4772 , n2395 );
not ( n4773 , n4558 );
or ( n4774 , n4772 , n4773 );
xor ( n4775 , n50 , n52 );
nand ( n4776 , n51 , n4775 );
nand ( n4777 , n4774 , n4776 );
xnor ( n4778 , n4771 , n4777 );
not ( n4779 , n4778 );
or ( n4780 , n4764 , n4779 );
or ( n4781 , n4763 , n4778 );
nand ( n4782 , n4780 , n4781 );
xnor ( n4783 , n4757 , n4782 );
not ( n4784 , n4783 );
not ( n4785 , n4784 );
or ( n4786 , n4752 , n4785 );
not ( n4787 , n4751 );
nand ( n4788 , n4787 , n4783 );
nand ( n4789 , n4786 , n4788 );
not ( n4790 , n4575 );
not ( n4791 , n4570 );
not ( n4792 , n4791 );
or ( n4793 , n4790 , n4792 );
not ( n4794 , n4566 );
nand ( n4795 , n4543 , n4794 );
nand ( n4796 , n4793 , n4795 );
and ( n4797 , n4789 , n4796 );
not ( n4798 , n4789 );
not ( n4799 , n4796 );
and ( n4800 , n4798 , n4799 );
nor ( n4801 , n4797 , n4800 );
not ( n4802 , n4801 );
nand ( n4803 , n4747 , n4802 );
nand ( n4804 , n4801 , n4746 );
nand ( n4805 , n4667 , n4803 , n4804 );
nand ( n4806 , n4659 , n4805 );
xor ( n4807 , n48 , n60 );
not ( n4808 , n4807 );
not ( n4809 , n2836 );
or ( n4810 , n4808 , n4809 );
nand ( n4811 , n2702 , n4253 );
nand ( n4812 , n4810 , n4811 );
not ( n4813 , n4812 );
not ( n4814 , n677 );
nand ( n4815 , n4814 , n64 );
not ( n4816 , n64 );
nand ( n4817 , n4816 , n688 );
nand ( n4818 , n4815 , n4817 );
not ( n4819 , n4818 );
not ( n4820 , n4302 );
or ( n4821 , n4819 , n4820 );
nand ( n4822 , n704 , n4296 );
nand ( n4823 , n4821 , n4822 );
nand ( n4824 , n67 , n638 );
and ( n4825 , n4823 , n4824 );
not ( n4826 , n4823 );
not ( n4827 , n67 );
nor ( n4828 , n4827 , n885 );
and ( n4829 , n4826 , n4828 );
nor ( n4830 , n4825 , n4829 );
not ( n4831 , n4830 );
not ( n4832 , n4831 );
or ( n4833 , n4813 , n4832 );
not ( n4834 , n4824 );
nand ( n4835 , n4834 , n4823 );
nand ( n4836 , n4833 , n4835 );
not ( n4837 , n4836 );
xor ( n4838 , n42 , n66 );
not ( n4839 , n4838 );
not ( n4840 , n4314 );
or ( n4841 , n4839 , n4840 );
not ( n4842 , n4317 );
or ( n4843 , n4842 , n4311 );
nand ( n4844 , n4841 , n4843 );
not ( n4845 , n4844 );
nand ( n4846 , n51 , n4289 );
xor ( n4847 , n50 , n58 );
nand ( n4848 , n4288 , n4847 );
and ( n4849 , n4846 , n4848 );
xor ( n4850 , n46 , n62 );
not ( n4851 , n4850 );
not ( n4852 , n4269 );
not ( n4853 , n4852 );
not ( n4854 , n4853 );
or ( n4855 , n4851 , n4854 );
nand ( n4856 , n2332 , n4619 );
nand ( n4857 , n4855 , n4856 );
xnor ( n4858 , n4849 , n4857 );
not ( n4859 , n4858 );
or ( n4860 , n4845 , n4859 );
not ( n4861 , n4849 );
nand ( n4862 , n4861 , n4857 );
nand ( n4863 , n4860 , n4862 );
not ( n4864 , n4863 );
not ( n4865 , n4864 );
or ( n4866 , n4837 , n4865 );
not ( n4867 , n4836 );
nand ( n4868 , n4867 , n4863 );
nand ( n4869 , n4866 , n4868 );
not ( n4870 , n4322 );
not ( n4871 , n4870 );
nand ( n4872 , n4871 , n4310 );
not ( n4873 , n4320 );
and ( n4874 , n4872 , n4873 );
not ( n4875 , n4872 );
and ( n4876 , n4875 , n4320 );
nor ( n4877 , n4874 , n4876 );
xor ( n4878 , n4869 , n4877 );
xor ( n4879 , n710 , n65 );
not ( n4880 , n4879 );
not ( n4881 , n4342 );
or ( n4882 , n4880 , n4881 );
nand ( n4883 , n1100 , n4818 );
nand ( n4884 , n4882 , n4883 );
not ( n4885 , n4884 );
not ( n4886 , n4885 );
not ( n4887 , n4886 );
not ( n4888 , n4288 );
xor ( n4889 , n50 , n59 );
not ( n4890 , n4889 );
or ( n4891 , n4888 , n4890 );
nand ( n4892 , n51 , n4847 );
nand ( n4893 , n4891 , n4892 );
not ( n4894 , n4893 );
not ( n4895 , n4894 );
xor ( n4896 , n42 , n67 );
not ( n4897 , n4896 );
not ( n4898 , n776 );
not ( n4899 , n4898 );
or ( n4900 , n4897 , n4899 );
nand ( n4901 , n788 , n4838 );
nand ( n4902 , n4900 , n4901 );
not ( n4903 , n4902 );
or ( n4904 , n4895 , n4903 );
or ( n4905 , n4894 , n4902 );
nand ( n4906 , n4904 , n4905 );
not ( n4907 , n4906 );
or ( n4908 , n4887 , n4907 );
not ( n4909 , n4894 );
nand ( n4910 , n4909 , n4902 );
nand ( n4911 , n4908 , n4910 );
not ( n4912 , n4911 );
not ( n4913 , n67 );
not ( n4914 , n4913 );
not ( n4915 , n2827 );
or ( n4916 , n4914 , n4915 );
nand ( n4917 , n4916 , n2823 );
nand ( n4918 , n42 , n4917 );
not ( n4919 , n4918 );
xor ( n4920 , n48 , n61 );
not ( n4921 , n4920 );
not ( n4922 , n2208 );
or ( n4923 , n4921 , n4922 );
nand ( n4924 , n1017 , n4807 );
nand ( n4925 , n4923 , n4924 );
nand ( n4926 , n4919 , n4925 );
not ( n4927 , n4926 );
not ( n4928 , n4830 );
not ( n4929 , n4928 );
not ( n4930 , n4812 );
not ( n4931 , n4930 );
or ( n4932 , n4929 , n4931 );
nand ( n4933 , n4812 , n4830 );
nand ( n4934 , n4932 , n4933 );
not ( n4935 , n4934 );
or ( n4936 , n4927 , n4935 );
or ( n4937 , n4926 , n4934 );
nand ( n4938 , n4936 , n4937 );
not ( n4939 , n4938 );
or ( n4940 , n4912 , n4939 );
not ( n4941 , n4926 );
nand ( n4942 , n4941 , n4934 );
nand ( n4943 , n4940 , n4942 );
not ( n4944 , n4943 );
not ( n4945 , n4609 );
and ( n4946 , n4630 , n4945 );
not ( n4947 , n4630 );
and ( n4948 , n4947 , n4609 );
nor ( n4949 , n4946 , n4948 );
not ( n4950 , n4949 );
and ( n4951 , n4944 , n4950 );
not ( n4952 , n4944 );
and ( n4953 , n4952 , n4949 );
nor ( n4954 , n4951 , n4953 );
not ( n4955 , n4954 );
and ( n4956 , n4878 , n4955 );
nor ( n4957 , n4949 , n4944 );
nor ( n4958 , n4956 , n4957 );
xor ( n4959 , n4650 , n4635 );
not ( n4960 , n4959 );
not ( n4961 , n4277 );
not ( n4962 , n4280 );
nand ( n4963 , n4961 , n4962 );
nor ( n4964 , n4963 , n4324 );
not ( n4965 , n4964 );
nand ( n4966 , n4281 , n4278 );
nand ( n4967 , n4324 , n4966 );
not ( n4968 , n4962 );
not ( n4969 , n4324 );
nand ( n4970 , n4968 , n4277 , n4969 );
nand ( n4971 , n4965 , n4967 , n4970 );
not ( n4972 , n4877 );
not ( n4973 , n4869 );
or ( n4974 , n4972 , n4973 );
not ( n4975 , n4864 );
nand ( n4976 , n4975 , n4836 );
nand ( n4977 , n4974 , n4976 );
xor ( n4978 , n4971 , n4977 );
nand ( n4979 , n4960 , n4978 );
not ( n4980 , n4979 );
not ( n4981 , n4959 );
nor ( n4982 , n4981 , n4978 );
nor ( n4983 , n4980 , n4982 );
nand ( n4984 , n4958 , n4983 );
not ( n4985 , n4984 );
nor ( n4986 , n4806 , n4985 );
xor ( n4987 , n4844 , n4858 );
and ( n4988 , n1130 , n66 );
not ( n4989 , n1130 );
and ( n4990 , n4989 , n4442 );
nor ( n4991 , n4988 , n4990 );
not ( n4992 , n4991 );
not ( n4993 , n4342 );
or ( n4994 , n4992 , n4993 );
nand ( n4995 , n1100 , n4879 );
nand ( n4996 , n4994 , n4995 );
not ( n4997 , n4996 );
not ( n4998 , n788 );
nor ( n4999 , n4998 , n4913 );
not ( n5000 , n1935 );
not ( n5001 , n5000 );
xor ( n5002 , n50 , n60 );
not ( n5003 , n5002 );
or ( n5004 , n5001 , n5003 );
nand ( n5005 , n51 , n4889 );
nand ( n5006 , n5004 , n5005 );
xnor ( n5007 , n4999 , n5006 );
not ( n5008 , n5007 );
not ( n5009 , n5008 );
or ( n5010 , n4997 , n5009 );
nand ( n5011 , n4999 , n5006 );
nand ( n5012 , n5010 , n5011 );
not ( n5013 , n5012 );
xor ( n5014 , n46 , n63 );
not ( n5015 , n5014 );
not ( n5016 , n4853 );
or ( n5017 , n5015 , n5016 );
nand ( n5018 , n2332 , n4850 );
nand ( n5019 , n5017 , n5018 );
not ( n5020 , n5019 );
not ( n5021 , n4918 );
not ( n5022 , n4925 );
and ( n5023 , n5021 , n5022 );
and ( n5024 , n4918 , n4925 );
nor ( n5025 , n5023 , n5024 );
not ( n5026 , n5025 );
or ( n5027 , n5020 , n5026 );
or ( n5028 , n5019 , n5025 );
nand ( n5029 , n5027 , n5028 );
not ( n5030 , n5029 );
or ( n5031 , n5013 , n5030 );
not ( n5032 , n5025 );
nand ( n5033 , n5019 , n5032 );
nand ( n5034 , n5031 , n5033 );
nand ( n5035 , n4987 , n5034 );
nor ( n5036 , n4987 , n5034 );
not ( n5037 , n5036 );
not ( n5038 , n4911 );
and ( n5039 , n4938 , n5038 );
not ( n5040 , n4938 );
and ( n5041 , n5040 , n4911 );
nor ( n5042 , n5039 , n5041 );
not ( n5043 , n5042 );
nand ( n5044 , n5037 , n5043 );
nand ( n5045 , n5035 , n5044 );
xnor ( n5046 , n4878 , n4954 );
and ( n5047 , n5045 , n5046 );
not ( n5048 , n3067 );
not ( n5049 , n67 );
nand ( n5050 , n5049 , n3061 );
not ( n5051 , n5050 );
or ( n5052 , n5048 , n5051 );
nand ( n5053 , n5052 , n1134 );
not ( n5054 , n5053 );
not ( n5055 , n2395 );
xor ( n5056 , n50 , n61 );
not ( n5057 , n5056 );
or ( n5058 , n5055 , n5057 );
nand ( n5059 , n51 , n5002 );
nand ( n5060 , n5058 , n5059 );
nand ( n5061 , n5054 , n5060 );
not ( n5062 , n5061 );
xor ( n5063 , n46 , n64 );
not ( n5064 , n4852 );
and ( n5065 , n5063 , n5064 );
not ( n5066 , n5014 );
nor ( n5067 , n746 , n5066 );
nor ( n5068 , n5065 , n5067 );
not ( n5069 , n5068 );
nand ( n5070 , n5062 , n5069 );
xor ( n5071 , n48 , n62 );
not ( n5072 , n5071 );
not ( n5073 , n3300 );
or ( n5074 , n5072 , n5073 );
nand ( n5075 , n3296 , n4920 );
nand ( n5076 , n5074 , n5075 );
nand ( n5077 , n5061 , n5068 );
nand ( n5078 , n5076 , n5077 );
nand ( n5079 , n5070 , n5078 );
not ( n5080 , n5079 );
not ( n5081 , n4884 );
not ( n5082 , n5081 );
not ( n5083 , n4906 );
or ( n5084 , n5082 , n5083 );
or ( n5085 , n4885 , n4906 );
nand ( n5086 , n5084 , n5085 );
not ( n5087 , n5086 );
nand ( n5088 , n5080 , n5087 );
not ( n5089 , n5088 );
not ( n5090 , n5029 );
not ( n5091 , n5012 );
not ( n5092 , n5091 );
and ( n5093 , n5090 , n5092 );
and ( n5094 , n5091 , n5029 );
nor ( n5095 , n5093 , n5094 );
not ( n5096 , n5095 );
not ( n5097 , n5096 );
or ( n5098 , n5089 , n5097 );
nand ( n5099 , n5079 , n5086 );
nand ( n5100 , n5098 , n5099 );
not ( n5101 , n5100 );
not ( n5102 , n5036 );
nand ( n5103 , n5102 , n5035 );
xnor ( n5104 , n5103 , n5042 );
nor ( n5105 , n5101 , n5104 );
nor ( n5106 , n5047 , n5105 );
not ( n5107 , n5100 );
nand ( n5108 , n5107 , n5104 );
not ( n5109 , n5076 );
nand ( n5110 , n5070 , n5077 );
not ( n5111 , n5110 );
or ( n5112 , n5109 , n5111 );
or ( n5113 , n5076 , n5110 );
nand ( n5114 , n5112 , n5113 );
not ( n5115 , n5114 );
not ( n5116 , n4996 );
not ( n5117 , n5007 );
and ( n5118 , n5116 , n5117 );
and ( n5119 , n4996 , n5007 );
nor ( n5120 , n5118 , n5119 );
not ( n5121 , n5120 );
not ( n5122 , n2182 );
not ( n5123 , n4991 );
or ( n5124 , n5122 , n5123 );
nand ( n5125 , n1134 , n67 );
or ( n5126 , n1107 , n67 );
nand ( n5127 , n5125 , n5126 , n4342 );
nand ( n5128 , n5124 , n5127 );
not ( n5129 , n5128 );
xor ( n5130 , n46 , n65 );
not ( n5131 , n5130 );
not ( n5132 , n4269 );
or ( n5133 , n5131 , n5132 );
nand ( n5134 , n755 , n5063 );
nand ( n5135 , n5133 , n5134 );
not ( n5136 , n5135 );
xor ( n5137 , n48 , n63 );
not ( n5138 , n5137 );
not ( n5139 , n2208 );
or ( n5140 , n5138 , n5139 );
nand ( n5141 , n800 , n5071 );
nand ( n5142 , n5140 , n5141 );
not ( n5143 , n5142 );
not ( n5144 , n5143 );
or ( n5145 , n5136 , n5144 );
not ( n5146 , n5142 );
or ( n5147 , n5146 , n5135 );
nand ( n5148 , n5145 , n5147 );
not ( n5149 , n5148 );
or ( n5150 , n5129 , n5149 );
not ( n5151 , n5146 );
nand ( n5152 , n5135 , n5151 );
nand ( n5153 , n5150 , n5152 );
not ( n5154 , n5153 );
and ( n5155 , n5121 , n5154 );
and ( n5156 , n5120 , n5153 );
nor ( n5157 , n5155 , n5156 );
not ( n5158 , n5157 );
not ( n5159 , n5158 );
or ( n5160 , n5115 , n5159 );
not ( n5161 , n5120 );
nand ( n5162 , n5161 , n5153 );
nand ( n5163 , n5160 , n5162 );
nand ( n5164 , n5099 , n5088 );
nand ( n5165 , n5096 , n5164 );
not ( n5166 , n5164 );
nand ( n5167 , n5166 , n5095 );
nand ( n5168 , n5165 , n5167 );
and ( n5169 , n5163 , n5168 );
xor ( n5170 , n5114 , n5157 );
not ( n5171 , n5054 );
not ( n5172 , n5060 );
not ( n5173 , n5172 );
and ( n5174 , n5171 , n5173 );
and ( n5175 , n5054 , n5172 );
nor ( n5176 , n5174 , n5175 );
not ( n5177 , n5176 );
not ( n5178 , n5177 );
nand ( n5179 , n67 , n705 );
xor ( n5180 , n50 , n62 );
and ( n5181 , n2395 , n5180 );
nand ( n5182 , n51 , n5056 );
not ( n5183 , n5182 );
nor ( n5184 , n5181 , n5183 );
nand ( n5185 , n5179 , n5184 );
not ( n5186 , n5185 );
xor ( n5187 , n48 , n64 );
not ( n5188 , n5187 );
not ( n5189 , n2498 );
or ( n5190 , n5188 , n5189 );
nand ( n5191 , n1018 , n5137 );
nand ( n5192 , n5190 , n5191 );
not ( n5193 , n5192 );
or ( n5194 , n5186 , n5193 );
nor ( n5195 , n5184 , n5179 );
not ( n5196 , n5195 );
nand ( n5197 , n5194 , n5196 );
not ( n5198 , n5197 );
or ( n5199 , n5178 , n5198 );
or ( n5200 , n5177 , n5197 );
not ( n5201 , n5128 );
not ( n5202 , n5201 );
not ( n5203 , n5148 );
and ( n5204 , n5202 , n5203 );
buf ( n5205 , n5148 );
and ( n5206 , n5201 , n5205 );
nor ( n5207 , n5204 , n5206 );
not ( n5208 , n5207 );
nand ( n5209 , n5200 , n5208 );
nand ( n5210 , n5199 , n5209 );
not ( n5211 , n5210 );
nor ( n5212 , n5170 , n5211 );
or ( n5213 , n5169 , n5212 );
or ( n5214 , n5163 , n5168 );
nand ( n5215 , n5213 , n5214 );
not ( n5216 , n51 );
not ( n5217 , n5180 );
or ( n5218 , n5216 , n5217 );
not ( n5219 , n51 );
not ( n5220 , n50 );
nand ( n5221 , n5220 , n63 );
not ( n5222 , n63 );
nand ( n5223 , n5222 , n50 );
nand ( n5224 , n5221 , n5223 );
nand ( n5225 , n5219 , n50 , n5224 );
nand ( n5226 , n5218 , n5225 );
not ( n5227 , n5226 );
not ( n5228 , n3279 );
not ( n5229 , n67 );
nand ( n5230 , n5229 , n3276 );
not ( n5231 , n5230 );
or ( n5232 , n5228 , n5231 );
nand ( n5233 , n5232 , n46 );
not ( n5234 , n5233 );
or ( n5235 , n5227 , n5234 );
or ( n5236 , n5233 , n5226 );
nand ( n5237 , n5235 , n5236 );
not ( n5238 , n5237 );
not ( n5239 , n2150 );
not ( n5240 , n5239 );
xor ( n5241 , n46 , n66 );
not ( n5242 , n5241 );
or ( n5243 , n5240 , n5242 );
xor ( n5244 , n46 , n67 );
nand ( n5245 , n5244 , n4269 );
nand ( n5246 , n5243 , n5245 );
not ( n5247 , n5246 );
xor ( n5248 , n48 , n65 );
not ( n5249 , n5248 );
not ( n5250 , n2498 );
or ( n5251 , n5249 , n5250 );
nand ( n5252 , n2507 , n5187 );
nand ( n5253 , n5251 , n5252 );
not ( n5254 , n5253 );
not ( n5255 , n5254 );
or ( n5256 , n5247 , n5255 );
or ( n5257 , n5246 , n5254 );
nand ( n5258 , n5256 , n5257 );
not ( n5259 , n5258 );
or ( n5260 , n5238 , n5259 );
nand ( n5261 , n5246 , n5253 );
nand ( n5262 , n5260 , n5261 );
not ( n5263 , n5241 );
not ( n5264 , n4269 );
or ( n5265 , n5263 , n5264 );
nand ( n5266 , n5239 , n5130 );
nand ( n5267 , n5265 , n5266 );
not ( n5268 , n5226 );
nor ( n5269 , n5268 , n5233 );
nor ( n5270 , n5267 , n5269 );
not ( n5271 , n5270 );
nand ( n5272 , n5269 , n5267 );
nand ( n5273 , n5271 , n5272 );
not ( n5274 , n5273 );
not ( n5275 , n5195 );
nand ( n5276 , n5275 , n5185 );
not ( n5277 , n5192 );
and ( n5278 , n5276 , n5277 );
not ( n5279 , n5276 );
and ( n5280 , n5279 , n5192 );
nor ( n5281 , n5278 , n5280 );
not ( n5282 , n5281 );
or ( n5283 , n5274 , n5282 );
or ( n5284 , n5273 , n5281 );
nand ( n5285 , n5283 , n5284 );
or ( n5286 , n5262 , n5285 );
not ( n5287 , n5286 );
not ( n5288 , n5176 );
not ( n5289 , n5197 );
or ( n5290 , n5288 , n5289 );
or ( n5291 , n5176 , n5197 );
nand ( n5292 , n5290 , n5291 );
not ( n5293 , n5292 );
not ( n5294 , n5293 );
not ( n5295 , n5208 );
or ( n5296 , n5294 , n5295 );
nand ( n5297 , n5292 , n5207 );
nand ( n5298 , n5296 , n5297 );
not ( n5299 , n5270 );
not ( n5300 , n5299 );
not ( n5301 , n5281 );
or ( n5302 , n5300 , n5301 );
nand ( n5303 , n5302 , n5272 );
nor ( n5304 , n5298 , n5303 );
nor ( n5305 , n5287 , n5304 );
not ( n5306 , n5305 );
nand ( n5307 , n67 , n745 );
not ( n5308 , n5307 );
not ( n5309 , n1935 );
not ( n5310 , n5309 );
xor ( n5311 , n50 , n64 );
not ( n5312 , n5311 );
or ( n5313 , n5310 , n5312 );
nand ( n5314 , n51 , n5224 );
nand ( n5315 , n5313 , n5314 );
nand ( n5316 , n5308 , n5315 );
xor ( n5317 , n48 , n66 );
not ( n5318 , n5317 );
not ( n5319 , n3215 );
or ( n5320 , n5318 , n5319 );
nand ( n5321 , n1018 , n5248 );
nand ( n5322 , n5320 , n5321 );
not ( n5323 , n5307 );
not ( n5324 , n5315 );
and ( n5325 , n5323 , n5324 );
and ( n5326 , n5307 , n5315 );
nor ( n5327 , n5325 , n5326 );
not ( n5328 , n5327 );
nand ( n5329 , n5322 , n5328 );
and ( n5330 , n5316 , n5329 );
not ( n5331 , n5237 );
nand ( n5332 , n5331 , n5258 );
not ( n5333 , n5332 );
not ( n5334 , n5237 );
nor ( n5335 , n5334 , n5258 );
nor ( n5336 , n5333 , n5335 );
nor ( n5337 , n5330 , n5336 );
not ( n5338 , n5337 );
nand ( n5339 , n5262 , n5285 );
nand ( n5340 , n5330 , n5336 );
not ( n5341 , n4913 );
not ( n5342 , n3459 );
or ( n5343 , n5341 , n5342 );
nand ( n5344 , n5343 , n3463 );
nand ( n5345 , n48 , n5344 );
not ( n5346 , n5345 );
not ( n5347 , n4288 );
xor ( n5348 , n50 , n65 );
not ( n5349 , n5348 );
or ( n5350 , n5347 , n5349 );
nand ( n5351 , n51 , n5311 );
nand ( n5352 , n5350 , n5351 );
nand ( n5353 , n5346 , n5352 );
not ( n5354 , n5353 );
not ( n5355 , n5354 );
not ( n5356 , n5322 );
not ( n5357 , n5327 );
or ( n5358 , n5356 , n5357 );
or ( n5359 , n5322 , n5327 );
nand ( n5360 , n5358 , n5359 );
not ( n5361 , n5360 );
or ( n5362 , n5355 , n5361 );
not ( n5363 , n5354 );
not ( n5364 , n5360 );
not ( n5365 , n5364 );
or ( n5366 , n5363 , n5365 );
nand ( n5367 , n5353 , n5360 );
nand ( n5368 , n5366 , n5367 );
not ( n5369 , n51 );
not ( n5370 , n5348 );
or ( n5371 , n5369 , n5370 );
or ( n5372 , n66 , n4287 );
nand ( n5373 , n5371 , n5372 );
not ( n5374 , n3160 );
and ( n5375 , n67 , n5374 );
not ( n5376 , n67 );
or ( n5377 , n4442 , n1937 );
nand ( n5378 , n5377 , n50 );
and ( n5379 , n5376 , n5378 );
nor ( n5380 , n5375 , n5379 );
nand ( n5381 , n5373 , n5380 );
and ( n5382 , n48 , n67 );
not ( n5383 , n48 );
and ( n5384 , n5383 , n4913 );
nor ( n5385 , n5382 , n5384 );
not ( n5386 , n5385 );
not ( n5387 , n3217 );
or ( n5388 , n5386 , n5387 );
nand ( n5389 , n3296 , n5317 );
nand ( n5390 , n5388 , n5389 );
not ( n5391 , n5346 );
not ( n5392 , n5352 );
not ( n5393 , n5392 );
or ( n5394 , n5391 , n5393 );
nand ( n5395 , n5345 , n5352 );
nand ( n5396 , n5394 , n5395 );
nor ( n5397 , n5390 , n5396 );
or ( n5398 , n5381 , n5397 );
nand ( n5399 , n5390 , n5396 );
nand ( n5400 , n5398 , n5399 );
nand ( n5401 , n5368 , n5400 );
nand ( n5402 , n5362 , n5401 );
nand ( n5403 , n5340 , n5402 );
nand ( n5404 , n5338 , n5339 , n5403 );
not ( n5405 , n5404 );
or ( n5406 , n5306 , n5405 );
nand ( n5407 , n5303 , n5298 );
nand ( n5408 , n5406 , n5407 );
not ( n5409 , n5210 );
nand ( n5410 , n5409 , n5170 );
not ( n5411 , n5163 );
nand ( n5412 , n5411 , n5165 , n5167 );
nand ( n5413 , n5408 , n5410 , n5412 );
nand ( n5414 , n5215 , n5413 );
nand ( n5415 , n5108 , n5414 );
and ( n5416 , n5106 , n5415 );
nor ( n5417 , n5045 , n5046 );
nor ( n5418 , n5416 , n5417 );
not ( n5419 , n5418 );
and ( n5420 , n4959 , n4978 );
and ( n5421 , n4971 , n4977 );
nor ( n5422 , n5420 , n5421 );
xor ( n5423 , n4596 , n4655 );
nand ( n5424 , n5422 , n5423 );
not ( n5425 , n5424 );
nor ( n5426 , n5419 , n5425 );
and ( n5427 , n4986 , n5426 );
nand ( n5428 , n4801 , n4747 );
nand ( n5429 , n4802 , n4746 );
and ( n5430 , n5428 , n5429 , n4666 );
nor ( n5431 , n5427 , n5430 );
not ( n5432 , n4806 );
nor ( n5433 , n5422 , n5423 );
not ( n5434 , n5433 );
nor ( n5435 , n4958 , n4983 );
nand ( n5436 , n5435 , n5424 );
nand ( n5437 , n5434 , n5436 );
and ( n5438 , n5432 , n5437 );
not ( n5439 , n4805 );
not ( n5440 , n4658 );
not ( n5441 , n4590 );
nand ( n5442 , n5440 , n5441 );
nor ( n5443 , n5439 , n5442 );
nor ( n5444 , n5438 , n5443 );
nand ( n5445 , n5431 , n5444 );
not ( n5446 , n5445 );
not ( n5447 , n4685 );
not ( n5448 , n4271 );
or ( n5449 , n5447 , n5448 );
xor ( n5450 , n46 , n55 );
nand ( n5451 , n3014 , n5450 );
nand ( n5452 , n5449 , n5451 );
not ( n5453 , n5452 );
not ( n5454 , n4761 );
not ( n5455 , n573 );
or ( n5456 , n5454 , n5455 );
xor ( n5457 , n38 , n63 );
nand ( n5458 , n1022 , n5457 );
nand ( n5459 , n5456 , n5458 );
not ( n5460 , n5459 );
or ( n5461 , n5453 , n5460 );
or ( n5462 , n5452 , n5459 );
not ( n5463 , n4696 );
not ( n5464 , n4153 );
or ( n5465 , n5463 , n5464 );
xor ( n5466 , n40 , n61 );
nand ( n5467 , n2742 , n5466 );
nand ( n5468 , n5465 , n5467 );
nand ( n5469 , n5462 , n5468 );
nand ( n5470 , n5461 , n5469 );
not ( n5471 , n5470 );
not ( n5472 , n4716 );
not ( n5473 , n51 );
nand ( n5474 , n5473 , n52 );
nand ( n5475 , n50 , n5474 );
not ( n5476 , n5475 );
not ( n5477 , n5476 );
or ( n5478 , n5472 , n5477 );
not ( n5479 , n4716 );
nand ( n5480 , n5479 , n5475 );
nand ( n5481 , n5478 , n5480 );
not ( n5482 , n5481 );
not ( n5483 , n4724 );
not ( n5484 , n3082 );
or ( n5485 , n5483 , n5484 );
xor ( n5486 , n48 , n53 );
nand ( n5487 , n3160 , n5486 );
nand ( n5488 , n5485 , n5487 );
not ( n5489 , n5488 );
or ( n5490 , n5482 , n5489 );
not ( n5491 , n4716 );
nand ( n5492 , n5491 , n5476 );
nand ( n5493 , n5490 , n5492 );
not ( n5494 , n5493 );
not ( n5495 , n5494 );
not ( n5496 , n4708 );
not ( n5497 , n4082 );
or ( n5498 , n5496 , n5497 );
xor ( n5499 , n36 , n65 );
nand ( n5500 , n477 , n5499 );
nand ( n5501 , n5498 , n5500 );
not ( n5502 , n4704 );
not ( n5503 , n4303 );
or ( n5504 , n5502 , n5503 );
not ( n5505 , n1102 );
not ( n5506 , n57 );
not ( n5507 , n5506 );
or ( n5508 , n5505 , n5507 );
not ( n5509 , n1129 );
nand ( n5510 , n5509 , n57 );
nand ( n5511 , n5508 , n5510 );
nand ( n5512 , n705 , n5511 );
nand ( n5513 , n5504 , n5512 );
nand ( n5514 , n5501 , n5513 );
or ( n5515 , n5513 , n5501 );
not ( n5516 , n4680 );
and ( n5517 , n2827 , n2823 );
nor ( n5518 , n5517 , n4676 );
not ( n5519 , n5518 );
or ( n5520 , n5516 , n5519 );
xor ( n5521 , n42 , n59 );
nand ( n5522 , n1903 , n5521 );
nand ( n5523 , n5520 , n5522 );
nand ( n5524 , n5515 , n5523 );
nand ( n5525 , n5514 , n5524 );
not ( n5526 , n5525 );
or ( n5527 , n5495 , n5526 );
nand ( n5528 , n5493 , n5514 , n5524 );
nand ( n5529 , n5527 , n5528 );
not ( n5530 , n5529 );
or ( n5531 , n5471 , n5530 );
not ( n5532 , n5494 );
nand ( n5533 , n5532 , n5525 );
nand ( n5534 , n5531 , n5533 );
not ( n5535 , n5534 );
xor ( n5536 , n42 , n58 );
not ( n5537 , n5536 );
not ( n5538 , n777 );
or ( n5539 , n5537 , n5538 );
xor ( n5540 , n42 , n57 );
nand ( n5541 , n2165 , n5540 );
nand ( n5542 , n5539 , n5541 );
nand ( n5543 , n36 , n65 );
not ( n5544 , n5543 );
xor ( n5545 , n46 , n54 );
not ( n5546 , n5545 );
not ( n5547 , n4268 );
or ( n5548 , n5546 , n5547 );
xor ( n5549 , n46 , n53 );
nand ( n5550 , n730 , n5549 );
nand ( n5551 , n5548 , n5550 );
not ( n5552 , n5551 );
or ( n5553 , n5544 , n5552 );
or ( n5554 , n5543 , n5551 );
nand ( n5555 , n5553 , n5554 );
xor ( n5556 , n5542 , n5555 );
not ( n5557 , n5556 );
xor ( n5558 , n36 , n64 );
not ( n5559 , n5558 );
not ( n5560 , n4082 );
or ( n5561 , n5559 , n5560 );
xor ( n5562 , n36 , n63 );
nand ( n5563 , n1472 , n5562 );
nand ( n5564 , n5561 , n5563 );
not ( n5565 , n5511 );
not ( n5566 , n4303 );
or ( n5567 , n5565 , n5566 );
and ( n5568 , n688 , n56 );
not ( n5569 , n688 );
and ( n5570 , n5569 , n4181 );
nor ( n5571 , n5568 , n5570 );
nand ( n5572 , n3189 , n5571 );
nand ( n5573 , n5567 , n5572 );
and ( n5574 , n5564 , n5573 );
not ( n5575 , n5564 );
not ( n5576 , n5573 );
and ( n5577 , n5575 , n5576 );
nor ( n5578 , n5574 , n5577 );
not ( n5579 , n5578 );
xor ( n5580 , n48 , n52 );
not ( n5581 , n5580 );
not ( n5582 , n3300 );
or ( n5583 , n5581 , n5582 );
nand ( n5584 , n5583 , n1019 );
not ( n5585 , n5584 );
and ( n5586 , n5579 , n5585 );
not ( n5587 , n5579 );
and ( n5588 , n5587 , n5584 );
nor ( n5589 , n5586 , n5588 );
not ( n5590 , n5589 );
or ( n5591 , n5557 , n5590 );
or ( n5592 , n5556 , n5589 );
nand ( n5593 , n5591 , n5592 );
not ( n5594 , n5593 );
not ( n5595 , n5594 );
or ( n5596 , n5535 , n5595 );
or ( n5597 , n5534 , n5594 );
nand ( n5598 , n5596 , n5597 );
xor ( n5599 , n5468 , n5459 );
not ( n5600 , n5452 );
not ( n5601 , n5600 );
xor ( n5602 , n5599 , n5601 );
not ( n5603 , n5602 );
xnor ( n5604 , n5488 , n5481 );
not ( n5605 , n5604 );
not ( n5606 , n5513 );
not ( n5607 , n5523 );
or ( n5608 , n5606 , n5607 );
or ( n5609 , n5513 , n5523 );
nand ( n5610 , n5608 , n5609 );
not ( n5611 , n5501 );
and ( n5612 , n5610 , n5611 );
not ( n5613 , n5610 );
not ( n5614 , n5611 );
and ( n5615 , n5613 , n5614 );
nor ( n5616 , n5612 , n5615 );
not ( n5617 , n5616 );
or ( n5618 , n5605 , n5617 );
or ( n5619 , n5604 , n5616 );
nand ( n5620 , n5618 , n5619 );
not ( n5621 , n5620 );
or ( n5622 , n5603 , n5621 );
not ( n5623 , n5604 );
nand ( n5624 , n5623 , n5616 );
nand ( n5625 , n5622 , n5624 );
not ( n5626 , n5625 );
xor ( n5627 , n5470 , n5529 );
not ( n5628 , n5466 );
not ( n5629 , n4155 );
or ( n5630 , n5628 , n5629 );
xor ( n5631 , n40 , n60 );
nand ( n5632 , n1519 , n5631 );
nand ( n5633 , n5630 , n5632 );
not ( n5634 , n5576 );
not ( n5635 , n5457 );
not ( n5636 , n1088 );
or ( n5637 , n5635 , n5636 );
xor ( n5638 , n38 , n62 );
nand ( n5639 , n1022 , n5638 );
nand ( n5640 , n5637 , n5639 );
not ( n5641 , n5640 );
not ( n5642 , n5641 );
or ( n5643 , n5634 , n5642 );
not ( n5644 , n5576 );
nand ( n5645 , n5644 , n5640 );
nand ( n5646 , n5643 , n5645 );
xnor ( n5647 , n5633 , n5646 );
xnor ( n5648 , n5627 , n5647 );
not ( n5649 , n5648 );
or ( n5650 , n5626 , n5649 );
not ( n5651 , n5647 );
xor ( n5652 , n5470 , n5529 );
nand ( n5653 , n5651 , n5652 );
nand ( n5654 , n5650 , n5653 );
xor ( n5655 , n5598 , n5654 );
not ( n5656 , n5655 );
not ( n5657 , n5633 );
not ( n5658 , n5646 );
or ( n5659 , n5657 , n5658 );
not ( n5660 , n5576 );
not ( n5661 , n5660 );
not ( n5662 , n5641 );
nand ( n5663 , n5661 , n5662 );
nand ( n5664 , n5659 , n5663 );
not ( n5665 , n50 );
nand ( n5666 , n36 , n66 );
not ( n5667 , n5666 );
not ( n5668 , n5667 );
or ( n5669 , n5665 , n5668 );
or ( n5670 , n50 , n5667 );
nand ( n5671 , n5669 , n5670 );
not ( n5672 , n5671 );
not ( n5673 , n5499 );
not ( n5674 , n4712 );
not ( n5675 , n5674 );
or ( n5676 , n5673 , n5675 );
nand ( n5677 , n477 , n5558 );
nand ( n5678 , n5676 , n5677 );
not ( n5679 , n5678 );
or ( n5680 , n5672 , n5679 );
nand ( n5681 , n1406 , n5667 );
nand ( n5682 , n5680 , n5681 );
not ( n5683 , n5682 );
not ( n5684 , n5571 );
not ( n5685 , n4302 );
or ( n5686 , n5684 , n5685 );
and ( n5687 , n688 , n55 );
not ( n5688 , n688 );
not ( n5689 , n55 );
and ( n5690 , n5688 , n5689 );
nor ( n5691 , n5687 , n5690 );
nand ( n5692 , n5691 , n704 );
nand ( n5693 , n5686 , n5692 );
not ( n5694 , n637 );
xor ( n5695 , n40 , n59 );
not ( n5696 , n5695 );
or ( n5697 , n5694 , n5696 );
nand ( n5698 , n5631 , n4152 );
nand ( n5699 , n5697 , n5698 );
xor ( n5700 , n5693 , n5699 );
not ( n5701 , n5638 );
not ( n5702 , n2433 );
or ( n5703 , n5701 , n5702 );
xor ( n5704 , n38 , n61 );
nand ( n5705 , n560 , n5704 );
nand ( n5706 , n5703 , n5705 );
xor ( n5707 , n5700 , n5706 );
xor ( n5708 , n5683 , n5707 );
not ( n5709 , n5450 );
not ( n5710 , n4271 );
or ( n5711 , n5709 , n5710 );
nand ( n5712 , n3312 , n5545 );
nand ( n5713 , n5711 , n5712 );
not ( n5714 , n5713 );
not ( n5715 , n5521 );
not ( n5716 , n5518 );
or ( n5717 , n5715 , n5716 );
nand ( n5718 , n788 , n5536 );
nand ( n5719 , n5717 , n5718 );
not ( n5720 , n5486 );
not ( n5721 , n2498 );
or ( n5722 , n5720 , n5721 );
nand ( n5723 , n2507 , n5580 );
nand ( n5724 , n5722 , n5723 );
xor ( n5725 , n5719 , n5724 );
not ( n5726 , n5725 );
or ( n5727 , n5714 , n5726 );
nand ( n5728 , n5719 , n5724 );
nand ( n5729 , n5727 , n5728 );
xnor ( n5730 , n5708 , n5729 );
xor ( n5731 , n5664 , n5730 );
not ( n5732 , n4683 );
and ( n5733 , n5732 , n4699 );
and ( n5734 , n4692 , n4698 );
nor ( n5735 , n5733 , n5734 );
not ( n5736 , n5735 );
not ( n5737 , n5736 );
nand ( n5738 , n4771 , n4777 );
not ( n5739 , n5738 );
not ( n5740 , n4706 );
not ( n5741 , n5740 );
nand ( n5742 , n4728 , n5741 );
not ( n5743 , n5740 );
not ( n5744 , n4727 );
or ( n5745 , n5743 , n5744 );
nand ( n5746 , n5745 , n4718 );
nand ( n5747 , n5742 , n5746 );
not ( n5748 , n5747 );
or ( n5749 , n5739 , n5748 );
not ( n5750 , n5738 );
nand ( n5751 , n5750 , n5742 , n5746 );
nand ( n5752 , n5749 , n5751 );
not ( n5753 , n5752 );
or ( n5754 , n5737 , n5753 );
not ( n5755 , n5738 );
nand ( n5756 , n5755 , n5747 );
nand ( n5757 , n5754 , n5756 );
not ( n5758 , n5757 );
not ( n5759 , n5725 );
xor ( n5760 , n5713 , n5759 );
xor ( n5761 , n5678 , n5671 );
xnor ( n5762 , n5760 , n5761 );
not ( n5763 , n5762 );
or ( n5764 , n5758 , n5763 );
not ( n5765 , n5713 );
nand ( n5766 , n5765 , n5725 );
not ( n5767 , n5766 );
nand ( n5768 , n5713 , n5759 );
not ( n5769 , n5768 );
or ( n5770 , n5767 , n5769 );
nand ( n5771 , n5770 , n5761 );
nand ( n5772 , n5764 , n5771 );
not ( n5773 , n5772 );
and ( n5774 , n5731 , n5773 );
not ( n5775 , n5731 );
and ( n5776 , n5775 , n5772 );
nor ( n5777 , n5774 , n5776 );
not ( n5778 , n5777 );
and ( n5779 , n5656 , n5778 );
and ( n5780 , n5655 , n5777 );
nor ( n5781 , n5779 , n5780 );
not ( n5782 , n5781 );
and ( n5783 , n5648 , n5625 );
not ( n5784 , n5648 );
not ( n5785 , n5625 );
and ( n5786 , n5784 , n5785 );
nor ( n5787 , n5783 , n5786 );
not ( n5788 , n5787 );
not ( n5789 , n4729 );
xor ( n5790 , n4699 , n5732 );
not ( n5791 , n5790 );
or ( n5792 , n5789 , n5791 );
nand ( n5793 , n4673 , n4730 );
nand ( n5794 , n5792 , n5793 );
not ( n5795 , n5794 );
not ( n5796 , n4757 );
not ( n5797 , n4782 );
or ( n5798 , n5796 , n5797 );
not ( n5799 , n4778 );
nand ( n5800 , n4763 , n5799 );
nand ( n5801 , n5798 , n5800 );
not ( n5802 , n5801 );
not ( n5803 , n5735 );
not ( n5804 , n5752 );
or ( n5805 , n5803 , n5804 );
or ( n5806 , n5735 , n5752 );
nand ( n5807 , n5805 , n5806 );
not ( n5808 , n5807 );
not ( n5809 , n5808 );
or ( n5810 , n5802 , n5809 );
not ( n5811 , n5801 );
nand ( n5812 , n5811 , n5807 );
nand ( n5813 , n5810 , n5812 );
not ( n5814 , n5813 );
or ( n5815 , n5795 , n5814 );
nand ( n5816 , n5801 , n5807 );
nand ( n5817 , n5815 , n5816 );
xnor ( n5818 , n5757 , n5762 );
not ( n5819 , n5818 );
and ( n5820 , n5817 , n5819 );
not ( n5821 , n5817 );
and ( n5822 , n5821 , n5818 );
nor ( n5823 , n5820 , n5822 );
not ( n5824 , n5823 );
or ( n5825 , n5788 , n5824 );
nand ( n5826 , n5819 , n5817 );
nand ( n5827 , n5825 , n5826 );
nor ( n5828 , n5782 , n5827 );
not ( n5829 , n5828 );
not ( n5830 , n5829 );
nor ( n5831 , n5446 , n5830 );
not ( n5832 , n5831 );
and ( n5833 , n42 , n4105 );
not ( n5834 , n42 );
and ( n5835 , n5834 , n53 );
nor ( n5836 , n5833 , n5835 );
not ( n5837 , n5836 );
nand ( n5838 , n5837 , n4317 );
not ( n5839 , n42 );
not ( n5840 , n54 );
and ( n5841 , n5839 , n5840 );
and ( n5842 , n42 , n54 );
nor ( n5843 , n5841 , n5842 );
nand ( n5844 , n5843 , n4314 );
and ( n5845 , n5838 , n5844 );
not ( n5846 , n5845 );
nand ( n5847 , n36 , n61 );
not ( n5848 , n5847 );
and ( n5849 , n40 , n56 );
not ( n5850 , n40 );
and ( n5851 , n5850 , n4181 );
nor ( n5852 , n5849 , n5851 );
not ( n5853 , n5852 );
not ( n5854 , n4154 );
not ( n5855 , n5854 );
or ( n5856 , n5853 , n5855 );
not ( n5857 , n640 );
xor ( n5858 , n40 , n55 );
nand ( n5859 , n5857 , n5858 );
nand ( n5860 , n5856 , n5859 );
not ( n5861 , n5860 );
and ( n5862 , n5848 , n5861 );
and ( n5863 , n5847 , n5860 );
nor ( n5864 , n5862 , n5863 );
not ( n5865 , n5864 );
not ( n5866 , n5865 );
or ( n5867 , n5846 , n5866 );
not ( n5868 , n5847 );
nand ( n5869 , n5868 , n5860 );
nand ( n5870 , n5867 , n5869 );
or ( n5871 , n4840 , n5836 );
not ( n5872 , n42 );
not ( n5873 , n52 );
and ( n5874 , n5872 , n5873 );
and ( n5875 , n42 , n52 );
nor ( n5876 , n5874 , n5875 );
not ( n5877 , n5876 );
or ( n5878 , n4842 , n5877 );
nand ( n5879 , n5871 , n5878 );
and ( n5880 , n38 , n57 );
not ( n5881 , n38 );
and ( n5882 , n5881 , n5506 );
nor ( n5883 , n5880 , n5882 );
not ( n5884 , n574 );
and ( n5885 , n5883 , n5884 );
xor ( n5886 , n38 , n56 );
and ( n5887 , n1022 , n5886 );
nor ( n5888 , n5885 , n5887 );
not ( n5889 , n1325 );
not ( n5890 , n5889 );
not ( n5891 , n4304 );
not ( n5892 , n5891 );
or ( n5893 , n5890 , n5892 );
not ( n5894 , n1650 );
not ( n5895 , n5894 );
nand ( n5896 , n5893 , n5895 );
not ( n5897 , n5896 );
and ( n5898 , n5888 , n5897 );
not ( n5899 , n5888 );
and ( n5900 , n5899 , n5896 );
nor ( n5901 , n5898 , n5900 );
xor ( n5902 , n5879 , n5901 );
xor ( n5903 , n5870 , n5902 );
not ( n5904 , n5858 );
not ( n5905 , n4155 );
or ( n5906 , n5904 , n5905 );
xor ( n5907 , n40 , n54 );
not ( n5908 , n5907 );
or ( n5909 , n1707 , n5908 );
nand ( n5910 , n5906 , n5909 );
nand ( n5911 , n36 , n60 );
not ( n5912 , n5911 );
xor ( n5913 , n36 , n59 );
not ( n5914 , n5913 );
not ( n5915 , n4084 );
or ( n5916 , n5914 , n5915 );
not ( n5917 , n479 );
and ( n5918 , n36 , n58 );
not ( n5919 , n36 );
not ( n5920 , n58 );
and ( n5921 , n5919 , n5920 );
nor ( n5922 , n5918 , n5921 );
nand ( n5923 , n5917 , n5922 );
nand ( n5924 , n5916 , n5923 );
not ( n5925 , n5924 );
and ( n5926 , n5912 , n5925 );
and ( n5927 , n5911 , n5924 );
nor ( n5928 , n5926 , n5927 );
xor ( n5929 , n5910 , n5928 );
not ( n5930 , n5929 );
not ( n5931 , n5845 );
and ( n5932 , n1107 , n52 );
not ( n5933 , n1107 );
and ( n5934 , n5933 , n4209 );
nor ( n5935 , n5932 , n5934 );
not ( n5936 , n5935 );
not ( n5937 , n4304 );
or ( n5938 , n5936 , n5937 );
nand ( n5939 , n5938 , n1651 );
not ( n5940 , n5939 );
xor ( n5941 , n36 , n60 );
not ( n5942 , n5941 );
not ( n5943 , n4083 );
not ( n5944 , n5943 );
or ( n5945 , n5942 , n5944 );
nand ( n5946 , n478 , n5913 );
nand ( n5947 , n5945 , n5946 );
not ( n5948 , n5947 );
or ( n5949 , n5940 , n5948 );
not ( n5950 , n5939 );
not ( n5951 , n5950 );
not ( n5952 , n5947 );
not ( n5953 , n5952 );
or ( n5954 , n5951 , n5953 );
and ( n5955 , n38 , n58 );
not ( n5956 , n38 );
and ( n5957 , n5956 , n5920 );
nor ( n5958 , n5955 , n5957 );
not ( n5959 , n5958 );
not ( n5960 , n1507 );
or ( n5961 , n5959 , n5960 );
nand ( n5962 , n1022 , n5883 );
nand ( n5963 , n5961 , n5962 );
nand ( n5964 , n5954 , n5963 );
nand ( n5965 , n5949 , n5964 );
not ( n5966 , n5965 );
or ( n5967 , n5931 , n5966 );
or ( n5968 , n5845 , n5965 );
nand ( n5969 , n5967 , n5968 );
not ( n5970 , n5969 );
or ( n5971 , n5930 , n5970 );
or ( n5972 , n5929 , n5969 );
nand ( n5973 , n5971 , n5972 );
xor ( n5974 , n5903 , n5973 );
not ( n5975 , n5845 );
not ( n5976 , n5975 );
not ( n5977 , n5865 );
or ( n5978 , n5976 , n5977 );
nand ( n5979 , n5845 , n5864 );
nand ( n5980 , n5978 , n5979 );
nand ( n5981 , n36 , n62 );
xor ( n5982 , n46 , n52 );
not ( n5983 , n5982 );
not ( n5984 , n4853 );
or ( n5985 , n5983 , n5984 );
nand ( n5986 , n5985 , n748 );
not ( n5987 , n5986 );
nand ( n5988 , n5981 , n5987 );
not ( n5989 , n5988 );
xor ( n5990 , n1129 , n54 );
not ( n5991 , n5990 );
not ( n5992 , n4303 );
or ( n5993 , n5991 , n5992 );
xor ( n5994 , n1102 , n53 );
nand ( n5995 , n2304 , n5994 );
nand ( n5996 , n5993 , n5995 );
not ( n5997 , n5996 );
not ( n5998 , n5997 );
not ( n5999 , n5998 );
xor ( n6000 , n38 , n60 );
not ( n6001 , n6000 );
not ( n6002 , n2433 );
or ( n6003 , n6001 , n6002 );
xor ( n6004 , n38 , n59 );
nand ( n6005 , n560 , n6004 );
nand ( n6006 , n6003 , n6005 );
not ( n6007 , n6006 );
not ( n6008 , n6007 );
not ( n6009 , n6008 );
or ( n6010 , n5999 , n6009 );
not ( n6011 , n5997 );
not ( n6012 , n6007 );
or ( n6013 , n6011 , n6012 );
xor ( n6014 , n40 , n58 );
not ( n6015 , n6014 );
not ( n6016 , n4153 );
or ( n6017 , n6015 , n6016 );
xor ( n6018 , n40 , n57 );
nand ( n6019 , n1074 , n6018 );
nand ( n6020 , n6017 , n6019 );
nand ( n6021 , n6013 , n6020 );
nand ( n6022 , n6010 , n6021 );
not ( n6023 , n6022 );
or ( n6024 , n5989 , n6023 );
not ( n6025 , n5981 );
nand ( n6026 , n6025 , n5986 );
nand ( n6027 , n6024 , n6026 );
xor ( n6028 , n5980 , n6027 );
not ( n6029 , n55 );
nor ( n6030 , n6029 , n42 );
not ( n6031 , n42 );
nor ( n6032 , n6031 , n55 );
nor ( n6033 , n6030 , n6032 );
not ( n6034 , n6033 );
not ( n6035 , n4840 );
and ( n6036 , n6034 , n6035 );
and ( n6037 , n4317 , n5843 );
nor ( n6038 , n6036 , n6037 );
xor ( n6039 , n36 , n61 );
not ( n6040 , n6039 );
not ( n6041 , n4084 );
or ( n6042 , n6040 , n6041 );
nand ( n6043 , n1059 , n5941 );
nand ( n6044 , n6042 , n6043 );
not ( n6045 , n6004 );
not ( n6046 , n1507 );
or ( n6047 , n6045 , n6046 );
nand ( n6048 , n562 , n5958 );
nand ( n6049 , n6047 , n6048 );
xor ( n6050 , n6044 , n6049 );
xnor ( n6051 , n6038 , n6050 );
not ( n6052 , n6051 );
xor ( n6053 , n36 , n62 );
not ( n6054 , n6053 );
not ( n6055 , n4085 );
or ( n6056 , n6054 , n6055 );
nand ( n6057 , n1751 , n6039 );
nand ( n6058 , n6056 , n6057 );
and ( n6059 , n36 , n63 );
xor ( n6060 , n42 , n56 );
not ( n6061 , n6060 );
not ( n6062 , n5518 );
or ( n6063 , n6061 , n6062 );
not ( n6064 , n6033 );
nand ( n6065 , n6064 , n2795 );
nand ( n6066 , n6063 , n6065 );
xor ( n6067 , n6059 , n6066 );
and ( n6068 , n6058 , n6067 );
and ( n6069 , n6059 , n6066 );
nor ( n6070 , n6068 , n6069 );
not ( n6071 , n6070 );
not ( n6072 , n6018 );
not ( n6073 , n4153 );
or ( n6074 , n6072 , n6073 );
nand ( n6075 , n4611 , n5852 );
nand ( n6076 , n6074 , n6075 );
not ( n6077 , n2718 );
not ( n6078 , n4270 );
or ( n6079 , n6077 , n6078 );
nand ( n6080 , n6079 , n46 );
not ( n6081 , n6080 );
not ( n6082 , n6081 );
not ( n6083 , n5994 );
not ( n6084 , n4342 );
or ( n6085 , n6083 , n6084 );
nand ( n6086 , n1100 , n5935 );
nand ( n6087 , n6085 , n6086 );
not ( n6088 , n6087 );
or ( n6089 , n6082 , n6088 );
or ( n6090 , n6081 , n6087 );
nand ( n6091 , n6089 , n6090 );
xor ( n6092 , n6076 , n6091 );
not ( n6093 , n6092 );
or ( n6094 , n6071 , n6093 );
or ( n6095 , n6070 , n6092 );
nand ( n6096 , n6094 , n6095 );
not ( n6097 , n6096 );
or ( n6098 , n6052 , n6097 );
not ( n6099 , n6070 );
nand ( n6100 , n6099 , n6092 );
nand ( n6101 , n6098 , n6100 );
and ( n6102 , n6028 , n6101 );
and ( n6103 , n5980 , n6027 );
nor ( n6104 , n6102 , n6103 );
not ( n6105 , n6038 );
and ( n6106 , n6105 , n6050 );
and ( n6107 , n6044 , n6049 );
nor ( n6108 , n6106 , n6107 );
not ( n6109 , n6108 );
not ( n6110 , n6109 );
not ( n6111 , n6076 );
not ( n6112 , n6091 );
or ( n6113 , n6111 , n6112 );
nand ( n6114 , n6080 , n6087 );
nand ( n6115 , n6113 , n6114 );
not ( n6116 , n6115 );
not ( n6117 , n5950 );
not ( n6118 , n5947 );
or ( n6119 , n6117 , n6118 );
or ( n6120 , n5950 , n5947 );
nand ( n6121 , n6119 , n6120 );
and ( n6122 , n6121 , n5963 );
not ( n6123 , n6121 );
not ( n6124 , n5963 );
and ( n6125 , n6123 , n6124 );
nor ( n6126 , n6122 , n6125 );
xnor ( n6127 , n6116 , n6126 );
not ( n6128 , n6127 );
or ( n6129 , n6110 , n6128 );
nand ( n6130 , n6115 , n6126 );
nand ( n6131 , n6129 , n6130 );
not ( n6132 , n6131 );
and ( n6133 , n6104 , n6132 );
not ( n6134 , n6104 );
and ( n6135 , n6134 , n6131 );
nor ( n6136 , n6133 , n6135 );
xor ( n6137 , n5974 , n6136 );
not ( n6138 , n6137 );
not ( n6139 , n6028 );
not ( n6140 , n6101 );
not ( n6141 , n6140 );
and ( n6142 , n6139 , n6141 );
and ( n6143 , n6028 , n6140 );
nor ( n6144 , n6142 , n6143 );
not ( n6145 , n6144 );
not ( n6146 , n6145 );
xor ( n6147 , n6108 , n6127 );
not ( n6148 , n6147 );
xor ( n6149 , n6067 , n6058 );
not ( n6150 , n6149 );
not ( n6151 , n6006 );
not ( n6152 , n5996 );
not ( n6153 , n6152 );
or ( n6154 , n6151 , n6153 );
or ( n6155 , n5997 , n6006 );
nand ( n6156 , n6154 , n6155 );
and ( n6157 , n6156 , n6020 );
not ( n6158 , n6156 );
not ( n6159 , n6020 );
and ( n6160 , n6158 , n6159 );
nor ( n6161 , n6157 , n6160 );
not ( n6162 , n5562 );
not ( n6163 , n5943 );
or ( n6164 , n6162 , n6163 );
nand ( n6165 , n1472 , n6053 );
nand ( n6166 , n6164 , n6165 );
not ( n6167 , n6166 );
not ( n6168 , n5704 );
not ( n6169 , n1506 );
or ( n6170 , n6168 , n6169 );
nand ( n6171 , n1022 , n6000 );
nand ( n6172 , n6170 , n6171 );
not ( n6173 , n6172 );
or ( n6174 , n6167 , n6173 );
or ( n6175 , n6166 , n6172 );
nand ( n6176 , n6175 , n5584 );
nand ( n6177 , n6174 , n6176 );
and ( n6178 , n6161 , n6177 );
not ( n6179 , n6161 );
not ( n6180 , n6177 );
and ( n6181 , n6179 , n6180 );
nor ( n6182 , n6178 , n6181 );
not ( n6183 , n6182 );
or ( n6184 , n6150 , n6183 );
not ( n6185 , n6180 );
nand ( n6186 , n6161 , n6185 );
nand ( n6187 , n6184 , n6186 );
not ( n6188 , n6187 );
xor ( n6189 , n5981 , n5987 );
xor ( n6190 , n6189 , n6022 );
not ( n6191 , n5540 );
not ( n6192 , n1051 );
or ( n6193 , n6191 , n6192 );
nand ( n6194 , n2165 , n6060 );
nand ( n6195 , n6193 , n6194 );
not ( n6196 , n3093 );
not ( n6197 , n3216 );
or ( n6198 , n6196 , n6197 );
nand ( n6199 , n6198 , n48 );
xor ( n6200 , n6195 , n6199 );
not ( n6201 , n5549 );
not ( n6202 , n4271 );
or ( n6203 , n6201 , n6202 );
nand ( n6204 , n2719 , n5982 );
nand ( n6205 , n6203 , n6204 );
and ( n6206 , n6200 , n6205 );
and ( n6207 , n6195 , n6199 );
or ( n6208 , n6206 , n6207 );
not ( n6209 , n6208 );
not ( n6210 , n5691 );
not ( n6211 , n4303 );
or ( n6212 , n6210 , n6211 );
nand ( n6213 , n3189 , n5990 );
nand ( n6214 , n6212 , n6213 );
not ( n6215 , n6214 );
nand ( n6216 , n36 , n64 );
not ( n6217 , n6216 );
and ( n6218 , n5695 , n4152 );
not ( n6219 , n637 );
not ( n6220 , n6014 );
nor ( n6221 , n6219 , n6220 );
nor ( n6222 , n6218 , n6221 );
not ( n6223 , n6222 );
not ( n6224 , n6223 );
or ( n6225 , n6217 , n6224 );
not ( n6226 , n6216 );
nand ( n6227 , n6226 , n6222 );
nand ( n6228 , n6225 , n6227 );
not ( n6229 , n6228 );
or ( n6230 , n6215 , n6229 );
not ( n6231 , n6216 );
nand ( n6232 , n6231 , n6223 );
nand ( n6233 , n6230 , n6232 );
and ( n6234 , n5987 , n6233 );
not ( n6235 , n5987 );
not ( n6236 , n6233 );
and ( n6237 , n6235 , n6236 );
nor ( n6238 , n6234 , n6237 );
not ( n6239 , n6238 );
or ( n6240 , n6209 , n6239 );
not ( n6241 , n6236 );
nand ( n6242 , n5987 , n6241 );
nand ( n6243 , n6240 , n6242 );
xor ( n6244 , n6190 , n6243 );
not ( n6245 , n6244 );
or ( n6246 , n6188 , n6245 );
nand ( n6247 , n6190 , n6243 );
nand ( n6248 , n6246 , n6247 );
not ( n6249 , n6248 );
or ( n6250 , n6148 , n6249 );
or ( n6251 , n6147 , n6248 );
nand ( n6252 , n6250 , n6251 );
not ( n6253 , n6252 );
or ( n6254 , n6146 , n6253 );
not ( n6255 , n6147 );
nand ( n6256 , n6255 , n6248 );
nand ( n6257 , n6254 , n6256 );
not ( n6258 , n6257 );
nand ( n6259 , n6138 , n6258 );
xnor ( n6260 , n5813 , n5794 );
not ( n6261 , n6260 );
and ( n6262 , n5620 , n5602 );
not ( n6263 , n5620 );
not ( n6264 , n5602 );
and ( n6265 , n6263 , n6264 );
nor ( n6266 , n6262 , n6265 );
not ( n6267 , n4796 );
not ( n6268 , n4789 );
or ( n6269 , n6267 , n6268 );
not ( n6270 , n4751 );
nand ( n6271 , n6270 , n4784 );
nand ( n6272 , n6269 , n6271 );
xor ( n6273 , n6266 , n6272 );
not ( n6274 , n6273 );
or ( n6275 , n6261 , n6274 );
or ( n6276 , n6260 , n6273 );
nand ( n6277 , n6275 , n6276 );
not ( n6278 , n6277 );
not ( n6279 , n4735 );
and ( n6280 , n6279 , n4802 );
nor ( n6281 , n6280 , n4742 );
nor ( n6282 , n4802 , n6279 );
nor ( n6283 , n6281 , n6282 );
nand ( n6284 , n6278 , n6283 );
not ( n6285 , n5817 );
xor ( n6286 , n5818 , n6285 );
xnor ( n6287 , n6286 , n5787 );
not ( n6288 , n6260 );
and ( n6289 , n6288 , n6273 );
and ( n6290 , n6266 , n6272 );
nor ( n6291 , n6289 , n6290 );
and ( n6292 , n6287 , n6291 );
not ( n6293 , n6292 );
and ( n6294 , n6259 , n6284 , n6293 );
not ( n6295 , n5777 );
and ( n6296 , n5655 , n6295 );
and ( n6297 , n5598 , n5654 );
nor ( n6298 , n6296 , n6297 );
xnor ( n6299 , n6228 , n6214 );
not ( n6300 , n6299 );
not ( n6301 , n5585 );
not ( n6302 , n5578 );
or ( n6303 , n6301 , n6302 );
nand ( n6304 , n5564 , n5660 );
nand ( n6305 , n6303 , n6304 );
not ( n6306 , n6305 );
or ( n6307 , n6300 , n6306 );
or ( n6308 , n6299 , n6305 );
nand ( n6309 , n6307 , n6308 );
not ( n6310 , n6309 );
xor ( n6311 , n6172 , n6166 );
and ( n6312 , n6311 , n5584 );
not ( n6313 , n6311 );
and ( n6314 , n6313 , n5585 );
nor ( n6315 , n6312 , n6314 );
not ( n6316 , n6315 );
not ( n6317 , n6316 );
or ( n6318 , n6310 , n6317 );
or ( n6319 , n6316 , n6309 );
nand ( n6320 , n6318 , n6319 );
not ( n6321 , n6320 );
and ( n6322 , n5731 , n5772 );
and ( n6323 , n5664 , n5730 );
nor ( n6324 , n6322 , n6323 );
not ( n6325 , n6324 );
or ( n6326 , n6321 , n6325 );
buf ( n6327 , n6320 );
or ( n6328 , n6327 , n6324 );
nand ( n6329 , n6326 , n6328 );
not ( n6330 , n6329 );
not ( n6331 , n5729 );
not ( n6332 , n5683 );
not ( n6333 , n5707 );
or ( n6334 , n6332 , n6333 );
or ( n6335 , n5683 , n5707 );
nand ( n6336 , n6334 , n6335 );
not ( n6337 , n6336 );
or ( n6338 , n6331 , n6337 );
not ( n6339 , n5683 );
nand ( n6340 , n6339 , n5707 );
nand ( n6341 , n6338 , n6340 );
not ( n6342 , n6341 );
and ( n6343 , n5542 , n5555 );
not ( n6344 , n5543 );
nand ( n6345 , n6344 , n5551 );
not ( n6346 , n6345 );
nor ( n6347 , n6343 , n6346 );
not ( n6348 , n5706 );
not ( n6349 , n5699 );
not ( n6350 , n5693 );
and ( n6351 , n6349 , n6350 );
not ( n6352 , n6349 );
and ( n6353 , n6352 , n5693 );
nor ( n6354 , n6351 , n6353 );
not ( n6355 , n6354 );
or ( n6356 , n6348 , n6355 );
not ( n6357 , n6349 );
nand ( n6358 , n5693 , n6357 );
nand ( n6359 , n6356 , n6358 );
not ( n6360 , n6359 );
xor ( n6361 , n6347 , n6360 );
xor ( n6362 , n6195 , n6199 );
xor ( n6363 , n6362 , n6205 );
xnor ( n6364 , n6361 , n6363 );
not ( n6365 , n6364 );
or ( n6366 , n6342 , n6365 );
or ( n6367 , n6341 , n6364 );
nand ( n6368 , n6366 , n6367 );
not ( n6369 , n5534 );
not ( n6370 , n5593 );
or ( n6371 , n6369 , n6370 );
not ( n6372 , n5589 );
nand ( n6373 , n5556 , n6372 );
nand ( n6374 , n6371 , n6373 );
not ( n6375 , n6374 );
and ( n6376 , n6368 , n6375 );
not ( n6377 , n6368 );
not ( n6378 , n6375 );
and ( n6379 , n6377 , n6378 );
nor ( n6380 , n6376 , n6379 );
not ( n6381 , n6380 );
and ( n6382 , n6330 , n6381 );
and ( n6383 , n6380 , n6329 );
nor ( n6384 , n6382 , n6383 );
nand ( n6385 , n6298 , n6384 );
not ( n6386 , n6385 );
not ( n6387 , n6386 );
not ( n6388 , n6380 );
not ( n6389 , n6388 );
not ( n6390 , n6329 );
or ( n6391 , n6389 , n6390 );
not ( n6392 , n6324 );
nand ( n6393 , n6327 , n6392 );
nand ( n6394 , n6391 , n6393 );
not ( n6395 , n6149 );
and ( n6396 , n6182 , n6395 );
not ( n6397 , n6182 );
and ( n6398 , n6397 , n6149 );
nor ( n6399 , n6396 , n6398 );
buf ( n6400 , n6399 );
not ( n6401 , n6400 );
xor ( n6402 , n6208 , n6238 );
not ( n6403 , n6402 );
not ( n6404 , n6363 );
not ( n6405 , n6360 );
not ( n6406 , n6347 );
and ( n6407 , n6405 , n6406 );
not ( n6408 , n6405 );
not ( n6409 , n6406 );
and ( n6410 , n6408 , n6409 );
nor ( n6411 , n6407 , n6410 );
not ( n6412 , n6411 );
or ( n6413 , n6404 , n6412 );
not ( n6414 , n6409 );
nand ( n6415 , n6414 , n6405 );
nand ( n6416 , n6413 , n6415 );
not ( n6417 , n6416 );
not ( n6418 , n6417 );
or ( n6419 , n6403 , n6418 );
not ( n6420 , n6402 );
nand ( n6421 , n6420 , n6416 );
nand ( n6422 , n6419 , n6421 );
not ( n6423 , n6422 );
and ( n6424 , n6401 , n6423 );
and ( n6425 , n6400 , n6422 );
nor ( n6426 , n6424 , n6425 );
not ( n6427 , n6426 );
not ( n6428 , n6315 );
not ( n6429 , n6309 );
or ( n6430 , n6428 , n6429 );
not ( n6431 , n6299 );
nand ( n6432 , n6431 , n6305 );
nand ( n6433 , n6430 , n6432 );
not ( n6434 , n6433 );
not ( n6435 , n6374 );
not ( n6436 , n6368 );
or ( n6437 , n6435 , n6436 );
not ( n6438 , n6364 );
nand ( n6439 , n6341 , n6438 );
nand ( n6440 , n6437 , n6439 );
not ( n6441 , n6440 );
not ( n6442 , n6441 );
or ( n6443 , n6434 , n6442 );
not ( n6444 , n6433 );
nand ( n6445 , n6444 , n6440 );
nand ( n6446 , n6443 , n6445 );
not ( n6447 , n6446 );
or ( n6448 , n6427 , n6447 );
or ( n6449 , n6426 , n6446 );
nand ( n6450 , n6448 , n6449 );
nor ( n6451 , n6394 , n6450 );
not ( n6452 , n6426 );
not ( n6453 , n6452 );
not ( n6454 , n6446 );
or ( n6455 , n6453 , n6454 );
nand ( n6456 , n6433 , n6440 );
nand ( n6457 , n6455 , n6456 );
not ( n6458 , n6051 );
xor ( n6459 , n6458 , n6096 );
not ( n6460 , n6459 );
not ( n6461 , n6187 );
not ( n6462 , n6461 );
not ( n6463 , n6244 );
or ( n6464 , n6462 , n6463 );
or ( n6465 , n6461 , n6244 );
nand ( n6466 , n6464 , n6465 );
not ( n6467 , n6466 );
or ( n6468 , n6460 , n6467 );
or ( n6469 , n6459 , n6466 );
nand ( n6470 , n6468 , n6469 );
not ( n6471 , n6470 );
not ( n6472 , n6400 );
not ( n6473 , n6472 );
not ( n6474 , n6422 );
or ( n6475 , n6473 , n6474 );
nand ( n6476 , n6402 , n6416 );
nand ( n6477 , n6475 , n6476 );
not ( n6478 , n6477 );
not ( n6479 , n6478 );
or ( n6480 , n6471 , n6479 );
or ( n6481 , n6478 , n6470 );
nand ( n6482 , n6480 , n6481 );
nor ( n6483 , n6457 , n6482 );
nor ( n6484 , n6451 , n6483 );
not ( n6485 , n6144 );
not ( n6486 , n6252 );
or ( n6487 , n6485 , n6486 );
or ( n6488 , n6144 , n6252 );
nand ( n6489 , n6487 , n6488 );
not ( n6490 , n6477 );
not ( n6491 , n6470 );
or ( n6492 , n6490 , n6491 );
not ( n6493 , n6459 );
nand ( n6494 , n6493 , n6466 );
nand ( n6495 , n6492 , n6494 );
nor ( n6496 , n6489 , n6495 );
not ( n6497 , n6496 );
nand ( n6498 , n6294 , n6387 , n6484 , n6497 );
not ( n6499 , n6498 );
not ( n6500 , n6499 );
or ( n6501 , n5832 , n6500 );
not ( n6502 , n5827 );
nor ( n6503 , n5781 , n6502 );
nand ( n6504 , n6503 , n6385 );
not ( n6505 , n6298 );
not ( n6506 , n6384 );
nand ( n6507 , n6505 , n6506 );
nand ( n6508 , n6504 , n6507 );
not ( n6509 , n6508 );
not ( n6510 , n6386 );
not ( n6511 , n6291 );
not ( n6512 , n6511 );
not ( n6513 , n6287 );
not ( n6514 , n6513 );
or ( n6515 , n6512 , n6514 );
not ( n6516 , n6283 );
nand ( n6517 , n6516 , n6277 );
nand ( n6518 , n6515 , n6517 );
nor ( n6519 , n6292 , n5828 );
nand ( n6520 , n6510 , n6518 , n6519 );
nand ( n6521 , n6457 , n6482 );
nand ( n6522 , n6137 , n6257 );
nand ( n6523 , n6489 , n6495 );
and ( n6524 , n6521 , n6522 , n6523 );
nand ( n6525 , n6394 , n6450 );
not ( n6526 , n6525 );
not ( n6527 , n6483 );
nand ( n6528 , n6526 , n6527 );
nand ( n6529 , n6509 , n6520 , n6524 , n6528 );
not ( n6530 , n6484 );
and ( n6531 , n6530 , n6524 );
nand ( n6532 , n6522 , n6523 );
nor ( n6533 , n6497 , n6532 );
nor ( n6534 , n6531 , n6533 );
nand ( n6535 , n6529 , n6259 , n6534 );
nand ( n6536 , n6501 , n6535 );
not ( n6537 , n6536 );
not ( n6538 , n6537 );
nand ( n6539 , n4237 , n4247 );
not ( n6540 , n5907 );
not ( n6541 , n4152 );
or ( n6542 , n6540 , n6541 );
not ( n6543 , n886 );
xor ( n6544 , n40 , n53 );
nand ( n6545 , n6543 , n6544 );
nand ( n6546 , n6542 , n6545 );
and ( n6547 , n5886 , n607 );
xor ( n6548 , n38 , n55 );
and ( n6549 , n562 , n6548 );
nor ( n6550 , n6547 , n6549 );
not ( n6551 , n6550 );
and ( n6552 , n6546 , n6551 );
not ( n6553 , n6546 );
and ( n6554 , n6553 , n6550 );
nor ( n6555 , n6552 , n6554 );
not ( n6556 , n5910 );
not ( n6557 , n5928 );
not ( n6558 , n6557 );
or ( n6559 , n6556 , n6558 );
not ( n6560 , n5911 );
nand ( n6561 , n6560 , n5924 );
nand ( n6562 , n6559 , n6561 );
nand ( n6563 , n6555 , n6562 );
not ( n6564 , n6563 );
not ( n6565 , n6555 );
not ( n6566 , n6562 );
and ( n6567 , n6565 , n6566 );
nor ( n6568 , n6564 , n6567 );
not ( n6569 , n5879 );
not ( n6570 , n5901 );
or ( n6571 , n6569 , n6570 );
not ( n6572 , n5888 );
nand ( n6573 , n5896 , n6572 );
nand ( n6574 , n6571 , n6573 );
not ( n6575 , n6574 );
and ( n6576 , n36 , n59 );
not ( n6577 , n5876 );
not ( n6578 , n4314 );
or ( n6579 , n6577 , n6578 );
nand ( n6580 , n6579 , n3859 );
xor ( n6581 , n6576 , n6580 );
not ( n6582 , n5922 );
not ( n6583 , n4085 );
or ( n6584 , n6582 , n6583 );
and ( n6585 , n36 , n57 );
not ( n6586 , n36 );
and ( n6587 , n6586 , n5506 );
nor ( n6588 , n6585 , n6587 );
nand ( n6589 , n1751 , n6588 );
nand ( n6590 , n6584 , n6589 );
not ( n6591 , n6590 );
and ( n6592 , n6581 , n6591 );
not ( n6593 , n6581 );
and ( n6594 , n6593 , n6590 );
nor ( n6595 , n6592 , n6594 );
and ( n6596 , n6575 , n6595 );
not ( n6597 , n6575 );
not ( n6598 , n6595 );
and ( n6599 , n6597 , n6598 );
nor ( n6600 , n6596 , n6599 );
not ( n6601 , n6600 );
or ( n6602 , n6568 , n6601 );
or ( n6603 , n6575 , n6595 );
nand ( n6604 , n6602 , n6603 );
or ( n6605 , n6555 , n6566 );
or ( n6606 , n6550 , n6546 );
nand ( n6607 , n6605 , n6606 );
not ( n6608 , n6607 );
nand ( n6609 , n36 , n58 );
not ( n6610 , n6609 );
not ( n6611 , n6546 );
and ( n6612 , n6610 , n6611 );
and ( n6613 , n6609 , n6546 );
nor ( n6614 , n6612 , n6613 );
not ( n6615 , n6614 );
not ( n6616 , n6548 );
not ( n6617 , n1507 );
or ( n6618 , n6616 , n6617 );
nand ( n6619 , n1022 , n4166 );
nand ( n6620 , n6618 , n6619 );
not ( n6621 , n6620 );
or ( n6622 , n6615 , n6621 );
or ( n6623 , n6620 , n6614 );
nand ( n6624 , n6622 , n6623 );
not ( n6625 , n6624 );
and ( n6626 , n6590 , n6581 );
and ( n6627 , n6576 , n6580 );
nor ( n6628 , n6626 , n6627 );
not ( n6629 , n6628 );
and ( n6630 , n6625 , n6629 );
and ( n6631 , n6628 , n6624 );
nor ( n6632 , n6630 , n6631 );
not ( n6633 , n6632 );
not ( n6634 , n6544 );
not ( n6635 , n6634 );
not ( n6636 , n4203 );
and ( n6637 , n6635 , n6636 );
not ( n6638 , n4202 );
and ( n6639 , n6638 , n4144 );
nor ( n6640 , n6637 , n6639 );
not ( n6641 , n6640 );
not ( n6642 , n6641 );
not ( n6643 , n6588 );
not ( n6644 , n4085 );
or ( n6645 , n6643 , n6644 );
nand ( n6646 , n1059 , n4183 );
nand ( n6647 , n6645 , n6646 );
not ( n6648 , n3823 );
and ( n6649 , n6647 , n6648 );
not ( n6650 , n6647 );
and ( n6651 , n6650 , n3823 );
nor ( n6652 , n6649 , n6651 );
not ( n6653 , n6652 );
not ( n6654 , n6653 );
or ( n6655 , n6642 , n6654 );
nand ( n6656 , n6640 , n6652 );
nand ( n6657 , n6655 , n6656 );
not ( n6658 , n6657 );
and ( n6659 , n6633 , n6658 );
and ( n6660 , n6657 , n6632 );
nor ( n6661 , n6659 , n6660 );
not ( n6662 , n6661 );
and ( n6663 , n6608 , n6662 );
and ( n6664 , n6607 , n6661 );
nor ( n6665 , n6663 , n6664 );
and ( n6666 , n6604 , n6665 );
not ( n6667 , n6604 );
not ( n6668 , n6665 );
and ( n6669 , n6667 , n6668 );
or ( n6670 , n6666 , n6669 );
not ( n6671 , n6568 );
not ( n6672 , n6600 );
or ( n6673 , n6671 , n6672 );
or ( n6674 , n6568 , n6600 );
nand ( n6675 , n6673 , n6674 );
not ( n6676 , n6675 );
not ( n6677 , n5929 );
and ( n6678 , n6677 , n5969 );
and ( n6679 , n5975 , n5965 );
nor ( n6680 , n6678 , n6679 );
not ( n6681 , n6680 );
and ( n6682 , n5903 , n5973 );
and ( n6683 , n5870 , n5902 );
nor ( n6684 , n6682 , n6683 );
not ( n6685 , n6684 );
not ( n6686 , n6685 );
or ( n6687 , n6681 , n6686 );
not ( n6688 , n6680 );
nand ( n6689 , n6688 , n6684 );
nand ( n6690 , n6687 , n6689 );
not ( n6691 , n6690 );
or ( n6692 , n6676 , n6691 );
not ( n6693 , n6680 );
nand ( n6694 , n6693 , n6685 );
nand ( n6695 , n6692 , n6694 );
nor ( n6696 , n6670 , n6695 );
not ( n6697 , n6696 );
xor ( n6698 , n6675 , n6690 );
not ( n6699 , n6698 );
not ( n6700 , n5974 );
not ( n6701 , n6136 );
or ( n6702 , n6700 , n6701 );
not ( n6703 , n6104 );
nand ( n6704 , n6131 , n6703 );
nand ( n6705 , n6702 , n6704 );
not ( n6706 , n6705 );
nand ( n6707 , n6699 , n6706 );
and ( n6708 , n6697 , n6707 );
xor ( n6709 , n4205 , n4206 );
xor ( n6710 , n6709 , n4214 );
and ( n6711 , n4138 , n4160 );
not ( n6712 , n4138 );
and ( n6713 , n6712 , n4159 );
nor ( n6714 , n6711 , n6713 );
xor ( n6715 , n6714 , n4198 );
xnor ( n6716 , n6710 , n6715 );
not ( n6717 , n6640 );
not ( n6718 , n6653 );
and ( n6719 , n6717 , n6718 );
and ( n6720 , n3824 , n6647 );
nor ( n6721 , n6719 , n6720 );
not ( n6722 , n6721 );
not ( n6723 , n4159 );
not ( n6724 , n4174 );
not ( n6725 , n4193 );
or ( n6726 , n6724 , n6725 );
or ( n6727 , n4174 , n4193 );
nand ( n6728 , n6726 , n6727 );
not ( n6729 , n6728 );
and ( n6730 , n6723 , n6729 );
and ( n6731 , n4159 , n6728 );
nor ( n6732 , n6730 , n6731 );
not ( n6733 , n6732 );
and ( n6734 , n6722 , n6733 );
and ( n6735 , n4160 , n6728 );
nor ( n6736 , n6734 , n6735 );
xor ( n6737 , n6716 , n6736 );
not ( n6738 , n6737 );
not ( n6739 , n6628 );
not ( n6740 , n6624 );
not ( n6741 , n6740 );
and ( n6742 , n6739 , n6741 );
not ( n6743 , n6632 );
and ( n6744 , n6657 , n6743 );
nor ( n6745 , n6742 , n6744 );
not ( n6746 , n6745 );
not ( n6747 , n6609 );
not ( n6748 , n6747 );
not ( n6749 , n6546 );
or ( n6750 , n6748 , n6749 );
not ( n6751 , n6620 );
or ( n6752 , n6751 , n6614 );
nand ( n6753 , n6750 , n6752 );
xor ( n6754 , n6721 , n6732 );
and ( n6755 , n6753 , n6754 );
not ( n6756 , n6753 );
not ( n6757 , n6754 );
and ( n6758 , n6756 , n6757 );
or ( n6759 , n6755 , n6758 );
not ( n6760 , n6759 );
and ( n6761 , n6746 , n6760 );
and ( n6762 , n6753 , n6754 );
nor ( n6763 , n6761 , n6762 );
nand ( n6764 , n6738 , n6763 );
not ( n6765 , n6604 );
not ( n6766 , n6668 );
or ( n6767 , n6765 , n6766 );
not ( n6768 , n6661 );
nand ( n6769 , n6768 , n6607 );
nand ( n6770 , n6767 , n6769 );
not ( n6771 , n6770 );
not ( n6772 , n6759 );
and ( n6773 , n6745 , n6772 );
not ( n6774 , n6745 );
and ( n6775 , n6774 , n6759 );
nor ( n6776 , n6773 , n6775 );
nand ( n6777 , n6771 , n6776 );
and ( n6778 , n6708 , n6764 , n6777 );
and ( n6779 , n6539 , n6778 );
xor ( n6780 , n4201 , n4217 );
xor ( n6781 , n6780 , n4234 );
or ( n6782 , n6736 , n6716 );
or ( n6783 , n6710 , n6715 );
nand ( n6784 , n6782 , n6783 );
not ( n6785 , n6784 );
nand ( n6786 , n6781 , n6785 );
nand ( n6787 , n6538 , n6779 , n6786 );
not ( n6788 , n6763 );
nand ( n6789 , n6737 , n6788 );
not ( n6790 , n6789 );
not ( n6791 , n6777 );
nand ( n6792 , n6698 , n6705 );
or ( n6793 , n6696 , n6792 );
nand ( n6794 , n6695 , n6670 );
nand ( n6795 , n6793 , n6794 );
not ( n6796 , n6795 );
or ( n6797 , n6791 , n6796 );
not ( n6798 , n6776 );
nand ( n6799 , n6770 , n6798 );
nand ( n6800 , n6797 , n6799 );
nand ( n6801 , n6800 , n6764 );
not ( n6802 , n6801 );
or ( n6803 , n6790 , n6802 );
nand ( n6804 , n6803 , n6786 );
not ( n6805 , n6781 );
nand ( n6806 , n6805 , n6784 );
nand ( n6807 , n6804 , n6806 );
nand ( n6808 , n6539 , n6807 );
nand ( n6809 , n4249 , n6787 , n6808 );
and ( n6810 , n4103 , n4117 );
not ( n6811 , n4103 );
and ( n6812 , n6811 , n4118 );
nor ( n6813 , n6810 , n6812 );
and ( n6814 , n4246 , n4245 );
and ( n6815 , n4232 , n4241 );
nor ( n6816 , n6814 , n6815 );
nand ( n6817 , n6813 , n6816 );
and ( n6818 , n6809 , n6817 );
nor ( n6819 , n6813 , n6816 );
nor ( n6820 , n6818 , n6819 );
not ( n6821 , n6820 );
not ( n6822 , n6821 );
or ( n6823 , n4127 , n6822 );
and ( n6824 , n4125 , n6820 );
nor ( n6825 , n6824 , n2 );
nand ( n6826 , n6823 , n6825 );
nand ( n6827 , n4071 , n6826 );
not ( n6828 , n6827 );
or ( n6829 , n474 , n6828 );
xor ( n6830 , n466 , n467 );
nand ( n6831 , n381 , n6830 );
nand ( n6832 , n6829 , n6831 );
not ( n6833 , n6832 );
xnor ( n6834 , n395 , n421 );
xnor ( n6835 , n443 , n463 );
or ( n6836 , n6834 , n6835 );
xor ( n6837 , n459 , n450 );
or ( n6838 , n73 , n84 );
nand ( n6839 , n6838 , n457 );
not ( n6840 , n310 );
or ( n6841 , n6839 , n6840 );
or ( n6842 , n346 , n453 );
nand ( n6843 , n6841 , n6842 );
not ( n6844 , n6843 );
xor ( n6845 , n91 , n92 );
not ( n6846 , n6845 );
not ( n6847 , n6846 );
not ( n6848 , n6847 );
not ( n6849 , n6848 );
not ( n6850 , n6849 );
not ( n6851 , n6850 );
not ( n6852 , n6851 );
not ( n6853 , n90 );
not ( n6854 , n91 );
or ( n6855 , n6853 , n6854 );
nor ( n6856 , n90 , n91 );
nor ( n6857 , n6856 , n6845 );
nand ( n6858 , n6855 , n6857 );
not ( n6859 , n6858 );
not ( n6860 , n6859 );
not ( n6861 , n6860 );
not ( n6862 , n6861 );
not ( n6863 , n6862 );
not ( n6864 , n6863 );
and ( n6865 , n6852 , n6864 );
not ( n6866 , n90 );
nor ( n6867 , n6865 , n6866 );
and ( n6868 , n389 , n419 );
and ( n6869 , n69 , n88 );
nor ( n6870 , n6868 , n6869 );
and ( n6871 , n6870 , n416 );
and ( n6872 , n405 , n429 );
nor ( n6873 , n6871 , n6872 );
xor ( n6874 , n6867 , n6873 );
not ( n6875 , n6874 );
or ( n6876 , n6844 , n6875 );
or ( n6877 , n6867 , n6873 );
nand ( n6878 , n6876 , n6877 );
xor ( n6879 , n6878 , n432 );
and ( n6880 , n6837 , n6879 );
and ( n6881 , n432 , n6878 );
nor ( n6882 , n6880 , n6881 );
and ( n6883 , n6836 , n6882 );
and ( n6884 , n6834 , n6835 );
nor ( n6885 , n6883 , n6884 , n1 );
not ( n6886 , n6885 );
nor ( n6887 , n6833 , n6886 );
not ( n6888 , n6887 );
or ( n6889 , n473 , n6888 );
nand ( n6890 , n388 , n470 );
nand ( n6891 , n6889 , n6890 );
not ( n6892 , n6891 );
not ( n6893 , n6892 );
and ( n6894 , n386 , n6893 );
xor ( n6895 , n6879 , n6837 );
not ( n6896 , n6895 );
nand ( n6897 , n74 , n84 );
and ( n6898 , n444 , n419 );
and ( n6899 , n70 , n88 );
nor ( n6900 , n6898 , n6899 );
not ( n6901 , n415 );
and ( n6902 , n6900 , n6901 );
and ( n6903 , n405 , n6870 );
nor ( n6904 , n6902 , n6903 );
xnor ( n6905 , n6897 , n6904 );
not ( n6906 , n71 );
and ( n6907 , n6906 , n358 );
and ( n6908 , n71 , n86 );
nor ( n6909 , n6907 , n6908 );
and ( n6910 , n6909 , n338 );
not ( n6911 , n328 );
and ( n6912 , n6911 , n447 );
nor ( n6913 , n6910 , n6912 );
xnor ( n6914 , n6905 , n6913 );
not ( n6915 , n6914 );
not ( n6916 , n6915 );
xor ( n6917 , n6874 , n6843 );
not ( n6918 , n6917 );
or ( n6919 , n6916 , n6918 );
or ( n6920 , n6915 , n6917 );
not ( n6921 , n90 );
and ( n6922 , n296 , n6921 );
and ( n6923 , n68 , n90 );
nor ( n6924 , n6922 , n6923 );
not ( n6925 , n6864 );
and ( n6926 , n6924 , n6925 );
not ( n6927 , n6852 );
and ( n6928 , n90 , n6927 );
nor ( n6929 , n6926 , n6928 );
nand ( n6930 , n75 , n84 );
or ( n6931 , n74 , n84 );
nand ( n6932 , n6931 , n6897 );
or ( n6933 , n6932 , n309 );
or ( n6934 , n346 , n6839 );
nand ( n6935 , n6933 , n6934 );
and ( n6936 , n6930 , n6935 );
not ( n6937 , n6930 );
not ( n6938 , n6935 );
and ( n6939 , n6937 , n6938 );
nor ( n6940 , n6936 , n6939 );
or ( n6941 , n6929 , n6940 );
or ( n6942 , n6930 , n6938 );
nand ( n6943 , n6941 , n6942 );
nand ( n6944 , n6920 , n6943 );
nand ( n6945 , n6919 , n6944 );
or ( n6946 , n6913 , n6905 );
or ( n6947 , n6897 , n6904 );
nand ( n6948 , n6946 , n6947 );
xnor ( n6949 , n6945 , n6948 );
or ( n6950 , n6896 , n6949 );
and ( n6951 , n6896 , n6949 );
nor ( n6952 , n6951 , n1 );
nand ( n6953 , n6950 , n6952 );
not ( n6954 , n72 );
and ( n6955 , n6954 , n358 );
and ( n6956 , n72 , n86 );
nor ( n6957 , n6955 , n6956 );
and ( n6958 , n6957 , n337 );
and ( n6959 , n327 , n6909 );
nor ( n6960 , n6958 , n6959 );
not ( n6961 , n6960 );
and ( n6962 , n6904 , n6961 );
not ( n6963 , n6904 );
and ( n6964 , n6963 , n6960 );
nor ( n6965 , n6962 , n6964 );
and ( n6966 , n71 , n88 );
nor ( n6967 , n71 , n88 );
nor ( n6968 , n6966 , n6967 );
and ( n6969 , n6968 , n414 );
and ( n6970 , n403 , n6900 );
nor ( n6971 , n6969 , n6970 );
nand ( n6972 , n76 , n84 );
not ( n6973 , n6972 );
not ( n6974 , n6930 );
nor ( n6975 , n75 , n84 );
nor ( n6976 , n6974 , n6975 );
not ( n6977 , n6976 );
not ( n6978 , n306 );
or ( n6979 , n6977 , n6978 );
or ( n6980 , n346 , n6932 );
nand ( n6981 , n6979 , n6980 );
not ( n6982 , n6981 );
and ( n6983 , n6973 , n6982 );
and ( n6984 , n6972 , n6981 );
nor ( n6985 , n6983 , n6984 );
or ( n6986 , n6971 , n6985 );
not ( n6987 , n6981 );
or ( n6988 , n6972 , n6987 );
nand ( n6989 , n6986 , n6988 );
and ( n6990 , n6965 , n6989 );
and ( n6991 , n6961 , n6904 );
nor ( n6992 , n6990 , n6991 );
xor ( n6993 , n6989 , n6965 );
xor ( n6994 , n6929 , n6940 );
and ( n6995 , n73 , n86 );
nor ( n6996 , n73 , n86 );
nor ( n6997 , n6995 , n6996 );
and ( n6998 , n6997 , n336 );
not ( n6999 , n326 );
and ( n7000 , n6999 , n6957 );
nor ( n7001 , n6998 , n7000 );
not ( n7002 , n69 );
not ( n7003 , n90 );
and ( n7004 , n7002 , n7003 );
and ( n7005 , n69 , n90 );
nor ( n7006 , n7004 , n7005 );
not ( n7007 , n7006 );
not ( n7008 , n7007 );
not ( n7009 , n6860 );
and ( n7010 , n7008 , n7009 );
and ( n7011 , n6924 , n6849 );
nor ( n7012 , n7010 , n7011 );
xor ( n7013 , n93 , n94 );
buf ( n7014 , n7013 );
not ( n7015 , n7014 );
not ( n7016 , n7015 );
not ( n7017 , n7016 );
not ( n7018 , n7017 );
not ( n7019 , n92 );
not ( n7020 , n93 );
or ( n7021 , n7019 , n7020 );
nor ( n7022 , n92 , n93 );
nor ( n7023 , n7022 , n7013 );
nand ( n7024 , n7021 , n7023 );
not ( n7025 , n7024 );
not ( n7026 , n7025 );
not ( n7027 , n7026 );
or ( n7028 , n7018 , n7027 );
nand ( n7029 , n7028 , n92 );
and ( n7030 , n7012 , n7029 );
not ( n7031 , n7012 );
not ( n7032 , n7029 );
and ( n7033 , n7031 , n7032 );
nor ( n7034 , n7030 , n7033 );
or ( n7035 , n7001 , n7034 );
or ( n7036 , n7032 , n7012 );
nand ( n7037 , n7035 , n7036 );
xor ( n7038 , n6994 , n7037 );
and ( n7039 , n6993 , n7038 );
and ( n7040 , n7037 , n6994 );
nor ( n7041 , n7039 , n7040 );
or ( n7042 , n6992 , n7041 );
not ( n7043 , n6917 );
not ( n7044 , n6943 );
not ( n7045 , n6914 );
and ( n7046 , n7044 , n7045 );
and ( n7047 , n6943 , n6914 );
nor ( n7048 , n7046 , n7047 );
not ( n7049 , n7048 );
and ( n7050 , n7043 , n7049 );
and ( n7051 , n6917 , n7048 );
nor ( n7052 , n7050 , n7051 );
xnor ( n7053 , n7041 , n6992 );
nor ( n7054 , n7052 , n7053 );
not ( n7055 , n7054 );
nand ( n7056 , n7042 , n7055 );
nand ( n7057 , n381 , n7056 );
and ( n7058 , n6953 , n7057 );
not ( n7059 , n4060 );
nand ( n7060 , n7059 , n3846 );
not ( n7061 , n7060 );
not ( n7062 , n4046 );
not ( n7063 , t_1 );
and ( n7064 , n7061 , n7063 );
and ( n7065 , n7060 , t_1 );
nor ( n7066 , n7064 , n7065 );
not ( n7067 , n2 );
nor ( n7068 , n7066 , n7067 );
not ( n7069 , n6537 );
nand ( n7070 , n7069 , n6778 );
not ( n7071 , n4248 );
nand ( n7072 , n7071 , n6539 );
not ( n7073 , n6807 );
nand ( n7074 , n7072 , n7073 );
and ( n7075 , n7070 , n7074 );
not ( n7076 , n7070 );
not ( n7077 , n7072 );
nand ( n7078 , n7077 , n6786 );
and ( n7079 , n7076 , n7078 );
nor ( n7080 , n7075 , n7079 );
nand ( n7081 , n7067 , n7072 , n6807 );
not ( n7082 , n6786 );
nand ( n7083 , n7082 , n7072 );
nand ( n7084 , n7083 , n7067 , n7073 );
and ( n7085 , n7081 , n7084 );
nor ( n7086 , n7080 , n7085 );
or ( n7087 , n7068 , n7086 );
nand ( n7088 , n7087 , n1 );
nand ( n7089 , n7058 , n7088 );
not ( n7090 , n6817 );
nor ( n7091 , n7090 , n6819 );
not ( n7092 , n7091 );
not ( n7093 , n6809 );
nand ( n7094 , n7092 , n7093 );
and ( n7095 , n7091 , n6809 );
nor ( n7096 , n7095 , n2 );
nand ( n7097 , n7094 , n7096 );
nand ( n7098 , n4064 , n634 );
not ( n7099 , n7098 );
not ( n7100 , t_0 );
or ( n7101 , n7099 , n7100 );
or ( n7102 , n7098 , t_0 );
nand ( n7103 , n7101 , n7102 );
nand ( n7104 , n7103 , n2 );
and ( n7105 , n7097 , n7104 );
nor ( n7106 , n7105 , n381 );
xnor ( n7107 , n6834 , n6835 );
and ( n7108 , n6882 , n7107 );
nor ( n7109 , n6882 , n7107 );
nor ( n7110 , n7108 , n7109 , n1 );
nor ( n7111 , n7106 , n7110 );
or ( n7112 , n6948 , n6895 );
and ( n7113 , n6948 , n6895 );
nor ( n7114 , n7113 , n6945 );
nor ( n7115 , n1 , n7114 );
nand ( n7116 , n7112 , n7115 );
nand ( n7117 , n7111 , n7116 );
and ( n7118 , n7089 , n7117 );
not ( n7119 , n7118 );
not ( n7120 , n7119 );
and ( n7121 , n3992 , n4045 );
not ( n7122 , n7121 );
nand ( n7123 , n4048 , n4003 );
nor ( n7124 , n7123 , n7067 );
not ( n7125 , n7124 );
buf ( n7126 , n4058 );
not ( n7127 , n7126 );
or ( n7128 , n7125 , n7127 );
nand ( n7129 , n7128 , n1 );
nor ( n7130 , n7122 , n7129 );
not ( n7131 , n7130 );
buf ( n7132 , n3704 );
not ( n7133 , n7132 );
or ( n7134 , n7131 , n7133 );
not ( n7135 , n7126 );
nand ( n7136 , n2 , n7123 , n7135 );
not ( n7137 , n7129 );
nand ( n7138 , n7136 , n7137 );
nand ( n7139 , n7134 , n7138 );
not ( n7140 , n7067 );
nand ( n7141 , n6789 , n6764 );
not ( n7142 , n7141 );
or ( n7143 , n7140 , n7142 );
not ( n7144 , n6800 );
nand ( n7145 , n7143 , n7144 );
or ( n7146 , n6777 , n7145 );
nor ( n7147 , n7141 , n2 );
or ( n7148 , n7144 , n7147 );
nand ( n7149 , n7146 , n7148 );
not ( n7150 , n7149 );
not ( n7151 , n6537 );
nand ( n7152 , n7151 , n6708 );
nand ( n7153 , n7150 , n7152 , n7145 );
not ( n7154 , n7147 );
nand ( n7155 , n7154 , n6777 );
not ( n7156 , n7152 );
not ( n7157 , n7149 );
nand ( n7158 , n7155 , n7156 , n7157 );
nand ( n7159 , n7139 , n7153 , n7158 );
and ( n7160 , n3705 , n7121 , n7124 );
or ( n7161 , n7159 , n7160 );
and ( n7162 , n72 , n88 );
nor ( n7163 , n72 , n88 );
nor ( n7164 , n7162 , n7163 );
and ( n7165 , n7164 , n414 );
and ( n7166 , n401 , n6968 );
nor ( n7167 , n7165 , n7166 );
nand ( n7168 , n77 , n84 );
xnor ( n7169 , n7167 , n7168 );
not ( n7170 , n70 );
not ( n7171 , n90 );
and ( n7172 , n7170 , n7171 );
and ( n7173 , n70 , n90 );
nor ( n7174 , n7172 , n7173 );
not ( n7175 , n7174 );
not ( n7176 , n7175 );
not ( n7177 , n6860 );
and ( n7178 , n7176 , n7177 );
not ( n7179 , n6846 );
and ( n7180 , n7006 , n7179 );
nor ( n7181 , n7178 , n7180 );
and ( n7182 , n7169 , n7181 );
not ( n7183 , n7169 );
not ( n7184 , n7181 );
and ( n7185 , n7183 , n7184 );
nor ( n7186 , n7182 , n7185 );
and ( n7187 , n78 , n84 );
xor ( n7188 , n95 , n96 );
buf ( n7189 , n7188 );
not ( n7190 , n7189 );
not ( n7191 , n7190 );
nand ( n7192 , n94 , n7191 );
not ( n7193 , n68 );
not ( n7194 , n94 );
and ( n7195 , n7193 , n7194 );
and ( n7196 , n68 , n94 );
nor ( n7197 , n7195 , n7196 );
not ( n7198 , n94 );
not ( n7199 , n95 );
or ( n7200 , n7198 , n7199 );
nor ( n7201 , n94 , n95 );
nor ( n7202 , n7201 , n7188 );
nand ( n7203 , n7200 , n7202 );
not ( n7204 , n7203 );
nand ( n7205 , n7197 , n7204 );
and ( n7206 , n7192 , n7205 );
not ( n7207 , n7206 );
and ( n7208 , n7187 , n7207 );
not ( n7209 , n7187 );
and ( n7210 , n7209 , n7206 );
nor ( n7211 , n7208 , n7210 );
not ( n7212 , n92 );
and ( n7213 , n444 , n7212 );
and ( n7214 , n70 , n92 );
nor ( n7215 , n7213 , n7214 );
not ( n7216 , n7026 );
and ( n7217 , n7215 , n7216 );
not ( n7218 , n7017 );
and ( n7219 , n389 , n7212 );
and ( n7220 , n69 , n92 );
nor ( n7221 , n7219 , n7220 );
and ( n7222 , n7218 , n7221 );
nor ( n7223 , n7217 , n7222 );
not ( n7224 , n7223 );
not ( n7225 , n7224 );
not ( n7226 , n76 );
not ( n7227 , n86 );
and ( n7228 , n7226 , n7227 );
and ( n7229 , n76 , n86 );
nor ( n7230 , n7228 , n7229 );
and ( n7231 , n7230 , n333 );
and ( n7232 , n75 , n86 );
nor ( n7233 , n75 , n86 );
nor ( n7234 , n7232 , n7233 );
and ( n7235 , n324 , n7234 );
nor ( n7236 , n7231 , n7235 );
and ( n7237 , n74 , n88 );
nor ( n7238 , n74 , n88 );
nor ( n7239 , n7237 , n7238 );
and ( n7240 , n7239 , n412 );
not ( n7241 , n73 );
not ( n7242 , n88 );
and ( n7243 , n7241 , n7242 );
and ( n7244 , n73 , n88 );
nor ( n7245 , n7243 , n7244 );
and ( n7246 , n401 , n7245 );
nor ( n7247 , n7240 , n7246 );
and ( n7248 , n7236 , n7247 );
not ( n7249 , n7236 );
not ( n7250 , n7247 );
and ( n7251 , n7249 , n7250 );
nor ( n7252 , n7248 , n7251 );
not ( n7253 , n7252 );
or ( n7254 , n7225 , n7253 );
not ( n7255 , n7236 );
nand ( n7256 , n7250 , n7255 );
nand ( n7257 , n7254 , n7256 );
and ( n7258 , n7211 , n7257 );
and ( n7259 , n7187 , n7207 );
nor ( n7260 , n7258 , n7259 );
xnor ( n7261 , n7186 , n7260 );
and ( n7262 , n7221 , n7216 );
and ( n7263 , n296 , n7212 );
and ( n7264 , n68 , n92 );
nor ( n7265 , n7263 , n7264 );
and ( n7266 , n7218 , n7265 );
nor ( n7267 , n7262 , n7266 );
not ( n7268 , n413 );
and ( n7269 , n7245 , n7268 );
not ( n7270 , n402 );
and ( n7271 , n7270 , n7164 );
nor ( n7272 , n7269 , n7271 );
not ( n7273 , n7191 );
not ( n7274 , n7273 );
not ( n7275 , n7203 );
or ( n7276 , n7274 , n7275 );
nand ( n7277 , n7276 , n94 );
and ( n7278 , n7272 , n7277 );
not ( n7279 , n7272 );
not ( n7280 , n7277 );
and ( n7281 , n7279 , n7280 );
nor ( n7282 , n7278 , n7281 );
xnor ( n7283 , n7267 , n7282 );
not ( n7284 , n7283 );
or ( n7285 , n77 , n84 );
nand ( n7286 , n7285 , n7168 );
or ( n7287 , n7286 , n307 );
or ( n7288 , n76 , n84 );
nand ( n7289 , n7288 , n6972 );
or ( n7290 , n346 , n7289 );
nand ( n7291 , n7287 , n7290 );
not ( n7292 , n74 );
not ( n7293 , n86 );
and ( n7294 , n7292 , n7293 );
and ( n7295 , n74 , n86 );
nor ( n7296 , n7294 , n7295 );
nand ( n7297 , n325 , n7296 );
nand ( n7298 , n7234 , n333 );
and ( n7299 , n7297 , n7298 );
nand ( n7300 , n7174 , n7179 );
not ( n7301 , n71 );
not ( n7302 , n90 );
or ( n7303 , n7301 , n7302 );
or ( n7304 , n71 , n90 );
nand ( n7305 , n7303 , n7304 );
not ( n7306 , n7305 );
nand ( n7307 , n7306 , n6859 );
and ( n7308 , n7300 , n7307 );
xor ( n7309 , n7299 , n7308 );
xor ( n7310 , n7291 , n7309 );
not ( n7311 , n7305 );
not ( n7312 , n6850 );
and ( n7313 , n7311 , n7312 );
not ( n7314 , n90 );
and ( n7315 , n6954 , n7314 );
and ( n7316 , n72 , n90 );
nor ( n7317 , n7315 , n7316 );
not ( n7318 , n6862 );
and ( n7319 , n7317 , n7318 );
nor ( n7320 , n7313 , n7319 );
nand ( n7321 , n79 , n84 );
xor ( n7322 , n78 , n84 );
not ( n7323 , n7322 );
not ( n7324 , n306 );
or ( n7325 , n7323 , n7324 );
or ( n7326 , n346 , n7286 );
nand ( n7327 , n7325 , n7326 );
and ( n7328 , n7321 , n7327 );
not ( n7329 , n7321 );
not ( n7330 , n7327 );
and ( n7331 , n7329 , n7330 );
nor ( n7332 , n7328 , n7331 );
or ( n7333 , n7320 , n7332 );
or ( n7334 , n7321 , n7330 );
nand ( n7335 , n7333 , n7334 );
xnor ( n7336 , n7310 , n7335 );
not ( n7337 , n7336 );
and ( n7338 , n7284 , n7337 );
and ( n7339 , n7335 , n7310 );
nor ( n7340 , n7338 , n7339 );
or ( n7341 , n7261 , n7340 );
or ( n7342 , n7186 , n7260 );
nand ( n7343 , n7341 , n7342 );
not ( n7344 , n7343 );
or ( n7345 , n7184 , n7169 );
or ( n7346 , n7168 , n7167 );
nand ( n7347 , n7345 , n7346 );
xor ( n7348 , n7001 , n7034 );
xnor ( n7349 , n7347 , n7348 );
xor ( n7350 , n6971 , n6985 );
not ( n7351 , n7026 );
and ( n7352 , n7265 , n7351 );
not ( n7353 , n7014 );
not ( n7354 , n7353 );
and ( n7355 , n92 , n7354 );
nor ( n7356 , n7352 , n7355 );
not ( n7357 , n7356 );
not ( n7358 , n7357 );
and ( n7359 , n7296 , n333 );
and ( n7360 , n324 , n6997 );
nor ( n7361 , n7359 , n7360 );
not ( n7362 , n7289 );
not ( n7363 , n7362 );
not ( n7364 , n306 );
or ( n7365 , n7363 , n7364 );
nand ( n7366 , n302 , n6976 );
nand ( n7367 , n7365 , n7366 );
xnor ( n7368 , n7361 , n7367 );
not ( n7369 , n7368 );
or ( n7370 , n7358 , n7369 );
not ( n7371 , n7361 );
nand ( n7372 , n7367 , n7371 );
nand ( n7373 , n7370 , n7372 );
and ( n7374 , n7373 , n7184 );
not ( n7375 , n7373 );
and ( n7376 , n7375 , n7181 );
nor ( n7377 , n7374 , n7376 );
xnor ( n7378 , n7350 , n7377 );
xnor ( n7379 , n7349 , n7378 );
or ( n7380 , n7267 , n7282 );
or ( n7381 , n7280 , n7272 );
nand ( n7382 , n7380 , n7381 );
not ( n7383 , n7291 );
not ( n7384 , n7309 );
or ( n7385 , n7383 , n7384 );
or ( n7386 , n7308 , n7299 );
nand ( n7387 , n7385 , n7386 );
and ( n7388 , n7368 , n7357 );
not ( n7389 , n7368 );
and ( n7390 , n7389 , n7356 );
nor ( n7391 , n7388 , n7390 );
xor ( n7392 , n7387 , n7391 );
and ( n7393 , n7382 , n7392 );
and ( n7394 , n7387 , n7391 );
nor ( n7395 , n7393 , n7394 );
xor ( n7396 , n7379 , n7395 );
not ( n7397 , n7396 );
or ( n7398 , n7344 , n7397 );
or ( n7399 , n7395 , n7379 );
nand ( n7400 , n7398 , n7399 );
nand ( n7401 , n381 , n7400 );
nand ( n7402 , n7161 , n7401 );
xnor ( n7403 , n7038 , n6993 );
not ( n7404 , n7349 );
not ( n7405 , n7378 );
and ( n7406 , n7404 , n7405 );
and ( n7407 , n7347 , n7348 );
nor ( n7408 , n7406 , n7407 );
and ( n7409 , n7350 , n7377 );
and ( n7410 , n7184 , n7373 );
nor ( n7411 , n7409 , n7410 );
xnor ( n7412 , n7408 , n7411 );
or ( n7413 , n7403 , n7412 );
and ( n7414 , n7403 , n7412 );
nor ( n7415 , n7414 , n1 );
nand ( n7416 , n7413 , n7415 );
not ( n7417 , n7416 );
and ( n7418 , n7402 , n7417 );
and ( n7419 , n7052 , n7053 );
nor ( n7420 , n7419 , n1 , n7054 );
not ( n7421 , n7420 );
and ( n7422 , n4047 , n3840 );
not ( n7423 , n7422 );
not ( n7424 , n7062 );
not ( n7425 , n7132 );
or ( n7426 , n7424 , n7425 );
not ( n7427 , n4048 );
not ( n7428 , n4059 );
nor ( n7429 , n7427 , n7428 );
nand ( n7430 , n7426 , n7429 );
not ( n7431 , n7430 );
or ( n7432 , n7423 , n7431 );
or ( n7433 , n7422 , n7430 );
nand ( n7434 , n7432 , n7433 );
nand ( n7435 , n2 , n7434 );
not ( n7436 , n6789 );
not ( n7437 , n7436 );
nand ( n7438 , n7437 , n7070 , n6801 );
nand ( n7439 , n6806 , n6786 );
and ( n7440 , n7438 , n7439 );
not ( n7441 , n7438 );
not ( n7442 , n7439 );
and ( n7443 , n7441 , n7442 );
nor ( n7444 , n7440 , n7443 );
nand ( n7445 , n7067 , n7444 );
nand ( n7446 , n7435 , n1 , n7445 );
or ( n7447 , n7411 , n7403 );
and ( n7448 , n7408 , n7447 );
and ( n7449 , n7411 , n7403 );
nor ( n7450 , n7448 , n7449 , n1 );
not ( n7451 , n7450 );
nand ( n7452 , n7421 , n7446 , n7451 );
nand ( n7453 , n7418 , n7452 );
not ( n7454 , n7420 );
not ( n7455 , n7454 );
not ( n7456 , n7446 );
or ( n7457 , n7455 , n7456 );
nand ( n7458 , n7457 , n7450 );
nand ( n7459 , n7453 , n7458 );
nand ( n7460 , n7120 , n7459 );
not ( n7461 , n7116 );
not ( n7462 , n7111 );
or ( n7463 , n7461 , n7462 );
and ( n7464 , n7088 , n6953 );
nor ( n7465 , n7464 , n7057 );
nand ( n7466 , n7463 , n7465 );
buf ( n7467 , n7466 );
not ( n7468 , n7110 );
not ( n7469 , n7468 );
not ( n7470 , n7106 );
not ( n7471 , n7470 );
or ( n7472 , n7469 , n7471 );
not ( n7473 , n7116 );
nand ( n7474 , n7472 , n7473 );
nand ( n7475 , n7460 , n7467 , n7474 );
nor ( n7476 , n6832 , n6885 );
nor ( n7477 , n7476 , n471 );
not ( n7478 , n7477 );
nor ( n7479 , n385 , n7478 );
and ( n7480 , n7475 , n7479 );
nor ( n7481 , n6894 , n7480 );
nand ( n7482 , n82 , n84 );
not ( n7483 , n7482 );
not ( n7484 , n7483 );
nand ( n7485 , n81 , n84 );
nor ( n7486 , n81 , n84 );
not ( n7487 , n7486 );
nand ( n7488 , n7485 , n7487 );
not ( n7489 , n7488 );
not ( n7490 , n305 );
and ( n7491 , n7489 , n7490 );
or ( n7492 , n80 , n84 );
nand ( n7493 , n80 , n84 );
nand ( n7494 , n7492 , n7493 );
nor ( n7495 , n346 , n7494 );
nor ( n7496 , n7491 , n7495 );
not ( n7497 , n7496 );
not ( n7498 , n7497 );
or ( n7499 , n7484 , n7498 );
and ( n7500 , n92 , n72 );
not ( n7501 , n92 );
and ( n7502 , n7501 , n6954 );
nor ( n7503 , n7500 , n7502 );
not ( n7504 , n7503 );
not ( n7505 , n7504 );
not ( n7506 , n7017 );
and ( n7507 , n7505 , n7506 );
not ( n7508 , n73 );
and ( n7509 , n7508 , n7212 );
and ( n7510 , n73 , n92 );
nor ( n7511 , n7509 , n7510 );
not ( n7512 , n7025 );
not ( n7513 , n7512 );
and ( n7514 , n7511 , n7513 );
nor ( n7515 , n7507 , n7514 );
and ( n7516 , n7496 , n7483 );
not ( n7517 , n7496 );
and ( n7518 , n7517 , n7482 );
nor ( n7519 , n7516 , n7518 );
or ( n7520 , n7515 , n7519 );
nand ( n7521 , n7499 , n7520 );
or ( n7522 , n7494 , n307 );
or ( n7523 , n79 , n84 );
nand ( n7524 , n7523 , n7321 );
or ( n7525 , n346 , n7524 );
nand ( n7526 , n7522 , n7525 );
not ( n7527 , n75 );
not ( n7528 , n90 );
and ( n7529 , n7527 , n7528 );
and ( n7530 , n75 , n90 );
nor ( n7531 , n7529 , n7530 );
and ( n7532 , n7531 , n6859 );
and ( n7533 , n90 , n74 );
not ( n7534 , n90 );
not ( n7535 , n74 );
and ( n7536 , n7534 , n7535 );
nor ( n7537 , n7533 , n7536 );
and ( n7538 , n7537 , n7179 );
nor ( n7539 , n7532 , n7538 );
nand ( n7540 , n98 , n7539 );
xor ( n7541 , n7526 , n7540 );
xor ( n7542 , n7521 , n7541 );
and ( n7543 , n79 , n86 );
not ( n7544 , n79 );
and ( n7545 , n7544 , n358 );
nor ( n7546 , n7543 , n7545 );
and ( n7547 , n7546 , n333 );
not ( n7548 , n78 );
and ( n7549 , n7548 , n358 );
and ( n7550 , n78 , n86 );
nor ( n7551 , n7549 , n7550 );
and ( n7552 , n325 , n7551 );
nor ( n7553 , n7547 , n7552 );
nand ( n7554 , n83 , n84 );
not ( n7555 , n99 );
nand ( n7556 , n98 , n7555 );
not ( n7557 , n7556 );
xor ( n7558 , n68 , n98 );
and ( n7559 , n7557 , n7558 );
and ( n7560 , n98 , n99 );
nor ( n7561 , n7559 , n7560 );
nor ( n7562 , n7554 , n7561 );
and ( n7563 , n7553 , n7562 );
not ( n7564 , n7553 );
not ( n7565 , n7562 );
and ( n7566 , n7564 , n7565 );
nor ( n7567 , n7563 , n7566 );
nand ( n7568 , n83 , n85 );
or ( n7569 , n83 , n85 );
nand ( n7570 , n7569 , n86 );
nand ( n7571 , n7568 , n84 , n7570 );
not ( n7572 , n7571 );
nand ( n7573 , n7572 , n4 );
not ( n7574 , n7573 );
and ( n7575 , n94 , n72 );
not ( n7576 , n94 );
and ( n7577 , n7576 , n6954 );
nor ( n7578 , n7575 , n7577 );
not ( n7579 , n7578 );
not ( n7580 , n7204 );
or ( n7581 , n7579 , n7580 );
not ( n7582 , n71 );
not ( n7583 , n94 );
and ( n7584 , n7582 , n7583 );
and ( n7585 , n71 , n94 );
nor ( n7586 , n7584 , n7585 );
nand ( n7587 , n7586 , n7189 );
nand ( n7588 , n7581 , n7587 );
not ( n7589 , n7588 );
not ( n7590 , n7589 );
and ( n7591 , n7574 , n7590 );
xor ( n7592 , n76 , n90 );
not ( n7593 , n7592 );
not ( n7594 , n6858 );
not ( n7595 , n7594 );
or ( n7596 , n7593 , n7595 );
not ( n7597 , n6846 );
nand ( n7598 , n7531 , n7597 );
nand ( n7599 , n7596 , n7598 );
not ( n7600 , n7573 );
nor ( n7601 , n7600 , n7588 );
not ( n7602 , n7601 );
and ( n7603 , n7599 , n7602 );
nor ( n7604 , n7591 , n7603 );
or ( n7605 , n7567 , n7604 );
or ( n7606 , n7565 , n7553 );
nand ( n7607 , n7605 , n7606 );
and ( n7608 , n7537 , n6861 );
not ( n7609 , n73 );
not ( n7610 , n90 );
and ( n7611 , n7609 , n7610 );
and ( n7612 , n73 , n90 );
nor ( n7613 , n7611 , n7612 );
not ( n7614 , n6848 );
and ( n7615 , n7613 , n7614 );
nor ( n7616 , n7608 , n7615 );
not ( n7617 , n7616 );
not ( n7618 , n7485 );
and ( n7619 , n76 , n88 );
nor ( n7620 , n76 , n88 );
nor ( n7621 , n7619 , n7620 );
not ( n7622 , n7621 );
nand ( n7623 , n398 , n400 );
not ( n7624 , n411 );
nor ( n7625 , n7623 , n7624 );
not ( n7626 , n7625 );
or ( n7627 , n7622 , n7626 );
not ( n7628 , n75 );
not ( n7629 , n88 );
and ( n7630 , n7628 , n7629 );
and ( n7631 , n75 , n88 );
nor ( n7632 , n7630 , n7631 );
nand ( n7633 , n401 , n7632 );
nand ( n7634 , n7627 , n7633 );
not ( n7635 , n7634 );
or ( n7636 , n7618 , n7635 );
or ( n7637 , n7485 , n7634 );
nand ( n7638 , n7636 , n7637 );
not ( n7639 , n7638 );
or ( n7640 , n7617 , n7639 );
or ( n7641 , n7616 , n7638 );
nand ( n7642 , n7640 , n7641 );
xor ( n7643 , n7607 , n7642 );
xnor ( n7644 , n7542 , n7643 );
and ( n7645 , n7519 , n7515 );
not ( n7646 , n7519 );
not ( n7647 , n7515 );
and ( n7648 , n7646 , n7647 );
nor ( n7649 , n7645 , n7648 );
or ( n7650 , n98 , n7539 );
nand ( n7651 , n7650 , n7540 );
xor ( n7652 , n7649 , n7651 );
not ( n7653 , n74 );
not ( n7654 , n92 );
and ( n7655 , n7653 , n7654 );
and ( n7656 , n74 , n92 );
nor ( n7657 , n7655 , n7656 );
and ( n7658 , n7657 , n7216 );
and ( n7659 , n7354 , n7511 );
nor ( n7660 , n7658 , n7659 );
not ( n7661 , n7660 );
not ( n7662 , n7661 );
xnor ( n7663 , n82 , n84 );
or ( n7664 , n7663 , n305 );
or ( n7665 , n346 , n7488 );
nand ( n7666 , n7664 , n7665 );
not ( n7667 , n7666 );
and ( n7668 , n96 , n70 );
not ( n7669 , n96 );
and ( n7670 , n7669 , n444 );
nor ( n7671 , n7668 , n7670 );
not ( n7672 , n7671 );
nor ( n7673 , n96 , n97 );
not ( n7674 , n7673 );
not ( n7675 , n97 );
not ( n7676 , n98 );
or ( n7677 , n7675 , n7676 );
or ( n7678 , n97 , n98 );
nand ( n7679 , n7677 , n7678 );
nand ( n7680 , n96 , n97 );
nand ( n7681 , n7674 , n7679 , n7680 );
not ( n7682 , n7681 );
not ( n7683 , n7682 );
or ( n7684 , n7672 , n7683 );
and ( n7685 , n96 , n69 );
not ( n7686 , n96 );
and ( n7687 , n7686 , n389 );
nor ( n7688 , n7685 , n7687 );
not ( n7689 , n7679 );
nand ( n7690 , n7688 , n7689 );
nand ( n7691 , n7684 , n7690 );
not ( n7692 , n7691 );
not ( n7693 , n7692 );
or ( n7694 , n7667 , n7693 );
or ( n7695 , n7666 , n7692 );
nand ( n7696 , n7694 , n7695 );
not ( n7697 , n7696 );
or ( n7698 , n7662 , n7697 );
not ( n7699 , n7666 );
or ( n7700 , n7699 , n7692 );
nand ( n7701 , n7698 , n7700 );
xor ( n7702 , n7652 , n7701 );
and ( n7703 , n7561 , n7554 );
not ( n7704 , n7561 );
not ( n7705 , n7554 );
and ( n7706 , n7704 , n7705 );
or ( n7707 , n7703 , n7706 );
not ( n7708 , n7707 );
and ( n7709 , n80 , n86 );
not ( n7710 , n80 );
and ( n7711 , n7710 , n358 );
nor ( n7712 , n7709 , n7711 );
not ( n7713 , n7712 );
not ( n7714 , n333 );
or ( n7715 , n7713 , n7714 );
nand ( n7716 , n324 , n7546 );
nand ( n7717 , n7715 , n7716 );
not ( n7718 , n7717 );
not ( n7719 , n78 );
not ( n7720 , n88 );
or ( n7721 , n7719 , n7720 );
or ( n7722 , n78 , n88 );
nand ( n7723 , n7721 , n7722 );
not ( n7724 , n7723 );
not ( n7725 , n7625 );
not ( n7726 , n7725 );
and ( n7727 , n7724 , n7726 );
nand ( n7728 , n398 , n400 );
xor ( n7729 , n77 , n88 );
and ( n7730 , n7728 , n7729 );
nor ( n7731 , n7727 , n7730 );
not ( n7732 , n7731 );
or ( n7733 , n7718 , n7732 );
or ( n7734 , n7731 , n7717 );
nand ( n7735 , n7733 , n7734 );
not ( n7736 , n7735 );
or ( n7737 , n7708 , n7736 );
or ( n7738 , n7707 , n7735 );
nand ( n7739 , n7737 , n7738 );
not ( n7740 , n7739 );
not ( n7741 , n7661 );
not ( n7742 , n7697 );
or ( n7743 , n7741 , n7742 );
nand ( n7744 , n7660 , n7696 );
nand ( n7745 , n7743 , n7744 );
not ( n7746 , n7745 );
or ( n7747 , n7740 , n7746 );
or ( n7748 , n7739 , n7745 );
and ( n7749 , n7599 , n7601 );
not ( n7750 , n7599 );
and ( n7751 , n7750 , n7573 , n7588 );
nor ( n7752 , n7749 , n7751 );
nor ( n7753 , n7573 , n7588 );
and ( n7754 , n7750 , n7753 );
and ( n7755 , n7599 , n7600 , n7588 );
nor ( n7756 , n7754 , n7755 );
nand ( n7757 , n7752 , n7756 );
nand ( n7758 , n7748 , n7757 );
nand ( n7759 , n7747 , n7758 );
xor ( n7760 , n7604 , n7567 );
xor ( n7761 , n7759 , n7760 );
and ( n7762 , n7702 , n7761 );
and ( n7763 , n7760 , n7759 );
nor ( n7764 , n7762 , n7763 );
or ( n7765 , n7644 , n7764 );
and ( n7766 , n7652 , n7701 );
and ( n7767 , n7651 , n7649 );
nor ( n7768 , n7766 , n7767 );
not ( n7769 , n68 );
not ( n7770 , n96 );
and ( n7771 , n7769 , n7770 );
and ( n7772 , n68 , n96 );
nor ( n7773 , n7771 , n7772 );
not ( n7774 , n7773 );
not ( n7775 , n7681 );
not ( n7776 , n7775 );
or ( n7777 , n7774 , n7776 );
nand ( n7778 , n96 , n7689 );
nand ( n7779 , n7777 , n7778 );
not ( n7780 , n7779 );
not ( n7781 , n69 );
not ( n7782 , n94 );
and ( n7783 , n7781 , n7782 );
and ( n7784 , n69 , n94 );
nor ( n7785 , n7783 , n7784 );
not ( n7786 , n7190 );
nand ( n7787 , n7785 , n7786 );
not ( n7788 , n70 );
not ( n7789 , n94 );
and ( n7790 , n7788 , n7789 );
and ( n7791 , n70 , n94 );
nor ( n7792 , n7790 , n7791 );
nand ( n7793 , n7792 , n7204 );
and ( n7794 , n7787 , n7793 );
nor ( n7795 , n7780 , n7794 );
not ( n7796 , n7795 );
nand ( n7797 , n7794 , n7780 );
nand ( n7798 , n7796 , n7797 );
not ( n7799 , n7503 );
not ( n7800 , n7025 );
or ( n7801 , n7799 , n7800 );
not ( n7802 , n7353 );
not ( n7803 , n71 );
not ( n7804 , n92 );
and ( n7805 , n7803 , n7804 );
and ( n7806 , n71 , n92 );
nor ( n7807 , n7805 , n7806 );
nand ( n7808 , n7802 , n7807 );
nand ( n7809 , n7801 , n7808 );
not ( n7810 , n325 );
not ( n7811 , n77 );
and ( n7812 , n7811 , n358 );
and ( n7813 , n77 , n86 );
nor ( n7814 , n7812 , n7813 );
not ( n7815 , n7814 );
or ( n7816 , n7810 , n7815 );
nand ( n7817 , n7551 , n334 );
nand ( n7818 , n7816 , n7817 );
xor ( n7819 , n7809 , n7818 );
xor ( n7820 , n7798 , n7819 );
and ( n7821 , n7586 , n7204 );
not ( n7822 , n7273 );
and ( n7823 , n7792 , n7822 );
nor ( n7824 , n7821 , n7823 );
not ( n7825 , n7688 );
not ( n7826 , n7775 );
or ( n7827 , n7825 , n7826 );
nand ( n7828 , n7773 , n7689 );
nand ( n7829 , n7827 , n7828 );
not ( n7830 , n7829 );
and ( n7831 , n7729 , n7268 );
and ( n7832 , n401 , n7621 );
nor ( n7833 , n7831 , n7832 );
xnor ( n7834 , n7830 , n7833 );
or ( n7835 , n7824 , n7834 );
or ( n7836 , n7830 , n7833 );
nand ( n7837 , n7835 , n7836 );
xnor ( n7838 , n7820 , n7837 );
xnor ( n7839 , n7768 , n7838 );
xor ( n7840 , n7834 , n7824 );
not ( n7841 , n7735 );
or ( n7842 , n7707 , n7841 );
not ( n7843 , n7717 );
or ( n7844 , n7731 , n7843 );
nand ( n7845 , n7842 , n7844 );
xor ( n7846 , n7840 , n7845 );
and ( n7847 , n94 , n73 );
not ( n7848 , n94 );
and ( n7849 , n7848 , n7508 );
nor ( n7850 , n7847 , n7849 );
and ( n7851 , n7850 , n7204 );
and ( n7852 , n7578 , n7191 );
nor ( n7853 , n7851 , n7852 );
xor ( n7854 , n81 , n86 );
and ( n7855 , n333 , n7854 );
and ( n7856 , n325 , n7712 );
nor ( n7857 , n7855 , n7856 );
or ( n7858 , n7663 , n346 );
or ( n7859 , n83 , n84 );
not ( n7860 , n305 );
nand ( n7861 , n7859 , n7554 , n7860 );
nand ( n7862 , n7858 , n7861 );
and ( n7863 , n7857 , n7862 );
not ( n7864 , n7857 );
not ( n7865 , n7862 );
and ( n7866 , n7864 , n7865 );
nor ( n7867 , n7863 , n7866 );
or ( n7868 , n7853 , n7867 );
or ( n7869 , n7865 , n7857 );
nand ( n7870 , n7868 , n7869 );
not ( n7871 , n75 );
and ( n7872 , n92 , n7871 );
not ( n7873 , n92 );
and ( n7874 , n7873 , n75 );
nor ( n7875 , n7872 , n7874 );
not ( n7876 , n7875 );
not ( n7877 , n7026 );
and ( n7878 , n7876 , n7877 );
not ( n7879 , n7017 );
and ( n7880 , n7879 , n7657 );
nor ( n7881 , n7878 , n7880 );
not ( n7882 , n7881 );
xor ( n7883 , n69 , n98 );
and ( n7884 , n7557 , n7883 );
and ( n7885 , n99 , n7558 );
nor ( n7886 , n7884 , n7885 );
xor ( n7887 , n7571 , n4 );
and ( n7888 , n7886 , n7887 );
not ( n7889 , n7888 );
and ( n7890 , n7882 , n7889 );
not ( n7891 , n7886 );
not ( n7892 , n7887 );
nand ( n7893 , n7891 , n7892 );
not ( n7894 , n7893 );
nor ( n7895 , n7890 , n7894 );
not ( n7896 , n7895 );
nand ( n7897 , n7671 , n7689 );
and ( n7898 , n96 , n71 );
not ( n7899 , n96 );
and ( n7900 , n7899 , n6906 );
nor ( n7901 , n7898 , n7900 );
not ( n7902 , n7681 );
nand ( n7903 , n7901 , n7902 );
and ( n7904 , n7897 , n7903 );
not ( n7905 , n77 );
not ( n7906 , n90 );
and ( n7907 , n7905 , n7906 );
and ( n7908 , n77 , n90 );
nor ( n7909 , n7907 , n7908 );
not ( n7910 , n7909 );
not ( n7911 , n7910 );
not ( n7912 , n6858 );
and ( n7913 , n7911 , n7912 );
not ( n7914 , n6846 );
and ( n7915 , n7592 , n7914 );
nor ( n7916 , n7913 , n7915 );
and ( n7917 , n79 , n88 );
not ( n7918 , n79 );
and ( n7919 , n7918 , n419 );
nor ( n7920 , n7917 , n7919 );
and ( n7921 , n7920 , n7625 );
not ( n7922 , n7728 );
nor ( n7923 , n7922 , n7723 );
nor ( n7924 , n7921 , n7923 );
not ( n7925 , n7924 );
and ( n7926 , n7916 , n7925 );
not ( n7927 , n7916 );
and ( n7928 , n7927 , n7924 );
nor ( n7929 , n7926 , n7928 );
or ( n7930 , n7904 , n7929 );
or ( n7931 , n7916 , n7924 );
nand ( n7932 , n7930 , n7931 );
not ( n7933 , n7932 );
or ( n7934 , n7896 , n7933 );
or ( n7935 , n7895 , n7932 );
nand ( n7936 , n7934 , n7935 );
and ( n7937 , n7870 , n7936 );
not ( n7938 , n7895 );
and ( n7939 , n7938 , n7932 );
nor ( n7940 , n7937 , n7939 );
not ( n7941 , n7940 );
and ( n7942 , n7846 , n7941 );
and ( n7943 , n7845 , n7840 );
nor ( n7944 , n7942 , n7943 );
xor ( n7945 , n7839 , n7944 );
xor ( n7946 , n7764 , n7644 );
nand ( n7947 , n7945 , n7946 );
nand ( n7948 , n7765 , n7947 );
nand ( n7949 , n381 , n7948 );
not ( n7950 , n2663 );
not ( n7951 , n1738 );
nand ( n7952 , n7950 , n7951 );
and ( n7953 , n2 , n7952 );
not ( n7954 , n3700 );
or ( n7955 , n7954 , n2690 );
nand ( n7956 , n7955 , n2633 );
not ( n7957 , n2629 );
not ( n7958 , n2473 );
or ( n7959 , n7957 , n7958 );
nand ( n7960 , n7959 , n2658 );
nor ( n7961 , n7956 , n7960 );
not ( n7962 , n7961 );
nand ( n7963 , n7962 , n3702 );
not ( n7964 , n7963 );
nand ( n7965 , n1 , n7953 , n7964 );
and ( n7966 , n7949 , n7965 );
not ( n7967 , n6530 );
not ( n7968 , n7967 );
not ( n7969 , n6520 );
nor ( n7970 , n7969 , n6508 );
nand ( n7971 , n6293 , n6284 );
nor ( n7972 , n7971 , n6386 );
nand ( n7973 , n7972 , n5445 , n5829 );
nand ( n7974 , n7970 , n7973 );
not ( n7975 , n7974 );
or ( n7976 , n7968 , n7975 );
and ( n7977 , n6521 , n6528 );
nand ( n7978 , n7976 , n7977 );
not ( n7979 , n6523 );
buf ( n7980 , n6497 );
not ( n7981 , n7980 );
nor ( n7982 , n2 , n7979 , n7981 );
nor ( n7983 , n7978 , n7982 );
not ( n7984 , n7983 );
not ( n7985 , n7067 );
not ( n7986 , n7980 );
not ( n7987 , n7986 );
nand ( n7988 , n6523 , n7987 );
not ( n7989 , n7988 );
or ( n7990 , n7985 , n7989 );
nand ( n7991 , n7990 , n7978 );
nand ( n7992 , n7984 , n1 , n7991 );
not ( n7993 , n2653 );
not ( n7994 , n7993 );
nand ( n7995 , n2637 , n7994 );
not ( n7996 , n2668 );
nand ( n7997 , n7995 , n7996 );
not ( n7998 , n7997 );
not ( n7999 , n7998 );
nand ( n8000 , n7953 , n7999 );
not ( n8001 , n8000 );
nor ( n8002 , n7997 , n7952 );
nand ( n8003 , n8002 , n2 , n7963 );
not ( n8004 , n8003 );
or ( n8005 , n8001 , n8004 );
nand ( n8006 , n8005 , n1 );
nand ( n8007 , n7966 , n7992 , n8006 );
and ( n8008 , n7785 , n7204 );
and ( n8009 , n7197 , n7191 );
nor ( n8010 , n8008 , n8009 );
not ( n8011 , n6860 );
not ( n8012 , n7613 );
not ( n8013 , n8012 );
and ( n8014 , n8011 , n8013 );
and ( n8015 , n7317 , n7179 );
nor ( n8016 , n8014 , n8015 );
not ( n8017 , n7679 );
not ( n8018 , n7775 );
not ( n8019 , n8018 );
or ( n8020 , n8017 , n8019 );
nand ( n8021 , n8020 , n96 );
and ( n8022 , n8016 , n8021 );
not ( n8023 , n8016 );
not ( n8024 , n8021 );
and ( n8025 , n8023 , n8024 );
nor ( n8026 , n8022 , n8025 );
xor ( n8027 , n8010 , n8026 );
not ( n8028 , n7634 );
or ( n8029 , n7485 , n8028 );
not ( n8030 , n7616 );
nand ( n8031 , n8030 , n7638 );
nand ( n8032 , n8029 , n8031 );
xor ( n8033 , n8032 , n7797 );
xnor ( n8034 , n8027 , n8033 );
and ( n8035 , n7837 , n7820 );
and ( n8036 , n7798 , n7819 );
nor ( n8037 , n8035 , n8036 );
xnor ( n8038 , n8034 , n8037 );
and ( n8039 , n7542 , n7643 );
and ( n8040 , n7642 , n7607 );
nor ( n8041 , n8039 , n8040 );
xor ( n8042 , n8038 , n8041 );
and ( n8043 , n7807 , n7351 );
and ( n8044 , n7354 , n7215 );
nor ( n8045 , n8043 , n8044 );
not ( n8046 , n7632 );
not ( n8047 , n412 );
or ( n8048 , n8046 , n8047 );
nand ( n8049 , n7728 , n7239 );
nand ( n8050 , n8048 , n8049 );
xor ( n8051 , n7493 , n8050 );
xnor ( n8052 , n8045 , n8051 );
and ( n8053 , n7541 , n7521 );
and ( n8054 , n7526 , n7540 );
nor ( n8055 , n8053 , n8054 );
xnor ( n8056 , n8052 , n8055 );
and ( n8057 , n7809 , n7818 );
not ( n8058 , n308 );
or ( n8059 , n7524 , n8058 );
not ( n8060 , n7322 );
or ( n8061 , n346 , n8060 );
nand ( n8062 , n8059 , n8061 );
and ( n8063 , n7814 , n336 );
and ( n8064 , n327 , n7230 );
nor ( n8065 , n8063 , n8064 );
not ( n8066 , n8065 );
and ( n8067 , n8062 , n8066 );
not ( n8068 , n8062 );
and ( n8069 , n8068 , n8065 );
nor ( n8070 , n8067 , n8069 );
xnor ( n8071 , n8057 , n8070 );
xnor ( n8072 , n8056 , n8071 );
not ( n8073 , n8072 );
or ( n8074 , n7839 , n7944 );
or ( n8075 , n7768 , n7838 );
nand ( n8076 , n8074 , n8075 );
not ( n8077 , n8076 );
or ( n8078 , n8073 , n8077 );
or ( n8079 , n8072 , n8076 );
nand ( n8080 , n8078 , n8079 );
or ( n8081 , n8042 , n8080 );
nand ( n8082 , n8042 , n8080 );
and ( n8083 , n8081 , n381 , n8082 );
nand ( n8084 , n8007 , n8083 );
not ( n8085 , n8084 );
not ( n8086 , n8085 );
buf ( n8087 , n2671 );
not ( n8088 , n8087 );
not ( n8089 , n7961 );
not ( n8090 , n8089 );
or ( n8091 , n8088 , n8090 );
not ( n8092 , n7994 );
nand ( n8093 , n8091 , n8092 );
not ( n8094 , n2637 );
not ( n8095 , n8094 );
nand ( n8096 , n8095 , n7996 );
not ( n8097 , n8096 );
and ( n8098 , n8093 , n8097 );
not ( n8099 , n8093 );
and ( n8100 , n8099 , n8096 );
or ( n8101 , n8098 , n8100 );
nor ( n8102 , n8101 , n7067 );
not ( n8103 , n7067 );
nand ( n8104 , n6521 , n6527 );
not ( n8105 , n8104 );
not ( n8106 , n6451 );
not ( n8107 , n8106 );
not ( n8108 , n7974 );
or ( n8109 , n8107 , n8108 );
nand ( n8110 , n8109 , n6525 );
not ( n8111 , n8110 );
or ( n8112 , n8105 , n8111 );
or ( n8113 , n8104 , n8110 );
nand ( n8114 , n8112 , n8113 );
not ( n8115 , n8114 );
or ( n8116 , n8103 , n8115 );
xor ( n8117 , n7761 , n7702 );
not ( n8118 , n7881 );
not ( n8119 , n7888 );
and ( n8120 , n7893 , n8119 );
not ( n8121 , n8120 );
and ( n8122 , n8118 , n8121 );
and ( n8123 , n7881 , n8120 );
nor ( n8124 , n8122 , n8123 );
not ( n8125 , n8124 );
not ( n8126 , n7904 );
not ( n8127 , n7929 );
not ( n8128 , n8127 );
or ( n8129 , n8126 , n8128 );
or ( n8130 , n7904 , n8127 );
nand ( n8131 , n8129 , n8130 );
not ( n8132 , n8131 );
not ( n8133 , n8132 );
and ( n8134 , n8125 , n8133 );
not ( n8135 , n8131 );
not ( n8136 , n8124 );
or ( n8137 , n8135 , n8136 );
or ( n8138 , n8124 , n8131 );
nand ( n8139 , n8137 , n8138 );
xor ( n8140 , n7867 , n7853 );
and ( n8141 , n8139 , n8140 );
nor ( n8142 , n8134 , n8141 );
not ( n8143 , n5 );
nand ( n8144 , n83 , n302 );
not ( n8145 , n8144 );
not ( n8146 , n8145 );
or ( n8147 , n8143 , n8146 );
and ( n8148 , n98 , n70 );
not ( n8149 , n98 );
and ( n8150 , n8149 , n444 );
nor ( n8151 , n8148 , n8150 );
and ( n8152 , n7557 , n8151 );
and ( n8153 , n99 , n7883 );
nor ( n8154 , n8152 , n8153 );
not ( n8155 , n8154 );
not ( n8156 , n5 );
not ( n8157 , n8144 );
or ( n8158 , n8156 , n8157 );
or ( n8159 , n5 , n8144 );
nand ( n8160 , n8158 , n8159 );
nand ( n8161 , n8155 , n8160 );
nand ( n8162 , n8147 , n8161 );
not ( n8163 , n90 );
and ( n8164 , n7548 , n8163 );
and ( n8165 , n78 , n90 );
nor ( n8166 , n8164 , n8165 );
not ( n8167 , n8166 );
not ( n8168 , n6859 );
or ( n8169 , n8167 , n8168 );
nand ( n8170 , n7909 , n7179 );
nand ( n8171 , n8169 , n8170 );
not ( n8172 , n8171 );
nand ( n8173 , n83 , n87 );
or ( n8174 , n83 , n87 );
nand ( n8175 , n8174 , n88 );
and ( n8176 , n8173 , n86 , n8175 );
and ( n8177 , n6 , n8176 );
and ( n8178 , n96 , n72 );
not ( n8179 , n96 );
and ( n8180 , n8179 , n6954 );
nor ( n8181 , n8178 , n8180 );
not ( n8182 , n8181 );
not ( n8183 , n7682 );
or ( n8184 , n8182 , n8183 );
nand ( n8185 , n7901 , n7689 );
nand ( n8186 , n8184 , n8185 );
xor ( n8187 , n8177 , n8186 );
not ( n8188 , n8187 );
or ( n8189 , n8172 , n8188 );
nand ( n8190 , n8177 , n8186 );
nand ( n8191 , n8189 , n8190 );
xor ( n8192 , n8162 , n8191 );
not ( n8193 , n7875 );
not ( n8194 , n7017 );
and ( n8195 , n8193 , n8194 );
and ( n8196 , n76 , n92 );
nor ( n8197 , n76 , n92 );
nor ( n8198 , n8196 , n8197 );
and ( n8199 , n8198 , n7351 );
nor ( n8200 , n8195 , n8199 );
and ( n8201 , n82 , n86 );
not ( n8202 , n82 );
and ( n8203 , n8202 , n358 );
nor ( n8204 , n8201 , n8203 );
buf ( n8205 , n333 );
and ( n8206 , n8204 , n8205 );
not ( n8207 , n323 );
and ( n8208 , n8207 , n7854 );
nor ( n8209 , n8206 , n8208 );
and ( n8210 , n74 , n94 );
nor ( n8211 , n74 , n94 );
nor ( n8212 , n8210 , n8211 );
not ( n8213 , n8212 );
not ( n8214 , n7204 );
or ( n8215 , n8213 , n8214 );
nand ( n8216 , n7850 , n7189 );
nand ( n8217 , n8215 , n8216 );
xor ( n8218 , n8209 , n8217 );
or ( n8219 , n8200 , n8218 );
not ( n8220 , n8217 );
or ( n8221 , n8220 , n8209 );
nand ( n8222 , n8219 , n8221 );
and ( n8223 , n8192 , n8222 );
and ( n8224 , n8162 , n8191 );
nor ( n8225 , n8223 , n8224 );
xnor ( n8226 , n8142 , n8225 );
xnor ( n8227 , n7936 , n7870 );
or ( n8228 , n8226 , n8227 );
or ( n8229 , n8225 , n8142 );
nand ( n8230 , n8228 , n8229 );
and ( n8231 , n7846 , n7941 );
not ( n8232 , n7846 );
and ( n8233 , n8232 , n7940 );
nor ( n8234 , n8231 , n8233 );
xor ( n8235 , n8230 , n8234 );
and ( n8236 , n8117 , n8235 );
and ( n8237 , n8234 , n8230 );
nor ( n8238 , n8236 , n8237 );
nor ( n8239 , n1 , n8238 );
not ( n8240 , n8239 );
nand ( n8241 , n8116 , n8240 );
or ( n8242 , n8102 , n8241 );
not ( n8243 , n7945 );
not ( n8244 , n7946 );
nand ( n8245 , n8243 , n8244 );
and ( n8246 , n8245 , n381 , n7947 );
nand ( n8247 , n8242 , n8246 );
and ( n8248 , n381 , n8240 );
nor ( n8249 , n8247 , n8248 );
not ( n8250 , n8249 );
buf ( n8251 , n8139 );
xnor ( n8252 , n8140 , n8251 );
nand ( n8253 , n325 , n8204 );
not ( n8254 , n83 );
or ( n8255 , n8254 , n358 );
or ( n8256 , n83 , n86 );
nand ( n8257 , n8255 , n8256 , n335 );
and ( n8258 , n8253 , n8257 );
not ( n8259 , n99 );
nand ( n8260 , n8259 , n98 );
not ( n8261 , n8260 );
not ( n8262 , n8261 );
not ( n8263 , n8262 );
and ( n8264 , n98 , n6906 );
not ( n8265 , n98 );
and ( n8266 , n8265 , n71 );
nor ( n8267 , n8264 , n8266 );
not ( n8268 , n8267 );
and ( n8269 , n8263 , n8268 );
and ( n8270 , n99 , n8151 );
nor ( n8271 , n8269 , n8270 );
xor ( n8272 , n6 , n8176 );
and ( n8273 , n8271 , n8272 );
not ( n8274 , n8271 );
not ( n8275 , n8272 );
and ( n8276 , n8274 , n8275 );
nor ( n8277 , n8273 , n8276 );
xor ( n8278 , n8258 , n8277 );
not ( n8279 , n8278 );
not ( n8280 , n8 );
nand ( n8281 , n83 , n89 );
or ( n8282 , n83 , n89 );
nand ( n8283 , n8282 , n90 );
nand ( n8284 , n8281 , n88 , n8283 );
or ( n8285 , n8280 , n8284 );
not ( n8286 , n8285 );
xnor ( n8287 , n94 , n76 );
not ( n8288 , n8287 );
not ( n8289 , n8288 );
not ( n8290 , n7204 );
or ( n8291 , n8289 , n8290 );
not ( n8292 , n75 );
not ( n8293 , n94 );
and ( n8294 , n8292 , n8293 );
and ( n8295 , n75 , n94 );
nor ( n8296 , n8294 , n8295 );
nand ( n8297 , n8296 , n7189 );
nand ( n8298 , n8291 , n8297 );
nand ( n8299 , n8286 , n8298 );
not ( n8300 , n7353 );
not ( n8301 , n77 );
not ( n8302 , n92 );
and ( n8303 , n8301 , n8302 );
and ( n8304 , n77 , n92 );
nor ( n8305 , n8303 , n8304 );
not ( n8306 , n8305 );
not ( n8307 , n8306 );
and ( n8308 , n8300 , n8307 );
and ( n8309 , n92 , n78 );
not ( n8310 , n92 );
and ( n8311 , n8310 , n7548 );
nor ( n8312 , n8309 , n8311 );
and ( n8313 , n8312 , n7025 );
nor ( n8314 , n8308 , n8313 );
not ( n8315 , n8314 );
not ( n8316 , n8298 );
nand ( n8317 , n8316 , n8285 );
nand ( n8318 , n8315 , n8317 );
nand ( n8319 , n8299 , n8318 );
and ( n8320 , n98 , n6954 );
not ( n8321 , n98 );
and ( n8322 , n8321 , n72 );
nor ( n8323 , n8320 , n8322 );
or ( n8324 , n8262 , n8323 );
or ( n8325 , n7555 , n8267 );
nand ( n8326 , n8324 , n8325 );
and ( n8327 , n83 , n322 );
and ( n8328 , n8327 , n7 );
not ( n8329 , n8327 );
and ( n8330 , n8329 , n2401 );
nor ( n8331 , n8328 , n8330 );
and ( n8332 , n8326 , n8331 );
and ( n8333 , n7 , n8327 );
nor ( n8334 , n8332 , n8333 );
xnor ( n8335 , n8319 , n8334 );
not ( n8336 , n8335 );
or ( n8337 , n8279 , n8336 );
not ( n8338 , n8319 );
or ( n8339 , n8334 , n8338 );
nand ( n8340 , n8337 , n8339 );
not ( n8341 , n79 );
not ( n8342 , n90 );
and ( n8343 , n8341 , n8342 );
and ( n8344 , n79 , n90 );
nor ( n8345 , n8343 , n8344 );
and ( n8346 , n8345 , n7594 );
and ( n8347 , n8166 , n6847 );
nor ( n8348 , n8346 , n8347 );
and ( n8349 , n81 , n88 );
nor ( n8350 , n81 , n88 );
nor ( n8351 , n8349 , n8350 );
not ( n8352 , n413 );
and ( n8353 , n8351 , n8352 );
not ( n8354 , n80 );
and ( n8355 , n8354 , n419 );
and ( n8356 , n80 , n88 );
nor ( n8357 , n8355 , n8356 );
and ( n8358 , n401 , n8357 );
nor ( n8359 , n8353 , n8358 );
xor ( n8360 , n8348 , n8359 );
not ( n8361 , n8360 );
not ( n8362 , n80 );
not ( n8363 , n90 );
and ( n8364 , n8362 , n8363 );
and ( n8365 , n80 , n90 );
nor ( n8366 , n8364 , n8365 );
and ( n8367 , n8366 , n6863 );
and ( n8368 , n8345 , n6851 );
nor ( n8369 , n8367 , n8368 );
and ( n8370 , n96 , n73 );
not ( n8371 , n96 );
and ( n8372 , n8371 , n7508 );
nor ( n8373 , n8370 , n8372 );
nand ( n8374 , n8373 , n7689 );
not ( n8375 , n74 );
not ( n8376 , n96 );
and ( n8377 , n8375 , n8376 );
and ( n8378 , n74 , n96 );
nor ( n8379 , n8377 , n8378 );
nand ( n8380 , n8379 , n7682 );
and ( n8381 , n8374 , n8380 );
not ( n8382 , n82 );
and ( n8383 , n8382 , n419 );
and ( n8384 , n82 , n88 );
nor ( n8385 , n8383 , n8384 );
and ( n8386 , n8385 , n7625 );
and ( n8387 , n401 , n8351 );
nor ( n8388 , n8386 , n8387 );
xnor ( n8389 , n8381 , n8388 );
or ( n8390 , n8369 , n8389 );
or ( n8391 , n8381 , n8388 );
nand ( n8392 , n8390 , n8391 );
not ( n8393 , n8392 );
or ( n8394 , n8361 , n8393 );
or ( n8395 , n8348 , n8359 );
nand ( n8396 , n8394 , n8395 );
xor ( n8397 , n8340 , n8396 );
and ( n8398 , n8373 , n7902 );
and ( n8399 , n8181 , n7689 );
nor ( n8400 , n8398 , n8399 );
not ( n8401 , n8296 );
not ( n8402 , n7204 );
or ( n8403 , n8401 , n8402 );
nand ( n8404 , n8212 , n7786 );
nand ( n8405 , n8403 , n8404 );
not ( n8406 , n8405 );
and ( n8407 , n8305 , n7513 );
not ( n8408 , n7015 );
and ( n8409 , n8408 , n8198 );
nor ( n8410 , n8407 , n8409 );
xnor ( n8411 , n8406 , n8410 );
or ( n8412 , n8400 , n8411 );
or ( n8413 , n8406 , n8410 );
nand ( n8414 , n8412 , n8413 );
not ( n8415 , n8357 );
not ( n8416 , n414 );
or ( n8417 , n8415 , n8416 );
not ( n8418 , n404 );
nand ( n8419 , n8418 , n7920 );
nand ( n8420 , n8417 , n8419 );
xor ( n8421 , n8414 , n8420 );
not ( n8422 , n8154 );
not ( n8423 , n8160 );
or ( n8424 , n8422 , n8423 );
or ( n8425 , n8154 , n8160 );
nand ( n8426 , n8424 , n8425 );
xor ( n8427 , n8421 , n8426 );
and ( n8428 , n8397 , n8427 );
and ( n8429 , n8396 , n8340 );
nor ( n8430 , n8428 , n8429 );
or ( n8431 , n8252 , n8430 );
and ( n8432 , n8192 , n8222 );
not ( n8433 , n8192 );
not ( n8434 , n8222 );
and ( n8435 , n8433 , n8434 );
nor ( n8436 , n8432 , n8435 );
xnor ( n8437 , n8187 , n8171 );
not ( n8438 , n8437 );
xnor ( n8439 , n8200 , n8218 );
not ( n8440 , n8439 );
nand ( n8441 , n8438 , n8440 );
not ( n8442 , n8437 );
not ( n8443 , n8439 );
or ( n8444 , n8442 , n8443 );
or ( n8445 , n8258 , n8277 );
or ( n8446 , n8271 , n8275 );
nand ( n8447 , n8445 , n8446 );
nand ( n8448 , n8444 , n8447 );
nand ( n8449 , n8441 , n8448 );
xor ( n8450 , n8436 , n8449 );
xor ( n8451 , n8414 , n8420 );
and ( n8452 , n8451 , n8426 );
and ( n8453 , n8414 , n8420 );
or ( n8454 , n8452 , n8453 );
xor ( n8455 , n8450 , n8454 );
xor ( n8456 , n8430 , n8252 );
nand ( n8457 , n8455 , n8456 );
nand ( n8458 , n8431 , n8457 );
nand ( n8459 , n381 , n8458 );
not ( n8460 , n7971 );
not ( n8461 , n8460 );
not ( n8462 , n5445 );
or ( n8463 , n8461 , n8462 );
nand ( n8464 , n6518 , n6293 );
nand ( n8465 , n8463 , n8464 );
not ( n8466 , n5830 );
nand ( n8467 , n8465 , n8466 );
not ( n8468 , n6503 );
not ( n8469 , n8468 );
not ( n8470 , n8469 );
and ( n8471 , n8467 , n8470 );
not ( n8472 , n6387 );
not ( n8473 , n8472 );
nand ( n8474 , n8473 , n6507 );
nand ( n8475 , n7067 , n8474 );
nor ( n8476 , n8471 , n8475 );
not ( n8477 , n8476 );
not ( n8478 , n2657 );
not ( n8479 , n8478 );
not ( n8480 , n2689 );
not ( n8481 , n8480 );
not ( n8482 , n2688 );
not ( n8483 , n3700 );
or ( n8484 , n8482 , n8483 );
not ( n8485 , n2474 );
not ( n8486 , n2686 );
nor ( n8487 , n8486 , n2478 );
not ( n8488 , n8487 );
nand ( n8489 , n8485 , n8488 );
not ( n8490 , n2472 );
nand ( n8491 , n8489 , n8490 );
nand ( n8492 , n8484 , n8491 );
nand ( n8493 , n8481 , n8492 );
not ( n8494 , n8493 );
or ( n8495 , n8479 , n8494 );
not ( n8496 , n2656 );
not ( n8497 , n2633 );
nor ( n8498 , n8496 , n8497 );
nor ( n8499 , n7067 , n8498 );
nand ( n8500 , n8495 , n8499 );
nand ( n8501 , n8477 , n8500 );
nor ( n8502 , n8474 , n8469 );
nand ( n8503 , n8502 , n7067 , n8467 );
and ( n8504 , n2 , n8478 );
nand ( n8505 , n8504 , n8493 , n8498 );
nand ( n8506 , n8503 , n8505 );
or ( n8507 , n8501 , n8506 );
nand ( n8508 , n8507 , n1 );
and ( n8509 , n8459 , n8508 );
xnor ( n8510 , n8226 , n8227 );
xor ( n8511 , n8436 , n8449 );
and ( n8512 , n8511 , n8454 );
and ( n8513 , n8436 , n8449 );
or ( n8514 , n8512 , n8513 );
and ( n8515 , n7745 , n7757 , n7739 );
nor ( n8516 , n7757 , n7740 , n7745 );
nor ( n8517 , n8515 , n8516 );
and ( n8518 , n7757 , n7740 , n7746 );
nor ( n8519 , n7757 , n7739 , n7746 );
nor ( n8520 , n8518 , n8519 );
nand ( n8521 , n8517 , n8520 );
xnor ( n8522 , n8514 , n8521 );
or ( n8523 , n8510 , n8522 );
and ( n8524 , n8510 , n8522 );
nor ( n8525 , n8524 , n1 );
nand ( n8526 , n8523 , n8525 );
nor ( n8527 , n8509 , n8526 );
not ( n8528 , n8527 );
and ( n8529 , n8521 , n8514 );
nor ( n8530 , n8510 , n8522 );
nor ( n8531 , n8529 , n8530 );
nor ( n8532 , n8531 , n1 );
not ( n8533 , n8532 );
not ( n8534 , n6451 );
nand ( n8535 , n8534 , n6525 );
not ( n8536 , n8535 );
not ( n8537 , n7974 );
or ( n8538 , n8536 , n8537 );
or ( n8539 , n8535 , n7974 );
nand ( n8540 , n8538 , n8539 );
nand ( n8541 , n8540 , n7067 );
not ( n8542 , n8541 );
nand ( n8543 , n7993 , n8087 );
not ( n8544 , n8543 );
not ( n8545 , n8544 );
not ( n8546 , n8089 );
or ( n8547 , n8545 , n8546 );
and ( n8548 , n7961 , n8543 );
nor ( n8549 , n8548 , n7067 );
nand ( n8550 , n8547 , n8549 );
not ( n8551 , n8550 );
or ( n8552 , n8542 , n8551 );
nand ( n8553 , n8552 , n1 );
not ( n8554 , n8117 );
not ( n8555 , n8235 );
or ( n8556 , n8554 , n8555 );
not ( n8557 , n8117 );
not ( n8558 , n8235 );
and ( n8559 , n8557 , n8558 );
nor ( n8560 , n8559 , n1 );
nand ( n8561 , n8556 , n8560 );
nand ( n8562 , n8533 , n8553 , n8561 );
not ( n8563 , n8562 );
or ( n8564 , n8528 , n8563 );
not ( n8565 , n8553 );
or ( n8566 , n8565 , n8532 );
not ( n8567 , n8561 );
nand ( n8568 , n8566 , n8567 );
nand ( n8569 , n8564 , n8568 );
not ( n8570 , n1 );
not ( n8571 , n7067 );
not ( n8572 , n8104 );
not ( n8573 , n8110 );
or ( n8574 , n8572 , n8573 );
or ( n8575 , n8104 , n8110 );
nand ( n8576 , n8574 , n8575 );
not ( n8577 , n8576 );
or ( n8578 , n8571 , n8577 );
nand ( n8579 , n8097 , n8093 );
not ( n8580 , n8093 );
and ( n8581 , n8580 , n8096 );
nor ( n8582 , n8581 , n7067 );
nand ( n8583 , n8579 , n8582 );
nand ( n8584 , n8578 , n8583 );
not ( n8585 , n8584 );
or ( n8586 , n8570 , n8585 );
nor ( n8587 , n8239 , n8246 );
nand ( n8588 , n8586 , n8587 );
nand ( n8589 , n8569 , n8588 );
nand ( n8590 , n8086 , n8250 , n8589 );
not ( n8591 , n8083 );
nand ( n8592 , n7992 , n8006 , n7966 , n8591 );
not ( n8593 , n2 );
not ( n8594 , n4044 );
nand ( n8595 , n4050 , n8594 );
not ( n8596 , n8595 );
not ( n8597 , n7132 );
or ( n8598 , n8596 , n8597 );
or ( n8599 , n8595 , n3705 );
nand ( n8600 , n8598 , n8599 );
not ( n8601 , n8600 );
or ( n8602 , n8593 , n8601 );
nand ( n8603 , n6792 , n6707 );
xor ( n8604 , n6537 , n8603 );
nand ( n8605 , n8604 , n7067 );
nand ( n8606 , n8602 , n8605 );
nand ( n8607 , n8606 , n1 );
or ( n8608 , n8071 , n8056 );
or ( n8609 , n8052 , n8055 );
nand ( n8610 , n8608 , n8609 );
or ( n8611 , n8026 , n8010 );
or ( n8612 , n8024 , n8016 );
nand ( n8613 , n8611 , n8612 );
or ( n8614 , n8045 , n8051 );
not ( n8615 , n8050 );
or ( n8616 , n7493 , n8615 );
nand ( n8617 , n8614 , n8616 );
xor ( n8618 , n7206 , n8617 );
xor ( n8619 , n8613 , n8618 );
and ( n8620 , n8027 , n8033 );
and ( n8621 , n7797 , n8032 );
nor ( n8622 , n8620 , n8621 );
not ( n8623 , n8622 );
and ( n8624 , n8619 , n8623 );
not ( n8625 , n8619 );
and ( n8626 , n8625 , n8622 );
nor ( n8627 , n8624 , n8626 );
and ( n8628 , n8610 , n8627 );
and ( n8629 , n8623 , n8619 );
nor ( n8630 , n8628 , n8629 );
xnor ( n8631 , n7320 , n7332 );
not ( n8632 , n8631 );
and ( n8633 , n7252 , n7223 );
not ( n8634 , n7252 );
and ( n8635 , n8634 , n7224 );
nor ( n8636 , n8633 , n8635 );
not ( n8637 , n8636 );
and ( n8638 , n8632 , n8637 );
and ( n8639 , n8631 , n8636 );
and ( n8640 , n8057 , n8070 );
and ( n8641 , n8062 , n8066 );
nor ( n8642 , n8640 , n8641 );
nor ( n8643 , n8639 , n8642 );
nor ( n8644 , n8638 , n8643 );
not ( n8645 , n7283 );
and ( n8646 , n7336 , n8645 );
not ( n8647 , n7336 );
and ( n8648 , n8647 , n7283 );
nor ( n8649 , n8646 , n8648 );
and ( n8650 , n8613 , n8618 );
and ( n8651 , n7206 , n8617 );
nor ( n8652 , n8650 , n8651 );
xnor ( n8653 , n7211 , n7257 );
not ( n8654 , n8653 );
and ( n8655 , n8652 , n8654 );
not ( n8656 , n8652 );
and ( n8657 , n8656 , n8653 );
nor ( n8658 , n8655 , n8657 );
xnor ( n8659 , n8649 , n8658 );
nor ( n8660 , n8644 , n8659 );
not ( n8661 , n8660 );
nand ( n8662 , n8644 , n8659 );
nand ( n8663 , n8661 , n8662 );
and ( n8664 , n8630 , n8663 );
or ( n8665 , n8663 , n8630 );
nand ( n8666 , n8665 , n381 );
nor ( n8667 , n8664 , n8666 );
not ( n8668 , n8667 );
nand ( n8669 , n8607 , n8668 );
xor ( n8670 , n8627 , n8610 );
or ( n8671 , n8038 , n8041 );
or ( n8672 , n8037 , n8034 );
nand ( n8673 , n8671 , n8672 );
xor ( n8674 , n8631 , n8642 );
xnor ( n8675 , n8636 , n8674 );
and ( n8676 , n8673 , n8675 );
not ( n8677 , n8673 );
not ( n8678 , n8675 );
and ( n8679 , n8677 , n8678 );
nor ( n8680 , n8676 , n8679 );
and ( n8681 , n8670 , n8680 );
and ( n8682 , n8675 , n8673 );
nor ( n8683 , n8681 , n8682 );
nor ( n8684 , n1 , n8683 );
nor ( n8685 , n8669 , n8684 );
not ( n8686 , n8685 );
nor ( n8687 , n381 , n7067 );
not ( n8688 , n8687 );
not ( n8689 , n1864 );
nand ( n8690 , n8689 , n2681 );
nor ( n8691 , n8688 , n8690 );
not ( n8692 , n8691 );
and ( n8693 , n7963 , n7998 );
buf ( n8694 , n2663 );
nor ( n8695 , n8693 , n8694 );
not ( n8696 , n7951 );
nor ( n8697 , n8695 , n8696 );
not ( n8698 , n8697 );
or ( n8699 , n8692 , n8698 );
nor ( n8700 , n381 , n2 );
nand ( n8701 , n6522 , n6259 );
not ( n8702 , n8701 );
not ( n8703 , n7967 );
nor ( n8704 , n8703 , n7986 );
nand ( n8705 , n7974 , n8704 );
not ( n8706 , n7977 );
and ( n8707 , n8706 , n7987 );
nor ( n8708 , n8707 , n7979 );
nand ( n8709 , n8700 , n8702 , n8705 , n8708 );
nand ( n8710 , n8699 , n8709 );
not ( n8711 , n8710 );
not ( n8712 , n8670 );
not ( n8713 , n8680 );
or ( n8714 , n8712 , n8713 );
not ( n8715 , n8670 );
not ( n8716 , n8680 );
and ( n8717 , n8715 , n8716 );
nor ( n8718 , n8717 , n1 );
nand ( n8719 , n8714 , n8718 );
nand ( n8720 , n2 , n8690 );
not ( n8721 , n8720 );
not ( n8722 , n8697 );
nand ( n8723 , n8721 , n8722 , n1 );
nor ( n8724 , n381 , n2 );
nand ( n8725 , n8705 , n8708 );
nand ( n8726 , n8724 , n8725 , n8701 );
not ( n8727 , n8076 );
or ( n8728 , n8072 , n8727 );
nand ( n8729 , n8728 , n8082 );
nand ( n8730 , n381 , n8729 );
nand ( n8731 , n8726 , n8730 );
not ( n8732 , n8731 );
nand ( n8733 , n8711 , n8719 , n8723 , n8732 );
nand ( n8734 , n8686 , n8733 );
xnor ( n8735 , n7392 , n7382 );
xnor ( n8736 , n7340 , n7261 );
and ( n8737 , n8735 , n8736 );
not ( n8738 , n8735 );
not ( n8739 , n8736 );
and ( n8740 , n8738 , n8739 );
or ( n8741 , n8649 , n8658 );
not ( n8742 , n8654 );
or ( n8743 , n8742 , n8652 );
nand ( n8744 , n8741 , n8743 );
nor ( n8745 , n8740 , n8744 );
nor ( n8746 , n8737 , n1 , n8745 );
and ( n8747 , n7343 , n7396 );
or ( n8748 , n7343 , n7396 );
nand ( n8749 , n8748 , n381 );
nor ( n8750 , n8747 , n8749 );
nor ( n8751 , n8746 , n8750 );
not ( n8752 , n8751 );
and ( n8753 , n6799 , n6777 );
nor ( n8754 , n2 , n8753 );
nand ( n8755 , n8754 , n6795 );
not ( n8756 , n6795 );
nand ( n8757 , n7067 , n8753 , n8756 );
nand ( n8758 , n8755 , n7152 , n8757 );
not ( n8759 , n8758 );
not ( n8760 , n8754 );
nand ( n8761 , n7156 , n8760 );
not ( n8762 , n8761 );
or ( n8763 , n8759 , n8762 );
nand ( n8764 , n4057 , n3992 );
not ( n8765 , n8764 );
not ( n8766 , n4045 );
not ( n8767 , n3704 );
or ( n8768 , n8766 , n8767 );
not ( n8769 , n4053 );
nand ( n8770 , n8768 , n8769 );
not ( n8771 , n8770 );
or ( n8772 , n8765 , n8771 );
or ( n8773 , n8770 , n8764 );
nand ( n8774 , n8772 , n8773 );
nand ( n8775 , n2 , n8774 );
nand ( n8776 , n8763 , n8775 );
nand ( n8777 , n1 , n8776 );
not ( n8778 , n8777 );
or ( n8779 , n8752 , n8778 );
and ( n8780 , n8594 , n3705 );
not ( n8781 , n4050 );
nor ( n8782 , n8780 , n8781 );
not ( n8783 , n8782 );
nor ( n8784 , n381 , n7067 );
not ( n8785 , n4052 );
nor ( n8786 , n8785 , n4036 );
not ( n8787 , n8786 );
and ( n8788 , n8783 , n8784 , n8787 );
not ( n8789 , n8630 );
or ( n8790 , n8789 , n8660 );
nand ( n8791 , n8790 , n381 , n8662 );
not ( n8792 , n8735 );
not ( n8793 , n8744 );
and ( n8794 , n8792 , n8793 );
and ( n8795 , n8735 , n8744 );
nor ( n8796 , n8794 , n8795 );
or ( n8797 , n8736 , n8796 );
and ( n8798 , n8736 , n8796 );
nor ( n8799 , n8798 , n1 );
nand ( n8800 , n8797 , n8799 );
nand ( n8801 , n8791 , n8800 );
nor ( n8802 , n8788 , n8801 );
not ( n8803 , n6707 );
not ( n8804 , n6536 );
or ( n8805 , n8803 , n8804 );
nand ( n8806 , n8805 , n6792 );
nand ( n8807 , n6794 , n6697 );
nand ( n8808 , n7067 , n8806 , n8807 );
nand ( n8809 , n2 , n8782 , n8786 );
nand ( n8810 , n8808 , n8809 );
not ( n8811 , n8806 );
not ( n8812 , n8807 );
and ( n8813 , n7067 , n8811 , n8812 );
or ( n8814 , n8810 , n8813 );
nand ( n8815 , n8814 , n1 );
nand ( n8816 , n8802 , n8815 );
nand ( n8817 , n8779 , n8816 );
nor ( n8818 , n8734 , n8817 );
nand ( n8819 , n8590 , n8592 , n8818 );
not ( n8820 , n8819 );
not ( n8821 , n8720 );
nand ( n8822 , n8821 , n1 , n8722 );
nand ( n8823 , n8822 , n8732 );
or ( n8824 , n8823 , n8710 );
not ( n8825 , n8719 );
nand ( n8826 , n8824 , n8825 );
not ( n8827 , n8684 );
and ( n8828 , n8827 , n8607 , n8668 );
or ( n8829 , n8826 , n8828 );
not ( n8830 , n8607 );
or ( n8831 , n8830 , n8667 );
nand ( n8832 , n8831 , n8684 );
nand ( n8833 , n8829 , n8832 );
not ( n8834 , n8833 );
buf ( n8835 , n8817 );
or ( n8836 , n8834 , n8835 );
nor ( n8837 , n8791 , n8800 );
not ( n8838 , n8837 );
nand ( n8839 , n8751 , n8777 );
not ( n8840 , n8839 );
or ( n8841 , n8838 , n8840 );
not ( n8842 , n8746 );
not ( n8843 , n8842 );
not ( n8844 , n8777 );
or ( n8845 , n8843 , n8844 );
nand ( n8846 , n8845 , n8750 );
nand ( n8847 , n8841 , n8846 );
not ( n8848 , n8847 );
nand ( n8849 , n8836 , n8848 );
nor ( n8850 , n8820 , n8849 );
not ( n8851 , n8818 );
not ( n8852 , n8851 );
not ( n8853 , n8447 );
not ( n8854 , n8437 );
or ( n8855 , n8853 , n8854 );
or ( n8856 , n8447 , n8437 );
nand ( n8857 , n8855 , n8856 );
xor ( n8858 , n8439 , n8857 );
xor ( n8859 , n8411 , n8400 );
not ( n8860 , n8859 );
not ( n8861 , n8860 );
not ( n8862 , n96 );
and ( n8863 , n7871 , n8862 );
and ( n8864 , n75 , n96 );
nor ( n8865 , n8863 , n8864 );
not ( n8866 , n8018 );
and ( n8867 , n8865 , n8866 );
and ( n8868 , n8379 , n7689 );
nor ( n8869 , n8867 , n8868 );
xor ( n8870 , n81 , n90 );
and ( n8871 , n8870 , n7594 );
not ( n8872 , n6846 );
and ( n8873 , n8366 , n8872 );
nor ( n8874 , n8871 , n8873 );
and ( n8875 , n79 , n92 );
nor ( n8876 , n79 , n92 );
nor ( n8877 , n8875 , n8876 );
not ( n8878 , n7512 );
and ( n8879 , n8877 , n8878 );
and ( n8880 , n7014 , n8312 );
nor ( n8881 , n8879 , n8880 );
xnor ( n8882 , n8874 , n8881 );
or ( n8883 , n8869 , n8882 );
or ( n8884 , n8874 , n8881 );
nand ( n8885 , n8883 , n8884 );
xor ( n8886 , n8326 , n8331 );
and ( n8887 , n94 , n77 );
not ( n8888 , n94 );
and ( n8889 , n8888 , n7811 );
nor ( n8890 , n8887 , n8889 );
not ( n8891 , n8890 );
not ( n8892 , n7204 );
or ( n8893 , n8891 , n8892 );
or ( n8894 , n8287 , n7190 );
nand ( n8895 , n8893 , n8894 );
not ( n8896 , n8895 );
and ( n8897 , n8284 , n8280 );
not ( n8898 , n8284 );
and ( n8899 , n8898 , n8 );
nor ( n8900 , n8897 , n8899 );
and ( n8901 , n98 , n7508 );
not ( n8902 , n98 );
and ( n8903 , n8902 , n73 );
nor ( n8904 , n8901 , n8903 );
or ( n8905 , n8262 , n8904 );
or ( n8906 , n7555 , n8323 );
nand ( n8907 , n8905 , n8906 );
xor ( n8908 , n8900 , n8907 );
not ( n8909 , n8908 );
or ( n8910 , n8896 , n8909 );
nand ( n8911 , n8907 , n8900 );
nand ( n8912 , n8910 , n8911 );
xor ( n8913 , n8886 , n8912 );
and ( n8914 , n8885 , n8913 );
and ( n8915 , n8886 , n8912 );
nor ( n8916 , n8914 , n8915 );
not ( n8917 , n8916 );
and ( n8918 , n8861 , n8917 );
xor ( n8919 , n8392 , n8360 );
not ( n8920 , n8859 );
not ( n8921 , n8916 );
or ( n8922 , n8920 , n8921 );
or ( n8923 , n8859 , n8916 );
nand ( n8924 , n8922 , n8923 );
and ( n8925 , n8919 , n8924 );
nor ( n8926 , n8918 , n8925 );
or ( n8927 , n8858 , n8926 );
xnor ( n8928 , n8397 , n8427 );
xnor ( n8929 , n8926 , n8858 );
nor ( n8930 , n8928 , n8929 );
not ( n8931 , n8930 );
nand ( n8932 , n8927 , n8931 );
nand ( n8933 , n381 , n8932 );
not ( n8934 , n8933 );
not ( n8935 , n8480 );
nand ( n8936 , n8935 , n8478 );
not ( n8937 , n8936 );
and ( n8938 , n8937 , n8492 );
not ( n8939 , n8936 );
not ( n8940 , n8492 );
not ( n8941 , n8940 );
or ( n8942 , n8939 , n8941 );
nand ( n8943 , n8942 , n2 );
or ( n8944 , n8938 , n8943 );
not ( n8945 , n5830 );
nand ( n8946 , n8945 , n8468 );
xnor ( n8947 , n8465 , n8946 );
nand ( n8948 , n7067 , n8947 );
nand ( n8949 , n8944 , n8948 );
nand ( n8950 , n1 , n8949 );
not ( n8951 , n8950 );
or ( n8952 , n8934 , n8951 );
not ( n8953 , n1 );
not ( n8954 , n84 );
or ( n8955 , n8953 , n8954 );
or ( n8956 , n8455 , n8456 );
nand ( n8957 , n8956 , n381 , n8457 );
nand ( n8958 , n8955 , n8957 );
nand ( n8959 , n8952 , n8958 );
not ( n8960 , n8959 );
not ( n8961 , n8960 );
not ( n8962 , n3677 );
not ( n8963 , n8962 );
not ( n8964 , n3505 );
not ( n8965 , n8964 );
not ( n8966 , n8965 );
or ( n8967 , n8963 , n8966 );
not ( n8968 , n3688 );
nand ( n8969 , n8967 , n8968 );
not ( n8970 , n8969 );
not ( n8971 , n3606 );
or ( n8972 , n8970 , n8971 );
not ( n8973 , n3693 );
not ( n8974 , n8973 );
nand ( n8975 , n8972 , n8974 );
not ( n8976 , n8975 );
nand ( n8977 , n3697 , n3619 );
not ( n8978 , n8977 );
not ( n8979 , n8978 );
or ( n8980 , n8976 , n8979 );
not ( n8981 , n8975 );
and ( n8982 , n8981 , n8977 );
nor ( n8983 , n8982 , n8688 );
nand ( n8984 , n8980 , n8983 );
not ( n8985 , n8984 );
not ( n8986 , n4659 );
nor ( n8987 , n4985 , n5425 );
not ( n8988 , n8987 );
buf ( n8989 , n5418 );
not ( n8990 , n8989 );
or ( n8991 , n8988 , n8990 );
not ( n8992 , n5437 );
nand ( n8993 , n8991 , n8992 );
not ( n8994 , n8993 );
or ( n8995 , n8986 , n8994 );
nand ( n8996 , n8995 , n5442 );
nor ( n8997 , n5430 , n5439 );
nor ( n8998 , n8996 , n8997 );
not ( n8999 , n8998 );
nor ( n9000 , n381 , n2 );
nand ( n9001 , n8996 , n8997 );
nand ( n9002 , n8999 , n9000 , n9001 );
not ( n9003 , n9002 );
nor ( n9004 , n8985 , n9003 );
and ( n9005 , n8354 , n7212 );
and ( n9006 , n80 , n92 );
nor ( n9007 , n9005 , n9006 );
and ( n9008 , n9007 , n7025 );
and ( n9009 , n7014 , n8877 );
nor ( n9010 , n9008 , n9009 );
and ( n9011 , n94 , n78 );
not ( n9012 , n94 );
and ( n9013 , n9012 , n7548 );
nor ( n9014 , n9011 , n9013 );
not ( n9015 , n9014 );
not ( n9016 , n9015 );
not ( n9017 , n7203 );
and ( n9018 , n9016 , n9017 );
and ( n9019 , n8890 , n7786 );
nor ( n9020 , n9018 , n9019 );
nand ( n9021 , n83 , n91 );
or ( n9022 , n83 , n91 );
nand ( n9023 , n9022 , n92 );
nand ( n9024 , n9021 , n90 , n9023 );
not ( n9025 , n9024 );
nand ( n9026 , n9025 , n10 );
not ( n9027 , n9026 );
and ( n9028 , n9020 , n9027 );
not ( n9029 , n9020 );
and ( n9030 , n9029 , n9026 );
nor ( n9031 , n9028 , n9030 );
or ( n9032 , n9010 , n9031 );
or ( n9033 , n9026 , n9020 );
nand ( n9034 , n9032 , n9033 );
not ( n9035 , n9 );
nand ( n9036 , n83 , n7728 );
not ( n9037 , n9036 );
not ( n9038 , n9037 );
or ( n9039 , n9035 , n9038 );
not ( n9040 , n7555 );
not ( n9041 , n8904 );
and ( n9042 , n9040 , n9041 );
and ( n9043 , n98 , n74 );
not ( n9044 , n98 );
and ( n9045 , n9044 , n7535 );
nor ( n9046 , n9043 , n9045 );
and ( n9047 , n7557 , n9046 );
nor ( n9048 , n9042 , n9047 );
not ( n9049 , n9 );
not ( n9050 , n9036 );
and ( n9051 , n9049 , n9050 );
and ( n9052 , n9 , n9036 );
nor ( n9053 , n9051 , n9052 );
or ( n9054 , n9048 , n9053 );
nand ( n9055 , n9039 , n9054 );
not ( n9056 , n403 );
not ( n9057 , n8385 );
or ( n9058 , n9056 , n9057 );
or ( n9059 , n8254 , n419 );
or ( n9060 , n83 , n88 );
nand ( n9061 , n9059 , n9060 , n412 );
nand ( n9062 , n9058 , n9061 );
xor ( n9063 , n9055 , n9062 );
xnor ( n9064 , n9034 , n9063 );
xnor ( n9065 , n9048 , n9053 );
not ( n9066 , n9065 );
not ( n9067 , n9031 );
not ( n9068 , n9010 );
not ( n9069 , n9068 );
and ( n9070 , n9067 , n9069 );
and ( n9071 , n9068 , n9031 );
nor ( n9072 , n9070 , n9071 );
not ( n9073 , n9072 );
and ( n9074 , n9066 , n9073 );
not ( n9075 , n81 );
and ( n9076 , n9075 , n7212 );
and ( n9077 , n81 , n92 );
nor ( n9078 , n9076 , n9077 );
and ( n9079 , n9078 , n7216 );
and ( n9080 , n7218 , n9007 );
nor ( n9081 , n9079 , n9080 );
and ( n9082 , n90 , n82 );
not ( n9083 , n90 );
and ( n9084 , n9083 , n8382 );
nor ( n9085 , n9082 , n9084 );
nand ( n9086 , n9085 , n6847 );
not ( n9087 , n90 );
or ( n9088 , n8254 , n9087 );
or ( n9089 , n83 , n90 );
not ( n9090 , n6858 );
nand ( n9091 , n9088 , n9089 , n9090 );
and ( n9092 , n9086 , n9091 );
and ( n9093 , n7811 , n8862 );
and ( n9094 , n77 , n96 );
nor ( n9095 , n9093 , n9094 );
and ( n9096 , n9095 , n7682 );
and ( n9097 , n76 , n96 );
not ( n9098 , n76 );
and ( n9099 , n9098 , n8862 );
nor ( n9100 , n9097 , n9099 );
and ( n9101 , n9100 , n7689 );
nor ( n9102 , n9096 , n9101 );
xnor ( n9103 , n9092 , n9102 );
or ( n9104 , n9081 , n9103 );
or ( n9105 , n9102 , n9092 );
nand ( n9106 , n9104 , n9105 );
xnor ( n9107 , n9065 , n9072 );
not ( n9108 , n9107 );
and ( n9109 , n9106 , n9108 );
nor ( n9110 , n9074 , n9109 );
or ( n9111 , n9064 , n9110 );
xnor ( n9112 , n8882 , n8869 );
xnor ( n9113 , n8908 , n8895 );
not ( n9114 , n9113 );
and ( n9115 , n9100 , n7902 );
and ( n9116 , n8865 , n7689 );
nor ( n9117 , n9115 , n9116 );
and ( n9118 , n9085 , n6859 );
and ( n9119 , n8870 , n6847 );
nor ( n9120 , n9118 , n9119 );
xor ( n9121 , n9117 , n9120 );
not ( n9122 , n9121 );
not ( n9123 , n94 );
and ( n9124 , n8341 , n9123 );
and ( n9125 , n79 , n94 );
nor ( n9126 , n9124 , n9125 );
and ( n9127 , n9126 , n7204 );
and ( n9128 , n9014 , n7822 );
nor ( n9129 , n9127 , n9128 );
not ( n9130 , n7556 );
and ( n9131 , n98 , n75 );
not ( n9132 , n98 );
and ( n9133 , n9132 , n7871 );
nor ( n9134 , n9131 , n9133 );
and ( n9135 , n9130 , n9134 );
and ( n9136 , n99 , n9046 );
nor ( n9137 , n9135 , n9136 );
not ( n9138 , n10 );
not ( n9139 , n9024 );
and ( n9140 , n9138 , n9139 );
and ( n9141 , n10 , n9024 );
nor ( n9142 , n9140 , n9141 );
xnor ( n9143 , n9137 , n9142 );
or ( n9144 , n9129 , n9143 );
or ( n9145 , n9137 , n9142 );
nand ( n9146 , n9144 , n9145 );
not ( n9147 , n9146 );
or ( n9148 , n9122 , n9147 );
or ( n9149 , n9120 , n9117 );
nand ( n9150 , n9148 , n9149 );
not ( n9151 , n9150 );
or ( n9152 , n9114 , n9151 );
or ( n9153 , n9113 , n9150 );
nand ( n9154 , n9152 , n9153 );
and ( n9155 , n9112 , n9154 );
nor ( n9156 , n9112 , n9154 );
nor ( n9157 , n9155 , n9156 );
xnor ( n9158 , n9110 , n9064 );
nor ( n9159 , n9157 , n9158 );
not ( n9160 , n9159 );
nand ( n9161 , n9111 , n9160 );
nand ( n9162 , n381 , n9161 );
and ( n9163 , n9004 , n9162 );
and ( n9164 , n9063 , n9034 );
and ( n9165 , n9062 , n9055 );
nor ( n9166 , n9164 , n9165 );
not ( n9167 , n9166 );
not ( n9168 , n8314 );
and ( n9169 , n8299 , n8317 );
not ( n9170 , n9169 );
and ( n9171 , n9168 , n9170 );
and ( n9172 , n8314 , n9169 );
nor ( n9173 , n9171 , n9172 );
xnor ( n9174 , n8369 , n8389 );
xor ( n9175 , n9173 , n9174 );
not ( n9176 , n9175 );
or ( n9177 , n9167 , n9176 );
or ( n9178 , n9166 , n9175 );
nand ( n9179 , n9177 , n9178 );
xor ( n9180 , n8913 , n8885 );
or ( n9181 , n9113 , n9112 );
not ( n9182 , n9113 );
not ( n9183 , n9112 );
or ( n9184 , n9182 , n9183 );
nand ( n9185 , n9184 , n9150 );
nand ( n9186 , n9181 , n9185 );
xor ( n9187 , n9180 , n9186 );
xor ( n9188 , n9179 , n9187 );
and ( n9189 , n381 , n9188 );
and ( n9190 , n1 , n87 );
nor ( n9191 , n9189 , n9190 );
nor ( n9192 , n9163 , n9191 );
not ( n9193 , n3700 );
not ( n9194 , n2687 );
not ( n9195 , n8487 );
nand ( n9196 , n9194 , n9195 );
not ( n9197 , n9196 );
not ( n9198 , n9197 );
or ( n9199 , n9193 , n9198 );
and ( n9200 , n7954 , n9196 );
nor ( n9201 , n9200 , n7067 );
nand ( n9202 , n9199 , n9201 );
not ( n9203 , n9202 );
buf ( n9204 , n6517 );
nand ( n9205 , n9204 , n6284 );
not ( n9206 , n9205 );
buf ( n9207 , n5445 );
not ( n9208 , n9207 );
or ( n9209 , n9206 , n9208 );
or ( n9210 , n9205 , n9207 );
nand ( n9211 , n9209 , n9210 );
nand ( n9212 , n7067 , n9211 );
not ( n9213 , n9212 );
or ( n9214 , n9203 , n9213 );
nand ( n9215 , n9214 , n1 );
and ( n9216 , n9180 , n9186 );
and ( n9217 , n9179 , n9187 );
or ( n9218 , n9216 , n9217 );
nand ( n9219 , n9218 , n381 );
and ( n9220 , n1 , n86 );
not ( n9221 , n1 );
not ( n9222 , n9173 );
not ( n9223 , n9174 );
and ( n9224 , n9222 , n9223 );
and ( n9225 , n9173 , n9174 );
nor ( n9226 , n9225 , n9166 );
nor ( n9227 , n9224 , n9226 );
xnor ( n9228 , n8278 , n8335 );
xnor ( n9229 , n9227 , n9228 );
xnor ( n9230 , n8924 , n8919 );
and ( n9231 , n9229 , n9230 );
nor ( n9232 , n9229 , n9230 );
nor ( n9233 , n9231 , n9232 );
and ( n9234 , n9221 , n9233 );
nor ( n9235 , n9220 , n9234 );
nand ( n9236 , n9215 , n9219 , n9235 );
nand ( n9237 , n9192 , n9236 );
not ( n9238 , n9237 );
not ( n9239 , n8490 );
not ( n9240 , n8485 );
nor ( n9241 , n9239 , n9240 );
or ( n9242 , n7954 , n2687 );
nand ( n9243 , n9242 , n9195 );
nor ( n9244 , n9241 , n9243 );
not ( n9245 , n9244 );
not ( n9246 , n9242 );
not ( n9247 , n9195 );
or ( n9248 , n9246 , n9247 );
nand ( n9249 , n9248 , n9241 );
nand ( n9250 , n9245 , n8687 , n9249 );
or ( n9251 , n9228 , n9227 );
not ( n9252 , n9232 );
nand ( n9253 , n9251 , n9252 );
nand ( n9254 , n381 , n9253 );
nand ( n9255 , n9250 , n9254 );
nand ( n9256 , n6511 , n6513 );
and ( n9257 , n9256 , n6293 );
not ( n9258 , n9257 );
not ( n9259 , n9258 );
not ( n9260 , n6284 );
not ( n9261 , n9207 );
or ( n9262 , n9260 , n9261 );
buf ( n9263 , n9204 );
nand ( n9264 , n9262 , n9263 );
not ( n9265 , n9264 );
not ( n9266 , n9265 );
and ( n9267 , n9259 , n9266 );
or ( n9268 , n9257 , n9264 );
nand ( n9269 , n1 , n7067 );
not ( n9270 , n9269 );
nand ( n9271 , n9268 , n9270 );
nor ( n9272 , n9267 , n9271 );
or ( n9273 , n9255 , n9272 );
and ( n9274 , n8928 , n8929 );
nor ( n9275 , n9274 , n8930 );
and ( n9276 , n9275 , n381 );
and ( n9277 , n1 , n85 );
nor ( n9278 , n9276 , n9277 );
not ( n9279 , n9278 );
nand ( n9280 , n9273 , n9279 );
not ( n9281 , n9219 );
not ( n9282 , n9215 );
or ( n9283 , n9281 , n9282 );
not ( n9284 , n9235 );
nand ( n9285 , n9283 , n9284 );
nand ( n9286 , n9280 , n9285 );
nor ( n9287 , n9238 , n9286 );
not ( n9288 , n9287 );
nor ( n9289 , n5433 , n5425 );
not ( n9290 , n9289 );
not ( n9291 , n4984 );
not ( n9292 , n8989 );
or ( n9293 , n9291 , n9292 );
not ( n9294 , n5435 );
nand ( n9295 , n9293 , n9294 );
not ( n9296 , n9295 );
nand ( n9297 , n9290 , n9296 );
and ( n9298 , n9295 , n9289 );
nor ( n9299 , n9298 , n9269 );
and ( n9300 , n9297 , n9299 );
xor ( n9301 , n9103 , n9081 );
not ( n9302 , n78 );
not ( n9303 , n96 );
and ( n9304 , n9302 , n9303 );
and ( n9305 , n78 , n96 );
nor ( n9306 , n9304 , n9305 );
and ( n9307 , n9306 , n8866 );
and ( n9308 , n9095 , n7689 );
nor ( n9309 , n9307 , n9308 );
xor ( n9310 , n76 , n98 );
and ( n9311 , n9130 , n9310 );
and ( n9312 , n99 , n9134 );
nor ( n9313 , n9311 , n9312 );
nand ( n9314 , n83 , n6845 );
and ( n9315 , n9314 , n11 );
not ( n9316 , n9314 );
not ( n9317 , n11 );
and ( n9318 , n9316 , n9317 );
nor ( n9319 , n9315 , n9318 );
xnor ( n9320 , n9313 , n9319 );
or ( n9321 , n9309 , n9320 );
not ( n9322 , n9309 );
not ( n9323 , n9320 );
or ( n9324 , n9322 , n9323 );
and ( n9325 , n94 , n80 );
not ( n9326 , n94 );
and ( n9327 , n9326 , n8354 );
nor ( n9328 , n9325 , n9327 );
not ( n9329 , n9328 );
not ( n9330 , n7189 );
or ( n9331 , n9329 , n9330 );
not ( n9332 , n81 );
not ( n9333 , n94 );
and ( n9334 , n9332 , n9333 );
and ( n9335 , n81 , n94 );
nor ( n9336 , n9334 , n9335 );
nand ( n9337 , n9336 , n7204 );
nand ( n9338 , n9331 , n9337 );
not ( n9339 , n9338 );
xor ( n9340 , n77 , n98 );
and ( n9341 , n9130 , n9340 );
and ( n9342 , n99 , n9310 );
nor ( n9343 , n9341 , n9342 );
not ( n9344 , n9343 );
nand ( n9345 , n83 , n93 );
or ( n9346 , n83 , n93 );
nand ( n9347 , n9346 , n94 );
nand ( n9348 , n9345 , n92 , n9347 );
xnor ( n9349 , n9348 , n12 );
not ( n9350 , n9349 );
or ( n9351 , n9344 , n9350 );
or ( n9352 , n9343 , n9349 );
nand ( n9353 , n9351 , n9352 );
not ( n9354 , n9353 );
or ( n9355 , n9339 , n9354 );
not ( n9356 , n9343 );
nand ( n9357 , n9356 , n9349 );
nand ( n9358 , n9355 , n9357 );
nand ( n9359 , n9324 , n9358 );
nand ( n9360 , n9321 , n9359 );
and ( n9361 , n9301 , n9360 );
and ( n9362 , n9328 , n7204 );
and ( n9363 , n9126 , n7822 );
nor ( n9364 , n9362 , n9363 );
and ( n9365 , n8382 , n7212 );
and ( n9366 , n82 , n92 );
nor ( n9367 , n9365 , n9366 );
not ( n9368 , n7026 );
and ( n9369 , n9367 , n9368 );
and ( n9370 , n7354 , n9078 );
nor ( n9371 , n9369 , n9370 );
not ( n9372 , n9348 );
nand ( n9373 , n9372 , n12 );
xnor ( n9374 , n9371 , n9373 );
or ( n9375 , n9364 , n9374 );
or ( n9376 , n9373 , n9371 );
nand ( n9377 , n9375 , n9376 );
or ( n9378 , n9313 , n9319 );
or ( n9379 , n9317 , n9314 );
nand ( n9380 , n9378 , n9379 );
xor ( n9381 , n9377 , n9380 );
xor ( n9382 , n9143 , n9129 );
xor ( n9383 , n9381 , n9382 );
xor ( n9384 , n9360 , n9301 );
and ( n9385 , n9383 , n9384 );
nor ( n9386 , n9361 , n9385 );
nor ( n9387 , n1 , n9386 );
nor ( n9388 , n9300 , n9387 );
xor ( n9389 , n9377 , n9380 );
and ( n9390 , n9389 , n9382 );
and ( n9391 , n9377 , n9380 );
or ( n9392 , n9390 , n9391 );
not ( n9393 , n9106 );
not ( n9394 , n9393 );
not ( n9395 , n9108 );
or ( n9396 , n9394 , n9395 );
nand ( n9397 , n9106 , n9107 );
nand ( n9398 , n9396 , n9397 );
xor ( n9399 , n9121 , n9146 );
xor ( n9400 , n9398 , n9399 );
xor ( n9401 , n9392 , n9400 );
and ( n9402 , n381 , n9401 );
and ( n9403 , n1 , n89 );
nor ( n9404 , n9402 , n9403 );
nor ( n9405 , n381 , n7067 );
not ( n9406 , n3676 );
not ( n9407 , n8964 );
not ( n9408 , n9407 );
or ( n9409 , n9406 , n9408 );
nand ( n9410 , n9409 , n3683 );
not ( n9411 , n9410 );
not ( n9412 , n3684 );
nor ( n9413 , n9412 , n3687 );
not ( n9414 , n9413 );
and ( n9415 , n9411 , n9414 );
and ( n9416 , n9410 , n9413 );
nor ( n9417 , n9415 , n9416 );
nand ( n9418 , n9405 , n9417 );
nand ( n9419 , n9388 , n9404 , n9418 );
nand ( n9420 , n9294 , n4984 );
and ( n9421 , n9420 , n8989 );
not ( n9422 , n9420 );
not ( n9423 , n8989 );
and ( n9424 , n9422 , n9423 );
nor ( n9425 , n9421 , n9424 );
nor ( n9426 , n2 , n9425 );
nand ( n9427 , n3676 , n3683 );
not ( n9428 , n9427 );
nor ( n9429 , n9428 , n9407 );
or ( n9430 , n9427 , n8964 );
nand ( n9431 , n9430 , n2 );
nor ( n9432 , n9429 , n9431 );
or ( n9433 , n9426 , n9432 );
nand ( n9434 , n9433 , n1 );
not ( n9435 , n9434 );
xnor ( n9436 , n9374 , n9364 );
not ( n9437 , n9309 );
not ( n9438 , n9358 );
and ( n9439 , n9437 , n9438 );
and ( n9440 , n9309 , n9358 );
nor ( n9441 , n9439 , n9440 );
xnor ( n9442 , n9441 , n9320 );
and ( n9443 , n9436 , n9442 );
not ( n9444 , n9436 );
not ( n9445 , n9442 );
and ( n9446 , n9444 , n9445 );
and ( n9447 , n83 , n7014 );
xor ( n9448 , n9447 , n13 );
and ( n9449 , n8382 , n9123 );
and ( n9450 , n82 , n94 );
nor ( n9451 , n9449 , n9450 );
not ( n9452 , n9451 );
not ( n9453 , n7204 );
or ( n9454 , n9452 , n9453 );
nand ( n9455 , n9336 , n7191 );
nand ( n9456 , n9454 , n9455 );
and ( n9457 , n9448 , n9456 );
and ( n9458 , n13 , n9447 );
nor ( n9459 , n9457 , n9458 );
nand ( n9460 , n7016 , n9367 );
or ( n9461 , n8254 , n7212 );
or ( n9462 , n83 , n92 );
nand ( n9463 , n9461 , n9462 , n7025 );
and ( n9464 , n9460 , n9463 );
nand ( n9465 , n9306 , n7689 );
not ( n9466 , n79 );
not ( n9467 , n96 );
and ( n9468 , n9466 , n9467 );
and ( n9469 , n79 , n96 );
nor ( n9470 , n9468 , n9469 );
nand ( n9471 , n9470 , n7775 );
and ( n9472 , n9465 , n9471 );
xnor ( n9473 , n9464 , n9472 );
or ( n9474 , n9459 , n9473 );
or ( n9475 , n9472 , n9464 );
nand ( n9476 , n9474 , n9475 );
nor ( n9477 , n9446 , n9476 );
nor ( n9478 , n9443 , n9477 , n1 );
or ( n9479 , n9435 , n9478 );
xor ( n9480 , n9383 , n9384 );
and ( n9481 , n381 , n9480 );
and ( n9482 , n1 , n90 );
nor ( n9483 , n9481 , n9482 );
not ( n9484 , n9483 );
nand ( n9485 , n9479 , n9484 );
not ( n9486 , n9478 );
nand ( n9487 , n9486 , n9483 , n9434 );
not ( n9488 , n9476 );
not ( n9489 , n9442 );
and ( n9490 , n9488 , n9489 );
and ( n9491 , n9476 , n9442 );
nor ( n9492 , n9490 , n9491 );
or ( n9493 , n9436 , n9492 );
and ( n9494 , n9436 , n9492 );
nor ( n9495 , n9494 , n1 );
and ( n9496 , n9493 , n9495 );
and ( n9497 , n1 , n91 );
nor ( n9498 , n9496 , n9497 );
not ( n9499 , n9498 );
xnor ( n9500 , n9353 , n9338 );
not ( n9501 , n9500 );
and ( n9502 , n8354 , n8862 );
and ( n9503 , n80 , n96 );
nor ( n9504 , n9502 , n9503 );
and ( n9505 , n9504 , n7902 );
and ( n9506 , n9470 , n7689 );
nor ( n9507 , n9505 , n9506 );
nand ( n9508 , n83 , n95 );
or ( n9509 , n83 , n95 );
nand ( n9510 , n9509 , n96 );
nand ( n9511 , n9508 , n94 , n9510 );
not ( n9512 , n9511 );
nand ( n9513 , n9512 , n14 );
nand ( n9514 , n99 , n9340 );
xor ( n9515 , n78 , n98 );
nand ( n9516 , n8261 , n9515 );
and ( n9517 , n9514 , n9516 );
xnor ( n9518 , n9513 , n9517 );
or ( n9519 , n9507 , n9518 );
or ( n9520 , n9513 , n9517 );
nand ( n9521 , n9519 , n9520 );
nand ( n9522 , n9501 , n9521 );
not ( n9523 , n9522 );
xnor ( n9524 , n9473 , n9459 );
and ( n9525 , n9521 , n9500 );
nor ( n9526 , n9521 , n9500 );
nor ( n9527 , n9525 , n9526 );
nor ( n9528 , n9524 , n9527 );
not ( n9529 , n9528 );
not ( n9530 , n9529 );
or ( n9531 , n9523 , n9530 );
nand ( n9532 , n9531 , n381 );
not ( n9533 , n5417 );
nand ( n9534 , n5045 , n5046 );
nand ( n9535 , n9533 , n9534 );
not ( n9536 , n9535 );
not ( n9537 , n5105 );
buf ( n9538 , n5414 );
nand ( n9539 , n5108 , n9538 );
nand ( n9540 , n7067 , n9536 , n9537 , n9539 );
not ( n9541 , n3143 );
not ( n9542 , n3495 );
or ( n9543 , n9542 , n3502 );
nand ( n9544 , n9543 , n3271 );
nand ( n9545 , n3274 , n9544 );
not ( n9546 , n9545 );
or ( n9547 , n9541 , n9546 );
not ( n9548 , n3048 );
not ( n9549 , n9548 );
nand ( n9550 , n3049 , n3051 );
nand ( n9551 , n9549 , n9550 );
not ( n9552 , n9551 );
nand ( n9553 , n9547 , n9552 );
nand ( n9554 , n9545 , n3143 , n9551 );
nand ( n9555 , n9553 , n2 , n9554 );
nand ( n9556 , n9537 , n9539 );
nand ( n9557 , n9556 , n7067 , n9535 );
nand ( n9558 , n9540 , n9555 , n9557 );
nand ( n9559 , n1 , n9558 );
nand ( n9560 , n9532 , n9559 );
and ( n9561 , n9499 , n9560 );
nand ( n9562 , n9487 , n9561 );
nand ( n9563 , n9485 , n9562 );
and ( n9564 , n9419 , n9563 );
and ( n9565 , n9418 , n9388 );
nor ( n9566 , n9565 , n9404 );
nor ( n9567 , n9564 , n9566 );
and ( n9568 , n9399 , n9398 );
and ( n9569 , n9392 , n9400 );
nor ( n9570 , n9568 , n9569 );
nor ( n9571 , n9570 , n1 );
or ( n9572 , n1 , n9571 );
not ( n9573 , n9572 );
not ( n9574 , n2 );
not ( n9575 , n8973 );
nand ( n9576 , n9575 , n3606 );
not ( n9577 , n9576 );
and ( n9578 , n8969 , n9577 );
not ( n9579 , n8969 );
and ( n9580 , n9579 , n9576 );
nor ( n9581 , n9578 , n9580 );
not ( n9582 , n9581 );
or ( n9583 , n9574 , n9582 );
not ( n9584 , n8993 );
nand ( n9585 , n5442 , n4659 );
not ( n9586 , n9585 );
or ( n9587 , n9584 , n9586 );
or ( n9588 , n8993 , n9585 );
nand ( n9589 , n9587 , n9588 );
and ( n9590 , n9589 , n7067 );
nor ( n9591 , n9590 , n9571 );
nand ( n9592 , n9583 , n9591 );
not ( n9593 , n9592 );
or ( n9594 , n9573 , n9593 );
and ( n9595 , n9157 , n9158 );
nor ( n9596 , n9595 , n9159 );
and ( n9597 , n381 , n9596 );
and ( n9598 , n1 , n88 );
nor ( n9599 , n9597 , n9598 );
nand ( n9600 , n9594 , n9599 );
not ( n9601 , n9600 );
or ( n9602 , n9567 , n9601 );
not ( n9603 , n9599 );
nand ( n9604 , n9603 , n9572 , n9592 );
nand ( n9605 , n9602 , n9604 );
not ( n9606 , n9605 );
nand ( n9607 , n83 , n7786 );
and ( n9608 , n9607 , n15 );
not ( n9609 , n9607 );
not ( n9610 , n15 );
and ( n9611 , n9609 , n9610 );
nor ( n9612 , n9608 , n9611 );
nand ( n9613 , n83 , n97 );
or ( n9614 , n83 , n97 );
nand ( n9615 , n9614 , n98 );
nand ( n9616 , n9613 , n96 , n9615 );
not ( n9617 , n9616 );
nand ( n9618 , n9617 , n16 );
xnor ( n9619 , n9612 , n9618 );
and ( n9620 , n8382 , n8862 );
and ( n9621 , n82 , n96 );
nor ( n9622 , n9620 , n9621 );
and ( n9623 , n9622 , n8866 );
and ( n9624 , n9075 , n8862 );
and ( n9625 , n81 , n96 );
nor ( n9626 , n9624 , n9625 );
and ( n9627 , n9626 , n7689 );
nor ( n9628 , n9623 , n9627 );
not ( n9629 , n98 );
and ( n9630 , n8354 , n9629 );
and ( n9631 , n80 , n98 );
nor ( n9632 , n9630 , n9631 );
and ( n9633 , n7557 , n9632 );
xor ( n9634 , n79 , n98 );
and ( n9635 , n99 , n9634 );
nor ( n9636 , n9633 , n9635 );
xnor ( n9637 , n9628 , n9636 );
or ( n9638 , n9619 , n9637 );
and ( n9639 , n9619 , n9637 );
nor ( n9640 , n9639 , n1 );
and ( n9641 , n9638 , n9640 );
and ( n9642 , n1 , n95 );
nor ( n9643 , n9641 , n9642 );
not ( n9644 , n99 );
not ( n9645 , n9632 );
or ( n9646 , n9644 , n9645 );
and ( n9647 , n9075 , n9629 );
and ( n9648 , n81 , n98 );
nor ( n9649 , n9647 , n9648 );
nand ( n9650 , n7557 , n9649 );
nand ( n9651 , n9646 , n9650 );
not ( n9652 , n16 );
not ( n9653 , n9616 );
or ( n9654 , n9652 , n9653 );
or ( n9655 , n16 , n9616 );
nand ( n9656 , n9654 , n9655 );
and ( n9657 , n9651 , n9656 );
not ( n9658 , n9622 );
not ( n9659 , n7689 );
or ( n9660 , n9658 , n9659 );
or ( n9661 , n8254 , n8862 );
or ( n9662 , n83 , n96 );
nand ( n9663 , n9661 , n9662 , n8866 );
nand ( n9664 , n9660 , n9663 );
xor ( n9665 , n9651 , n9656 );
and ( n9666 , n9664 , n9665 );
or ( n9667 , n9657 , n9666 );
nand ( n9668 , n9667 , n381 );
not ( n9669 , n3494 );
nor ( n9670 , n9669 , n3368 );
not ( n9671 , n3355 );
not ( n9672 , n9671 );
nand ( n9673 , n3416 , n3488 );
not ( n9674 , n9673 );
or ( n9675 , n9672 , n9674 );
nand ( n9676 , n9675 , n3419 );
and ( n9677 , n9670 , n9676 );
or ( n9678 , n9670 , n9676 );
nand ( n9679 , n9678 , n2 );
or ( n9680 , n9677 , n9679 );
not ( n9681 , n5304 );
nand ( n9682 , n9681 , n5407 );
not ( n9683 , n9682 );
not ( n9684 , n5286 );
nand ( n9685 , n5338 , n5403 );
not ( n9686 , n9685 );
or ( n9687 , n9684 , n9686 );
nand ( n9688 , n9687 , n5339 );
not ( n9689 , n9688 );
or ( n9690 , n9683 , n9689 );
or ( n9691 , n9682 , n9688 );
nand ( n9692 , n9690 , n9691 );
nand ( n9693 , n7067 , n9692 );
nand ( n9694 , n9680 , n9693 );
nand ( n9695 , n1 , n9694 );
nand ( n9696 , n9668 , n9695 );
not ( n9697 , n9696 );
nand ( n9698 , n9643 , n9697 );
nand ( n9699 , n83 , n99 );
and ( n9700 , n98 , n9699 );
not ( n9701 , n9700 );
nand ( n9702 , n9701 , n1187 );
and ( n9703 , n18 , n9700 );
nor ( n9704 , n9703 , n1 );
and ( n9705 , n9702 , n9704 );
and ( n9706 , n1 , n98 );
nor ( n9707 , n9705 , n9706 );
not ( n9708 , n9707 );
buf ( n9709 , n3474 );
not ( n9710 , n9709 );
not ( n9711 , n3486 );
nor ( n9712 , n9711 , n3484 );
not ( n9713 , n9712 );
or ( n9714 , n9710 , n9713 );
buf ( n9715 , n9709 );
or ( n9716 , n9715 , n9712 );
nand ( n9717 , n9714 , n9716 );
and ( n9718 , n8687 , n9717 );
not ( n9719 , n381 );
not ( n9720 , n99 );
and ( n9721 , n8382 , n9629 );
and ( n9722 , n82 , n98 );
nor ( n9723 , n9721 , n9722 );
not ( n9724 , n9723 );
or ( n9725 , n9720 , n9724 );
not ( n9726 , n7557 );
or ( n9727 , n83 , n9726 );
nand ( n9728 , n9725 , n9727 );
not ( n9729 , n9728 );
or ( n9730 , n9719 , n9729 );
nor ( n9731 , n5400 , n5368 );
not ( n9732 , n9731 );
nor ( n9733 , n381 , n2 );
nand ( n9734 , n9732 , n9733 , n5401 );
nand ( n9735 , n9730 , n9734 );
nor ( n9736 , n9718 , n9735 );
not ( n9737 , n9736 );
nand ( n9738 , n9708 , n9737 );
or ( n9739 , n1 , n9699 );
or ( n9740 , n381 , n7555 );
nand ( n9741 , n9739 , n9740 );
not ( n9742 , n3441 );
not ( n9743 , n3470 );
nor ( n9744 , n9743 , n3473 );
not ( n9745 , n9744 );
nand ( n9746 , n9742 , n9745 );
and ( n9747 , n3441 , n9744 );
nor ( n9748 , n9747 , n7067 );
and ( n9749 , n9746 , n9748 );
not ( n9750 , n5397 );
nand ( n9751 , n9750 , n5399 );
xnor ( n9752 , n9751 , n5381 );
nor ( n9753 , n2 , n9752 );
nor ( n9754 , n9749 , n9753 );
or ( n9755 , n381 , n9754 );
nand ( n9756 , n19 , n381 );
nand ( n9757 , n9755 , n9756 );
and ( n9758 , n9741 , n9757 );
nand ( n9759 , n9707 , n9736 );
nand ( n9760 , n9758 , n9759 );
nand ( n9761 , n9738 , n9760 );
not ( n9762 , n3487 );
not ( n9763 , n3416 );
not ( n9764 , n3421 );
nor ( n9765 , n9763 , n9764 );
and ( n9766 , n9762 , n9765 );
nor ( n9767 , n9766 , n7067 );
not ( n9768 , n9762 );
not ( n9769 , n9765 );
nand ( n9770 , n9768 , n9769 );
and ( n9771 , n9767 , n9770 );
not ( n9772 , n5337 );
nand ( n9773 , n9772 , n5340 );
not ( n9774 , n5402 );
and ( n9775 , n9773 , n9774 );
not ( n9776 , n9773 );
and ( n9777 , n9776 , n5402 );
nor ( n9778 , n9775 , n9777 );
nor ( n9779 , n2 , n9778 );
nor ( n9780 , n9771 , n9779 );
and ( n9781 , n9780 , n1 );
not ( n9782 , n9726 );
and ( n9783 , n9782 , n9723 );
and ( n9784 , n99 , n9649 );
nor ( n9785 , n9783 , n9784 );
nor ( n9786 , n1 , n9785 );
nor ( n9787 , n9781 , n9786 );
nand ( n9788 , n18 , n9700 );
nand ( n9789 , n83 , n7689 );
and ( n9790 , n9789 , n17 );
not ( n9791 , n9789 );
not ( n9792 , n17 );
and ( n9793 , n9791 , n9792 );
nor ( n9794 , n9790 , n9793 );
or ( n9795 , n9788 , n9794 );
and ( n9796 , n9788 , n9794 );
nor ( n9797 , n9796 , n1 );
and ( n9798 , n9795 , n9797 );
and ( n9799 , n1 , n97 );
nor ( n9800 , n9798 , n9799 );
nor ( n9801 , n9787 , n9800 );
or ( n9802 , n9761 , n9801 );
nand ( n9803 , n9800 , n9787 );
nand ( n9804 , n9802 , n9803 );
xor ( n9805 , n9664 , n9665 );
and ( n9806 , n381 , n9805 );
and ( n9807 , n1 , n96 );
nor ( n9808 , n9806 , n9807 );
not ( n9809 , n9808 );
not ( n9810 , n381 );
or ( n9811 , n9788 , n9794 );
or ( n9812 , n9792 , n9789 );
nand ( n9813 , n9811 , n9812 );
not ( n9814 , n9813 );
or ( n9815 , n9810 , n9814 );
nand ( n9816 , n5339 , n5286 );
not ( n9817 , n9816 );
not ( n9818 , n9685 );
or ( n9819 , n9817 , n9818 );
or ( n9820 , n9816 , n9685 );
nand ( n9821 , n9819 , n9820 );
nand ( n9822 , n7067 , n9821 );
not ( n9823 , n9822 );
not ( n9824 , n3355 );
nand ( n9825 , n9824 , n3419 );
not ( n9826 , n9825 );
nand ( n9827 , n9673 , n9826 );
not ( n9828 , n9673 );
nand ( n9829 , n9828 , n9825 );
nand ( n9830 , n9827 , n2 , n9829 );
not ( n9831 , n9830 );
or ( n9832 , n9823 , n9831 );
nand ( n9833 , n9832 , n1 );
nand ( n9834 , n9815 , n9833 );
nand ( n9835 , n9809 , n9834 );
and ( n9836 , n9804 , n9835 );
not ( n9837 , n9808 );
nor ( n9838 , n9837 , n9834 );
nor ( n9839 , n9836 , n9838 );
or ( n9840 , n9618 , n9612 );
or ( n9841 , n9610 , n9607 );
nand ( n9842 , n9840 , n9841 );
not ( n9843 , n9626 );
not ( n9844 , n8866 );
or ( n9845 , n9843 , n9844 );
nand ( n9846 , n9504 , n7689 );
nand ( n9847 , n9845 , n9846 );
nand ( n9848 , n83 , n94 );
and ( n9849 , n8254 , n9123 );
nor ( n9850 , n9849 , n7203 );
and ( n9851 , n9848 , n9850 );
and ( n9852 , n9451 , n7191 );
nor ( n9853 , n9851 , n9852 );
not ( n9854 , n9853 );
and ( n9855 , n8261 , n9634 );
and ( n9856 , n99 , n9515 );
nor ( n9857 , n9855 , n9856 );
xor ( n9858 , n9511 , n14 );
nand ( n9859 , n9857 , n9858 );
not ( n9860 , n9859 );
nor ( n9861 , n9857 , n9858 );
nor ( n9862 , n9860 , n9861 );
not ( n9863 , n9862 );
or ( n9864 , n9854 , n9863 );
or ( n9865 , n9853 , n9862 );
nand ( n9866 , n9864 , n9865 );
xor ( n9867 , n9847 , n9866 );
xor ( n9868 , n9842 , n9867 );
and ( n9869 , n381 , n9868 );
and ( n9870 , n1 , n94 );
nor ( n9871 , n9869 , n9870 );
or ( n9872 , n9619 , n9637 );
or ( n9873 , n9636 , n9628 );
nand ( n9874 , n9872 , n9873 );
nand ( n9875 , n381 , n9874 );
not ( n9876 , n5212 );
nand ( n9877 , n9876 , n5410 );
not ( n9878 , n5408 );
and ( n9879 , n9877 , n9878 );
not ( n9880 , n9877 );
not ( n9881 , n9878 );
and ( n9882 , n9880 , n9881 );
nor ( n9883 , n9879 , n9882 );
nand ( n9884 , n7067 , n9883 );
not ( n9885 , n9884 );
not ( n9886 , n3252 );
not ( n9887 , n9886 );
nand ( n9888 , n9887 , n3501 );
or ( n9889 , n9888 , n9542 );
nand ( n9890 , n9888 , n9542 );
nand ( n9891 , n9889 , n9890 , n2 );
not ( n9892 , n9891 );
or ( n9893 , n9885 , n9892 );
nand ( n9894 , n9893 , n1 );
nand ( n9895 , n9871 , n9875 , n9894 );
nand ( n9896 , n9698 , n9839 , n9895 );
not ( n9897 , n9896 );
and ( n9898 , n9524 , n9527 );
nor ( n9899 , n9898 , n9528 );
and ( n9900 , n381 , n9899 );
and ( n9901 , n1 , n92 );
nor ( n9902 , n9900 , n9901 );
xnor ( n9903 , n9448 , n9456 );
xnor ( n9904 , n9507 , n9518 );
nand ( n9905 , n9903 , n9904 );
or ( n9906 , n9903 , n9904 );
not ( n9907 , n9853 );
and ( n9908 , n9907 , n9859 );
nor ( n9909 , n9908 , n9861 );
nand ( n9910 , n9906 , n9909 );
nand ( n9911 , n9905 , n381 , n9910 );
not ( n9912 , n3273 );
nand ( n9913 , n9912 , n3143 );
not ( n9914 , n9913 );
not ( n9915 , n9544 );
not ( n9916 , n9915 );
nor ( n9917 , n9914 , n9916 );
or ( n9918 , n9913 , n9915 );
nand ( n9919 , n9918 , n2 );
or ( n9920 , n9917 , n9919 );
not ( n9921 , n5105 );
nand ( n9922 , n9921 , n5108 );
not ( n9923 , n9922 );
not ( n9924 , n9538 );
or ( n9925 , n9923 , n9924 );
or ( n9926 , n9922 , n9538 );
nand ( n9927 , n9925 , n9926 );
nand ( n9928 , n7067 , n9927 );
nand ( n9929 , n9920 , n9928 );
nand ( n9930 , n1 , n9929 );
nand ( n9931 , n9902 , n9911 , n9930 );
xnor ( n9932 , n9904 , n9909 );
or ( n9933 , n9903 , n9932 );
and ( n9934 , n9903 , n9932 );
nor ( n9935 , n9934 , n1 );
and ( n9936 , n9933 , n9935 );
and ( n9937 , n1 , n93 );
nor ( n9938 , n9936 , n9937 );
and ( n9939 , n9847 , n9866 );
and ( n9940 , n9842 , n9867 );
or ( n9941 , n9939 , n9940 );
nand ( n9942 , n9941 , n381 );
nor ( n9943 , n381 , n7067 );
not ( n9944 , n3501 );
not ( n9945 , n3495 );
or ( n9946 , n9944 , n9945 );
nand ( n9947 , n9946 , n3252 );
not ( n9948 , n3270 );
not ( n9949 , n9948 );
nand ( n9950 , n9949 , n3265 );
not ( n9951 , n9950 );
and ( n9952 , n9947 , n9951 );
not ( n9953 , n9947 );
and ( n9954 , n9953 , n9950 );
nor ( n9955 , n9952 , n9954 );
and ( n9956 , n9943 , n9955 );
not ( n9957 , n5212 );
not ( n9958 , n5410 );
nand ( n9959 , n9957 , n9958 );
not ( n9960 , n9959 );
not ( n9961 , n9881 );
nand ( n9962 , n9957 , n9961 );
not ( n9963 , n9962 );
or ( n9964 , n9960 , n9963 );
not ( n9965 , n5169 );
not ( n9966 , n9965 );
not ( n9967 , n5214 );
nor ( n9968 , n9966 , n9967 );
not ( n9969 , n9968 );
nand ( n9970 , n9964 , n9969 );
nor ( n9971 , n381 , n2 );
nand ( n9972 , n9962 , n9959 , n9968 );
and ( n9973 , n9970 , n9971 , n9972 );
nor ( n9974 , n9956 , n9973 );
nand ( n9975 , n9942 , n9974 );
not ( n9976 , n9975 );
nand ( n9977 , n9938 , n9976 );
nand ( n9978 , n9897 , n9931 , n9977 );
not ( n9979 , n9875 );
not ( n9980 , n9894 );
or ( n9981 , n9979 , n9980 );
not ( n9982 , n9871 );
nand ( n9983 , n9981 , n9982 );
not ( n9984 , n9983 );
not ( n9985 , n9984 );
not ( n9986 , n9643 );
nand ( n9987 , n9696 , n9986 );
not ( n9988 , n9987 );
nand ( n9989 , n9988 , n9895 );
nand ( n9990 , n9985 , n9989 );
nand ( n9991 , n9977 , n9931 , n9990 );
nand ( n9992 , n9978 , n9991 );
not ( n9993 , n9992 );
nand ( n9994 , n9902 , n9911 , n9930 );
not ( n9995 , n9975 );
nor ( n9996 , n9995 , n9938 );
and ( n9997 , n9994 , n9996 );
and ( n9998 , n9911 , n9930 );
nor ( n9999 , n9998 , n9902 );
nor ( n10000 , n9997 , n9999 );
nand ( n10001 , n9993 , n10000 );
nand ( n10002 , n9532 , n9498 , n9559 );
and ( n10003 , n9487 , n10002 );
and ( n10004 , n9419 , n10003 , n9600 );
nand ( n10005 , n10001 , n10004 );
nand ( n10006 , n9606 , n10005 );
and ( n10007 , n9162 , n9191 );
not ( n10008 , n10007 );
and ( n10009 , n8984 , n9002 );
not ( n10010 , n10009 );
or ( n10011 , n10008 , n10010 );
nand ( n10012 , n9235 , n9219 , n9215 );
nand ( n10013 , n10011 , n10012 );
not ( n10014 , n10013 );
nand ( n10015 , n10006 , n10014 );
not ( n10016 , n10015 );
or ( n10017 , n9288 , n10016 );
not ( n10018 , n9272 );
not ( n10019 , n9241 );
not ( n10020 , n9247 );
nand ( n10021 , n10019 , n10020 );
not ( n10022 , n10021 );
not ( n10023 , n9246 );
nand ( n10024 , n10022 , n10023 );
nand ( n10025 , n10024 , n8687 , n9249 );
nand ( n10026 , n10018 , n10025 , n9254 , n9278 );
not ( n10027 , n8958 );
nand ( n10028 , n10027 , n8933 , n8950 );
nand ( n10029 , n10026 , n10028 );
not ( n10030 , n10029 );
nand ( n10031 , n10017 , n10030 );
nand ( n10032 , n8961 , n10031 );
not ( n10033 , n1 );
not ( n10034 , n8584 );
or ( n10035 , n10033 , n10034 );
nand ( n10036 , n10035 , n8587 );
nand ( n10037 , n7953 , n7964 );
not ( n10038 , n7983 );
nand ( n10039 , n10038 , n7991 );
nand ( n10040 , n10037 , n10039 , n8000 , n8003 );
and ( n10041 , n10040 , n1 );
nor ( n10042 , n10041 , n8083 );
nand ( n10043 , n7949 , n10042 );
not ( n10044 , n8532 );
nand ( n10045 , n8553 , n10044 , n8561 );
not ( n10046 , n10045 );
and ( n10047 , n8459 , n8508 , n8526 );
nor ( n10048 , n10046 , n10047 );
nand ( n10049 , n10036 , n10043 , n10048 );
not ( n10050 , n10049 );
nand ( n10051 , n8852 , n10032 , n10050 );
and ( n10052 , n8850 , n10051 );
not ( n10053 , n10052 );
or ( n10054 , n7159 , n7160 );
nand ( n10055 , n10054 , n7416 , n7401 );
and ( n10056 , n10055 , n7452 );
nand ( n10057 , n7118 , n10056 );
not ( n10058 , n10057 );
nand ( n10059 , n7479 , n10053 , n10058 );
nand ( n10060 , n384 , n7481 , n10059 );
and ( n10061 , n298 , n316 );
not ( n10062 , n298 );
and ( n10063 , n10062 , n319 );
nor ( n10064 , n10061 , n10063 );
not ( n10065 , n312 );
and ( n10066 , n346 , n10065 );
nor ( n10067 , n10066 , n297 );
or ( n10068 , n10064 , n10067 );
and ( n10069 , n10064 , n10067 );
nor ( n10070 , n10069 , n1 );
nand ( n10071 , n10068 , n10070 );
or ( n10072 , n321 , n353 );
or ( n10073 , n319 , n315 );
nand ( n10074 , n10072 , n10073 );
nand ( n10075 , n381 , n10074 );
nor ( n10076 , n10071 , n10075 );
not ( n10077 , n10076 );
nand ( n10078 , n10071 , n10075 );
nand ( n10079 , n10077 , n10078 );
not ( n10080 , n10079 );
and ( n10081 , n10060 , n10080 );
not ( n10082 , n10060 );
and ( n10083 , n10082 , n10079 );
nor ( n10084 , n10081 , n10083 );
not ( n10085 , n10057 );
and ( n10086 , n7477 , n10085 );
not ( n10087 , n10051 );
buf ( n10088 , n10087 );
and ( n10089 , n10086 , n10088 );
nor ( n10090 , n10089 , n6891 );
not ( n10091 , n8850 );
buf ( n10092 , n10091 );
nand ( n10093 , n10092 , n10086 );
nand ( n10094 , n7475 , n7477 );
nand ( n10095 , n10090 , n10093 , n10094 );
nor ( n10096 , n385 , n383 );
and ( n10097 , n10095 , n10096 );
not ( n10098 , n10095 );
not ( n10099 , n10096 );
and ( n10100 , n10098 , n10099 );
nor ( n10101 , n10097 , n10100 );
and ( n10102 , n472 , n6890 );
not ( n10103 , n10102 );
not ( n10104 , n10032 );
not ( n10105 , n10104 );
not ( n10106 , n8851 );
nand ( n10107 , n10105 , n10106 , n10056 , n10050 );
not ( n10108 , n7459 );
and ( n10109 , n7466 , n7474 );
nand ( n10110 , n10107 , n10108 , n10109 );
not ( n10111 , n10110 );
nand ( n10112 , n7119 , n7474 , n7466 );
not ( n10113 , n10112 );
or ( n10114 , n10111 , n10113 );
not ( n10115 , n8849 );
not ( n10116 , n10115 );
not ( n10117 , n8819 );
or ( n10118 , n10116 , n10117 );
nand ( n10119 , n10118 , n10058 );
nand ( n10120 , n10114 , n10119 );
not ( n10121 , n7476 );
and ( n10122 , n10120 , n10121 );
not ( n10123 , n6887 );
not ( n10124 , n10123 );
nor ( n10125 , n10122 , n10124 );
not ( n10126 , n10125 );
or ( n10127 , n10103 , n10126 );
or ( n10128 , n10102 , n10125 );
nand ( n10129 , n10127 , n10128 );
nand ( n10130 , n10101 , n10129 );
not ( n10131 , n10130 );
not ( n10132 , n7089 );
not ( n10133 , n10056 );
nor ( n10134 , n10132 , n10133 );
not ( n10135 , n10134 );
not ( n10136 , n10091 );
or ( n10137 , n10135 , n10136 );
not ( n10138 , n7465 );
nand ( n10139 , n10137 , n10138 );
not ( n10140 , n10134 );
not ( n10141 , n10087 );
or ( n10142 , n10140 , n10141 );
nand ( n10143 , n7459 , n7089 );
nand ( n10144 , n10142 , n10143 );
nor ( n10145 , n10139 , n10144 );
not ( n10146 , n7474 );
not ( n10147 , n10146 );
nand ( n10148 , n10147 , n7117 );
not ( n10149 , n10148 );
and ( n10150 , n10145 , n10149 );
not ( n10151 , n10145 );
and ( n10152 , n10151 , n10148 );
nor ( n10153 , n10150 , n10152 );
not ( n10154 , n10110 );
not ( n10155 , n10112 );
or ( n10156 , n10154 , n10155 );
nand ( n10157 , n10156 , n10119 );
nand ( n10158 , n10123 , n10121 );
and ( n10159 , n10157 , n10158 );
not ( n10160 , n10157 );
not ( n10161 , n10158 );
and ( n10162 , n10160 , n10161 );
nor ( n10163 , n10159 , n10162 );
nor ( n10164 , n10153 , n10163 );
buf ( n10165 , n10164 );
nand ( n10166 , n10084 , n10131 , n10165 );
nand ( n10167 , n7458 , n7452 );
not ( n10168 , n10167 );
or ( n10169 , n7159 , n7160 );
nand ( n10170 , n7401 , n7416 , n10169 );
not ( n10171 , n10170 );
not ( n10172 , n10043 );
nand ( n10173 , n10029 , n8959 );
not ( n10174 , n10047 );
and ( n10175 , n10173 , n10174 , n10045 );
not ( n10176 , n10006 );
not ( n10177 , n10014 );
or ( n10178 , n10176 , n10177 );
not ( n10179 , n9237 );
nor ( n10180 , n10179 , n8960 , n9286 );
nand ( n10181 , n10178 , n10180 );
nand ( n10182 , n10175 , n10181 , n10036 );
or ( n10183 , n10172 , n10182 );
nand ( n10184 , n8569 , n8588 , n8592 );
and ( n10185 , n8249 , n10043 );
nor ( n10186 , n10185 , n8085 );
nand ( n10187 , n10184 , n10186 );
not ( n10188 , n10187 );
nand ( n10189 , n10183 , n10188 );
not ( n10190 , n10189 );
not ( n10191 , n10106 );
or ( n10192 , n10190 , n10191 );
nand ( n10193 , n10192 , n10115 );
not ( n10194 , n10193 );
or ( n10195 , n10171 , n10194 );
not ( n10196 , n7418 );
nand ( n10197 , n10195 , n10196 );
not ( n10198 , n10197 );
or ( n10199 , n10168 , n10198 );
or ( n10200 , n10197 , n10167 );
nand ( n10201 , n10199 , n10200 );
and ( n10202 , n7089 , n10138 );
not ( n10203 , n10202 );
not ( n10204 , n10187 );
not ( n10205 , n8734 );
not ( n10206 , n10205 );
or ( n10207 , n10204 , n10206 );
nand ( n10208 , n10207 , n8834 );
not ( n10209 , n8835 );
and ( n10210 , n10208 , n10209 );
nor ( n10211 , n10210 , n8847 );
or ( n10212 , n10211 , n10133 );
nand ( n10213 , n10212 , n10108 );
not ( n10214 , n10104 );
and ( n10215 , n10056 , n10214 , n10106 , n10050 );
nor ( n10216 , n10213 , n10215 );
not ( n10217 , n10216 );
or ( n10218 , n10203 , n10217 );
or ( n10219 , n10216 , n10202 );
nand ( n10220 , n10218 , n10219 );
nand ( n10221 , n10201 , n10220 );
not ( n10222 , n10221 );
buf ( n10223 , n8250 );
nand ( n10224 , n10223 , n8589 );
not ( n10225 , n10224 );
nand ( n10226 , n10225 , n10182 );
not ( n10227 , n10172 );
nand ( n10228 , n10227 , n8086 );
not ( n10229 , n10228 );
and ( n10230 , n10226 , n10229 );
not ( n10231 , n10226 );
and ( n10232 , n10231 , n10228 );
nor ( n10233 , n10230 , n10232 );
not ( n10234 , n10233 );
buf ( n10235 , n10189 );
not ( n10236 , n10235 );
not ( n10237 , n8733 );
not ( n10238 , n10237 );
buf ( n10239 , n8826 );
nand ( n10240 , n10238 , n10239 );
not ( n10241 , n10240 );
and ( n10242 , n10236 , n10241 );
buf ( n10243 , n10235 );
and ( n10244 , n10243 , n10240 );
nor ( n10245 , n10242 , n10244 );
nor ( n10246 , n10234 , n10245 );
and ( n10247 , n10174 , n10173 );
not ( n10248 , n10247 );
not ( n10249 , n10181 );
or ( n10250 , n10248 , n10249 );
not ( n10251 , n8527 );
nand ( n10252 , n10250 , n10251 );
nand ( n10253 , n10045 , n8568 );
xnor ( n10254 , n10252 , n10253 );
buf ( n10255 , n10032 );
not ( n10256 , n10255 );
nand ( n10257 , n10174 , n10251 );
not ( n10258 , n10257 );
or ( n10259 , n10256 , n10258 );
buf ( n10260 , n10255 );
or ( n10261 , n10260 , n10257 );
nand ( n10262 , n10259 , n10261 );
not ( n10263 , n10006 );
not ( n10264 , n10263 );
not ( n10265 , n9191 );
nand ( n10266 , n9162 , n8984 , n9002 );
nor ( n10267 , n10265 , n10266 );
not ( n10268 , n10267 );
buf ( n10269 , n9192 );
not ( n10270 , n10269 );
nand ( n10271 , n10268 , n10270 );
not ( n10272 , n10271 );
not ( n10273 , n10272 );
or ( n10274 , n10264 , n10273 );
nand ( n10275 , n10006 , n10271 );
nand ( n10276 , n10274 , n10275 );
not ( n10277 , n9419 );
and ( n10278 , n10000 , n9978 , n9991 );
not ( n10279 , n10003 );
or ( n10280 , n10278 , n10279 );
not ( n10281 , n9563 );
nand ( n10282 , n10280 , n10281 );
not ( n10283 , n10282 );
or ( n10284 , n10277 , n10283 );
not ( n10285 , n9566 );
nand ( n10286 , n10284 , n10285 );
not ( n10287 , n10286 );
not ( n10288 , n9601 );
nand ( n10289 , n10288 , n9604 );
not ( n10290 , n10289 );
or ( n10291 , n10287 , n10290 );
or ( n10292 , n10286 , n10289 );
nand ( n10293 , n10291 , n10292 );
not ( n10294 , n10293 );
not ( n10295 , n16 );
nand ( n10296 , n9499 , n9560 );
and ( n10297 , n10296 , n10002 );
and ( n10298 , n10297 , n10278 );
not ( n10299 , n10297 );
and ( n10300 , n10299 , n10001 );
nor ( n10301 , n10298 , n10300 );
nand ( n10302 , n10295 , n10301 );
not ( n10303 , n10302 );
not ( n10304 , n18 );
nand ( n10305 , n9668 , n9643 , n9695 );
not ( n10306 , n10305 );
not ( n10307 , n9839 );
or ( n10308 , n10306 , n10307 );
nand ( n10309 , n10308 , n9987 );
not ( n10310 , n10309 );
nand ( n10311 , n9983 , n9895 );
not ( n10312 , n10311 );
or ( n10313 , n10310 , n10312 );
or ( n10314 , n10309 , n10311 );
nand ( n10315 , n10313 , n10314 );
and ( n10316 , n19 , n10315 );
not ( n10317 , n10316 );
or ( n10318 , n10304 , n10317 );
and ( n10319 , n10316 , n18 );
not ( n10320 , n10316 );
and ( n10321 , n10320 , n1187 );
nor ( n10322 , n10319 , n10321 );
not ( n10323 , n9990 );
nand ( n10324 , n9896 , n10323 );
not ( n10325 , n10324 );
not ( n10326 , n9996 );
nand ( n10327 , n10326 , n9977 );
not ( n10328 , n10327 );
or ( n10329 , n10325 , n10328 );
or ( n10330 , n10324 , n10327 );
nand ( n10331 , n10329 , n10330 );
nand ( n10332 , n10322 , n10331 );
nand ( n10333 , n10318 , n10332 );
not ( n10334 , n10333 );
nand ( n10335 , n9977 , n9897 );
not ( n10336 , n10335 );
not ( n10337 , n9977 );
not ( n10338 , n9990 );
or ( n10339 , n10337 , n10338 );
not ( n10340 , n9996 );
nand ( n10341 , n10339 , n10340 );
or ( n10342 , n10336 , n10341 );
not ( n10343 , n9994 );
nor ( n10344 , n10343 , n9999 );
not ( n10345 , n10344 );
nand ( n10346 , n10342 , n10345 );
not ( n10347 , n10341 );
nand ( n10348 , n10347 , n10344 , n10335 );
nand ( n10349 , n9792 , n10346 , n10348 );
not ( n10350 , n10349 );
or ( n10351 , n10334 , n10350 );
nand ( n10352 , n10346 , n10348 );
nand ( n10353 , n17 , n10352 );
nand ( n10354 , n10351 , n10353 );
not ( n10355 , n10354 );
or ( n10356 , n10303 , n10355 );
not ( n10357 , n10301 );
nand ( n10358 , n16 , n10357 );
nand ( n10359 , n10356 , n10358 );
nand ( n10360 , n10285 , n9419 );
not ( n10361 , n10360 );
not ( n10362 , n10282 );
or ( n10363 , n10361 , n10362 );
not ( n10364 , n10360 );
not ( n10365 , n10282 );
nand ( n10366 , n10364 , n10365 );
nand ( n10367 , n10363 , n10366 );
not ( n10368 , n10001 );
not ( n10369 , n10002 );
or ( n10370 , n10368 , n10369 );
nand ( n10371 , n10370 , n10296 );
nand ( n10372 , n9485 , n9487 );
not ( n10373 , n10372 );
and ( n10374 , n10371 , n10373 );
not ( n10375 , n10371 );
and ( n10376 , n10375 , n10372 );
nor ( n10377 , n10374 , n10376 );
nand ( n10378 , n10359 , n10367 , n10377 );
nor ( n10379 , n10294 , n10378 );
and ( n10380 , n10276 , n10379 );
not ( n10381 , n9255 );
and ( n10382 , n10018 , n9278 );
nand ( n10383 , n10381 , n10382 );
and ( n10384 , n10383 , n10014 );
buf ( n10385 , n9605 );
buf ( n10386 , n10385 );
and ( n10387 , n10384 , n10386 );
not ( n10388 , n9280 );
nor ( n10389 , n10387 , n10388 );
nand ( n10390 , n9237 , n9285 );
nand ( n10391 , n10390 , n10383 );
not ( n10392 , n10005 );
nand ( n10393 , n10384 , n10392 );
nand ( n10394 , n10389 , n10391 , n10393 );
not ( n10395 , n10028 );
not ( n10396 , n10395 );
nand ( n10397 , n10396 , n8959 );
not ( n10398 , n10397 );
and ( n10399 , n10394 , n10398 );
not ( n10400 , n10394 );
and ( n10401 , n10400 , n10397 );
nor ( n10402 , n10399 , n10401 );
not ( n10403 , n10267 );
not ( n10404 , n10004 );
not ( n10405 , n10404 );
nand ( n10406 , n10403 , n10405 , n10001 );
not ( n10407 , n10269 );
and ( n10408 , n10406 , n10407 );
not ( n10409 , n10408 );
not ( n10410 , n10267 );
nand ( n10411 , n10385 , n10410 );
not ( n10412 , n10012 );
not ( n10413 , n9285 );
nor ( n10414 , n10412 , n10413 );
and ( n10415 , n10411 , n10414 );
not ( n10416 , n10415 );
or ( n10417 , n10409 , n10416 );
nand ( n10418 , n10406 , n10411 , n10407 );
not ( n10419 , n10414 );
nand ( n10420 , n10418 , n10419 );
nand ( n10421 , n10417 , n10420 );
not ( n10422 , n10421 );
nor ( n10423 , n10013 , n10278 , n10404 );
not ( n10424 , n10423 );
not ( n10425 , n10390 );
nand ( n10426 , n10410 , n10385 , n10012 );
nand ( n10427 , n10424 , n10425 , n10426 );
nand ( n10428 , n9280 , n10383 );
and ( n10429 , n10427 , n10428 );
not ( n10430 , n10427 );
not ( n10431 , n10428 );
and ( n10432 , n10430 , n10431 );
nor ( n10433 , n10429 , n10432 );
nor ( n10434 , n10422 , n10433 );
nand ( n10435 , n10380 , n10402 , n10434 );
not ( n10436 , n10435 );
and ( n10437 , n10254 , n10262 , n10436 );
not ( n10438 , n10048 );
not ( n10439 , n10173 );
nor ( n10440 , n10438 , n10439 );
not ( n10441 , n10440 );
not ( n10442 , n10181 );
or ( n10443 , n10441 , n10442 );
not ( n10444 , n8569 );
nand ( n10445 , n10443 , n10444 );
not ( n10446 , n10445 );
not ( n10447 , n10036 );
not ( n10448 , n10447 );
nand ( n10449 , n10448 , n10223 );
not ( n10450 , n10449 );
or ( n10451 , n10446 , n10450 );
or ( n10452 , n10445 , n10449 );
nand ( n10453 , n10451 , n10452 );
and ( n10454 , n10246 , n10437 , n10453 );
not ( n10455 , n10255 );
not ( n10456 , n10205 );
not ( n10457 , n10050 );
nor ( n10458 , n10456 , n10457 );
not ( n10459 , n10458 );
or ( n10460 , n10455 , n10459 );
not ( n10461 , n10208 );
nand ( n10462 , n10460 , n10461 );
not ( n10463 , n8816 );
not ( n10464 , n10463 );
not ( n10465 , n8837 );
nand ( n10466 , n10464 , n10465 );
not ( n10467 , n10466 );
and ( n10468 , n10462 , n10467 );
not ( n10469 , n10462 );
and ( n10470 , n10469 , n10466 );
nor ( n10471 , n10468 , n10470 );
not ( n10472 , n10471 );
not ( n10473 , n8832 );
nor ( n10474 , n10473 , n8828 );
not ( n10475 , n10237 );
not ( n10476 , n10475 );
not ( n10477 , n10032 );
not ( n10478 , n10050 );
or ( n10479 , n10477 , n10478 );
nand ( n10480 , n10479 , n10188 );
not ( n10481 , n10480 );
or ( n10482 , n10476 , n10481 );
buf ( n10483 , n10239 );
nand ( n10484 , n10482 , n10483 );
not ( n10485 , n10484 );
and ( n10486 , n10474 , n10485 );
not ( n10487 , n10474 );
and ( n10488 , n10487 , n10484 );
nor ( n10489 , n10486 , n10488 );
nor ( n10490 , n10472 , n10489 );
buf ( n10491 , n10490 );
nand ( n10492 , n10454 , n10491 );
not ( n10493 , n10492 );
nand ( n10494 , n10196 , n10170 );
buf ( n10495 , n10494 );
not ( n10496 , n10495 );
and ( n10497 , n10052 , n10496 );
not ( n10498 , n10052 );
and ( n10499 , n10498 , n10495 );
nor ( n10500 , n10497 , n10499 );
nand ( n10501 , n10187 , n10205 );
not ( n10502 , n10501 );
not ( n10503 , n8834 );
or ( n10504 , n10502 , n10503 );
nand ( n10505 , n10504 , n10464 );
and ( n10506 , n10205 , n10050 );
not ( n10507 , n10463 );
nand ( n10508 , n10506 , n10255 , n10507 );
nand ( n10509 , n10505 , n10508 , n10465 );
nand ( n10510 , n8846 , n8839 );
and ( n10511 , n10509 , n10510 );
not ( n10512 , n10509 );
not ( n10513 , n10510 );
and ( n10514 , n10512 , n10513 );
nor ( n10515 , n10511 , n10514 );
buf ( n10516 , n10515 );
nor ( n10517 , n10500 , n10516 );
nand ( n10518 , n10222 , n10493 , n10517 );
nor ( n10519 , n10166 , n10518 );
and ( n10520 , n3 , n1 );
not ( n10521 , n3 );
and ( n10522 , n10521 , n381 );
nor ( n10523 , n10520 , n10522 );
xnor ( n10524 , n7067 , n10523 );
buf ( n10525 , n10524 );
buf ( n10526 , n10525 );
not ( n10527 , n385 );
nand ( n10528 , n10527 , n10078 );
nor ( n10529 , n10528 , n7478 );
not ( n10530 , n10529 );
or ( n10531 , n10119 , n10530 );
not ( n10532 , n381 );
not ( n10533 , n10064 );
not ( n10534 , n10067 );
and ( n10535 , n10533 , n10534 );
and ( n10536 , n298 , n319 );
nor ( n10537 , n10535 , n10536 );
nor ( n10538 , n10532 , n10537 );
nor ( n10539 , n10538 , n1 );
nand ( n10540 , n10531 , n10539 );
not ( n10541 , n10528 );
not ( n10542 , n10541 );
not ( n10543 , n6891 );
or ( n10544 , n10542 , n10543 );
and ( n10545 , n10078 , n383 );
nor ( n10546 , n10545 , n10076 );
nand ( n10547 , n10544 , n10546 );
not ( n10548 , n10547 );
buf ( n10549 , n10088 );
nand ( n10550 , n10549 , n10058 , n10529 );
nand ( n10551 , n7475 , n10529 );
nand ( n10552 , n10548 , n10550 , n10551 );
nor ( n10553 , n10540 , n10552 );
nand ( n10554 , n10526 , n10553 );
or ( n10555 , n10519 , n10554 );
not ( n10556 , n1503 );
not ( n10557 , n10556 );
not ( n10558 , n3898 );
not ( n10559 , n3853 );
not ( n10560 , n10559 );
or ( n10561 , n10558 , n10560 );
not ( n10562 , n1499 );
not ( n10563 , n1665 );
and ( n10564 , n10562 , n10563 );
not ( n10565 , n2721 );
not ( n10566 , n2769 );
and ( n10567 , n10565 , n10566 );
and ( n10568 , n1759 , n2769 );
nor ( n10569 , n10567 , n10568 );
nor ( n10570 , n10564 , n10569 );
nand ( n10571 , n10561 , n10570 );
buf ( n10572 , n10571 );
not ( n10573 , n10572 );
not ( n10574 , n10573 );
not ( n10575 , n10574 );
and ( n10576 , n10557 , n10575 );
not ( n10577 , n3898 );
not ( n10578 , n10577 );
not ( n10579 , n37 );
and ( n10580 , n10578 , n10579 );
not ( n10581 , n10578 );
and ( n10582 , n10581 , n37 );
nor ( n10583 , n10580 , n10582 );
buf ( n10584 , n10569 );
buf ( n10585 , n10584 );
not ( n10586 , n10585 );
not ( n10587 , n10586 );
and ( n10588 , n10583 , n10587 );
nor ( n10589 , n10576 , n10588 );
not ( n10590 , n10589 );
not ( n10591 , n1521 );
not ( n10592 , n3752 );
not ( n10593 , n10592 );
not ( n10594 , n1820 );
not ( n10595 , n10594 );
nand ( n10596 , n10593 , n10595 );
nand ( n10597 , n10594 , n3753 );
not ( n10598 , n1499 );
not ( n10599 , n3752 );
or ( n10600 , n10598 , n10599 );
not ( n10601 , n1499 );
nand ( n10602 , n10601 , n3751 );
nand ( n10603 , n10600 , n10602 );
and ( n10604 , n10596 , n10597 , n10603 );
not ( n10605 , n10604 );
or ( n10606 , n10591 , n10605 );
buf ( n10607 , n3774 );
buf ( n10608 , n10607 );
and ( n10609 , n39 , n10608 );
not ( n10610 , n39 );
not ( n10611 , n1820 );
not ( n10612 , n10611 );
not ( n10613 , n10612 );
not ( n10614 , n10613 );
and ( n10615 , n10610 , n10614 );
nor ( n10616 , n10609 , n10615 );
not ( n10617 , n10603 );
not ( n10618 , n10617 );
not ( n10619 , n10618 );
nand ( n10620 , n10616 , n10619 );
nand ( n10621 , n10606 , n10620 );
not ( n10622 , n506 );
not ( n10623 , n10622 );
nand ( n10624 , n10623 , n45 );
xor ( n10625 , n10621 , n10624 );
or ( n10626 , n10590 , n10625 );
not ( n10627 , n10621 );
or ( n10628 , n10624 , n10627 );
nand ( n10629 , n10626 , n10628 );
not ( n10630 , n10583 );
not ( n10631 , n10571 );
not ( n10632 , n10631 );
or ( n10633 , n10630 , n10632 );
not ( n10634 , n3900 );
not ( n10635 , n3898 );
not ( n10636 , n10635 );
and ( n10637 , n497 , n10636 );
nor ( n10638 , n10634 , n10637 );
nand ( n10639 , n10638 , n10585 );
nand ( n10640 , n10633 , n10639 );
not ( n10641 , n1061 );
not ( n10642 , n10641 );
not ( n10643 , n2892 );
and ( n10644 , n10642 , n10643 );
and ( n10645 , n1686 , n970 );
nor ( n10646 , n10644 , n10645 );
buf ( n10647 , n10646 );
not ( n10648 , n10647 );
not ( n10649 , n10648 );
buf ( n10650 , n2721 );
not ( n10651 , n10650 );
not ( n10652 , n1688 );
or ( n10653 , n10651 , n10652 );
not ( n10654 , n10650 );
and ( n10655 , n10654 , n1687 );
nor ( n10656 , n10655 , n10646 );
nand ( n10657 , n10653 , n10656 );
not ( n10658 , n10657 );
not ( n10659 , n10658 );
not ( n10660 , n10659 );
or ( n10661 , n10649 , n10660 );
not ( n10662 , n10650 );
buf ( n10663 , n10662 );
not ( n10664 , n10663 );
nand ( n10665 , n10661 , n10664 );
xor ( n10666 , n10640 , n10665 );
and ( n10667 , n41 , n557 );
not ( n10668 , n41 );
not ( n10669 , n556 );
not ( n10670 , n10669 );
and ( n10671 , n10668 , n10670 );
nor ( n10672 , n10667 , n10671 );
or ( n10673 , n591 , n605 );
nand ( n10674 , n591 , n605 );
not ( n10675 , n605 );
nand ( n10676 , n10675 , n1820 );
nand ( n10677 , n3708 , n10611 );
nand ( n10678 , n10676 , n10677 );
and ( n10679 , n10673 , n10674 , n10678 );
buf ( n10680 , n10679 );
and ( n10681 , n10672 , n10680 );
and ( n10682 , n40 , n557 );
and ( n10683 , n647 , n592 );
nor ( n10684 , n10682 , n10683 );
not ( n10685 , n10684 );
not ( n10686 , n10678 );
buf ( n10687 , n10686 );
not ( n10688 , n10687 );
nor ( n10689 , n10685 , n10688 );
nor ( n10690 , n10681 , n10689 );
not ( n10691 , n10690 );
and ( n10692 , n10666 , n10691 );
not ( n10693 , n10666 );
and ( n10694 , n10693 , n10690 );
nor ( n10695 , n10692 , n10694 );
xnor ( n10696 , n10629 , n10695 );
not ( n10697 , n10696 );
or ( n10698 , n43 , n610 );
not ( n10699 , n10622 );
nand ( n10700 , n10699 , n43 );
nand ( n10701 , n10698 , n10700 );
nor ( n10702 , n519 , n10622 );
not ( n10703 , n10702 );
not ( n10704 , n506 );
nand ( n10705 , n519 , n10704 );
not ( n10706 , n3737 );
not ( n10707 , n10706 );
not ( n10708 , n556 );
or ( n10709 , n10707 , n10708 );
or ( n10710 , n3738 , n556 );
nand ( n10711 , n10709 , n10710 );
nand ( n10712 , n10703 , n10705 , n10711 );
not ( n10713 , n10712 );
not ( n10714 , n10713 );
or ( n10715 , n10701 , n10714 );
not ( n10716 , n532 );
xor ( n10717 , n10716 , n42 );
not ( n10718 , n10711 );
buf ( n10719 , n10718 );
not ( n10720 , n10719 );
or ( n10721 , n10717 , n10720 );
nand ( n10722 , n10715 , n10721 );
not ( n10723 , n10616 );
not ( n10724 , n10604 );
or ( n10725 , n10723 , n10724 );
and ( n10726 , n609 , n10608 );
not ( n10727 , n10608 );
and ( n10728 , n38 , n10727 );
nor ( n10729 , n10726 , n10728 );
not ( n10730 , n10729 );
buf ( n10731 , n10617 );
nand ( n10732 , n10730 , n10731 );
nand ( n10733 , n10725 , n10732 );
xor ( n10734 , n10722 , n10733 );
not ( n10735 , n5894 );
not ( n10736 , n533 );
not ( n10737 , n10736 );
not ( n10738 , n10737 );
not ( n10739 , n10738 );
not ( n10740 , n10739 );
and ( n10741 , n10735 , n10740 );
xnor ( n10742 , n10734 , n10741 );
not ( n10743 , n10742 );
not ( n10744 , n10590 );
not ( n10745 , n1478 );
not ( n10746 , n10659 );
not ( n10747 , n10746 );
or ( n10748 , n10745 , n10747 );
not ( n10749 , n10664 );
not ( n10750 , n10648 );
not ( n10751 , n10750 );
or ( n10752 , n10749 , n10751 );
nand ( n10753 , n10748 , n10752 );
not ( n10754 , n10753 );
not ( n10755 , n10701 );
not ( n10756 , n10719 );
not ( n10757 , n10756 );
and ( n10758 , n10755 , n10757 );
not ( n10759 , n10735 );
not ( n10760 , n533 );
or ( n10761 , n10759 , n10760 );
nand ( n10762 , n10761 , n1529 );
not ( n10763 , n10712 );
and ( n10764 , n10762 , n10763 );
nor ( n10765 , n10758 , n10764 );
not ( n10766 , n42 );
not ( n10767 , n10766 );
not ( n10768 , n10669 );
not ( n10769 , n10768 );
not ( n10770 , n10769 );
or ( n10771 , n10767 , n10770 );
nand ( n10772 , n10771 , n1487 );
not ( n10773 , n10772 );
not ( n10774 , n10679 );
or ( n10775 , n10773 , n10774 );
nand ( n10776 , n10672 , n10687 );
nand ( n10777 , n10775 , n10776 );
xnor ( n10778 , n10765 , n10777 );
not ( n10779 , n10778 );
or ( n10780 , n10754 , n10779 );
not ( n10781 , n10765 );
nand ( n10782 , n10781 , n10777 );
nand ( n10783 , n10780 , n10782 );
not ( n10784 , n10783 );
not ( n10785 , n10784 );
or ( n10786 , n10744 , n10785 );
nand ( n10787 , n10589 , n10783 );
nand ( n10788 , n10786 , n10787 );
not ( n10789 , n10788 );
or ( n10790 , n10743 , n10789 );
or ( n10791 , n10742 , n10788 );
nand ( n10792 , n10790 , n10791 );
not ( n10793 , n10792 );
not ( n10794 , n10793 );
and ( n10795 , n10697 , n10794 );
and ( n10796 , n10629 , n10695 );
nor ( n10797 , n10795 , n10796 );
not ( n10798 , n10589 );
not ( n10799 , n10784 );
and ( n10800 , n10798 , n10799 );
not ( n10801 , n10742 );
and ( n10802 , n10801 , n10788 );
nor ( n10803 , n10800 , n10802 );
and ( n10804 , n10741 , n10734 );
and ( n10805 , n10722 , n10733 );
nor ( n10806 , n10804 , n10805 );
and ( n10807 , n10684 , n10680 );
and ( n10808 , n39 , n10769 );
and ( n10809 , n10610 , n10670 );
nor ( n10810 , n10808 , n10809 );
not ( n10811 , n10688 );
and ( n10812 , n10810 , n10811 );
nor ( n10813 , n10807 , n10812 );
not ( n10814 , n10729 );
not ( n10815 , n10604 );
not ( n10816 , n10815 );
and ( n10817 , n10814 , n10816 );
not ( n10818 , n10727 );
and ( n10819 , n37 , n10818 );
and ( n10820 , n10579 , n10727 );
nor ( n10821 , n10819 , n10820 );
not ( n10822 , n10731 );
not ( n10823 , n10822 );
and ( n10824 , n10821 , n10823 );
nor ( n10825 , n10817 , n10824 );
and ( n10826 , n10813 , n10825 );
not ( n10827 , n10813 );
not ( n10828 , n10825 );
and ( n10829 , n10827 , n10828 );
nor ( n10830 , n10826 , n10829 );
xnor ( n10831 , n10806 , n10830 );
not ( n10832 , n10638 );
or ( n10833 , n10832 , n10572 );
buf ( n10834 , n10636 );
buf ( n10835 , n10584 );
not ( n10836 , n10835 );
or ( n10837 , n10834 , n10836 );
nand ( n10838 , n10833 , n10837 );
not ( n10839 , n10717 );
not ( n10840 , n10839 );
not ( n10841 , n10763 );
or ( n10842 , n10840 , n10841 );
not ( n10843 , n532 );
nor ( n10844 , n669 , n10843 );
not ( n10845 , n10844 );
nand ( n10846 , n669 , n10704 );
nand ( n10847 , n10845 , n10846 );
not ( n10848 , n10847 );
nand ( n10849 , n10848 , n10719 );
nand ( n10850 , n10842 , n10849 );
not ( n10851 , n10700 );
and ( n10852 , n10850 , n10851 );
not ( n10853 , n10850 );
and ( n10854 , n10853 , n10700 );
nor ( n10855 , n10852 , n10854 );
xor ( n10856 , n10838 , n10855 );
not ( n10857 , n10691 );
not ( n10858 , n10666 );
or ( n10859 , n10857 , n10858 );
nand ( n10860 , n10665 , n10640 );
nand ( n10861 , n10859 , n10860 );
not ( n10862 , n10861 );
and ( n10863 , n10856 , n10862 );
not ( n10864 , n10856 );
and ( n10865 , n10864 , n10861 );
nor ( n10866 , n10863 , n10865 );
not ( n10867 , n10866 );
and ( n10868 , n10831 , n10867 );
not ( n10869 , n10831 );
and ( n10870 , n10869 , n10866 );
nor ( n10871 , n10868 , n10870 );
xnor ( n10872 , n10803 , n10871 );
xnor ( n10873 , n10797 , n10872 );
xor ( n10874 , n10778 , n10753 );
not ( n10875 , n4300 );
not ( n10876 , n10716 );
or ( n10877 , n10875 , n10876 );
nand ( n10878 , n10877 , n10624 );
not ( n10879 , n10763 );
or ( n10880 , n10878 , n10879 );
not ( n10881 , n10762 );
or ( n10882 , n10881 , n10720 );
nand ( n10883 , n10880 , n10882 );
not ( n10884 , n10883 );
not ( n10885 , n10556 );
not ( n10886 , n10586 );
and ( n10887 , n10885 , n10886 );
and ( n10888 , n10610 , n3898 );
not ( n10889 , n10610 );
not ( n10890 , n3898 );
and ( n10891 , n10889 , n10890 );
nor ( n10892 , n10888 , n10891 );
and ( n10893 , n10892 , n10573 );
nor ( n10894 , n10887 , n10893 );
not ( n10895 , n10894 );
not ( n10896 , n43 );
not ( n10897 , n10768 );
and ( n10898 , n10896 , n10897 );
and ( n10899 , n43 , n10670 );
nor ( n10900 , n10898 , n10899 );
not ( n10901 , n10900 );
not ( n10902 , n10901 );
not ( n10903 , n10680 );
or ( n10904 , n10902 , n10903 );
nand ( n10905 , n10772 , n10687 );
nand ( n10906 , n10904 , n10905 );
not ( n10907 , n10906 );
or ( n10908 , n10895 , n10907 );
or ( n10909 , n10894 , n10906 );
nand ( n10910 , n10908 , n10909 );
not ( n10911 , n10910 );
or ( n10912 , n10884 , n10911 );
not ( n10913 , n10894 );
nand ( n10914 , n10913 , n10906 );
nand ( n10915 , n10912 , n10914 );
not ( n10916 , n3774 );
not ( n10917 , n10916 );
and ( n10918 , n41 , n10917 );
and ( n10919 , n669 , n10614 );
nor ( n10920 , n10918 , n10919 );
buf ( n10921 , n10604 );
and ( n10922 , n10920 , n10921 );
and ( n10923 , n1521 , n10823 );
nor ( n10924 , n10922 , n10923 );
not ( n10925 , n987 );
not ( n10926 , n10925 );
not ( n10927 , n3100 );
not ( n10928 , n10927 );
or ( n10929 , n10926 , n10928 );
not ( n10930 , n987 );
or ( n10931 , n10930 , n3374 );
nand ( n10932 , n10929 , n10931 );
not ( n10933 , n10932 );
buf ( n10934 , n10933 );
not ( n10935 , n10934 );
nor ( n10936 , n2892 , n10930 );
not ( n10937 , n10936 );
nand ( n10938 , n970 , n10930 );
nand ( n10939 , n10937 , n10932 , n10938 );
not ( n10940 , n10939 );
not ( n10941 , n10940 );
and ( n10942 , n10935 , n10941 );
not ( n10943 , n1575 );
not ( n10944 , n10943 );
nor ( n10945 , n10942 , n10944 );
and ( n10946 , n10663 , n10579 );
not ( n10947 , n10663 );
and ( n10948 , n10947 , n37 );
nor ( n10949 , n10946 , n10948 );
and ( n10950 , n10949 , n10746 );
not ( n10951 , n10647 );
nor ( n10952 , n10745 , n10951 );
nor ( n10953 , n10950 , n10952 );
xnor ( n10954 , n10945 , n10953 );
or ( n10955 , n10924 , n10954 );
or ( n10956 , n10945 , n10953 );
nand ( n10957 , n10955 , n10956 );
xor ( n10958 , n10915 , n10957 );
and ( n10959 , n10874 , n10958 );
and ( n10960 , n10957 , n10915 );
nor ( n10961 , n10959 , n10960 );
not ( n10962 , n10961 );
and ( n10963 , n10696 , n10792 );
not ( n10964 , n10696 );
and ( n10965 , n10964 , n10793 );
nor ( n10966 , n10963 , n10965 );
not ( n10967 , n10966 );
and ( n10968 , n10962 , n10967 );
and ( n10969 , n10625 , n10589 );
not ( n10970 , n10625 );
and ( n10971 , n10970 , n10590 );
nor ( n10972 , n10969 , n10971 );
and ( n10973 , n46 , n10738 );
not ( n10974 , n975 );
not ( n10975 , n10939 );
not ( n10976 , n10975 );
or ( n10977 , n10974 , n10976 );
buf ( n10978 , n10933 );
not ( n10979 , n10978 );
or ( n10980 , n10944 , n10979 );
nand ( n10981 , n10977 , n10980 );
not ( n10982 , n10981 );
and ( n10983 , n10973 , n10982 );
not ( n10984 , n10973 );
and ( n10985 , n10984 , n10981 );
nor ( n10986 , n10983 , n10985 );
not ( n10987 , n10986 );
not ( n10988 , n556 );
and ( n10989 , n10735 , n10988 );
and ( n10990 , n5894 , n592 );
nor ( n10991 , n10989 , n10990 );
not ( n10992 , n10991 );
not ( n10993 , n10679 );
or ( n10994 , n10992 , n10993 );
not ( n10995 , n10687 );
or ( n10996 , n10900 , n10995 );
nand ( n10997 , n10994 , n10996 );
not ( n10998 , n1030 );
not ( n10999 , n10659 );
not ( n11000 , n10999 );
or ( n11001 , n10998 , n11000 );
not ( n11002 , n10647 );
not ( n11003 , n11002 );
nand ( n11004 , n10949 , n11003 );
nand ( n11005 , n11001 , n11004 );
not ( n11006 , n10916 );
xor ( n11007 , n11006 , n42 );
not ( n11008 , n11007 );
not ( n11009 , n10921 );
or ( n11010 , n11008 , n11009 );
nand ( n11011 , n10920 , n10731 );
nand ( n11012 , n11010 , n11011 );
xor ( n11013 , n11005 , n11012 );
and ( n11014 , n10997 , n11013 );
and ( n11015 , n11005 , n11012 );
nor ( n11016 , n11014 , n11015 );
not ( n11017 , n11016 );
and ( n11018 , n10987 , n11017 );
and ( n11019 , n10973 , n10981 );
nor ( n11020 , n11018 , n11019 );
xnor ( n11021 , n10972 , n11020 );
xor ( n11022 , n10954 , n10924 );
or ( n11023 , n4266 , n10622 );
not ( n11024 , n40 );
not ( n11025 , n3898 );
or ( n11026 , n11024 , n11025 );
nand ( n11027 , n11026 , n648 );
and ( n11028 , n11027 , n10631 );
and ( n11029 , n10892 , n10835 );
nor ( n11030 , n11028 , n11029 );
not ( n11031 , n11030 );
not ( n11032 , n742 );
not ( n11033 , n10763 );
or ( n11034 , n11032 , n11033 );
not ( n11035 , n10878 );
nand ( n11036 , n11035 , n10719 );
nand ( n11037 , n11034 , n11036 );
not ( n11038 , n11037 );
and ( n11039 , n11031 , n11038 );
and ( n11040 , n11030 , n11037 );
nor ( n11041 , n11039 , n11040 );
or ( n11042 , n11023 , n11041 );
not ( n11043 , n11037 );
or ( n11044 , n11030 , n11043 );
nand ( n11045 , n11042 , n11044 );
xor ( n11046 , n10883 , n10910 );
xor ( n11047 , n11045 , n11046 );
and ( n11048 , n11022 , n11047 );
and ( n11049 , n11045 , n11046 );
nor ( n11050 , n11048 , n11049 );
or ( n11051 , n11021 , n11050 );
or ( n11052 , n10972 , n11020 );
nand ( n11053 , n11051 , n11052 );
xor ( n11054 , n10961 , n10966 );
and ( n11055 , n11053 , n11054 );
nor ( n11056 , n10968 , n11055 );
nand ( n11057 , n10873 , n11056 );
not ( n11058 , n11053 );
and ( n11059 , n11054 , n11058 );
not ( n11060 , n11054 );
and ( n11061 , n11060 , n11053 );
nor ( n11062 , n11059 , n11061 );
xnor ( n11063 , n10874 , n10958 );
not ( n11064 , n11063 );
not ( n11065 , n11050 );
and ( n11066 , n11021 , n11065 );
not ( n11067 , n11021 );
and ( n11068 , n11067 , n11050 );
nor ( n11069 , n11066 , n11068 );
not ( n11070 , n11069 );
and ( n11071 , n11064 , n11070 );
xor ( n11072 , n11013 , n10997 );
or ( n11073 , n47 , n610 );
nand ( n11074 , n11073 , n11023 );
or ( n11075 , n11074 , n10879 );
not ( n11076 , n742 );
or ( n11077 , n11076 , n10720 );
nand ( n11078 , n11075 , n11077 );
not ( n11079 , n11078 );
nand ( n11080 , n1030 , n11003 );
and ( n11081 , n10663 , n10610 );
not ( n11082 , n10663 );
and ( n11083 , n11082 , n39 );
nor ( n11084 , n11081 , n11083 );
buf ( n11085 , n10658 );
nand ( n11086 , n11084 , n11085 );
and ( n11087 , n11080 , n11086 );
and ( n11088 , n45 , n557 );
and ( n11089 , n4300 , n592 );
nor ( n11090 , n11088 , n11089 );
not ( n11091 , n11090 );
and ( n11092 , n10673 , n10674 , n10678 );
not ( n11093 , n11092 );
or ( n11094 , n11091 , n11093 );
nand ( n11095 , n10991 , n10687 );
nand ( n11096 , n11094 , n11095 );
xor ( n11097 , n11087 , n11096 );
or ( n11098 , n11079 , n11097 );
not ( n11099 , n11096 );
or ( n11100 , n11087 , n11099 );
nand ( n11101 , n11098 , n11100 );
xor ( n11102 , n11041 , n11023 );
xor ( n11103 , n11101 , n11102 );
and ( n11104 , n11072 , n11103 );
and ( n11105 , n11101 , n11102 );
nor ( n11106 , n11104 , n11105 );
not ( n11107 , n11016 );
and ( n11108 , n10986 , n11107 );
not ( n11109 , n10986 );
and ( n11110 , n11109 , n11016 );
nor ( n11111 , n11108 , n11110 );
not ( n11112 , n2790 );
buf ( n11113 , n11112 );
not ( n11114 , n11113 );
and ( n11115 , n2790 , n3377 );
not ( n11116 , n11115 );
and ( n11117 , n11114 , n11116 );
buf ( n11118 , n3377 );
buf ( n11119 , n11118 );
not ( n11120 , n11119 );
nor ( n11121 , n11117 , n11120 );
not ( n11122 , n10974 );
not ( n11123 , n10979 );
and ( n11124 , n11122 , n11123 );
not ( n11125 , n1575 );
and ( n11126 , n10579 , n11125 );
not ( n11127 , n10579 );
buf ( n11128 , n970 );
not ( n11129 , n11128 );
and ( n11130 , n11127 , n11129 );
nor ( n11131 , n11126 , n11130 );
not ( n11132 , n11131 );
and ( n11133 , n11132 , n10940 );
nor ( n11134 , n11124 , n11133 );
nand ( n11135 , n11121 , n11134 );
and ( n11136 , n11135 , n10982 );
not ( n11137 , n11135 );
and ( n11138 , n11137 , n10981 );
nor ( n11139 , n11136 , n11138 );
and ( n11140 , n43 , n10917 );
and ( n11141 , n10896 , n10916 );
nor ( n11142 , n11140 , n11141 );
and ( n11143 , n11142 , n10921 );
and ( n11144 , n11007 , n10731 );
nor ( n11145 , n11143 , n11144 );
nand ( n11146 , n48 , n10736 );
and ( n11147 , n3898 , n669 );
not ( n11148 , n3898 );
and ( n11149 , n11148 , n41 );
nor ( n11150 , n11147 , n11149 );
and ( n11151 , n11150 , n10573 );
and ( n11152 , n11027 , n10835 );
nor ( n11153 , n11151 , n11152 );
not ( n11154 , n11153 );
and ( n11155 , n11146 , n11154 );
not ( n11156 , n11146 );
and ( n11157 , n11156 , n11153 );
nor ( n11158 , n11155 , n11157 );
or ( n11159 , n11145 , n11158 );
or ( n11160 , n11146 , n11153 );
nand ( n11161 , n11159 , n11160 );
and ( n11162 , n11139 , n11161 );
and ( n11163 , n10982 , n11135 );
nor ( n11164 , n11162 , n11163 );
not ( n11165 , n11164 );
and ( n11166 , n11111 , n11165 );
not ( n11167 , n11111 );
and ( n11168 , n11167 , n11164 );
nor ( n11169 , n11166 , n11168 );
or ( n11170 , n11106 , n11169 );
or ( n11171 , n11164 , n11111 );
nand ( n11172 , n11170 , n11171 );
xor ( n11173 , n11069 , n11063 );
and ( n11174 , n11172 , n11173 );
nor ( n11175 , n11071 , n11174 );
nor ( n11176 , n11062 , n11175 );
and ( n11177 , n11057 , n11176 );
nor ( n11178 , n10873 , n11056 );
nor ( n11179 , n11177 , n11178 );
not ( n11180 , n10831 );
not ( n11181 , n10866 );
and ( n11182 , n11180 , n11181 );
and ( n11183 , n10856 , n10861 );
nor ( n11184 , n11182 , n11183 );
and ( n11185 , n10810 , n10680 );
or ( n11186 , n609 , n10769 );
nand ( n11187 , n11186 , n3732 );
and ( n11188 , n11187 , n10687 );
nor ( n11189 , n11185 , n11188 );
not ( n11190 , n10739 );
nand ( n11191 , n42 , n11190 );
xor ( n11192 , n11189 , n11191 );
and ( n11193 , n11192 , n10825 );
not ( n11194 , n11192 );
and ( n11195 , n11194 , n10828 );
nor ( n11196 , n11193 , n11195 );
not ( n11197 , n10838 );
not ( n11198 , n10855 );
or ( n11199 , n11197 , n11198 );
nand ( n11200 , n10851 , n10850 );
nand ( n11201 , n11199 , n11200 );
not ( n11202 , n11201 );
not ( n11203 , n10821 );
not ( n11204 , n10921 );
or ( n11205 , n11203 , n11204 );
xor ( n11206 , n36 , n3774 );
nand ( n11207 , n11206 , n10731 );
nand ( n11208 , n11205 , n11207 );
not ( n11209 , n10586 );
not ( n11210 , n10572 );
or ( n11211 , n11209 , n11210 );
not ( n11212 , n10834 );
nand ( n11213 , n11211 , n11212 );
xor ( n11214 , n11208 , n11213 );
or ( n11215 , n10847 , n10879 );
or ( n11216 , n3717 , n10720 );
nand ( n11217 , n11215 , n11216 );
xnor ( n11218 , n11214 , n11217 );
not ( n11219 , n11218 );
or ( n11220 , n11202 , n11219 );
or ( n11221 , n11201 , n11218 );
nand ( n11222 , n11220 , n11221 );
and ( n11223 , n11196 , n11222 );
not ( n11224 , n11196 );
not ( n11225 , n11222 );
and ( n11226 , n11224 , n11225 );
or ( n11227 , n11223 , n11226 );
or ( n11228 , n10830 , n10806 );
or ( n11229 , n10828 , n10813 );
nand ( n11230 , n11228 , n11229 );
xnor ( n11231 , n11227 , n11230 );
xnor ( n11232 , n11184 , n11231 );
or ( n11233 , n10797 , n10872 );
or ( n11234 , n10803 , n10871 );
nand ( n11235 , n11233 , n11234 );
not ( n11236 , n11235 );
and ( n11237 , n11232 , n11236 );
or ( n11238 , n11179 , n11237 );
not ( n11239 , n11232 );
nand ( n11240 , n11239 , n11235 );
nand ( n11241 , n11238 , n11240 );
not ( n11242 , n11241 );
not ( n11243 , n11237 );
nand ( n11244 , n11243 , n11057 );
not ( n11245 , n11244 );
xor ( n11246 , n11158 , n11145 );
or ( n11247 , n11121 , n11134 );
nand ( n11248 , n11247 , n11135 );
not ( n11249 , n11248 );
not ( n11250 , n11249 );
and ( n11251 , n11097 , n11078 );
not ( n11252 , n11097 );
and ( n11253 , n11252 , n11079 );
nor ( n11254 , n11251 , n11253 );
not ( n11255 , n11254 );
not ( n11256 , n11255 );
or ( n11257 , n11250 , n11256 );
nand ( n11258 , n11248 , n11254 );
nand ( n11259 , n11257 , n11258 );
and ( n11260 , n11246 , n11259 );
and ( n11261 , n11248 , n11255 );
nor ( n11262 , n11260 , n11261 );
xnor ( n11263 , n11139 , n11161 );
nand ( n11264 , n11084 , n11003 );
not ( n11265 , n882 );
not ( n11266 , n11265 );
not ( n11267 , n10657 );
nand ( n11268 , n11266 , n11267 );
and ( n11269 , n11264 , n11268 );
and ( n11270 , n46 , n557 );
and ( n11271 , n763 , n592 );
nor ( n11272 , n11270 , n11271 );
not ( n11273 , n11272 );
not ( n11274 , n10679 );
or ( n11275 , n11273 , n11274 );
nand ( n11276 , n11090 , n10687 );
nand ( n11277 , n11275 , n11276 );
not ( n11278 , n11277 );
or ( n11279 , n11269 , n11278 );
not ( n11280 , n11074 );
not ( n11281 , n10720 );
and ( n11282 , n11280 , n11281 );
xnor ( n11283 , n533 , n48 );
not ( n11284 , n10714 );
and ( n11285 , n11283 , n11284 );
nor ( n11286 , n11282 , n11285 );
not ( n11287 , n11286 );
not ( n11288 , n11269 );
not ( n11289 , n11277 );
or ( n11290 , n11288 , n11289 );
or ( n11291 , n11269 , n11277 );
nand ( n11292 , n11290 , n11291 );
nand ( n11293 , n11287 , n11292 );
nand ( n11294 , n11279 , n11293 );
or ( n11295 , n5894 , n3774 );
nand ( n11296 , n11295 , n941 );
not ( n11297 , n11296 );
not ( n11298 , n10921 );
or ( n11299 , n11297 , n11298 );
nand ( n11300 , n11142 , n10731 );
nand ( n11301 , n11299 , n11300 );
not ( n11302 , n11301 );
not ( n11303 , n854 );
not ( n11304 , n10571 );
not ( n11305 , n11304 );
or ( n11306 , n11303 , n11305 );
nand ( n11307 , n11150 , n10584 );
nand ( n11308 , n11306 , n11307 );
nand ( n11309 , n49 , n506 );
not ( n11310 , n11309 );
and ( n11311 , n11308 , n11310 );
not ( n11312 , n11308 );
not ( n11313 , n11310 );
and ( n11314 , n11312 , n11313 );
nor ( n11315 , n11311 , n11314 );
not ( n11316 , n11315 );
or ( n11317 , n11302 , n11316 );
nand ( n11318 , n11310 , n11308 );
nand ( n11319 , n11317 , n11318 );
not ( n11320 , n1335 );
or ( n11321 , n11116 , n11320 );
not ( n11322 , n11113 );
or ( n11323 , n11120 , n11322 );
nand ( n11324 , n11321 , n11323 );
not ( n11325 , n925 );
or ( n11326 , n11325 , n10976 );
or ( n11327 , n11131 , n10979 );
nand ( n11328 , n11326 , n11327 );
and ( n11329 , n11324 , n11328 );
xor ( n11330 , n11319 , n11329 );
and ( n11331 , n11294 , n11330 );
and ( n11332 , n11329 , n11319 );
nor ( n11333 , n11331 , n11332 );
xnor ( n11334 , n11263 , n11333 );
or ( n11335 , n11262 , n11334 );
or ( n11336 , n11263 , n11333 );
nand ( n11337 , n11335 , n11336 );
and ( n11338 , n11169 , n11106 );
not ( n11339 , n11169 );
not ( n11340 , n11106 );
and ( n11341 , n11339 , n11340 );
nor ( n11342 , n11338 , n11341 );
xor ( n11343 , n11022 , n11047 );
xor ( n11344 , n11342 , n11343 );
and ( n11345 , n11337 , n11344 );
and ( n11346 , n11343 , n11342 );
nor ( n11347 , n11345 , n11346 );
xnor ( n11348 , n11172 , n11173 );
nand ( n11349 , n11347 , n11348 );
xor ( n11350 , n11334 , n11262 );
xor ( n11351 , n11103 , n11072 );
xor ( n11352 , n11324 , n11328 );
not ( n11353 , n11352 );
and ( n11354 , n50 , n532 );
and ( n11355 , n11129 , n10610 );
not ( n11356 , n11129 );
and ( n11357 , n11356 , n39 );
nor ( n11358 , n11355 , n11357 );
not ( n11359 , n11358 );
not ( n11360 , n10940 );
or ( n11361 , n11359 , n11360 );
nand ( n11362 , n925 , n10934 );
nand ( n11363 , n11361 , n11362 );
nand ( n11364 , n11354 , n11363 );
and ( n11365 , n3898 , n43 );
not ( n11366 , n3898 );
and ( n11367 , n11366 , n10896 );
nor ( n11368 , n11365 , n11367 );
or ( n11369 , n11368 , n10572 );
not ( n11370 , n854 );
or ( n11371 , n11370 , n10586 );
nand ( n11372 , n11369 , n11371 );
and ( n11373 , n11363 , n11354 );
not ( n11374 , n11363 );
not ( n11375 , n11354 );
and ( n11376 , n11374 , n11375 );
nor ( n11377 , n11373 , n11376 );
nand ( n11378 , n11372 , n11377 );
and ( n11379 , n11364 , n11378 );
nor ( n11380 , n11353 , n11379 );
not ( n11381 , n11380 );
not ( n11382 , n11294 );
not ( n11383 , n11382 );
not ( n11384 , n11330 );
or ( n11385 , n11383 , n11384 );
not ( n11386 , n11330 );
nand ( n11387 , n11294 , n11386 );
nand ( n11388 , n11385 , n11387 );
not ( n11389 , n11388 );
or ( n11390 , n11381 , n11389 );
xor ( n11391 , n11315 , n11301 );
not ( n11392 , n10662 );
and ( n11393 , n41 , n11392 );
not ( n11394 , n41 );
and ( n11395 , n11394 , n10663 );
nor ( n11396 , n11393 , n11395 );
not ( n11397 , n11396 );
not ( n11398 , n10657 );
not ( n11399 , n11398 );
or ( n11400 , n11397 , n11399 );
nand ( n11401 , n882 , n10647 );
nand ( n11402 , n11400 , n11401 );
not ( n11403 , n11402 );
and ( n11404 , n45 , n10613 );
not ( n11405 , n3774 );
and ( n11406 , n4300 , n11405 );
nor ( n11407 , n11404 , n11406 );
not ( n11408 , n11407 );
not ( n11409 , n10604 );
or ( n11410 , n11408 , n11409 );
nand ( n11411 , n11296 , n10617 );
nand ( n11412 , n11410 , n11411 );
not ( n11413 , n11412 );
or ( n11414 , n11403 , n11413 );
and ( n11415 , n47 , n557 );
not ( n11416 , n47 );
not ( n11417 , n10988 );
and ( n11418 , n11416 , n11417 );
nor ( n11419 , n11415 , n11418 );
and ( n11420 , n11419 , n10680 );
and ( n11421 , n11272 , n10687 );
nor ( n11422 , n11420 , n11421 );
not ( n11423 , n11422 );
not ( n11424 , n11402 );
not ( n11425 , n11413 );
or ( n11426 , n11424 , n11425 );
or ( n11427 , n11402 , n11413 );
nand ( n11428 , n11426 , n11427 );
nand ( n11429 , n11423 , n11428 );
nand ( n11430 , n11414 , n11429 );
xnor ( n11431 , n11286 , n11292 );
xor ( n11432 , n11430 , n11431 );
and ( n11433 , n11391 , n11432 );
and ( n11434 , n11430 , n11431 );
nor ( n11435 , n11433 , n11434 );
not ( n11436 , n11435 );
and ( n11437 , n11388 , n11380 );
not ( n11438 , n11388 );
not ( n11439 , n11380 );
and ( n11440 , n11438 , n11439 );
nor ( n11441 , n11437 , n11440 );
nand ( n11442 , n11436 , n11441 );
nand ( n11443 , n11390 , n11442 );
xor ( n11444 , n11351 , n11443 );
and ( n11445 , n11350 , n11444 );
and ( n11446 , n11351 , n11443 );
nor ( n11447 , n11445 , n11446 );
xnor ( n11448 , n11337 , n11344 );
nor ( n11449 , n11447 , n11448 );
not ( n11450 , n11449 );
not ( n11451 , n11444 );
and ( n11452 , n11350 , n11451 );
not ( n11453 , n11350 );
and ( n11454 , n11453 , n11444 );
nor ( n11455 , n11452 , n11454 );
not ( n11456 , n11435 );
not ( n11457 , n11441 );
or ( n11458 , n11456 , n11457 );
or ( n11459 , n11435 , n11441 );
nand ( n11460 , n11458 , n11459 );
not ( n11461 , n11352 );
not ( n11462 , n11379 );
and ( n11463 , n11461 , n11462 );
and ( n11464 , n11352 , n11379 );
nor ( n11465 , n11463 , n11464 );
and ( n11466 , n10579 , n11119 );
buf ( n11467 , n3377 );
not ( n11468 , n11467 );
and ( n11469 , n37 , n11468 );
nor ( n11470 , n11466 , n11469 );
or ( n11471 , n11116 , n11470 );
or ( n11472 , n11322 , n11320 );
nand ( n11473 , n11471 , n11472 );
not ( n11474 , n11473 );
not ( n11475 , n11283 );
not ( n11476 , n10719 );
or ( n11477 , n11475 , n11476 );
not ( n11478 , n49 );
not ( n11479 , n11478 );
not ( n11480 , n532 );
not ( n11481 , n11480 );
or ( n11482 , n11479 , n11481 );
nand ( n11483 , n11482 , n11309 );
not ( n11484 , n11483 );
nand ( n11485 , n11484 , n10713 );
nand ( n11486 , n11477 , n11485 );
not ( n11487 , n11486 );
or ( n11488 , n11474 , n11487 );
not ( n11489 , n1258 );
not ( n11490 , n10940 );
or ( n11491 , n11489 , n11490 );
nand ( n11492 , n11358 , n10934 );
nand ( n11493 , n11491 , n11492 );
not ( n11494 , n1281 );
or ( n11495 , n11116 , n11494 );
not ( n11496 , n11113 );
or ( n11497 , n11496 , n11470 );
nand ( n11498 , n11495 , n11497 );
and ( n11499 , n51 , n610 );
and ( n11500 , n11498 , n11499 );
not ( n11501 , n11498 );
not ( n11502 , n11499 );
and ( n11503 , n11501 , n11502 );
nor ( n11504 , n11500 , n11503 );
and ( n11505 , n11493 , n11504 );
and ( n11506 , n11499 , n11498 );
nor ( n11507 , n11505 , n11506 );
xnor ( n11508 , n11486 , n11473 );
or ( n11509 , n11507 , n11508 );
nand ( n11510 , n11488 , n11509 );
and ( n11511 , n11465 , n11510 );
not ( n11512 , n11465 );
not ( n11513 , n11510 );
and ( n11514 , n11512 , n11513 );
nor ( n11515 , n11511 , n11514 );
xor ( n11516 , n11372 , n11377 );
not ( n11517 , n11516 );
not ( n11518 , n11422 );
not ( n11519 , n11428 );
and ( n11520 , n11518 , n11519 );
and ( n11521 , n11422 , n11428 );
nor ( n11522 , n11520 , n11521 );
not ( n11523 , n11396 );
not ( n11524 , n10750 );
or ( n11525 , n11523 , n11524 );
not ( n11526 , n1153 );
or ( n11527 , n11526 , n10659 );
nand ( n11528 , n11525 , n11527 );
not ( n11529 , n11528 );
buf ( n11530 , n1877 );
not ( n11531 , n11530 );
and ( n11532 , n10596 , n10597 , n10603 );
not ( n11533 , n11532 );
or ( n11534 , n11531 , n11533 );
nand ( n11535 , n11407 , n10619 );
nand ( n11536 , n11534 , n11535 );
not ( n11537 , n1144 );
not ( n11538 , n10631 );
or ( n11539 , n11537 , n11538 );
not ( n11540 , n11368 );
nand ( n11541 , n11540 , n10585 );
nand ( n11542 , n11539 , n11541 );
xor ( n11543 , n11536 , n11542 );
not ( n11544 , n11543 );
or ( n11545 , n11529 , n11544 );
nand ( n11546 , n11542 , n11536 );
nand ( n11547 , n11545 , n11546 );
not ( n11548 , n11547 );
and ( n11549 , n11522 , n11548 );
not ( n11550 , n11522 );
and ( n11551 , n11550 , n11547 );
nor ( n11552 , n11549 , n11551 );
not ( n11553 , n11552 );
or ( n11554 , n11517 , n11553 );
not ( n11555 , n11522 );
nand ( n11556 , n11547 , n11555 );
nand ( n11557 , n11554 , n11556 );
not ( n11558 , n11557 );
or ( n11559 , n11515 , n11558 );
or ( n11560 , n11513 , n11465 );
nand ( n11561 , n11559 , n11560 );
xor ( n11562 , n11259 , n11246 );
xor ( n11563 , n11561 , n11562 );
and ( n11564 , n11460 , n11563 );
and ( n11565 , n11562 , n11561 );
nor ( n11566 , n11564 , n11565 );
nand ( n11567 , n11455 , n11566 );
xnor ( n11568 , n11563 , n11460 );
xnor ( n11569 , n11507 , n11508 );
and ( n11570 , n51 , n520 );
not ( n11571 , n51 );
and ( n11572 , n11571 , n518 );
or ( n11573 , n556 , n11572 );
nand ( n11574 , n11573 , n532 );
nor ( n11575 , n11570 , n11574 );
and ( n11576 , n10610 , n11118 );
and ( n11577 , n39 , n11468 );
nor ( n11578 , n11576 , n11577 );
or ( n11579 , n11116 , n11578 );
or ( n11580 , n11496 , n11494 );
nand ( n11581 , n11579 , n11580 );
nand ( n11582 , n11575 , n11581 );
not ( n11583 , n1237 );
not ( n11584 , n11092 );
not ( n11585 , n11584 );
and ( n11586 , n11583 , n11585 );
and ( n11587 , n11419 , n10687 );
nor ( n11588 , n11586 , n11587 );
not ( n11589 , n11483 );
not ( n11590 , n10756 );
and ( n11591 , n11589 , n11590 );
xor ( n11592 , n50 , n532 );
and ( n11593 , n11592 , n10713 );
nor ( n11594 , n11591 , n11593 );
not ( n11595 , n11594 );
and ( n11596 , n11588 , n11595 );
not ( n11597 , n11588 );
and ( n11598 , n11597 , n11594 );
nor ( n11599 , n11596 , n11598 );
or ( n11600 , n11582 , n11599 );
or ( n11601 , n11594 , n11588 );
nand ( n11602 , n11600 , n11601 );
and ( n11603 , n11569 , n11602 );
not ( n11604 , n11569 );
not ( n11605 , n11602 );
and ( n11606 , n11604 , n11605 );
nor ( n11607 , n11603 , n11606 );
xor ( n11608 , n11504 , n11493 );
not ( n11609 , n11530 );
not ( n11610 , n10731 );
or ( n11611 , n11609 , n11610 );
and ( n11612 , n4266 , n3774 );
and ( n11613 , n47 , n10612 );
nor ( n11614 , n11612 , n11613 );
not ( n11615 , n11614 );
nand ( n11616 , n11615 , n10604 );
nand ( n11617 , n11611 , n11616 );
and ( n11618 , n3898 , n4300 );
not ( n11619 , n3898 );
and ( n11620 , n11619 , n45 );
nor ( n11621 , n11618 , n11620 );
not ( n11622 , n11621 );
not ( n11623 , n10631 );
or ( n11624 , n11622 , n11623 );
nand ( n11625 , n1144 , n10585 );
nand ( n11626 , n11624 , n11625 );
and ( n11627 , n41 , n1575 );
not ( n11628 , n41 );
and ( n11629 , n11628 , n11128 );
nor ( n11630 , n11627 , n11629 );
or ( n11631 , n11630 , n10976 );
not ( n11632 , n1258 );
or ( n11633 , n11632 , n10979 );
nand ( n11634 , n11631 , n11633 );
xor ( n11635 , n11626 , n11634 );
and ( n11636 , n11617 , n11635 );
and ( n11637 , n11626 , n11634 );
nor ( n11638 , n11636 , n11637 );
not ( n11639 , n11638 );
not ( n11640 , n11592 );
not ( n11641 , n10756 );
not ( n11642 , n11641 );
or ( n11643 , n11640 , n11642 );
or ( n11644 , n51 , n10738 );
nor ( n11645 , n11499 , n10712 );
nand ( n11646 , n11644 , n11645 );
nand ( n11647 , n11643 , n11646 );
not ( n11648 , n11647 );
not ( n11649 , n11526 );
not ( n11650 , n10648 );
and ( n11651 , n11649 , n11650 );
not ( n11652 , n10650 );
buf ( n11653 , n11652 );
and ( n11654 , n11653 , n10896 );
not ( n11655 , n11653 );
and ( n11656 , n11655 , n43 );
nor ( n11657 , n11654 , n11656 );
and ( n11658 , n11657 , n11085 );
nor ( n11659 , n11651 , n11658 );
not ( n11660 , n11659 );
and ( n11661 , n49 , n10769 );
not ( n11662 , n49 );
and ( n11663 , n11662 , n10670 );
nor ( n11664 , n11661 , n11663 );
not ( n11665 , n11664 );
not ( n11666 , n11092 );
or ( n11667 , n11665 , n11666 );
not ( n11668 , n1237 );
nand ( n11669 , n11668 , n10687 );
nand ( n11670 , n11667 , n11669 );
not ( n11671 , n11670 );
or ( n11672 , n11660 , n11671 );
or ( n11673 , n11659 , n11670 );
nand ( n11674 , n11672 , n11673 );
not ( n11675 , n11674 );
or ( n11676 , n11648 , n11675 );
not ( n11677 , n11659 );
nand ( n11678 , n11677 , n11670 );
nand ( n11679 , n11676 , n11678 );
not ( n11680 , n11679 );
or ( n11681 , n11639 , n11680 );
or ( n11682 , n11638 , n11679 );
nand ( n11683 , n11681 , n11682 );
and ( n11684 , n11608 , n11683 );
not ( n11685 , n11638 );
and ( n11686 , n11685 , n11679 );
nor ( n11687 , n11684 , n11686 );
or ( n11688 , n11607 , n11687 );
or ( n11689 , n11605 , n11569 );
nand ( n11690 , n11688 , n11689 );
and ( n11691 , n11515 , n11558 );
not ( n11692 , n11515 );
and ( n11693 , n11692 , n11557 );
nor ( n11694 , n11691 , n11693 );
xor ( n11695 , n11391 , n11432 );
xor ( n11696 , n11694 , n11695 );
and ( n11697 , n11690 , n11696 );
and ( n11698 , n11695 , n11694 );
nor ( n11699 , n11697 , n11698 );
nor ( n11700 , n11568 , n11699 );
and ( n11701 , n11567 , n11700 );
nor ( n11702 , n11455 , n11566 );
nor ( n11703 , n11701 , n11702 );
not ( n11704 , n11703 );
nand ( n11705 , n11447 , n11448 );
nand ( n11706 , n11704 , n11705 );
nand ( n11707 , n11450 , n11706 );
nand ( n11708 , n11349 , n11707 );
or ( n11709 , n11347 , n11348 );
nand ( n11710 , n11349 , n11705 );
not ( n11711 , n11710 );
xnor ( n11712 , n11696 , n11690 );
xor ( n11713 , n11687 , n11607 );
xor ( n11714 , n11581 , n11575 );
not ( n11715 , n2147 );
not ( n11716 , n11304 );
or ( n11717 , n11715 , n11716 );
nand ( n11718 , n11621 , n10585 );
nand ( n11719 , n11717 , n11718 );
not ( n11720 , n11719 );
and ( n11721 , n51 , n10718 );
xnor ( n11722 , n1575 , n42 );
not ( n11723 , n11722 );
not ( n11724 , n10939 );
not ( n11725 , n11724 );
or ( n11726 , n11723 , n11725 );
not ( n11727 , n11630 );
nand ( n11728 , n11727 , n10978 );
nand ( n11729 , n11726 , n11728 );
xor ( n11730 , n11721 , n11729 );
not ( n11731 , n11730 );
or ( n11732 , n11720 , n11731 );
nand ( n11733 , n11721 , n11729 );
nand ( n11734 , n11732 , n11733 );
nand ( n11735 , n11714 , n11734 );
not ( n11736 , n2216 );
not ( n11737 , n10679 );
or ( n11738 , n11736 , n11737 );
nand ( n11739 , n11664 , n10687 );
nand ( n11740 , n11738 , n11739 );
not ( n11741 , n2349 );
or ( n11742 , n11116 , n11741 );
or ( n11743 , n11114 , n11578 );
nand ( n11744 , n11742 , n11743 );
not ( n11745 , n11744 );
not ( n11746 , n2206 );
not ( n11747 , n10604 );
or ( n11748 , n11746 , n11747 );
not ( n11749 , n11614 );
not ( n11750 , n10618 );
nand ( n11751 , n11749 , n11750 );
nand ( n11752 , n11748 , n11751 );
not ( n11753 , n11752 );
not ( n11754 , n11753 );
or ( n11755 , n11745 , n11754 );
not ( n11756 , n11744 );
nand ( n11757 , n11756 , n11752 );
nand ( n11758 , n11755 , n11757 );
and ( n11759 , n11740 , n11758 );
and ( n11760 , n11744 , n11752 );
nor ( n11761 , n11759 , n11760 );
not ( n11762 , n11761 );
xor ( n11763 , n11714 , n11734 );
nand ( n11764 , n11762 , n11763 );
and ( n11765 , n11735 , n11764 );
xnor ( n11766 , n11582 , n11599 );
not ( n11767 , n11528 );
and ( n11768 , n11543 , n11767 );
not ( n11769 , n11543 );
and ( n11770 , n11769 , n11528 );
nor ( n11771 , n11768 , n11770 );
not ( n11772 , n11771 );
and ( n11773 , n11766 , n11772 );
not ( n11774 , n11766 );
and ( n11775 , n11774 , n11771 );
nor ( n11776 , n11773 , n11775 );
or ( n11777 , n11765 , n11776 );
or ( n11778 , n11766 , n11771 );
nand ( n11779 , n11777 , n11778 );
xor ( n11780 , n11552 , n11516 );
xor ( n11781 , n11779 , n11780 );
and ( n11782 , n11713 , n11781 );
and ( n11783 , n11780 , n11779 );
nor ( n11784 , n11782 , n11783 );
nor ( n11785 , n11712 , n11784 );
not ( n11786 , n11785 );
xnor ( n11787 , n11713 , n11781 );
and ( n11788 , n51 , n10676 );
nand ( n11789 , n10988 , n10677 );
nor ( n11790 , n11788 , n11789 );
and ( n11791 , n11129 , n10896 );
not ( n11792 , n11129 );
and ( n11793 , n11792 , n43 );
nor ( n11794 , n11791 , n11793 );
and ( n11795 , n11794 , n10940 );
and ( n11796 , n11722 , n10934 );
nor ( n11797 , n11795 , n11796 );
not ( n11798 , n11797 );
and ( n11799 , n11790 , n11798 );
not ( n11800 , n2179 );
not ( n11801 , n11085 );
or ( n11802 , n11800 , n11801 );
nand ( n11803 , n11657 , n11003 );
nand ( n11804 , n11802 , n11803 );
xor ( n11805 , n11799 , n11804 );
and ( n11806 , n41 , n11118 );
not ( n11807 , n41 );
and ( n11808 , n11807 , n11468 );
nor ( n11809 , n11806 , n11808 );
and ( n11810 , n11115 , n11809 );
not ( n11811 , n11114 );
not ( n11812 , n11741 );
and ( n11813 , n11811 , n11812 );
nor ( n11814 , n11810 , n11813 );
not ( n11815 , n11814 );
not ( n11816 , n11815 );
and ( n11817 , n4266 , n3898 );
not ( n11818 , n4266 );
not ( n11819 , n3898 );
and ( n11820 , n11818 , n11819 );
nor ( n11821 , n11817 , n11820 );
and ( n11822 , n11821 , n10631 );
and ( n11823 , n2147 , n10584 );
nor ( n11824 , n11822 , n11823 );
not ( n11825 , n11824 );
not ( n11826 , n11825 );
not ( n11827 , n1820 );
xor ( n11828 , n11827 , n49 );
not ( n11829 , n11828 );
not ( n11830 , n11532 );
or ( n11831 , n11829 , n11830 );
nand ( n11832 , n2206 , n10619 );
nand ( n11833 , n11831 , n11832 );
not ( n11834 , n11833 );
not ( n11835 , n11834 );
or ( n11836 , n11826 , n11835 );
nand ( n11837 , n11824 , n11833 );
nand ( n11838 , n11836 , n11837 );
not ( n11839 , n11838 );
or ( n11840 , n11816 , n11839 );
or ( n11841 , n11824 , n11834 );
nand ( n11842 , n11840 , n11841 );
and ( n11843 , n11805 , n11842 );
and ( n11844 , n11804 , n11799 );
nor ( n11845 , n11843 , n11844 );
not ( n11846 , n11647 );
and ( n11847 , n11674 , n11846 );
not ( n11848 , n11674 );
and ( n11849 , n11848 , n11647 );
nor ( n11850 , n11847 , n11849 );
xor ( n11851 , n11635 , n11617 );
and ( n11852 , n11850 , n11851 );
not ( n11853 , n11850 );
not ( n11854 , n11851 );
and ( n11855 , n11853 , n11854 );
nor ( n11856 , n11852 , n11855 );
or ( n11857 , n11845 , n11856 );
or ( n11858 , n11854 , n11850 );
nand ( n11859 , n11857 , n11858 );
xor ( n11860 , n11776 , n11765 );
xor ( n11861 , n11608 , n11683 );
xor ( n11862 , n11860 , n11861 );
and ( n11863 , n11859 , n11862 );
and ( n11864 , n11861 , n11860 );
nor ( n11865 , n11863 , n11864 );
nand ( n11866 , n11787 , n11865 );
xor ( n11867 , n11845 , n11856 );
not ( n11868 , n11790 );
not ( n11869 , n11797 );
and ( n11870 , n11868 , n11869 );
and ( n11871 , n11790 , n11797 );
nor ( n11872 , n11870 , n11871 );
not ( n11873 , n2179 );
not ( n11874 , n11873 );
not ( n11875 , n10648 );
and ( n11876 , n11874 , n11875 );
and ( n11877 , n4300 , n11653 );
not ( n11878 , n4300 );
and ( n11879 , n11878 , n11392 );
nor ( n11880 , n11877 , n11879 );
and ( n11881 , n11880 , n11085 );
nor ( n11882 , n11876 , n11881 );
not ( n11883 , n2216 );
not ( n11884 , n10687 );
or ( n11885 , n11883 , n11884 );
not ( n11886 , n10988 );
not ( n11887 , n11886 );
or ( n11888 , n51 , n11887 );
nand ( n11889 , n51 , n11887 );
nand ( n11890 , n11888 , n11889 , n11092 );
nand ( n11891 , n11885 , n11890 );
and ( n11892 , n11882 , n11891 );
not ( n11893 , n11882 );
not ( n11894 , n11891 );
and ( n11895 , n11893 , n11894 );
nor ( n11896 , n11892 , n11895 );
or ( n11897 , n11872 , n11896 );
or ( n11898 , n11882 , n11894 );
nand ( n11899 , n11897 , n11898 );
not ( n11900 , n11899 );
xnor ( n11901 , n11730 , n11719 );
xor ( n11902 , n11740 , n11758 );
not ( n11903 , n11902 );
and ( n11904 , n11901 , n11903 );
not ( n11905 , n11901 );
and ( n11906 , n11905 , n11902 );
nor ( n11907 , n11904 , n11906 );
not ( n11908 , n11907 );
or ( n11909 , n11900 , n11908 );
not ( n11910 , n11901 );
nand ( n11911 , n11910 , n11902 );
nand ( n11912 , n11909 , n11911 );
and ( n11913 , n11763 , n11762 );
not ( n11914 , n11763 );
and ( n11915 , n11914 , n11761 );
nor ( n11916 , n11913 , n11915 );
and ( n11917 , n11912 , n11916 );
not ( n11918 , n11912 );
not ( n11919 , n11916 );
and ( n11920 , n11918 , n11919 );
nor ( n11921 , n11917 , n11920 );
and ( n11922 , n11867 , n11921 );
and ( n11923 , n11916 , n11912 );
nor ( n11924 , n11922 , n11923 );
not ( n11925 , n11924 );
xnor ( n11926 , n11862 , n11859 );
not ( n11927 , n11926 );
nand ( n11928 , n11925 , n11927 );
and ( n11929 , n4266 , n10662 );
not ( n11930 , n4266 );
not ( n11931 , n11652 );
and ( n11932 , n11930 , n11931 );
nor ( n11933 , n11929 , n11932 );
and ( n11934 , n11933 , n11267 );
and ( n11935 , n763 , n11653 );
not ( n11936 , n763 );
and ( n11937 , n11936 , n11392 );
nor ( n11938 , n11935 , n11937 );
and ( n11939 , n11938 , n11003 );
nor ( n11940 , n11934 , n11939 );
nand ( n11941 , n51 , n10635 );
not ( n11942 , n51 );
nand ( n11943 , n11942 , n3898 );
nand ( n11944 , n3753 , n11943 );
and ( n11945 , n11941 , n11006 , n11944 );
not ( n11946 , n11945 );
and ( n11947 , n45 , n1575 );
not ( n11948 , n45 );
and ( n11949 , n11948 , n1576 );
or ( n11950 , n11947 , n11949 );
not ( n11951 , n11950 );
not ( n11952 , n11724 );
or ( n11953 , n11951 , n11952 );
nand ( n11954 , n2490 , n10978 );
nand ( n11955 , n11953 , n11954 );
not ( n11956 , n11955 );
not ( n11957 , n11956 );
and ( n11958 , n11946 , n11957 );
and ( n11959 , n11945 , n11956 );
nor ( n11960 , n11958 , n11959 );
not ( n11961 , n11960 );
and ( n11962 , n11940 , n11961 );
not ( n11963 , n11940 );
and ( n11964 , n11963 , n11960 );
nor ( n11965 , n11962 , n11964 );
xnor ( n11966 , n10562 , n49 );
not ( n11967 , n11966 );
not ( n11968 , n10836 );
and ( n11969 , n11967 , n11968 );
and ( n11970 , n2763 , n11304 );
nor ( n11971 , n11969 , n11970 );
not ( n11972 , n11971 );
not ( n11973 , n11115 );
not ( n11974 , n2783 );
or ( n11975 , n11973 , n11974 );
not ( n11976 , n11467 );
and ( n11977 , n10896 , n11976 );
not ( n11978 , n10896 );
and ( n11979 , n11978 , n11118 );
nor ( n11980 , n11977 , n11979 );
nand ( n11981 , n11113 , n11980 );
nand ( n11982 , n11975 , n11981 );
and ( n11983 , n51 , n10617 );
not ( n11984 , n11983 );
and ( n11985 , n11982 , n11984 );
not ( n11986 , n11982 );
and ( n11987 , n11986 , n11983 );
nor ( n11988 , n11985 , n11987 );
not ( n11989 , n11988 );
and ( n11990 , n11972 , n11989 );
and ( n11991 , n11983 , n11982 );
nor ( n11992 , n11990 , n11991 );
xor ( n11993 , n11965 , n11992 );
not ( n11994 , n11966 );
not ( n11995 , n11994 );
not ( n11996 , n11304 );
or ( n11997 , n11995 , n11996 );
not ( n11998 , n48 );
and ( n11999 , n3898 , n11998 );
not ( n12000 , n3898 );
and ( n12001 , n12000 , n48 );
nor ( n12002 , n11999 , n12001 );
nand ( n12003 , n12002 , n10584 );
nand ( n12004 , n11997 , n12003 );
not ( n12005 , n12004 );
not ( n12006 , n12005 );
not ( n12007 , n2940 );
not ( n12008 , n10619 );
or ( n12009 , n12007 , n12008 );
not ( n12010 , n51 );
nand ( n12011 , n12010 , n10916 );
nand ( n12012 , n51 , n10607 );
nand ( n12013 , n12011 , n12012 , n11532 );
nand ( n12014 , n12009 , n12013 );
not ( n12015 , n12014 );
or ( n12016 , n12006 , n12015 );
or ( n12017 , n12005 , n12014 );
nand ( n12018 , n12016 , n12017 );
not ( n12019 , n11980 );
or ( n12020 , n11116 , n12019 );
not ( n12021 , n42 );
and ( n12022 , n11118 , n12021 );
not ( n12023 , n11118 );
and ( n12024 , n12023 , n42 );
nor ( n12025 , n12022 , n12024 );
or ( n12026 , n11114 , n12025 );
nand ( n12027 , n12020 , n12026 );
and ( n12028 , n12018 , n12027 );
not ( n12029 , n12018 );
not ( n12030 , n12027 );
and ( n12031 , n12029 , n12030 );
nor ( n12032 , n12028 , n12031 );
not ( n12033 , n10662 );
not ( n12034 , n51 );
not ( n12035 , n3853 );
nand ( n12036 , n12034 , n12035 );
and ( n12037 , n12033 , n12036 );
not ( n12038 , n12035 );
and ( n12039 , n51 , n12038 );
not ( n12040 , n10890 );
nor ( n12041 , n12037 , n12039 , n12040 );
and ( n12042 , n4300 , n11976 );
not ( n12043 , n4300 );
and ( n12044 , n12043 , n11118 );
nor ( n12045 , n12042 , n12044 );
not ( n12046 , n12045 );
or ( n12047 , n11116 , n12046 );
not ( n12048 , n2783 );
or ( n12049 , n11322 , n12048 );
nand ( n12050 , n12047 , n12049 );
and ( n12051 , n12041 , n12050 );
not ( n12052 , n12051 );
xor ( n12053 , n11931 , n48 );
and ( n12054 , n12053 , n11267 );
not ( n12055 , n11933 );
nor ( n12056 , n12055 , n11002 );
nor ( n12057 , n12054 , n12056 );
not ( n12058 , n3017 );
not ( n12059 , n12058 );
not ( n12060 , n10976 );
and ( n12061 , n12059 , n12060 );
and ( n12062 , n11950 , n10934 );
nor ( n12063 , n12061 , n12062 );
and ( n12064 , n12057 , n12063 );
not ( n12065 , n12057 );
not ( n12066 , n12063 );
and ( n12067 , n12065 , n12066 );
nor ( n12068 , n12064 , n12067 );
not ( n12069 , n12068 );
or ( n12070 , n12052 , n12069 );
or ( n12071 , n12057 , n12063 );
nand ( n12072 , n12070 , n12071 );
and ( n12073 , n12032 , n12072 );
not ( n12074 , n12032 );
not ( n12075 , n12072 );
and ( n12076 , n12074 , n12075 );
nor ( n12077 , n12073 , n12076 );
and ( n12078 , n11993 , n12077 );
and ( n12079 , n12072 , n12032 );
nor ( n12080 , n12078 , n12079 );
and ( n12081 , n11938 , n11398 );
and ( n12082 , n11880 , n10647 );
nor ( n12083 , n12081 , n12082 );
not ( n12084 , n12083 );
not ( n12085 , n2940 );
not ( n12086 , n11532 );
or ( n12087 , n12085 , n12086 );
nand ( n12088 , n11828 , n10617 );
nand ( n12089 , n12087 , n12088 );
not ( n12090 , n12089 );
not ( n12091 , n12025 );
and ( n12092 , n11115 , n12091 );
not ( n12093 , n11322 );
and ( n12094 , n12093 , n11809 );
nor ( n12095 , n12092 , n12094 );
and ( n12096 , n12090 , n12095 );
not ( n12097 , n12090 );
not ( n12098 , n12095 );
and ( n12099 , n12097 , n12098 );
nor ( n12100 , n12096 , n12099 );
not ( n12101 , n12100 );
or ( n12102 , n12084 , n12101 );
or ( n12103 , n12083 , n12100 );
nand ( n12104 , n12102 , n12103 );
or ( n12105 , n11992 , n11965 );
or ( n12106 , n11940 , n11960 );
nand ( n12107 , n12105 , n12106 );
xor ( n12108 , n12104 , n12107 );
not ( n12109 , n2490 );
not ( n12110 , n11724 );
or ( n12111 , n12109 , n12110 );
nand ( n12112 , n11794 , n10934 );
nand ( n12113 , n12111 , n12112 );
and ( n12114 , n51 , n10686 );
and ( n12115 , n12113 , n12114 );
not ( n12116 , n12113 );
not ( n12117 , n12114 );
and ( n12118 , n12116 , n12117 );
nor ( n12119 , n12115 , n12118 );
not ( n12120 , n12119 );
and ( n12121 , n12002 , n10631 );
and ( n12122 , n11821 , n10835 );
nor ( n12123 , n12121 , n12122 );
xor ( n12124 , n12120 , n12123 );
not ( n12125 , n11945 );
nor ( n12126 , n12125 , n11956 );
not ( n12127 , n12126 );
not ( n12128 , n12027 );
not ( n12129 , n12018 );
or ( n12130 , n12128 , n12129 );
not ( n12131 , n12005 );
nand ( n12132 , n12131 , n12014 );
nand ( n12133 , n12130 , n12132 );
not ( n12134 , n12133 );
not ( n12135 , n12134 );
or ( n12136 , n12127 , n12135 );
not ( n12137 , n12126 );
nand ( n12138 , n12137 , n12133 );
nand ( n12139 , n12136 , n12138 );
not ( n12140 , n12139 );
and ( n12141 , n12124 , n12140 );
not ( n12142 , n12124 );
and ( n12143 , n12142 , n12139 );
nor ( n12144 , n12141 , n12143 );
and ( n12145 , n12108 , n12144 );
not ( n12146 , n12108 );
not ( n12147 , n12144 );
and ( n12148 , n12146 , n12147 );
nor ( n12149 , n12145 , n12148 );
nor ( n12150 , n12080 , n12149 );
xor ( n12151 , n12068 , n12051 );
not ( n12152 , n49 );
and ( n12153 , n12152 , n10662 );
not ( n12154 , n12152 );
and ( n12155 , n12154 , n12033 );
nor ( n12156 , n12153 , n12155 );
not ( n12157 , n12156 );
not ( n12158 , n12157 );
not ( n12159 , n10657 );
and ( n12160 , n12158 , n12159 );
and ( n12161 , n12053 , n10647 );
nor ( n12162 , n12160 , n12161 );
not ( n12163 , n12162 );
not ( n12164 , n12163 );
not ( n12165 , n2763 );
not ( n12166 , n10835 );
or ( n12167 , n12165 , n12166 );
nand ( n12168 , n51 , n10577 );
not ( n12169 , n51 );
nand ( n12170 , n12169 , n12040 );
not ( n12171 , n10571 );
nand ( n12172 , n12168 , n12170 , n12171 );
nand ( n12173 , n12167 , n12172 );
not ( n12174 , n12173 );
and ( n12175 , n4266 , n1576 );
not ( n12176 , n4266 );
and ( n12177 , n12176 , n11129 );
or ( n12178 , n12175 , n12177 );
and ( n12179 , n12178 , n11724 );
not ( n12180 , n10933 );
nor ( n12181 , n12058 , n12180 );
nor ( n12182 , n12179 , n12181 );
not ( n12183 , n12182 );
or ( n12184 , n12174 , n12183 );
or ( n12185 , n12173 , n12182 );
nand ( n12186 , n12184 , n12185 );
not ( n12187 , n12186 );
or ( n12188 , n12164 , n12187 );
not ( n12189 , n12182 );
nand ( n12190 , n12189 , n12173 );
nand ( n12191 , n12188 , n12190 );
and ( n12192 , n11988 , n11971 );
not ( n12193 , n11988 );
not ( n12194 , n11971 );
and ( n12195 , n12193 , n12194 );
nor ( n12196 , n12192 , n12195 );
and ( n12197 , n12191 , n12196 );
not ( n12198 , n12191 );
not ( n12199 , n12196 );
and ( n12200 , n12198 , n12199 );
nor ( n12201 , n12197 , n12200 );
not ( n12202 , n12201 );
not ( n12203 , n12202 );
and ( n12204 , n12151 , n12203 );
and ( n12205 , n12196 , n12191 );
nor ( n12206 , n12204 , n12205 );
xnor ( n12207 , n12077 , n11993 );
nor ( n12208 , n12206 , n12207 );
nor ( n12209 , n12150 , n12208 );
nand ( n12210 , n12206 , n12207 );
not ( n12211 , n3090 );
not ( n12212 , n10975 );
or ( n12213 , n12211 , n12212 );
nand ( n12214 , n12178 , n10978 );
nand ( n12215 , n12213 , n12214 );
not ( n12216 , n12215 );
not ( n12217 , n11115 );
not ( n12218 , n3104 );
or ( n12219 , n12217 , n12218 );
nand ( n12220 , n11113 , n12045 );
nand ( n12221 , n12219 , n12220 );
and ( n12222 , n51 , n10584 );
and ( n12223 , n12221 , n12222 );
not ( n12224 , n12221 );
not ( n12225 , n12222 );
and ( n12226 , n12224 , n12225 );
nor ( n12227 , n12223 , n12226 );
not ( n12228 , n12227 );
or ( n12229 , n12216 , n12228 );
nand ( n12230 , n12222 , n12221 );
nand ( n12231 , n12229 , n12230 );
xor ( n12232 , n12041 , n12050 );
and ( n12233 , n12231 , n12232 );
not ( n12234 , n12231 );
not ( n12235 , n12232 );
and ( n12236 , n12234 , n12235 );
nor ( n12237 , n12233 , n12236 );
and ( n12238 , n12186 , n12163 );
not ( n12239 , n12186 );
and ( n12240 , n12239 , n12162 );
nor ( n12241 , n12238 , n12240 );
and ( n12242 , n12237 , n12241 );
and ( n12243 , n12232 , n12231 );
nor ( n12244 , n12242 , n12243 );
not ( n12245 , n12244 );
not ( n12246 , n12151 );
not ( n12247 , n12202 );
or ( n12248 , n12246 , n12247 );
not ( n12249 , n12151 );
nand ( n12250 , n12249 , n12201 );
nand ( n12251 , n12248 , n12250 );
not ( n12252 , n12251 );
or ( n12253 , n12245 , n12252 );
or ( n12254 , n12244 , n12251 );
nand ( n12255 , n12253 , n12254 );
not ( n12256 , n12255 );
nand ( n12257 , n51 , n1576 );
or ( n12258 , n51 , n11128 );
nand ( n12259 , n12258 , n1688 );
and ( n12260 , n12257 , n11392 , n12259 );
and ( n12261 , n11976 , n47 );
not ( n12262 , n11976 );
and ( n12263 , n12262 , n4266 );
nor ( n12264 , n12261 , n12263 );
or ( n12265 , n11116 , n12264 );
not ( n12266 , n3104 );
or ( n12267 , n11496 , n12266 );
nand ( n12268 , n12265 , n12267 );
nand ( n12269 , n12260 , n12268 );
and ( n12270 , n50 , n12033 );
not ( n12271 , n50 );
and ( n12272 , n12271 , n11653 );
nor ( n12273 , n12270 , n12272 );
and ( n12274 , n12273 , n11398 );
and ( n12275 , n12156 , n10647 );
nor ( n12276 , n12274 , n12275 );
xnor ( n12277 , n12269 , n12276 );
not ( n12278 , n12215 );
and ( n12279 , n12227 , n12278 );
not ( n12280 , n12227 );
and ( n12281 , n12280 , n12215 );
nor ( n12282 , n12279 , n12281 );
or ( n12283 , n12277 , n12282 );
or ( n12284 , n12269 , n12276 );
nand ( n12285 , n12283 , n12284 );
not ( n12286 , n12285 );
not ( n12287 , n12241 );
and ( n12288 , n12237 , n12287 );
not ( n12289 , n12237 );
and ( n12290 , n12289 , n12241 );
nor ( n12291 , n12288 , n12290 );
nand ( n12292 , n12286 , n12291 );
not ( n12293 , n12292 );
and ( n12294 , n12268 , n12260 );
not ( n12295 , n12268 );
not ( n12296 , n12260 );
and ( n12297 , n12295 , n12296 );
nor ( n12298 , n12294 , n12297 );
not ( n12299 , n12273 );
not ( n12300 , n10647 );
or ( n12301 , n12299 , n12300 );
nand ( n12302 , n51 , n11392 );
not ( n12303 , n51 );
nand ( n12304 , n12303 , n11653 );
not ( n12305 , n10657 );
nand ( n12306 , n12302 , n12304 , n12305 );
nand ( n12307 , n12301 , n12306 );
not ( n12308 , n12307 );
not ( n12309 , n49 );
not ( n12310 , n1575 );
or ( n12311 , n12309 , n12310 );
or ( n12312 , n49 , n1575 );
nand ( n12313 , n12311 , n12312 );
not ( n12314 , n12313 );
not ( n12315 , n12314 );
not ( n12316 , n10975 );
not ( n12317 , n12316 );
and ( n12318 , n12315 , n12317 );
and ( n12319 , n3090 , n10934 );
nor ( n12320 , n12318 , n12319 );
not ( n12321 , n12320 );
or ( n12322 , n12308 , n12321 );
or ( n12323 , n12307 , n12320 );
nand ( n12324 , n12322 , n12323 );
and ( n12325 , n12298 , n12324 );
not ( n12326 , n12320 );
and ( n12327 , n12307 , n12326 );
nor ( n12328 , n12325 , n12327 );
xnor ( n12329 , n12277 , n12282 );
nand ( n12330 , n12328 , n12329 );
not ( n12331 , n12330 );
nand ( n12332 , n51 , n10933 );
not ( n12333 , n12332 );
not ( n12334 , n11113 );
and ( n12335 , n49 , n11118 );
not ( n12336 , n49 );
not ( n12337 , n11467 );
and ( n12338 , n12336 , n12337 );
nor ( n12339 , n12335 , n12338 );
not ( n12340 , n12339 );
or ( n12341 , n12334 , n12340 );
not ( n12342 , n3380 );
nand ( n12343 , n11115 , n12342 );
nand ( n12344 , n12341 , n12343 );
nand ( n12345 , n12333 , n12344 );
nand ( n12346 , n51 , n11112 );
and ( n12347 , n11119 , n12346 );
not ( n12348 , n51 );
not ( n12349 , n12348 );
not ( n12350 , n11115 );
or ( n12351 , n12349 , n12350 );
nand ( n12352 , n11113 , n12342 );
nand ( n12353 , n12351 , n12352 );
and ( n12354 , n12347 , n12353 );
not ( n12355 , n12344 );
nand ( n12356 , n12355 , n12332 );
nand ( n12357 , n12354 , n12356 );
nand ( n12358 , n12345 , n12357 );
and ( n12359 , n50 , n11128 );
not ( n12360 , n50 );
and ( n12361 , n12360 , n1575 );
nor ( n12362 , n12359 , n12361 );
not ( n12363 , n12362 );
not ( n12364 , n10934 );
or ( n12365 , n12363 , n12364 );
or ( n12366 , n51 , n10943 );
not ( n12367 , n51 );
or ( n12368 , n12367 , n11129 );
nand ( n12369 , n12366 , n12368 , n10975 );
nand ( n12370 , n12365 , n12369 );
nand ( n12371 , n51 , n11118 );
or ( n12372 , n51 , n11467 );
nand ( n12373 , n12372 , n10930 );
and ( n12374 , n12371 , n10943 , n12373 );
not ( n12375 , n11115 );
not ( n12376 , n12339 );
or ( n12377 , n12375 , n12376 );
not ( n12378 , n3173 );
or ( n12379 , n11496 , n12378 );
nand ( n12380 , n12377 , n12379 );
xor ( n12381 , n12374 , n12380 );
xor ( n12382 , n12370 , n12381 );
and ( n12383 , n12358 , n12382 );
and ( n12384 , n12370 , n12381 );
nor ( n12385 , n12383 , n12384 );
not ( n12386 , n12385 );
not ( n12387 , n12386 );
and ( n12388 , n12374 , n12380 );
not ( n12389 , n12388 );
not ( n12390 , n11116 );
not ( n12391 , n12378 );
and ( n12392 , n12390 , n12391 );
not ( n12393 , n12264 );
and ( n12394 , n12093 , n12393 );
nor ( n12395 , n12392 , n12394 );
not ( n12396 , n12395 );
and ( n12397 , n51 , n10646 );
not ( n12398 , n12397 );
not ( n12399 , n12362 );
not ( n12400 , n10939 );
not ( n12401 , n12400 );
or ( n12402 , n12399 , n12401 );
nand ( n12403 , n12313 , n10933 );
nand ( n12404 , n12402 , n12403 );
not ( n12405 , n12404 );
not ( n12406 , n12405 );
or ( n12407 , n12398 , n12406 );
not ( n12408 , n12397 );
nand ( n12409 , n12408 , n12404 );
nand ( n12410 , n12407 , n12409 );
not ( n12411 , n12410 );
or ( n12412 , n12396 , n12411 );
or ( n12413 , n12395 , n12410 );
nand ( n12414 , n12412 , n12413 );
not ( n12415 , n12414 );
not ( n12416 , n12415 );
or ( n12417 , n12389 , n12416 );
not ( n12418 , n12388 );
nand ( n12419 , n12418 , n12414 );
nand ( n12420 , n12417 , n12419 );
not ( n12421 , n12420 );
or ( n12422 , n12387 , n12421 );
nand ( n12423 , n12388 , n12414 );
nand ( n12424 , n12422 , n12423 );
not ( n12425 , n12424 );
not ( n12426 , n12395 );
and ( n12427 , n12426 , n12410 );
and ( n12428 , n12397 , n12404 );
nor ( n12429 , n12427 , n12428 );
not ( n12430 , n12429 );
not ( n12431 , n12324 );
and ( n12432 , n12298 , n12431 );
not ( n12433 , n12298 );
and ( n12434 , n12433 , n12324 );
nor ( n12435 , n12432 , n12434 );
not ( n12436 , n12435 );
not ( n12437 , n12436 );
or ( n12438 , n12430 , n12437 );
not ( n12439 , n12429 );
nand ( n12440 , n12439 , n12435 );
nand ( n12441 , n12438 , n12440 );
not ( n12442 , n12441 );
or ( n12443 , n12425 , n12442 );
not ( n12444 , n12429 );
nand ( n12445 , n12444 , n12436 );
nand ( n12446 , n12443 , n12445 );
not ( n12447 , n12446 );
or ( n12448 , n12331 , n12447 );
not ( n12449 , n12328 );
not ( n12450 , n12329 );
nand ( n12451 , n12449 , n12450 );
nand ( n12452 , n12448 , n12451 );
not ( n12453 , n12452 );
or ( n12454 , n12293 , n12453 );
not ( n12455 , n12291 );
nand ( n12456 , n12285 , n12455 );
nand ( n12457 , n12454 , n12456 );
not ( n12458 , n12457 );
or ( n12459 , n12256 , n12458 );
not ( n12460 , n12244 );
nand ( n12461 , n12460 , n12251 );
nand ( n12462 , n12459 , n12461 );
nand ( n12463 , n12210 , n12462 );
and ( n12464 , n12209 , n12463 );
and ( n12465 , n12080 , n12149 );
nor ( n12466 , n12464 , n12465 );
not ( n12467 , n12466 );
and ( n12468 , n12108 , n12147 );
and ( n12469 , n12104 , n12107 );
nor ( n12470 , n12468 , n12469 );
and ( n12471 , n11838 , n11814 );
not ( n12472 , n11838 );
and ( n12473 , n12472 , n11815 );
nor ( n12474 , n12471 , n12473 );
nand ( n12475 , n12098 , n12089 );
not ( n12476 , n12083 );
nand ( n12477 , n12476 , n12100 );
nand ( n12478 , n12475 , n12477 );
not ( n12479 , n12114 );
not ( n12480 , n12113 );
or ( n12481 , n12479 , n12480 );
not ( n12482 , n12123 );
nand ( n12483 , n12482 , n12119 );
nand ( n12484 , n12481 , n12483 );
not ( n12485 , n12484 );
and ( n12486 , n12478 , n12485 );
not ( n12487 , n12478 );
and ( n12488 , n12487 , n12484 );
nor ( n12489 , n12486 , n12488 );
not ( n12490 , n12489 );
and ( n12491 , n12474 , n12490 );
not ( n12492 , n12474 );
and ( n12493 , n12492 , n12489 );
nor ( n12494 , n12491 , n12493 );
xnor ( n12495 , n11872 , n11896 );
not ( n12496 , n12495 );
and ( n12497 , n12494 , n12496 );
not ( n12498 , n12494 );
and ( n12499 , n12498 , n12495 );
nor ( n12500 , n12497 , n12499 );
and ( n12501 , n12124 , n12139 );
and ( n12502 , n12126 , n12133 );
nor ( n12503 , n12501 , n12502 );
xnor ( n12504 , n12500 , n12503 );
nand ( n12505 , n12470 , n12504 );
not ( n12506 , n12505 );
or ( n12507 , n12467 , n12506 );
or ( n12508 , n12470 , n12504 );
nand ( n12509 , n12507 , n12508 );
or ( n12510 , n12503 , n12500 );
or ( n12511 , n12495 , n12494 );
nand ( n12512 , n12510 , n12511 );
not ( n12513 , n12512 );
xnor ( n12514 , n11907 , n11899 );
not ( n12515 , n12474 );
not ( n12516 , n12489 );
and ( n12517 , n12515 , n12516 );
and ( n12518 , n12484 , n12478 );
nor ( n12519 , n12517 , n12518 );
xor ( n12520 , n11842 , n11805 );
and ( n12521 , n12519 , n12520 );
not ( n12522 , n12519 );
not ( n12523 , n12520 );
and ( n12524 , n12522 , n12523 );
nor ( n12525 , n12521 , n12524 );
xnor ( n12526 , n12514 , n12525 );
nand ( n12527 , n12513 , n12526 );
and ( n12528 , n12509 , n12527 );
not ( n12529 , n12526 );
and ( n12530 , n12512 , n12529 );
nor ( n12531 , n12528 , n12530 );
xor ( n12532 , n11921 , n11867 );
or ( n12533 , n12514 , n12525 );
or ( n12534 , n12523 , n12519 );
nand ( n12535 , n12533 , n12534 );
nor ( n12536 , n12532 , n12535 );
nor ( n12537 , n12531 , n12536 );
and ( n12538 , n12535 , n12532 );
or ( n12539 , n12537 , n12538 );
nand ( n12540 , n11924 , n11926 );
nand ( n12541 , n12539 , n12540 );
nand ( n12542 , n11928 , n12541 );
nand ( n12543 , n11866 , n12542 );
not ( n12544 , n12543 );
not ( n12545 , n11787 );
not ( n12546 , n11865 );
nand ( n12547 , n12545 , n12546 );
not ( n12548 , n12547 );
or ( n12549 , n12544 , n12548 );
nand ( n12550 , n11712 , n11784 );
nand ( n12551 , n12549 , n12550 );
nand ( n12552 , n11786 , n12551 );
nand ( n12553 , n11568 , n11699 );
nand ( n12554 , n12553 , n11567 );
not ( n12555 , n12554 );
nand ( n12556 , n11711 , n12552 , n12555 );
nand ( n12557 , n11708 , n11709 , n12556 );
nand ( n12558 , n11062 , n11175 );
nand ( n12559 , n11245 , n12557 , n12558 );
nand ( n12560 , n11242 , n12559 );
not ( n12561 , n11206 );
not ( n12562 , n10921 );
or ( n12563 , n12561 , n12562 );
buf ( n12564 , n10818 );
nand ( n12565 , n12564 , n10731 );
nand ( n12566 , n12563 , n12565 );
not ( n12567 , n12566 );
not ( n12568 , n11217 );
not ( n12569 , n11214 );
or ( n12570 , n12568 , n12569 );
nand ( n12571 , n11213 , n11208 );
nand ( n12572 , n12570 , n12571 );
not ( n12573 , n12572 );
or ( n12574 , n12567 , n12573 );
or ( n12575 , n12566 , n12572 );
nand ( n12576 , n12574 , n12575 );
not ( n12577 , n11187 );
not ( n12578 , n10680 );
or ( n12579 , n12577 , n12578 );
and ( n12580 , n11886 , n37 );
not ( n12581 , n11886 );
and ( n12582 , n12581 , n10579 );
nor ( n12583 , n12580 , n12582 );
not ( n12584 , n12583 );
nand ( n12585 , n12584 , n10811 );
nand ( n12586 , n12579 , n12585 );
xor ( n12587 , n10844 , n12586 );
not ( n12588 , n10879 );
not ( n12589 , n12588 );
or ( n12590 , n3717 , n12589 );
or ( n12591 , n39 , n610 );
nand ( n12592 , n39 , n610 );
nand ( n12593 , n12591 , n12592 );
not ( n12594 , n11641 );
or ( n12595 , n12593 , n12594 );
nand ( n12596 , n12590 , n12595 );
xor ( n12597 , n12587 , n12596 );
and ( n12598 , n12576 , n12597 );
not ( n12599 , n12576 );
not ( n12600 , n12597 );
and ( n12601 , n12599 , n12600 );
nor ( n12602 , n12598 , n12601 );
not ( n12603 , n10828 );
not ( n12604 , n11192 );
or ( n12605 , n12603 , n12604 );
or ( n12606 , n11191 , n11189 );
nand ( n12607 , n12605 , n12606 );
xor ( n12608 , n12602 , n12607 );
or ( n12609 , n11196 , n11225 );
not ( n12610 , n11201 );
or ( n12611 , n12610 , n11218 );
nand ( n12612 , n12609 , n12611 );
xor ( n12613 , n12608 , n12612 );
not ( n12614 , n12613 );
not ( n12615 , n11230 );
not ( n12616 , n11227 );
or ( n12617 , n12615 , n12616 );
or ( n12618 , n11184 , n11231 );
nand ( n12619 , n12617 , n12618 );
not ( n12620 , n12619 );
nand ( n12621 , n12614 , n12620 );
nand ( n12622 , n12560 , n12621 );
and ( n12623 , n12597 , n12576 );
not ( n12624 , n12566 );
and ( n12625 , n12624 , n12572 );
nor ( n12626 , n12623 , n12625 );
and ( n12627 , n10822 , n10815 );
not ( n12628 , n12564 );
nor ( n12629 , n12627 , n12628 );
not ( n12630 , n12583 );
not ( n12631 , n10679 );
not ( n12632 , n12631 );
and ( n12633 , n12630 , n12632 );
and ( n12634 , n497 , n11886 );
not ( n12635 , n558 );
nor ( n12636 , n12634 , n12635 );
and ( n12637 , n12636 , n10811 );
nor ( n12638 , n12633 , n12637 );
xnor ( n12639 , n12629 , n12638 );
nand ( n12640 , n40 , n10740 );
xor ( n12641 , n12639 , n12640 );
not ( n12642 , n12566 );
not ( n12643 , n12593 );
and ( n12644 , n12643 , n11284 );
xor ( n12645 , n38 , n10736 );
and ( n12646 , n12645 , n11641 );
nor ( n12647 , n12644 , n12646 );
not ( n12648 , n12647 );
and ( n12649 , n12642 , n12648 );
and ( n12650 , n12566 , n12647 );
nor ( n12651 , n12649 , n12650 );
and ( n12652 , n12596 , n12587 );
and ( n12653 , n10844 , n12586 );
nor ( n12654 , n12652 , n12653 );
xor ( n12655 , n12651 , n12654 );
xnor ( n12656 , n12641 , n12655 );
xnor ( n12657 , n12626 , n12656 );
and ( n12658 , n12612 , n12608 );
and ( n12659 , n12607 , n12602 );
nor ( n12660 , n12658 , n12659 );
and ( n12661 , n12657 , n12660 );
or ( n12662 , n12622 , n12661 );
not ( n12663 , n12661 );
nand ( n12664 , n12613 , n12619 );
not ( n12665 , n12664 );
and ( n12666 , n12663 , n12665 );
nor ( n12667 , n12657 , n12660 );
nor ( n12668 , n12666 , n12667 );
nand ( n12669 , n12662 , n12668 );
buf ( n12670 , n12669 );
and ( n12671 , n12645 , n11284 );
and ( n12672 , n10579 , n10737 );
and ( n12673 , n37 , n10736 );
nor ( n12674 , n12672 , n12673 );
and ( n12675 , n12674 , n11641 );
nor ( n12676 , n12671 , n12675 );
xnor ( n12677 , n12592 , n12676 );
not ( n12678 , n12636 );
not ( n12679 , n10680 );
or ( n12680 , n12678 , n12679 );
not ( n12681 , n11887 );
not ( n12682 , n10811 );
or ( n12683 , n12681 , n12682 );
nand ( n12684 , n12680 , n12683 );
and ( n12685 , n12677 , n12684 );
not ( n12686 , n12677 );
not ( n12687 , n12684 );
and ( n12688 , n12686 , n12687 );
nor ( n12689 , n12685 , n12688 );
or ( n12690 , n12640 , n12639 );
or ( n12691 , n12629 , n12638 );
nand ( n12692 , n12690 , n12691 );
xor ( n12693 , n12689 , n12692 );
xnor ( n12694 , t_2 , n12693 );
not ( n12695 , n12626 );
not ( n12696 , n12656 );
and ( n12697 , n12695 , n12696 );
and ( n12698 , n12641 , n12655 );
nor ( n12699 , n12697 , n12698 );
nor ( n12700 , n12694 , n12699 );
or ( n12701 , n12684 , n12677 );
or ( n12702 , n12592 , n12676 );
nand ( n12703 , n12701 , n12702 );
not ( n12704 , n12682 );
not ( n12705 , n12679 );
or ( n12706 , n12704 , n12705 );
not ( n12707 , n12681 );
nand ( n12708 , n12706 , n12707 );
not ( n12709 , n12674 );
not ( n12710 , n12588 );
or ( n12711 , n12709 , n12710 );
or ( n12712 , n536 , n12594 );
nand ( n12713 , n12711 , n12712 );
xor ( n12714 , n12708 , n12713 );
and ( n12715 , n38 , n10736 );
xor ( n12716 , n12714 , n12715 );
and ( n12717 , n12716 , n12684 );
not ( n12718 , n12716 );
and ( n12719 , n12718 , n12687 );
nor ( n12720 , n12717 , n12719 );
xnor ( n12721 , n12703 , n12720 );
and ( n12722 , t_3 , n12693 );
and ( n12723 , n12692 , n12689 );
nor ( n12724 , n12722 , n12723 );
nand ( n12725 , n12721 , n12724 );
not ( n12726 , n12725 );
nor ( n12727 , n12721 , n12724 );
nor ( n12728 , n12726 , n12727 );
or ( n12729 , n12700 , n12728 );
or ( n12730 , n12670 , n12729 );
and ( n12731 , n12700 , n12728 );
nand ( n12732 , n12694 , n12699 );
nor ( n12733 , n12732 , n12729 );
nor ( n12734 , n12731 , n12733 , n10526 );
nand ( n12735 , n12730 , n12734 );
not ( n12736 , n12670 );
nand ( n12737 , n12732 , n12728 );
nor ( n12738 , n12736 , n12737 );
or ( n12739 , n12735 , n12738 );
nand ( n12740 , n10555 , n12739 );
and ( n12741 , n10437 , n10246 , n10453 );
not ( n12742 , n12741 );
not ( n12743 , n12742 );
not ( n12744 , n12743 );
not ( n12745 , n10221 );
nor ( n12746 , n10500 , n10515 );
nand ( n12747 , n10490 , n12746 );
not ( n12748 , n12747 );
nand ( n12749 , n12745 , n12748 , n10164 );
nor ( n12750 , n10130 , n12749 );
not ( n12751 , n12750 );
or ( n12752 , n12744 , n12751 );
nand ( n12753 , n12752 , n10526 );
not ( n12754 , n10084 );
or ( n12755 , n12753 , n12754 );
not ( n12756 , n12742 );
nand ( n12757 , n12750 , n10526 , n12756 , n12754 );
not ( n12758 , n12670 );
not ( n12759 , n12700 );
nand ( n12760 , n12759 , n12732 );
not ( n12761 , n12760 );
not ( n12762 , n12761 );
or ( n12763 , n12758 , n12762 );
not ( n12764 , n12670 );
and ( n12765 , n12764 , n12760 );
nor ( n12766 , n12765 , n10526 );
nand ( n12767 , n12763 , n12766 );
nand ( n12768 , n12755 , n12757 , n12767 );
not ( n12769 , n10526 );
buf ( n12770 , n10101 );
nor ( n12771 , n12769 , n12770 );
not ( n12772 , n10129 );
not ( n12773 , n12741 );
nor ( n12774 , n12772 , n12773 );
not ( n12775 , n12749 );
nand ( n12776 , n12771 , n12774 , n12775 );
nand ( n12777 , n12774 , n12775 );
buf ( n12778 , n12770 );
nand ( n12779 , n12777 , n10526 , n12778 );
nand ( n12780 , n12664 , n12622 );
not ( n12781 , n12780 );
nor ( n12782 , n12667 , n12661 );
not ( n12783 , n12782 );
or ( n12784 , n12781 , n12783 );
not ( n12785 , n12780 );
not ( n12786 , n12782 );
and ( n12787 , n12785 , n12786 );
nor ( n12788 , n12787 , n10526 );
nand ( n12789 , n12784 , n12788 );
nand ( n12790 , n12776 , n12779 , n12789 );
not ( n12791 , n12756 );
not ( n12792 , n12791 );
nand ( n12793 , n12792 , n12775 );
nand ( n12794 , n10526 , n10131 , n10084 , n10553 );
or ( n12795 , n12793 , n12794 );
not ( n12796 , n12673 );
not ( n12797 , n12589 );
and ( n12798 , n535 , n12797 );
not ( n12799 , n12594 );
and ( n12800 , n10740 , n12799 );
nor ( n12801 , n12798 , n12800 );
and ( n12802 , n12796 , n12801 );
nor ( n12803 , n12796 , n12801 );
nor ( n12804 , n12802 , n12803 );
and ( n12805 , n12715 , n12714 );
and ( n12806 , n12708 , n12713 );
nor ( n12807 , n12805 , n12806 );
xnor ( n12808 , n12804 , n12807 );
and ( n12809 , n12703 , n12720 );
and ( n12810 , n12684 , n12716 );
nor ( n12811 , n12809 , n12810 );
nor ( n12812 , n12808 , n12811 );
not ( n12813 , n12812 );
nand ( n12814 , n12808 , n12811 );
nand ( n12815 , n12813 , n12814 );
not ( n12816 , n12815 );
and ( n12817 , n12725 , n12732 );
not ( n12818 , n12817 );
not ( n12819 , n12669 );
or ( n12820 , n12818 , n12819 );
and ( n12821 , n12725 , n12700 );
nor ( n12822 , n12821 , n12727 );
nand ( n12823 , n12820 , n12822 );
not ( n12824 , n12823 );
and ( n12825 , n12816 , n12824 );
and ( n12826 , n12815 , n12823 );
nor ( n12827 , n12825 , n12826 );
or ( n12828 , n10526 , n12827 );
nand ( n12829 , n12795 , n12828 );
and ( n12830 , n10526 , n10129 );
nor ( n12831 , n12742 , n12749 );
not ( n12832 , n12560 );
not ( n12833 , n12832 );
nand ( n12834 , n12664 , n12621 );
not ( n12835 , n12834 );
and ( n12836 , n12833 , n12835 );
not ( n12837 , n12834 );
or ( n12838 , n12560 , n12837 );
not ( n12839 , n10526 );
nand ( n12840 , n12838 , n12839 );
nor ( n12841 , n12836 , n12840 );
nor ( n12842 , n12830 , n12831 , n12841 );
not ( n12843 , n12775 );
not ( n12844 , n10526 );
nor ( n12845 , n12844 , n10129 );
nor ( n12846 , n12843 , n12845 , n12841 , n12742 );
nor ( n12847 , n12842 , n12846 );
not ( n12848 , n10221 );
nand ( n12849 , n12848 , n10454 , n12748 );
buf ( n12850 , n10153 );
nor ( n12851 , n12849 , n12850 );
not ( n12852 , n10163 );
nand ( n12853 , n10526 , n12852 );
or ( n12854 , n12851 , n12853 );
not ( n12855 , n10526 );
nor ( n12856 , n12855 , n12852 );
not ( n12857 , n12849 );
not ( n12858 , n12850 );
nand ( n12859 , n12856 , n12857 , n12858 );
not ( n12860 , n10526 );
and ( n12861 , n12557 , n12558 );
nor ( n12862 , n12861 , n11176 );
not ( n12863 , n11057 );
not ( n12864 , n11240 );
nor ( n12865 , n12864 , n11237 );
or ( n12866 , n12862 , n12863 , n12865 );
not ( n12867 , n11178 );
or ( n12868 , n12867 , n12865 );
and ( n12869 , n12867 , n12865 );
nand ( n12870 , n12862 , n12869 );
nand ( n12871 , n12868 , n12870 );
and ( n12872 , n12863 , n12867 , n12865 );
nor ( n12873 , n12871 , n12872 );
nand ( n12874 , n12866 , n12873 );
nand ( n12875 , n12860 , n12874 );
nand ( n12876 , n12854 , n12859 , n12875 );
not ( n12877 , n10526 );
not ( n12878 , n12877 );
nand ( n12879 , n12878 , n12849 );
or ( n12880 , n12879 , n12850 );
nand ( n12881 , n12850 , n10526 , n12857 );
nand ( n12882 , n12867 , n11057 );
or ( n12883 , n12862 , n12882 );
and ( n12884 , n12862 , n12882 );
nor ( n12885 , n12884 , n10526 );
nand ( n12886 , n12883 , n12885 );
nand ( n12887 , n12880 , n12881 , n12886 );
not ( n12888 , n10500 );
not ( n12889 , n12888 );
buf ( n12890 , n10516 );
not ( n12891 , n12890 );
nand ( n12892 , n12889 , n10526 , n12891 , n10493 );
not ( n12893 , n12890 );
nand ( n12894 , n12893 , n10493 );
not ( n12895 , n10526 );
nor ( n12896 , n12895 , n12889 );
and ( n12897 , n12894 , n12896 );
not ( n12898 , n11705 );
nor ( n12899 , n12898 , n11449 );
not ( n12900 , n12552 );
or ( n12901 , n12900 , n12554 );
nand ( n12902 , n12901 , n11703 );
and ( n12903 , n12899 , n12902 );
nor ( n12904 , n12899 , n12902 );
nor ( n12905 , n12903 , n12904 , n10526 );
nor ( n12906 , n12897 , n12905 );
nand ( n12907 , n12892 , n12906 );
buf ( n12908 , n10220 );
nor ( n12909 , n12742 , n12908 );
not ( n12910 , n10526 );
buf ( n12911 , n10201 );
not ( n12912 , n12911 );
nor ( n12913 , n12910 , n12912 );
nand ( n12914 , n12909 , n12748 , n12913 );
not ( n12915 , n12557 );
not ( n12916 , n11176 );
nand ( n12917 , n12916 , n12558 );
or ( n12918 , n12915 , n12917 );
nand ( n12919 , n12915 , n12917 );
not ( n12920 , n10526 );
nand ( n12921 , n12918 , n12919 , n12920 );
not ( n12922 , n12773 );
nand ( n12923 , n12922 , n12748 , n12911 );
not ( n12924 , n10526 );
not ( n12925 , n12908 );
nor ( n12926 , n12924 , n12925 );
nand ( n12927 , n12923 , n12926 );
nand ( n12928 , n12914 , n12921 , n12927 );
nand ( n12929 , n10493 , n10517 );
nand ( n12930 , n12913 , n12929 );
not ( n12931 , n12911 );
nand ( n12932 , n12931 , n10526 , n10493 , n10517 );
and ( n12933 , n12902 , n11705 );
nor ( n12934 , n12933 , n11449 );
nand ( n12935 , n11709 , n11349 );
or ( n12936 , n12934 , n12935 );
and ( n12937 , n12934 , n12935 );
nor ( n12938 , n12937 , n10526 );
nand ( n12939 , n12936 , n12938 );
nand ( n12940 , n12930 , n12932 , n12939 );
nand ( n12941 , n12891 , n10526 , n10492 );
not ( n12942 , n11702 );
nand ( n12943 , n12942 , n11567 );
and ( n12944 , n12553 , n12552 );
nor ( n12945 , n12944 , n11700 );
or ( n12946 , n12943 , n12945 );
and ( n12947 , n12943 , n12945 );
nor ( n12948 , n12947 , n10526 );
nand ( n12949 , n12946 , n12948 );
not ( n12950 , n12891 );
nand ( n12951 , n12950 , n10526 , n10493 );
nand ( n12952 , n12941 , n12949 , n12951 );
buf ( n12953 , n10471 );
not ( n12954 , n12742 );
not ( n12955 , n10489 );
nand ( n12956 , n12954 , n10526 , n12955 );
or ( n12957 , n12953 , n12956 );
not ( n12958 , n11700 );
nand ( n12959 , n12958 , n12553 );
or ( n12960 , n12900 , n12959 );
and ( n12961 , n12900 , n12959 );
nor ( n12962 , n12961 , n10526 );
nand ( n12963 , n12960 , n12962 );
not ( n12964 , n12773 );
nand ( n12965 , n12964 , n12955 );
nand ( n12966 , n12953 , n10526 , n12965 );
nand ( n12967 , n12957 , n12963 , n12966 );
not ( n12968 , n12791 );
not ( n12969 , n10485 );
not ( n12970 , n12969 );
not ( n12971 , n10474 );
and ( n12972 , n12970 , n12971 );
and ( n12973 , n12969 , n10474 );
nor ( n12974 , n12972 , n12973 );
not ( n12975 , n12974 );
not ( n12976 , n12975 );
or ( n12977 , n12968 , n12976 );
and ( n12978 , n12922 , n12974 );
not ( n12979 , n10526 );
nor ( n12980 , n12978 , n12979 );
nand ( n12981 , n12977 , n12980 );
not ( n12982 , n10526 );
not ( n12983 , n12550 );
nor ( n12984 , n12983 , n11785 );
not ( n12985 , n12984 );
and ( n12986 , n12543 , n12547 );
not ( n12987 , n12986 );
or ( n12988 , n12985 , n12987 );
or ( n12989 , n12984 , n12986 );
nand ( n12990 , n12988 , n12989 );
nand ( n12991 , n12982 , n12990 );
nand ( n12992 , n12981 , n12991 );
not ( n12993 , n10526 );
not ( n12994 , n12993 );
or ( n12995 , n12537 , n12538 );
not ( n12996 , n12995 );
nand ( n12997 , n11928 , n12540 );
not ( n12998 , n12997 );
or ( n12999 , n12996 , n12998 );
or ( n13000 , n12995 , n12997 );
nand ( n13001 , n12999 , n13000 );
not ( n13002 , n13001 );
or ( n13003 , n12994 , n13002 );
not ( n13004 , n10254 );
not ( n13005 , n10262 );
nor ( n13006 , n13004 , n13005 );
not ( n13007 , n10380 );
not ( n13008 , n10433 );
nand ( n13009 , n10402 , n10421 , n13008 );
nor ( n13010 , n13007 , n13009 );
nand ( n13011 , n10453 , n13006 , n13010 );
not ( n13012 , n13011 );
nor ( n13013 , n10233 , n13012 );
not ( n13014 , n13013 );
not ( n13015 , n10233 );
nor ( n13016 , n13015 , n13011 );
not ( n13017 , n13016 );
nand ( n13018 , n13014 , n10526 , n13017 );
nand ( n13019 , n13003 , n13018 );
not ( n13020 , n10245 );
not ( n13021 , n13020 );
nand ( n13022 , n13021 , n10526 , n13016 );
not ( n13023 , n10526 );
not ( n13024 , n13020 );
nor ( n13025 , n13023 , n13024 );
nand ( n13026 , n13017 , n13025 );
nand ( n13027 , n12547 , n11866 );
not ( n13028 , n12542 );
or ( n13029 , n13027 , n13028 );
and ( n13030 , n13027 , n13028 );
nor ( n13031 , n13030 , n10526 );
nand ( n13032 , n13029 , n13031 );
nand ( n13033 , n13022 , n13026 , n13032 );
not ( n13034 , n10526 );
not ( n13035 , n13034 );
not ( n13036 , n12531 );
not ( n13037 , n13036 );
or ( n13038 , n12538 , n12536 );
not ( n13039 , n13038 );
or ( n13040 , n13037 , n13039 );
or ( n13041 , n13036 , n13038 );
nand ( n13042 , n13040 , n13041 );
not ( n13043 , n13042 );
or ( n13044 , n13035 , n13043 );
not ( n13045 , n13006 );
not ( n13046 , n13010 );
nor ( n13047 , n13045 , n13046 );
nor ( n13048 , n13047 , n10453 );
not ( n13049 , n13048 );
nand ( n13050 , n13049 , n10526 , n13011 );
nand ( n13051 , n13044 , n13050 );
not ( n13052 , n10526 );
not ( n13053 , n13052 );
not ( n13054 , n12509 );
not ( n13055 , n12530 );
nand ( n13056 , n13055 , n12527 );
not ( n13057 , n13056 );
or ( n13058 , n13054 , n13057 );
or ( n13059 , n12509 , n13056 );
nand ( n13060 , n13058 , n13059 );
not ( n13061 , n13060 );
or ( n13062 , n13053 , n13061 );
not ( n13063 , n10437 );
not ( n13064 , n10254 );
not ( n13065 , n13005 );
not ( n13066 , n10435 );
nand ( n13067 , n13065 , n13066 );
nand ( n13068 , n13064 , n13067 );
nand ( n13069 , n13063 , n13068 , n10526 );
nand ( n13070 , n13062 , n13069 );
nand ( n13071 , n13005 , n10525 , n13066 );
not ( n13072 , n12466 );
nand ( n13073 , n12508 , n12505 );
or ( n13074 , n13072 , n13073 );
nand ( n13075 , n13072 , n13073 );
not ( n13076 , n10525 );
nand ( n13077 , n13074 , n13075 , n13076 );
not ( n13078 , n13066 );
nand ( n13079 , n13078 , n10525 , n10262 );
nand ( n13080 , n13071 , n13077 , n13079 );
not ( n13081 , n12796 );
not ( n13082 , n13081 );
or ( n13083 , n12799 , n12797 );
nand ( n13084 , n13083 , n10740 );
not ( n13085 , n13084 );
and ( n13086 , n13082 , n13085 );
and ( n13087 , n13081 , n13084 );
nor ( n13088 , n13086 , n13087 );
not ( n13089 , n13088 );
not ( n13090 , n508 );
or ( n13091 , n12804 , n12807 );
or ( n13092 , n13081 , n12801 );
nand ( n13093 , n13091 , n13092 );
not ( n13094 , n13093 );
or ( n13095 , n13090 , n13094 );
or ( n13096 , n508 , n13093 );
nand ( n13097 , n13095 , n13096 );
not ( n13098 , n13097 );
or ( n13099 , n13089 , n13098 );
or ( n13100 , n13088 , n13097 );
nand ( n13101 , n13099 , n13100 );
not ( n13102 , n13101 );
not ( n13103 , n12661 );
nand ( n13104 , n12817 , n13103 , n12814 , n12621 );
buf ( n13105 , n12559 );
or ( n13106 , n13104 , n13105 );
not ( n13107 , n13104 );
and ( n13108 , n13107 , n11241 );
not ( n13109 , n12817 );
or ( n13110 , n13109 , n12668 );
nand ( n13111 , n13110 , n12822 );
and ( n13112 , n12814 , n13111 );
nor ( n13113 , n13108 , n13112 , n12812 );
nand ( n13114 , n13106 , n13113 );
not ( n13115 , n13114 );
and ( n13116 , n13102 , n13115 );
and ( n13117 , n13101 , n13114 );
nor ( n13118 , n13116 , n13117 );
nor ( n13119 , n10525 , n13118 );
nand ( n13120 , n10380 , n10434 );
not ( n13121 , n13120 );
nor ( n13122 , n13121 , n10402 );
not ( n13123 , n10402 );
or ( n13124 , n13120 , n13123 );
nand ( n13125 , n13124 , n10525 );
or ( n13126 , n13122 , n13125 );
nor ( n13127 , n12150 , n12465 );
not ( n13128 , n13127 );
not ( n13129 , n12463 );
nor ( n13130 , n13129 , n12208 );
not ( n13131 , n13130 );
and ( n13132 , n13128 , n13131 );
and ( n13133 , n13127 , n13130 );
nor ( n13134 , n13132 , n13133 );
or ( n13135 , n10525 , n13134 );
nand ( n13136 , n13126 , n13135 );
not ( n13137 , n10421 );
nor ( n13138 , n13137 , n13007 );
not ( n13139 , n13138 );
nand ( n13140 , n13139 , n10433 );
nand ( n13141 , n13138 , n13008 );
nand ( n13142 , n13140 , n10525 , n13141 );
not ( n13143 , n10525 );
not ( n13144 , n12210 );
nor ( n13145 , n13144 , n12208 );
xor ( n13146 , n13145 , n12462 );
nand ( n13147 , n13143 , n13146 );
nand ( n13148 , n13142 , n13147 );
not ( n13149 , n13137 );
not ( n13150 , n13007 );
or ( n13151 , n13149 , n13150 );
nand ( n13152 , n13151 , n10525 );
or ( n13153 , n13138 , n13152 );
xnor ( n13154 , n12457 , n12255 );
or ( n13155 , n10525 , n13154 );
nand ( n13156 , n13153 , n13155 );
nand ( n13157 , n10525 , n10276 );
or ( n13158 , n13157 , n10379 );
nand ( n13159 , n12456 , n12292 );
not ( n13160 , n12452 );
or ( n13161 , n13159 , n13160 );
and ( n13162 , n13159 , n13160 );
nor ( n13163 , n13162 , n10525 );
nand ( n13164 , n13161 , n13163 );
not ( n13165 , n10525 );
nor ( n13166 , n13165 , n10276 );
nand ( n13167 , n13166 , n10379 );
nand ( n13168 , n13158 , n13164 , n13167 );
not ( n13169 , n10379 );
not ( n13170 , n10293 );
nand ( n13171 , n13170 , n10378 );
nand ( n13172 , n13169 , n13171 );
and ( n13173 , n10525 , n13172 );
and ( n13174 , n12451 , n12330 );
not ( n13175 , n13174 );
nand ( n13176 , n13175 , n12446 );
not ( n13177 , n12446 );
and ( n13178 , n13174 , n13177 );
nor ( n13179 , n13178 , n10525 );
and ( n13180 , n13176 , n13179 );
nor ( n13181 , n13173 , n13180 );
buf ( n13182 , n10359 );
nand ( n13183 , n10377 , n13182 );
not ( n13184 , n13183 );
nor ( n13185 , n10367 , n13184 );
not ( n13186 , n10367 );
or ( n13187 , n13186 , n13183 );
nand ( n13188 , n13187 , n10525 );
or ( n13189 , n13185 , n13188 );
xnor ( n13190 , n12424 , n12441 );
or ( n13191 , n10525 , n13190 );
nand ( n13192 , n13189 , n13191 );
not ( n13193 , n10377 );
not ( n13194 , n13182 );
nor ( n13195 , n13193 , n13194 );
or ( n13196 , n10377 , n13182 );
nand ( n13197 , n13196 , n10525 );
or ( n13198 , n13195 , n13197 );
not ( n13199 , n12385 );
not ( n13200 , n12420 );
and ( n13201 , n13199 , n13200 );
and ( n13202 , n12385 , n12420 );
nor ( n13203 , n13201 , n13202 );
or ( n13204 , n10525 , n13203 );
nand ( n13205 , n13198 , n13204 );
nand ( n13206 , n10358 , n10302 );
not ( n13207 , n13206 );
not ( n13208 , n10354 );
not ( n13209 , n13208 );
nor ( n13210 , n13207 , n13209 );
or ( n13211 , n13206 , n13208 );
nand ( n13212 , n13211 , n10525 );
or ( n13213 , n13210 , n13212 );
xnor ( n13214 , n12358 , n12382 );
or ( n13215 , n10525 , n13214 );
nand ( n13216 , n13213 , n13215 );
and ( n13217 , n10353 , n10349 );
nor ( n13218 , n10333 , n13217 );
not ( n13219 , n10333 );
not ( n13220 , n13217 );
or ( n13221 , n13219 , n13220 );
nand ( n13222 , n13221 , n10524 );
or ( n13223 , n13218 , n13222 );
not ( n13224 , n12354 );
nand ( n13225 , n12345 , n12356 );
not ( n13226 , n13225 );
and ( n13227 , n13224 , n13226 );
and ( n13228 , n12354 , n13225 );
nor ( n13229 , n13227 , n13228 );
or ( n13230 , n10525 , n13229 );
nand ( n13231 , n13223 , n13230 );
nor ( n13232 , n12347 , n12353 );
or ( n13233 , n13232 , n10524 , n12354 );
not ( n13234 , n10332 );
or ( n13235 , n10322 , n10331 );
nand ( n13236 , n13235 , n10524 );
or ( n13237 , n13234 , n13236 );
nand ( n13238 , n13233 , n13237 );
or ( n13239 , n19 , n10315 );
nand ( n13240 , n13239 , n10524 );
or ( n13241 , n10316 , n13240 );
or ( n13242 , n12346 , n10524 );
nand ( n13243 , n13241 , n13242 );
not ( n13244 , n9839 );
nand ( n13245 , n9987 , n10305 );
not ( n13246 , n13245 );
or ( n13247 , n13244 , n13246 );
or ( n13248 , n9839 , n13245 );
nand ( n13249 , n13247 , n13248 );
not ( n13250 , n9761 );
not ( n13251 , n13250 );
not ( n13252 , n9803 );
not ( n13253 , n13252 );
and ( n13254 , n13251 , n13253 );
nor ( n13255 , n13254 , n9801 );
not ( n13256 , n13255 );
not ( n13257 , n9835 );
nor ( n13258 , n13257 , n9838 );
not ( n13259 , n13258 );
or ( n13260 , n13256 , n13259 );
or ( n13261 , n13255 , n13258 );
nand ( n13262 , n13260 , n13261 );
not ( n13263 , n13250 );
nor ( n13264 , n9801 , n13252 );
not ( n13265 , n13264 );
or ( n13266 , n13263 , n13265 );
or ( n13267 , n13250 , n13264 );
nand ( n13268 , n13266 , n13267 );
xor ( n13269 , n9707 , n9737 );
or ( n13270 , n9758 , n13269 );
not ( n13271 , n9738 );
not ( n13272 , n9759 );
or ( n13273 , n13271 , n13272 );
nand ( n13274 , n13273 , n9758 );
nand ( n13275 , n13270 , n13274 );
not ( n13276 , n9741 );
not ( n13277 , n9757 );
not ( n13278 , n13277 );
or ( n13279 , n13276 , n13278 );
or ( n13280 , n9741 , n13277 );
nand ( n13281 , n13279 , n13280 );
not ( n13282 , n12850 );
not ( n13283 , n12931 );
endmodule
