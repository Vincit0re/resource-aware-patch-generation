module top (out_0, out_1, out_2, out_3, out_4, out_5, out_6, out_7, out_8, out_9, out_10, out_11, out_12, out_13, out_14, out_15, out_16, out_17, out_18, out_19, out_20, out_21, in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, in_17, in_18, in_19, in_20, in_21);
	input in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, in_17, in_18, in_19, in_20, in_21;
	output out_0, out_1, out_2, out_3, out_4, out_5, out_6, out_7, out_8, out_9, out_10, out_11, out_12, out_13, out_14, out_15, out_16, out_17, out_18, out_19, out_20, out_21;
	wire gm_n100, gm_n1000, gm_n10000, gm_n10001, gm_n10002, gm_n10003, gm_n10004, gm_n10005, gm_n10006, gm_n10007, gm_n10008, gm_n10009, gm_n1001, gm_n10010, gm_n10011, gm_n10012, gm_n10013, gm_n10014, gm_n10015, gm_n10016, gm_n10017, gm_n10018, gm_n10019, gm_n1002, gm_n10020, gm_n10021, gm_n10022, gm_n10023, gm_n10024, gm_n10025, gm_n10026, gm_n10027, gm_n10028, gm_n10029, gm_n1003, gm_n10030, gm_n10031, gm_n10032, gm_n10033, gm_n10034, gm_n10035, gm_n10036, gm_n10037, gm_n10038, gm_n10039, gm_n1004, gm_n10040, gm_n10041, gm_n10042, gm_n10043, gm_n10044, gm_n10045, gm_n10046, gm_n10047, gm_n10048, gm_n10049, gm_n1005, gm_n10050, gm_n10051, gm_n10052, gm_n10053, gm_n10054, gm_n10055, gm_n10056, gm_n10057, gm_n10058, gm_n10059, gm_n1006, gm_n10060, gm_n10061, gm_n10062, gm_n10063, gm_n10064, gm_n10065, gm_n10066, gm_n10067, gm_n10068, gm_n10069, gm_n1007, gm_n10070, gm_n10071, gm_n10072, gm_n10073, gm_n10074, gm_n10075, gm_n10076, gm_n10077, gm_n10078, gm_n10079, gm_n1008, gm_n10080, gm_n10081, gm_n10082, gm_n10083, gm_n10084, gm_n10085, gm_n10086, gm_n10087, gm_n10088, gm_n10089, gm_n1009, gm_n10090, gm_n10091, gm_n10092, gm_n10093, gm_n10094, gm_n10095, gm_n10096, gm_n10097, gm_n10098, gm_n10099, gm_n101, gm_n1010, gm_n10100, gm_n10101, gm_n10102, gm_n10103, gm_n10104, gm_n10105, gm_n10106, gm_n10107, gm_n10108, gm_n10109, gm_n1011, gm_n10110, gm_n10111, gm_n10112, gm_n10113, gm_n10114, gm_n10115, gm_n10116, gm_n10117, gm_n10118, gm_n10119, gm_n1012, gm_n10120, gm_n10121, gm_n10122, gm_n10123, gm_n10124, gm_n10125, gm_n10126, gm_n10127, gm_n10128, gm_n10129, gm_n1013, gm_n10130, gm_n10131, gm_n10132, gm_n10133, gm_n10134, gm_n10135, gm_n10136, gm_n10137, gm_n10138, gm_n10139, gm_n1014, gm_n10140, gm_n10141, gm_n10142, gm_n10143, gm_n10144, gm_n10145, gm_n10146, gm_n10147, gm_n10148, gm_n10149, gm_n1015, gm_n10150, gm_n10151, gm_n10152, gm_n10153, gm_n10154, gm_n10155, gm_n10156, gm_n10157, gm_n10158, gm_n10159, gm_n1016, gm_n10160, gm_n10161, gm_n10162, gm_n10163, gm_n10164, gm_n10165, gm_n10166, gm_n10167, gm_n10168, gm_n10169, gm_n1017, gm_n10170, gm_n10171, gm_n10172, gm_n10173, gm_n10174, gm_n10175, gm_n10176, gm_n10177, gm_n10178, gm_n10179, gm_n1018, gm_n10180, gm_n10181, gm_n10182, gm_n10183, gm_n10184, gm_n10185, gm_n10186, gm_n10187, gm_n10188, gm_n10189, gm_n1019, gm_n10190, gm_n10191, gm_n10192, gm_n10193, gm_n10194, gm_n10195, gm_n10196, gm_n10197, gm_n10198, gm_n10199, gm_n102, gm_n1020, gm_n10200, gm_n10201, gm_n10202, gm_n10203, gm_n10204, gm_n10205, gm_n10206, gm_n10207, gm_n10208, gm_n10209, gm_n1021, gm_n10210, gm_n10211, gm_n10212, gm_n10213, gm_n10214, gm_n10215, gm_n10216, gm_n10217, gm_n10218, gm_n10219, gm_n1022, gm_n10220, gm_n10221, gm_n10222, gm_n10223, gm_n10224, gm_n10225, gm_n10226, gm_n10227, gm_n10228, gm_n10229, gm_n1023, gm_n10230, gm_n10231, gm_n10232, gm_n10233, gm_n10234, gm_n10235, gm_n10236, gm_n10237, gm_n10238, gm_n10239, gm_n1024, gm_n10240, gm_n10241, gm_n10242, gm_n10243, gm_n10244, gm_n10245, gm_n10246, gm_n10247, gm_n10248, gm_n10249, gm_n1025, gm_n10250, gm_n10251, gm_n10252, gm_n10253, gm_n10254, gm_n10255, gm_n10256, gm_n10257, gm_n10258, gm_n10259, gm_n1026, gm_n10260, gm_n10261, gm_n10262, gm_n10263, gm_n10264, gm_n10265, gm_n10266, gm_n10267, gm_n10268, gm_n10269, gm_n1027, gm_n10270, gm_n10271, gm_n10272, gm_n10273, gm_n10274, gm_n10275, gm_n10276, gm_n10277, gm_n10278, gm_n10279, gm_n1028, gm_n10280, gm_n10281, gm_n10282, gm_n10283, gm_n10284, gm_n10285, gm_n10286, gm_n10287, gm_n10288, gm_n10289, gm_n1029, gm_n10290, gm_n10291, gm_n10292, gm_n10293, gm_n10294, gm_n10295, gm_n10296, gm_n10297, gm_n10298, gm_n10299, gm_n103, gm_n1030, gm_n10300, gm_n10301, gm_n10302, gm_n10303, gm_n10304, gm_n10305, gm_n10306, gm_n10307, gm_n10308, gm_n10309, gm_n1031, gm_n10310, gm_n10311, gm_n10312, gm_n10313, gm_n10314, gm_n10315, gm_n10316, gm_n10317, gm_n10318, gm_n10319, gm_n1032, gm_n10320, gm_n10321, gm_n10322, gm_n10323, gm_n10324, gm_n10325, gm_n10326, gm_n10327, gm_n10328, gm_n10329, gm_n1033, gm_n10330, gm_n10331, gm_n10332, gm_n10333, gm_n10334, gm_n10335, gm_n10336, gm_n10337, gm_n10338, gm_n10339, gm_n1034, gm_n10340, gm_n10341, gm_n10342, gm_n10343, gm_n10344, gm_n10345, gm_n10346, gm_n10347, gm_n10348, gm_n10349, gm_n1035, gm_n10350, gm_n10351, gm_n10352, gm_n10353, gm_n10354, gm_n10355, gm_n10356, gm_n10357, gm_n10358, gm_n10359, gm_n1036, gm_n10360, gm_n10361, gm_n10362, gm_n10363, gm_n10364, gm_n10365, gm_n10366, gm_n10367, gm_n10368, gm_n10369, gm_n1037, gm_n10370, gm_n10371, gm_n10372, gm_n10373, gm_n10374, gm_n10375, gm_n10376, gm_n10377, gm_n10378, gm_n10379, gm_n1038, gm_n10380, gm_n10381, gm_n10382, gm_n10383, gm_n10384, gm_n10385, gm_n10386, gm_n10387, gm_n10388, gm_n10389, gm_n1039, gm_n10390, gm_n10391, gm_n10392, gm_n10393, gm_n10394, gm_n10395, gm_n10396, gm_n10397, gm_n10398, gm_n10399, gm_n104, gm_n1040, gm_n10400, gm_n10401, gm_n10402, gm_n10403, gm_n10404, gm_n10405, gm_n10406, gm_n10407, gm_n10408, gm_n10409, gm_n1041, gm_n10410, gm_n10411, gm_n10412, gm_n10413, gm_n10414, gm_n10415, gm_n10416, gm_n10417, gm_n10418, gm_n10419, gm_n1042, gm_n10420, gm_n10421, gm_n10422, gm_n10423, gm_n10424, gm_n10425, gm_n10426, gm_n10427, gm_n10428, gm_n10429, gm_n1043, gm_n10430, gm_n10431, gm_n10432, gm_n10433, gm_n10434, gm_n10435, gm_n10436, gm_n10437, gm_n10438, gm_n10439, gm_n1044, gm_n10440, gm_n10441, gm_n10442, gm_n10443, gm_n10444, gm_n10445, gm_n10446, gm_n10447, gm_n10448, gm_n10449, gm_n1045, gm_n10450, gm_n10451, gm_n10452, gm_n10453, gm_n10454, gm_n10455, gm_n10456, gm_n10457, gm_n10458, gm_n10459, gm_n1046, gm_n10460, gm_n10461, gm_n10462, gm_n10463, gm_n10464, gm_n10465, gm_n10466, gm_n10467, gm_n10468, gm_n10469, gm_n1047, gm_n10470, gm_n10471, gm_n10472, gm_n10473, gm_n10474, gm_n10475, gm_n10476, gm_n10477, gm_n10478, gm_n10479, gm_n1048, gm_n10480, gm_n10481, gm_n10482, gm_n10483, gm_n10484, gm_n10485, gm_n10486, gm_n10487, gm_n10488, gm_n10489, gm_n1049, gm_n10490, gm_n10492, gm_n10493, gm_n10494, gm_n10495, gm_n10496, gm_n10497, gm_n10498, gm_n10499, gm_n105, gm_n1050, gm_n10500, gm_n10501, gm_n10502, gm_n10503, gm_n10504, gm_n10505, gm_n10506, gm_n10507, gm_n10508, gm_n10509, gm_n1051, gm_n10510, gm_n10511, gm_n10512, gm_n10513, gm_n10514, gm_n10515, gm_n10516, gm_n10517, gm_n10518, gm_n10519, gm_n1052, gm_n10520, gm_n10521, gm_n10522, gm_n10523, gm_n10524, gm_n10525, gm_n10526, gm_n10527, gm_n10528, gm_n10529, gm_n1053, gm_n10530, gm_n10531, gm_n10532, gm_n10533, gm_n10534, gm_n10535, gm_n10536, gm_n10537, gm_n10538, gm_n10539, gm_n1054, gm_n10540, gm_n10541, gm_n10542, gm_n10543, gm_n10544, gm_n10545, gm_n10546, gm_n10547, gm_n10548, gm_n10549, gm_n1055, gm_n10550, gm_n10551, gm_n10552, gm_n10553, gm_n10554, gm_n10555, gm_n10556, gm_n10557, gm_n10558, gm_n10559, gm_n1056, gm_n10560, gm_n10561, gm_n10562, gm_n10563, gm_n10564, gm_n10565, gm_n10566, gm_n10567, gm_n10568, gm_n10569, gm_n1057, gm_n10570, gm_n10571, gm_n10572, gm_n10573, gm_n10574, gm_n10575, gm_n10576, gm_n10577, gm_n10578, gm_n10579, gm_n1058, gm_n10580, gm_n10581, gm_n10582, gm_n10583, gm_n10584, gm_n10585, gm_n10586, gm_n10587, gm_n10588, gm_n10589, gm_n1059, gm_n10590, gm_n10591, gm_n10592, gm_n10593, gm_n10594, gm_n10595, gm_n10596, gm_n10597, gm_n10598, gm_n10599, gm_n106, gm_n1060, gm_n10600, gm_n10601, gm_n10602, gm_n10603, gm_n10604, gm_n10605, gm_n10606, gm_n10607, gm_n10608, gm_n10609, gm_n1061, gm_n10610, gm_n10611, gm_n10612, gm_n10613, gm_n10614, gm_n10615, gm_n10616, gm_n10617, gm_n10618, gm_n10619, gm_n1062, gm_n10620, gm_n10621, gm_n10622, gm_n10623, gm_n10624, gm_n10625, gm_n10626, gm_n10627, gm_n10628, gm_n10629, gm_n1063, gm_n10630, gm_n10631, gm_n10632, gm_n10633, gm_n10634, gm_n10635, gm_n10636, gm_n10637, gm_n10638, gm_n10639, gm_n1064, gm_n10640, gm_n10641, gm_n10642, gm_n10643, gm_n10644, gm_n10645, gm_n10646, gm_n10647, gm_n10648, gm_n10649, gm_n1065, gm_n10650, gm_n10651, gm_n10652, gm_n10653, gm_n10654, gm_n10655, gm_n10656, gm_n10657, gm_n10658, gm_n10659, gm_n1066, gm_n10660, gm_n10661, gm_n10662, gm_n10663, gm_n10664, gm_n10665, gm_n10666, gm_n10667, gm_n10668, gm_n10669, gm_n1067, gm_n10670, gm_n10671, gm_n10672, gm_n10673, gm_n10674, gm_n10675, gm_n10676, gm_n10677, gm_n10678, gm_n10679, gm_n1068, gm_n10680, gm_n10681, gm_n10682, gm_n10683, gm_n10684, gm_n10685, gm_n10686, gm_n10687, gm_n10688, gm_n10689, gm_n1069, gm_n10690, gm_n10691, gm_n10692, gm_n10693, gm_n10694, gm_n10695, gm_n10696, gm_n10697, gm_n10698, gm_n10699, gm_n107, gm_n1070, gm_n10700, gm_n10701, gm_n10702, gm_n10703, gm_n10704, gm_n10705, gm_n10706, gm_n10707, gm_n10708, gm_n10709, gm_n1071, gm_n10710, gm_n10711, gm_n10712, gm_n10713, gm_n10714, gm_n10715, gm_n10716, gm_n10717, gm_n10718, gm_n10719, gm_n1072, gm_n10720, gm_n10721, gm_n10722, gm_n10723, gm_n10724, gm_n10725, gm_n10726, gm_n10727, gm_n10728, gm_n10729, gm_n1073, gm_n10730, gm_n10731, gm_n10732, gm_n10733, gm_n10734, gm_n10735, gm_n10736, gm_n10737, gm_n10738, gm_n10739, gm_n1074, gm_n10740, gm_n10741, gm_n10742, gm_n10743, gm_n10744, gm_n10745, gm_n10746, gm_n10747, gm_n10748, gm_n10749, gm_n1075, gm_n10750, gm_n10751, gm_n10752, gm_n10753, gm_n10754, gm_n10755, gm_n10756, gm_n10757, gm_n10758, gm_n10759, gm_n1076, gm_n10760, gm_n10761, gm_n10762, gm_n10763, gm_n10764, gm_n10765, gm_n10766, gm_n10767, gm_n10768, gm_n10769, gm_n1077, gm_n10770, gm_n10771, gm_n10772, gm_n10773, gm_n10774, gm_n10775, gm_n10776, gm_n10777, gm_n10778, gm_n10779, gm_n1078, gm_n10780, gm_n10781, gm_n10782, gm_n10783, gm_n10784, gm_n10785, gm_n10786, gm_n10787, gm_n10788, gm_n10789, gm_n1079, gm_n10790, gm_n10791, gm_n10792, gm_n10793, gm_n10794, gm_n10795, gm_n10796, gm_n10797, gm_n10798, gm_n10799, gm_n108, gm_n1080, gm_n10800, gm_n10801, gm_n10802, gm_n10803, gm_n10804, gm_n10805, gm_n10806, gm_n10807, gm_n10808, gm_n10809, gm_n1081, gm_n10810, gm_n10811, gm_n10812, gm_n10813, gm_n10814, gm_n10815, gm_n10816, gm_n10817, gm_n10818, gm_n10819, gm_n1082, gm_n10820, gm_n10821, gm_n10822, gm_n10823, gm_n10824, gm_n10825, gm_n10826, gm_n10827, gm_n10828, gm_n10829, gm_n1083, gm_n10830, gm_n10831, gm_n10832, gm_n10833, gm_n10834, gm_n10835, gm_n10836, gm_n10837, gm_n10838, gm_n10839, gm_n1084, gm_n10840, gm_n10841, gm_n10842, gm_n10843, gm_n10844, gm_n10845, gm_n10846, gm_n10847, gm_n10848, gm_n10849, gm_n1085, gm_n10850, gm_n10851, gm_n10852, gm_n10853, gm_n10854, gm_n10855, gm_n10856, gm_n10857, gm_n10858, gm_n10859, gm_n1086, gm_n10860, gm_n10861, gm_n10862, gm_n10863, gm_n10864, gm_n10865, gm_n10866, gm_n10867, gm_n10868, gm_n10869, gm_n1087, gm_n10870, gm_n10871, gm_n10872, gm_n10873, gm_n10874, gm_n10875, gm_n10876, gm_n10877, gm_n10878, gm_n10879, gm_n1088, gm_n10880, gm_n10881, gm_n10882, gm_n10883, gm_n10884, gm_n10885, gm_n10886, gm_n10887, gm_n10888, gm_n10889, gm_n1089, gm_n10890, gm_n10891, gm_n10892, gm_n10893, gm_n10894, gm_n10895, gm_n10896, gm_n10897, gm_n10898, gm_n10899, gm_n109, gm_n1090, gm_n10900, gm_n10901, gm_n10902, gm_n10903, gm_n10904, gm_n10905, gm_n10906, gm_n10907, gm_n10908, gm_n10909, gm_n1091, gm_n10910, gm_n10911, gm_n10912, gm_n10913, gm_n10914, gm_n10915, gm_n10916, gm_n10917, gm_n10918, gm_n10919, gm_n1092, gm_n10920, gm_n10921, gm_n10922, gm_n10923, gm_n10924, gm_n10925, gm_n10926, gm_n10927, gm_n10928, gm_n10929, gm_n1093, gm_n10930, gm_n10931, gm_n10932, gm_n10933, gm_n10934, gm_n10935, gm_n10936, gm_n10937, gm_n10938, gm_n10939, gm_n1094, gm_n10940, gm_n10941, gm_n10942, gm_n10943, gm_n10944, gm_n10945, gm_n10946, gm_n10947, gm_n10948, gm_n10949, gm_n1095, gm_n10950, gm_n10951, gm_n10952, gm_n10953, gm_n10954, gm_n10955, gm_n10956, gm_n10957, gm_n10958, gm_n10959, gm_n1096, gm_n10960, gm_n10961, gm_n10962, gm_n10963, gm_n10964, gm_n10965, gm_n10966, gm_n10967, gm_n10968, gm_n10969, gm_n1097, gm_n10970, gm_n10971, gm_n10972, gm_n10973, gm_n10974, gm_n10975, gm_n10976, gm_n10977, gm_n10978, gm_n10979, gm_n1098, gm_n10980, gm_n10981, gm_n10982, gm_n10983, gm_n10984, gm_n10985, gm_n10986, gm_n10987, gm_n10988, gm_n10989, gm_n1099, gm_n10990, gm_n10991, gm_n10992, gm_n10993, gm_n10994, gm_n10995, gm_n10996, gm_n10997, gm_n10998, gm_n10999, gm_n110, gm_n1100, gm_n11000, gm_n11001, gm_n11002, gm_n11004, gm_n11005, gm_n11006, gm_n11007, gm_n11008, gm_n11009, gm_n1101, gm_n11010, gm_n11011, gm_n11012, gm_n11013, gm_n11014, gm_n11015, gm_n11016, gm_n11017, gm_n11018, gm_n11019, gm_n1102, gm_n11020, gm_n11021, gm_n11022, gm_n11023, gm_n11024, gm_n11025, gm_n11026, gm_n11027, gm_n11028, gm_n11029, gm_n1103, gm_n11030, gm_n11031, gm_n11032, gm_n11033, gm_n11034, gm_n11035, gm_n11036, gm_n11037, gm_n11038, gm_n11039, gm_n1104, gm_n11040, gm_n11041, gm_n11042, gm_n11043, gm_n11044, gm_n11045, gm_n11046, gm_n11047, gm_n11048, gm_n11049, gm_n1105, gm_n11050, gm_n11051, gm_n11052, gm_n11053, gm_n11054, gm_n11055, gm_n11056, gm_n11057, gm_n11058, gm_n11059, gm_n1106, gm_n11060, gm_n11061, gm_n11062, gm_n11063, gm_n11064, gm_n11065, gm_n11066, gm_n11067, gm_n11068, gm_n11069, gm_n1107, gm_n11070, gm_n11071, gm_n11072, gm_n11073, gm_n11074, gm_n11075, gm_n11076, gm_n11077, gm_n11078, gm_n11079, gm_n1108, gm_n11080, gm_n11081, gm_n11082, gm_n11083, gm_n11084, gm_n11085, gm_n11086, gm_n11087, gm_n11088, gm_n11089, gm_n1109, gm_n11090, gm_n11091, gm_n11092, gm_n11093, gm_n11094, gm_n11095, gm_n11096, gm_n11097, gm_n11098, gm_n11099, gm_n111, gm_n1110, gm_n11100, gm_n11101, gm_n11102, gm_n11103, gm_n11104, gm_n11105, gm_n11106, gm_n11107, gm_n11108, gm_n11109, gm_n1111, gm_n11110, gm_n11111, gm_n11112, gm_n11113, gm_n11114, gm_n11115, gm_n11116, gm_n11117, gm_n11118, gm_n11119, gm_n1112, gm_n11120, gm_n11121, gm_n11122, gm_n11123, gm_n11124, gm_n11125, gm_n11126, gm_n11127, gm_n11128, gm_n11129, gm_n1113, gm_n11130, gm_n11131, gm_n11132, gm_n11133, gm_n11134, gm_n11135, gm_n11136, gm_n11137, gm_n11138, gm_n11139, gm_n1114, gm_n11140, gm_n11141, gm_n11142, gm_n11143, gm_n11144, gm_n11145, gm_n11146, gm_n11147, gm_n11148, gm_n11149, gm_n1115, gm_n11150, gm_n11151, gm_n11152, gm_n11153, gm_n11154, gm_n11155, gm_n11156, gm_n11157, gm_n11158, gm_n11159, gm_n1116, gm_n11160, gm_n11161, gm_n11162, gm_n11163, gm_n11164, gm_n11165, gm_n11166, gm_n11167, gm_n11168, gm_n11169, gm_n1117, gm_n11170, gm_n11171, gm_n11172, gm_n11173, gm_n11174, gm_n11175, gm_n11176, gm_n11177, gm_n11178, gm_n11179, gm_n1118, gm_n11180, gm_n11181, gm_n11182, gm_n11183, gm_n11184, gm_n11185, gm_n11186, gm_n11187, gm_n11188, gm_n11189, gm_n1119, gm_n11190, gm_n11191, gm_n11192, gm_n11193, gm_n11194, gm_n11195, gm_n11196, gm_n11197, gm_n11198, gm_n11199, gm_n112, gm_n1120, gm_n11200, gm_n11201, gm_n11202, gm_n11203, gm_n11204, gm_n11205, gm_n11206, gm_n11207, gm_n11208, gm_n11209, gm_n1121, gm_n11210, gm_n11211, gm_n11212, gm_n11213, gm_n11214, gm_n11215, gm_n11216, gm_n11217, gm_n11218, gm_n11219, gm_n1122, gm_n11220, gm_n11221, gm_n11222, gm_n11223, gm_n11224, gm_n11225, gm_n11226, gm_n11227, gm_n11228, gm_n11229, gm_n1123, gm_n11230, gm_n11231, gm_n11232, gm_n11233, gm_n11234, gm_n11235, gm_n11236, gm_n11237, gm_n11238, gm_n11239, gm_n1124, gm_n11240, gm_n11241, gm_n11242, gm_n11243, gm_n11244, gm_n11245, gm_n11246, gm_n11247, gm_n11248, gm_n11249, gm_n1125, gm_n11250, gm_n11251, gm_n11252, gm_n11253, gm_n11254, gm_n11255, gm_n11256, gm_n11257, gm_n11258, gm_n11259, gm_n1126, gm_n11260, gm_n11261, gm_n11262, gm_n11263, gm_n11264, gm_n11265, gm_n11266, gm_n11267, gm_n11268, gm_n11269, gm_n1127, gm_n11270, gm_n11271, gm_n11272, gm_n11273, gm_n11274, gm_n11275, gm_n11276, gm_n11277, gm_n11278, gm_n11279, gm_n1128, gm_n11280, gm_n11281, gm_n11282, gm_n11283, gm_n11284, gm_n11285, gm_n11286, gm_n11287, gm_n11288, gm_n11289, gm_n1129, gm_n11290, gm_n11291, gm_n11292, gm_n11293, gm_n11294, gm_n11295, gm_n11296, gm_n11297, gm_n11298, gm_n11299, gm_n113, gm_n1130, gm_n11300, gm_n11301, gm_n11302, gm_n11303, gm_n11304, gm_n11305, gm_n11306, gm_n11307, gm_n11308, gm_n11309, gm_n1131, gm_n11310, gm_n11311, gm_n11312, gm_n11313, gm_n11314, gm_n11315, gm_n11316, gm_n11317, gm_n11318, gm_n11319, gm_n1132, gm_n11320, gm_n11321, gm_n11322, gm_n11323, gm_n11324, gm_n11325, gm_n11326, gm_n11327, gm_n11328, gm_n11329, gm_n1133, gm_n11330, gm_n11331, gm_n11332, gm_n11333, gm_n11334, gm_n11335, gm_n11336, gm_n11337, gm_n11338, gm_n11339, gm_n1134, gm_n11340, gm_n11341, gm_n11342, gm_n11343, gm_n11344, gm_n11345, gm_n11346, gm_n11347, gm_n11348, gm_n11349, gm_n1135, gm_n11350, gm_n11351, gm_n11352, gm_n11353, gm_n11354, gm_n11355, gm_n11356, gm_n11357, gm_n11358, gm_n11359, gm_n1136, gm_n11360, gm_n11361, gm_n11362, gm_n11363, gm_n11364, gm_n11365, gm_n11366, gm_n11367, gm_n11368, gm_n11369, gm_n1137, gm_n11370, gm_n11371, gm_n11372, gm_n11373, gm_n11374, gm_n11375, gm_n11376, gm_n11377, gm_n11378, gm_n11379, gm_n1138, gm_n11380, gm_n11381, gm_n11382, gm_n11383, gm_n11384, gm_n11385, gm_n11386, gm_n11387, gm_n11388, gm_n11389, gm_n1139, gm_n11390, gm_n11391, gm_n11392, gm_n11393, gm_n11394, gm_n11395, gm_n11396, gm_n11397, gm_n11398, gm_n11399, gm_n114, gm_n1140, gm_n11400, gm_n11401, gm_n11402, gm_n11403, gm_n11404, gm_n11405, gm_n11406, gm_n11407, gm_n11408, gm_n11409, gm_n1141, gm_n11410, gm_n11411, gm_n11412, gm_n11413, gm_n11414, gm_n11415, gm_n11416, gm_n11417, gm_n11418, gm_n11419, gm_n1142, gm_n11420, gm_n11421, gm_n11422, gm_n11423, gm_n11424, gm_n11425, gm_n11426, gm_n11427, gm_n11428, gm_n11429, gm_n1143, gm_n11430, gm_n11431, gm_n11432, gm_n11433, gm_n11434, gm_n11435, gm_n11436, gm_n11437, gm_n11438, gm_n11439, gm_n1144, gm_n11440, gm_n11441, gm_n11442, gm_n11443, gm_n11444, gm_n11445, gm_n11446, gm_n11447, gm_n11448, gm_n11449, gm_n1145, gm_n11450, gm_n11451, gm_n11452, gm_n11453, gm_n11454, gm_n11455, gm_n11456, gm_n11457, gm_n11458, gm_n11459, gm_n1146, gm_n11460, gm_n11461, gm_n11462, gm_n11463, gm_n11464, gm_n11465, gm_n11466, gm_n11467, gm_n11468, gm_n11469, gm_n1147, gm_n11470, gm_n11471, gm_n11472, gm_n11473, gm_n11474, gm_n11475, gm_n11476, gm_n11477, gm_n11478, gm_n11479, gm_n1148, gm_n11480, gm_n11481, gm_n11482, gm_n11483, gm_n11484, gm_n11485, gm_n11486, gm_n11487, gm_n11488, gm_n11489, gm_n1149, gm_n11490, gm_n11491, gm_n11492, gm_n11493, gm_n11494, gm_n11495, gm_n11496, gm_n11497, gm_n11498, gm_n11499, gm_n115, gm_n1150, gm_n11500, gm_n11502, gm_n11503, gm_n11504, gm_n11505, gm_n11506, gm_n11507, gm_n11508, gm_n11509, gm_n1151, gm_n11510, gm_n11511, gm_n11512, gm_n11513, gm_n11514, gm_n11515, gm_n11516, gm_n11517, gm_n11518, gm_n11519, gm_n1152, gm_n11520, gm_n11521, gm_n11522, gm_n11523, gm_n11524, gm_n11525, gm_n11526, gm_n11527, gm_n11528, gm_n11529, gm_n1153, gm_n11530, gm_n11531, gm_n11532, gm_n11533, gm_n11534, gm_n11535, gm_n11536, gm_n11537, gm_n11538, gm_n11539, gm_n1154, gm_n11540, gm_n11541, gm_n11542, gm_n11543, gm_n11544, gm_n11545, gm_n11546, gm_n11547, gm_n11548, gm_n11549, gm_n1155, gm_n11550, gm_n11551, gm_n11552, gm_n11553, gm_n11554, gm_n11555, gm_n11556, gm_n11557, gm_n11558, gm_n11559, gm_n1156, gm_n11560, gm_n11561, gm_n11562, gm_n11563, gm_n11564, gm_n11565, gm_n11566, gm_n11567, gm_n11568, gm_n11569, gm_n1157, gm_n11570, gm_n11571, gm_n11572, gm_n11573, gm_n11574, gm_n11575, gm_n11576, gm_n11577, gm_n11578, gm_n11579, gm_n1158, gm_n11580, gm_n11581, gm_n11582, gm_n11583, gm_n11584, gm_n11585, gm_n11586, gm_n11587, gm_n11588, gm_n11589, gm_n1159, gm_n11590, gm_n11591, gm_n11592, gm_n11593, gm_n11594, gm_n11595, gm_n11596, gm_n11597, gm_n11598, gm_n11599, gm_n116, gm_n1160, gm_n11600, gm_n11601, gm_n11602, gm_n11603, gm_n11604, gm_n11605, gm_n11606, gm_n11607, gm_n11608, gm_n11609, gm_n1161, gm_n11610, gm_n11611, gm_n11612, gm_n11613, gm_n11614, gm_n11615, gm_n11616, gm_n11617, gm_n11618, gm_n11619, gm_n1162, gm_n11620, gm_n11621, gm_n11622, gm_n11623, gm_n11624, gm_n11625, gm_n11626, gm_n11627, gm_n11628, gm_n11629, gm_n1163, gm_n11630, gm_n11631, gm_n11632, gm_n11633, gm_n11634, gm_n11635, gm_n11636, gm_n11637, gm_n11638, gm_n11639, gm_n1164, gm_n11640, gm_n11641, gm_n11642, gm_n11643, gm_n11644, gm_n11645, gm_n11646, gm_n11647, gm_n11648, gm_n11649, gm_n1165, gm_n11650, gm_n11651, gm_n11652, gm_n11653, gm_n11654, gm_n11655, gm_n11656, gm_n11657, gm_n11658, gm_n11659, gm_n1166, gm_n11660, gm_n11661, gm_n11662, gm_n11663, gm_n11664, gm_n11665, gm_n11666, gm_n11667, gm_n11668, gm_n11669, gm_n1167, gm_n11670, gm_n11671, gm_n11672, gm_n11673, gm_n11674, gm_n11675, gm_n11676, gm_n11677, gm_n11678, gm_n11679, gm_n1168, gm_n11680, gm_n11681, gm_n11682, gm_n11683, gm_n11684, gm_n11685, gm_n11686, gm_n11687, gm_n11688, gm_n11689, gm_n1169, gm_n11690, gm_n11691, gm_n11692, gm_n11693, gm_n11694, gm_n11695, gm_n11696, gm_n11697, gm_n11698, gm_n11699, gm_n117, gm_n1170, gm_n11700, gm_n11701, gm_n11702, gm_n11703, gm_n11704, gm_n11705, gm_n11706, gm_n11707, gm_n11708, gm_n11709, gm_n1171, gm_n11710, gm_n11711, gm_n11712, gm_n11713, gm_n11714, gm_n11715, gm_n11716, gm_n11717, gm_n11718, gm_n11719, gm_n1172, gm_n11720, gm_n11721, gm_n11722, gm_n11723, gm_n11724, gm_n11725, gm_n11726, gm_n11727, gm_n11728, gm_n11729, gm_n1173, gm_n11730, gm_n11731, gm_n11732, gm_n11733, gm_n11734, gm_n11735, gm_n11736, gm_n11737, gm_n11738, gm_n11739, gm_n1174, gm_n11740, gm_n11741, gm_n11742, gm_n11743, gm_n11744, gm_n11745, gm_n11746, gm_n11747, gm_n11748, gm_n11749, gm_n1175, gm_n11750, gm_n11751, gm_n11752, gm_n11753, gm_n11754, gm_n11755, gm_n11756, gm_n11757, gm_n11758, gm_n11759, gm_n1176, gm_n11760, gm_n11761, gm_n11762, gm_n11763, gm_n11764, gm_n11765, gm_n11766, gm_n11767, gm_n11768, gm_n11769, gm_n1177, gm_n11770, gm_n11771, gm_n11772, gm_n11773, gm_n11774, gm_n11775, gm_n11776, gm_n11777, gm_n11778, gm_n11779, gm_n1178, gm_n11780, gm_n11781, gm_n11782, gm_n11783, gm_n11784, gm_n11785, gm_n11786, gm_n11787, gm_n11788, gm_n11789, gm_n1179, gm_n11790, gm_n11791, gm_n11792, gm_n11793, gm_n11794, gm_n11795, gm_n11796, gm_n11797, gm_n11798, gm_n11799, gm_n118, gm_n1180, gm_n11800, gm_n11801, gm_n11802, gm_n11803, gm_n11804, gm_n11805, gm_n11806, gm_n11807, gm_n11808, gm_n11809, gm_n1181, gm_n11810, gm_n11811, gm_n11812, gm_n11813, gm_n11814, gm_n11815, gm_n11816, gm_n11817, gm_n11818, gm_n11819, gm_n1182, gm_n11820, gm_n11821, gm_n11822, gm_n11823, gm_n11824, gm_n11825, gm_n11826, gm_n11827, gm_n11828, gm_n11829, gm_n1183, gm_n11830, gm_n11831, gm_n11832, gm_n11833, gm_n11834, gm_n11835, gm_n11836, gm_n11837, gm_n11838, gm_n11839, gm_n1184, gm_n11840, gm_n11841, gm_n11842, gm_n11843, gm_n11844, gm_n11845, gm_n11846, gm_n11847, gm_n11848, gm_n11849, gm_n1185, gm_n11850, gm_n11851, gm_n11852, gm_n11853, gm_n11854, gm_n11855, gm_n11856, gm_n11857, gm_n11858, gm_n11859, gm_n1186, gm_n11860, gm_n11861, gm_n11862, gm_n11863, gm_n11864, gm_n11865, gm_n11866, gm_n11867, gm_n11868, gm_n11869, gm_n1187, gm_n11870, gm_n11871, gm_n11872, gm_n11873, gm_n11874, gm_n11875, gm_n11876, gm_n11877, gm_n11878, gm_n11879, gm_n1188, gm_n11880, gm_n11881, gm_n11882, gm_n11883, gm_n11884, gm_n11885, gm_n11886, gm_n11887, gm_n11888, gm_n11889, gm_n1189, gm_n11890, gm_n11891, gm_n11892, gm_n11893, gm_n11894, gm_n11895, gm_n11896, gm_n11897, gm_n11898, gm_n11899, gm_n119, gm_n1190, gm_n11900, gm_n11901, gm_n11902, gm_n11903, gm_n11904, gm_n11905, gm_n11906, gm_n11907, gm_n11908, gm_n11909, gm_n1191, gm_n11910, gm_n11911, gm_n11912, gm_n11913, gm_n11914, gm_n11915, gm_n11916, gm_n11917, gm_n11918, gm_n11919, gm_n1192, gm_n11920, gm_n11921, gm_n11922, gm_n11923, gm_n11924, gm_n11925, gm_n11926, gm_n11927, gm_n11928, gm_n11929, gm_n1193, gm_n11930, gm_n11931, gm_n11932, gm_n11933, gm_n11934, gm_n11935, gm_n11936, gm_n11937, gm_n11938, gm_n11939, gm_n1194, gm_n11940, gm_n11941, gm_n11942, gm_n11943, gm_n11944, gm_n11945, gm_n11946, gm_n11947, gm_n11948, gm_n11949, gm_n1195, gm_n11950, gm_n11951, gm_n11952, gm_n11953, gm_n11954, gm_n11955, gm_n11956, gm_n11957, gm_n11958, gm_n11959, gm_n1196, gm_n11960, gm_n11961, gm_n11962, gm_n11963, gm_n11964, gm_n11965, gm_n11966, gm_n11967, gm_n11968, gm_n11969, gm_n1197, gm_n11970, gm_n11971, gm_n11972, gm_n11973, gm_n11974, gm_n11975, gm_n11976, gm_n11977, gm_n11978, gm_n11979, gm_n1198, gm_n11980, gm_n11981, gm_n11982, gm_n11983, gm_n11984, gm_n11985, gm_n11986, gm_n11987, gm_n11988, gm_n11989, gm_n1199, gm_n11990, gm_n11991, gm_n11992, gm_n11993, gm_n11994, gm_n11995, gm_n11997, gm_n11998, gm_n11999, gm_n120, gm_n1200, gm_n12000, gm_n12001, gm_n12002, gm_n12003, gm_n12004, gm_n12005, gm_n12006, gm_n12007, gm_n12008, gm_n12009, gm_n1201, gm_n12010, gm_n12011, gm_n12012, gm_n12013, gm_n12014, gm_n12015, gm_n12016, gm_n12017, gm_n12018, gm_n12019, gm_n1202, gm_n12020, gm_n12021, gm_n12022, gm_n12023, gm_n12024, gm_n12025, gm_n12026, gm_n12027, gm_n12028, gm_n12029, gm_n1203, gm_n12030, gm_n12031, gm_n12032, gm_n12033, gm_n12034, gm_n12035, gm_n12036, gm_n12037, gm_n12038, gm_n12039, gm_n1204, gm_n12040, gm_n12041, gm_n12042, gm_n12043, gm_n12044, gm_n12045, gm_n12046, gm_n12047, gm_n12048, gm_n12049, gm_n1205, gm_n12050, gm_n12051, gm_n12052, gm_n12053, gm_n12054, gm_n12055, gm_n12056, gm_n12057, gm_n12058, gm_n12059, gm_n1206, gm_n12060, gm_n12061, gm_n12062, gm_n12063, gm_n12064, gm_n12065, gm_n12066, gm_n12067, gm_n12068, gm_n12069, gm_n1207, gm_n12070, gm_n12071, gm_n12072, gm_n12073, gm_n12074, gm_n12075, gm_n12076, gm_n12077, gm_n12078, gm_n12079, gm_n1208, gm_n12080, gm_n12081, gm_n12082, gm_n12083, gm_n12084, gm_n12085, gm_n12086, gm_n12087, gm_n12088, gm_n12089, gm_n1209, gm_n12090, gm_n12091, gm_n12092, gm_n12093, gm_n12094, gm_n12095, gm_n12096, gm_n12097, gm_n12098, gm_n12099, gm_n121, gm_n1210, gm_n12100, gm_n12101, gm_n12102, gm_n12103, gm_n12104, gm_n12105, gm_n12106, gm_n12107, gm_n12108, gm_n12109, gm_n1211, gm_n12110, gm_n12111, gm_n12112, gm_n12113, gm_n12114, gm_n12115, gm_n12116, gm_n12117, gm_n12118, gm_n12119, gm_n1212, gm_n12120, gm_n12121, gm_n12122, gm_n12123, gm_n12124, gm_n12125, gm_n12126, gm_n12127, gm_n12128, gm_n12129, gm_n1213, gm_n12130, gm_n12131, gm_n12132, gm_n12133, gm_n12134, gm_n12135, gm_n12136, gm_n12137, gm_n12138, gm_n12139, gm_n1214, gm_n12140, gm_n12141, gm_n12142, gm_n12143, gm_n12144, gm_n12145, gm_n12146, gm_n12147, gm_n12148, gm_n12149, gm_n1215, gm_n12150, gm_n12151, gm_n12152, gm_n12153, gm_n12154, gm_n12155, gm_n12156, gm_n12157, gm_n12158, gm_n12159, gm_n1216, gm_n12160, gm_n12161, gm_n12162, gm_n12163, gm_n12164, gm_n12165, gm_n12166, gm_n12167, gm_n12168, gm_n12169, gm_n1217, gm_n12170, gm_n12171, gm_n12172, gm_n12173, gm_n12174, gm_n12175, gm_n12176, gm_n12177, gm_n12178, gm_n12179, gm_n1218, gm_n12180, gm_n12181, gm_n12182, gm_n12183, gm_n12184, gm_n12185, gm_n12186, gm_n12187, gm_n12188, gm_n12189, gm_n1219, gm_n12190, gm_n12191, gm_n12192, gm_n12193, gm_n12194, gm_n12195, gm_n12196, gm_n12197, gm_n12198, gm_n12199, gm_n122, gm_n1220, gm_n12200, gm_n12201, gm_n12202, gm_n12203, gm_n12204, gm_n12205, gm_n12206, gm_n12207, gm_n12208, gm_n12209, gm_n1221, gm_n12210, gm_n12211, gm_n12212, gm_n12213, gm_n12214, gm_n12215, gm_n12216, gm_n12217, gm_n12218, gm_n12219, gm_n1222, gm_n12220, gm_n12221, gm_n12222, gm_n12223, gm_n12224, gm_n12225, gm_n12226, gm_n12227, gm_n12228, gm_n12229, gm_n1223, gm_n12230, gm_n12231, gm_n12232, gm_n12233, gm_n12234, gm_n12235, gm_n12236, gm_n12237, gm_n12238, gm_n12239, gm_n1224, gm_n12240, gm_n12241, gm_n12242, gm_n12243, gm_n12244, gm_n12245, gm_n12246, gm_n12247, gm_n12248, gm_n12249, gm_n1225, gm_n12250, gm_n12251, gm_n12252, gm_n12253, gm_n12254, gm_n12255, gm_n12256, gm_n12257, gm_n12258, gm_n12259, gm_n1226, gm_n12260, gm_n12261, gm_n12262, gm_n12263, gm_n12264, gm_n12265, gm_n12266, gm_n12267, gm_n12268, gm_n12269, gm_n1227, gm_n12270, gm_n12271, gm_n12272, gm_n12273, gm_n12274, gm_n12275, gm_n12276, gm_n12277, gm_n12278, gm_n12279, gm_n1228, gm_n12280, gm_n12281, gm_n12282, gm_n12283, gm_n12284, gm_n12285, gm_n12286, gm_n12287, gm_n12288, gm_n12289, gm_n1229, gm_n12290, gm_n12291, gm_n12292, gm_n12293, gm_n12294, gm_n12295, gm_n12296, gm_n12297, gm_n12298, gm_n12299, gm_n123, gm_n1230, gm_n12300, gm_n12301, gm_n12302, gm_n12303, gm_n12304, gm_n12305, gm_n12306, gm_n12307, gm_n12308, gm_n12309, gm_n1231, gm_n12310, gm_n12311, gm_n12312, gm_n12313, gm_n12314, gm_n12315, gm_n12316, gm_n12317, gm_n12318, gm_n12319, gm_n1232, gm_n12320, gm_n12321, gm_n12322, gm_n12323, gm_n12324, gm_n12325, gm_n12326, gm_n12327, gm_n12328, gm_n12329, gm_n1233, gm_n12330, gm_n12331, gm_n12332, gm_n12333, gm_n12334, gm_n12335, gm_n12336, gm_n12337, gm_n12338, gm_n12339, gm_n1234, gm_n12340, gm_n12341, gm_n12342, gm_n12343, gm_n12344, gm_n12345, gm_n12346, gm_n12347, gm_n12348, gm_n12349, gm_n1235, gm_n12350, gm_n12351, gm_n12352, gm_n12353, gm_n12354, gm_n12355, gm_n12356, gm_n12357, gm_n12358, gm_n12359, gm_n1236, gm_n12360, gm_n12361, gm_n12362, gm_n12363, gm_n12364, gm_n12365, gm_n12366, gm_n12367, gm_n12368, gm_n12369, gm_n1237, gm_n12370, gm_n12371, gm_n12372, gm_n12373, gm_n12374, gm_n12375, gm_n12376, gm_n12377, gm_n12378, gm_n12379, gm_n1238, gm_n12380, gm_n12381, gm_n12382, gm_n12383, gm_n12384, gm_n12385, gm_n12386, gm_n12387, gm_n12388, gm_n12389, gm_n1239, gm_n12390, gm_n12391, gm_n12392, gm_n12393, gm_n12394, gm_n12395, gm_n12396, gm_n12397, gm_n12398, gm_n12399, gm_n124, gm_n1240, gm_n12400, gm_n12401, gm_n12402, gm_n12403, gm_n12404, gm_n12405, gm_n12406, gm_n12407, gm_n12408, gm_n12409, gm_n1241, gm_n12410, gm_n12411, gm_n12412, gm_n12413, gm_n12414, gm_n12415, gm_n12416, gm_n12417, gm_n12418, gm_n12419, gm_n1242, gm_n12420, gm_n12421, gm_n12422, gm_n12423, gm_n12424, gm_n12425, gm_n12426, gm_n12427, gm_n12428, gm_n12429, gm_n1243, gm_n12430, gm_n12431, gm_n12432, gm_n12433, gm_n12434, gm_n12435, gm_n12436, gm_n12437, gm_n12438, gm_n12439, gm_n1244, gm_n12440, gm_n12441, gm_n12442, gm_n12443, gm_n12444, gm_n12445, gm_n12446, gm_n12447, gm_n12448, gm_n12449, gm_n1245, gm_n12450, gm_n12451, gm_n12452, gm_n12453, gm_n12454, gm_n12455, gm_n12456, gm_n12457, gm_n12458, gm_n12459, gm_n1246, gm_n12460, gm_n12461, gm_n12462, gm_n12463, gm_n12464, gm_n12465, gm_n12466, gm_n12467, gm_n12468, gm_n12469, gm_n1247, gm_n12470, gm_n12471, gm_n12472, gm_n12473, gm_n12474, gm_n12475, gm_n12476, gm_n12477, gm_n12478, gm_n12479, gm_n1248, gm_n12480, gm_n12481, gm_n1249, gm_n125, gm_n1250, gm_n1251, gm_n1252, gm_n1253, gm_n1254, gm_n1255, gm_n1256, gm_n1257, gm_n1258, gm_n1259, gm_n126, gm_n1260, gm_n1261, gm_n1262, gm_n1263, gm_n1264, gm_n1265, gm_n1266, gm_n1267, gm_n1268, gm_n1269, gm_n127, gm_n1270, gm_n1271, gm_n1272, gm_n1273, gm_n1274, gm_n1275, gm_n1276, gm_n1277, gm_n1278, gm_n1279, gm_n128, gm_n1280, gm_n1281, gm_n1282, gm_n1283, gm_n1284, gm_n1285, gm_n1286, gm_n1287, gm_n1288, gm_n1289, gm_n129, gm_n1290, gm_n1291, gm_n1292, gm_n1293, gm_n1294, gm_n1295, gm_n1296, gm_n1297, gm_n1298, gm_n1299, gm_n130, gm_n1300, gm_n1301, gm_n1302, gm_n1303, gm_n1304, gm_n1305, gm_n1306, gm_n1307, gm_n1308, gm_n1309, gm_n131, gm_n1310, gm_n1311, gm_n1312, gm_n1313, gm_n1314, gm_n1315, gm_n1316, gm_n1317, gm_n1318, gm_n1319, gm_n132, gm_n1320, gm_n1321, gm_n1322, gm_n1323, gm_n1324, gm_n1325, gm_n1326, gm_n1327, gm_n1328, gm_n1329, gm_n133, gm_n1330, gm_n1331, gm_n1332, gm_n1333, gm_n1334, gm_n1335, gm_n1336, gm_n1337, gm_n1338, gm_n1339, gm_n134, gm_n1340, gm_n1341, gm_n1342, gm_n1343, gm_n1344, gm_n1345, gm_n1346, gm_n1347, gm_n1348, gm_n1349, gm_n135, gm_n1350, gm_n1351, gm_n1352, gm_n1353, gm_n1354, gm_n1355, gm_n1356, gm_n1357, gm_n1358, gm_n1359, gm_n136, gm_n1360, gm_n1361, gm_n1362, gm_n1363, gm_n1364, gm_n1365, gm_n1366, gm_n1367, gm_n1368, gm_n1369, gm_n137, gm_n1370, gm_n1371, gm_n1372, gm_n1373, gm_n1374, gm_n1375, gm_n1376, gm_n1377, gm_n1378, gm_n1379, gm_n138, gm_n1380, gm_n1381, gm_n1382, gm_n1383, gm_n1384, gm_n1385, gm_n1386, gm_n1387, gm_n1388, gm_n1389, gm_n139, gm_n1390, gm_n1391, gm_n1392, gm_n1393, gm_n1394, gm_n1395, gm_n1396, gm_n1397, gm_n1398, gm_n1399, gm_n140, gm_n1400, gm_n1401, gm_n1402, gm_n1403, gm_n1404, gm_n1405, gm_n1406, gm_n1407, gm_n1408, gm_n1409, gm_n141, gm_n1410, gm_n1411, gm_n1412, gm_n1413, gm_n1414, gm_n1415, gm_n1416, gm_n1417, gm_n1418, gm_n1419, gm_n142, gm_n1420, gm_n1421, gm_n1422, gm_n1423, gm_n1424, gm_n1425, gm_n1426, gm_n1427, gm_n1428, gm_n1429, gm_n143, gm_n1430, gm_n1431, gm_n1432, gm_n1433, gm_n1434, gm_n1435, gm_n1436, gm_n1437, gm_n1438, gm_n1439, gm_n144, gm_n1440, gm_n1441, gm_n1442, gm_n1443, gm_n1444, gm_n1445, gm_n1446, gm_n1447, gm_n1448, gm_n1449, gm_n145, gm_n1450, gm_n1451, gm_n1452, gm_n1453, gm_n1454, gm_n1455, gm_n1456, gm_n1457, gm_n1458, gm_n1459, gm_n146, gm_n1460, gm_n1461, gm_n1462, gm_n1463, gm_n1464, gm_n1465, gm_n1466, gm_n1467, gm_n1468, gm_n1469, gm_n147, gm_n1470, gm_n1471, gm_n1472, gm_n1473, gm_n1474, gm_n1475, gm_n1476, gm_n1477, gm_n1478, gm_n1479, gm_n148, gm_n1480, gm_n1481, gm_n1482, gm_n1483, gm_n1484, gm_n1485, gm_n1486, gm_n1487, gm_n1488, gm_n1489, gm_n149, gm_n1490, gm_n1491, gm_n1492, gm_n1493, gm_n1494, gm_n1495, gm_n1496, gm_n1497, gm_n1498, gm_n1499, gm_n150, gm_n1500, gm_n1501, gm_n1502, gm_n1503, gm_n1504, gm_n1505, gm_n1506, gm_n1507, gm_n1508, gm_n1509, gm_n151, gm_n1510, gm_n1511, gm_n1512, gm_n1513, gm_n1514, gm_n1515, gm_n1516, gm_n1517, gm_n1518, gm_n1519, gm_n152, gm_n1520, gm_n1521, gm_n1522, gm_n1524, gm_n1525, gm_n1526, gm_n1527, gm_n1528, gm_n1529, gm_n153, gm_n1530, gm_n1531, gm_n1532, gm_n1533, gm_n1534, gm_n1535, gm_n1536, gm_n1537, gm_n1538, gm_n1539, gm_n154, gm_n1540, gm_n1541, gm_n1542, gm_n1543, gm_n1544, gm_n1545, gm_n1546, gm_n1547, gm_n1548, gm_n1549, gm_n155, gm_n1550, gm_n1551, gm_n1552, gm_n1553, gm_n1554, gm_n1555, gm_n1556, gm_n1557, gm_n1558, gm_n1559, gm_n156, gm_n1560, gm_n1561, gm_n1562, gm_n1563, gm_n1564, gm_n1565, gm_n1566, gm_n1567, gm_n1568, gm_n1569, gm_n157, gm_n1570, gm_n1571, gm_n1572, gm_n1573, gm_n1574, gm_n1575, gm_n1576, gm_n1577, gm_n1578, gm_n1579, gm_n158, gm_n1580, gm_n1581, gm_n1582, gm_n1583, gm_n1584, gm_n1585, gm_n1586, gm_n1587, gm_n1588, gm_n1589, gm_n159, gm_n1590, gm_n1591, gm_n1592, gm_n1593, gm_n1594, gm_n1595, gm_n1596, gm_n1597, gm_n1598, gm_n1599, gm_n160, gm_n1600, gm_n1601, gm_n1602, gm_n1603, gm_n1604, gm_n1605, gm_n1606, gm_n1607, gm_n1608, gm_n1609, gm_n161, gm_n1610, gm_n1611, gm_n1612, gm_n1613, gm_n1614, gm_n1615, gm_n1616, gm_n1617, gm_n1618, gm_n1619, gm_n162, gm_n1620, gm_n1621, gm_n1622, gm_n1623, gm_n1624, gm_n1625, gm_n1626, gm_n1627, gm_n1628, gm_n1629, gm_n163, gm_n1630, gm_n1631, gm_n1632, gm_n1633, gm_n1634, gm_n1635, gm_n1636, gm_n1637, gm_n1638, gm_n1639, gm_n164, gm_n1640, gm_n1641, gm_n1642, gm_n1643, gm_n1644, gm_n1645, gm_n1646, gm_n1647, gm_n1648, gm_n1649, gm_n165, gm_n1650, gm_n1651, gm_n1652, gm_n1653, gm_n1654, gm_n1655, gm_n1656, gm_n1657, gm_n1658, gm_n1659, gm_n166, gm_n1660, gm_n1661, gm_n1662, gm_n1663, gm_n1664, gm_n1665, gm_n1666, gm_n1667, gm_n1668, gm_n1669, gm_n167, gm_n1670, gm_n1671, gm_n1672, gm_n1673, gm_n1674, gm_n1675, gm_n1676, gm_n1677, gm_n1678, gm_n1679, gm_n168, gm_n1680, gm_n1681, gm_n1682, gm_n1683, gm_n1684, gm_n1685, gm_n1686, gm_n1687, gm_n1688, gm_n1689, gm_n169, gm_n1690, gm_n1691, gm_n1692, gm_n1693, gm_n1694, gm_n1695, gm_n1696, gm_n1697, gm_n1698, gm_n1699, gm_n170, gm_n1700, gm_n1701, gm_n1702, gm_n1703, gm_n1704, gm_n1705, gm_n1706, gm_n1707, gm_n1708, gm_n1709, gm_n171, gm_n1710, gm_n1711, gm_n1712, gm_n1713, gm_n1714, gm_n1715, gm_n1716, gm_n1717, gm_n1718, gm_n1719, gm_n172, gm_n1720, gm_n1721, gm_n1722, gm_n1723, gm_n1724, gm_n1725, gm_n1726, gm_n1727, gm_n1728, gm_n1729, gm_n173, gm_n1730, gm_n1731, gm_n1732, gm_n1733, gm_n1734, gm_n1735, gm_n1736, gm_n1737, gm_n1738, gm_n1739, gm_n174, gm_n1740, gm_n1741, gm_n1742, gm_n1743, gm_n1744, gm_n1745, gm_n1746, gm_n1747, gm_n1748, gm_n1749, gm_n175, gm_n1750, gm_n1751, gm_n1752, gm_n1753, gm_n1754, gm_n1755, gm_n1756, gm_n1757, gm_n1758, gm_n1759, gm_n176, gm_n1760, gm_n1761, gm_n1762, gm_n1763, gm_n1764, gm_n1765, gm_n1766, gm_n1767, gm_n1768, gm_n1769, gm_n177, gm_n1770, gm_n1771, gm_n1772, gm_n1773, gm_n1774, gm_n1775, gm_n1776, gm_n1777, gm_n1778, gm_n1779, gm_n178, gm_n1780, gm_n1781, gm_n1782, gm_n1783, gm_n1784, gm_n1785, gm_n1786, gm_n1787, gm_n1788, gm_n1789, gm_n179, gm_n1790, gm_n1791, gm_n1792, gm_n1793, gm_n1794, gm_n1795, gm_n1796, gm_n1797, gm_n1798, gm_n1799, gm_n180, gm_n1800, gm_n1801, gm_n1802, gm_n1803, gm_n1804, gm_n1805, gm_n1806, gm_n1807, gm_n1808, gm_n1809, gm_n181, gm_n1810, gm_n1811, gm_n1812, gm_n1813, gm_n1814, gm_n1815, gm_n1816, gm_n1817, gm_n1818, gm_n1819, gm_n182, gm_n1820, gm_n1821, gm_n1822, gm_n1823, gm_n1824, gm_n1825, gm_n1826, gm_n1827, gm_n1828, gm_n1829, gm_n183, gm_n1830, gm_n1831, gm_n1832, gm_n1833, gm_n1834, gm_n1835, gm_n1836, gm_n1837, gm_n1838, gm_n1839, gm_n184, gm_n1840, gm_n1841, gm_n1842, gm_n1843, gm_n1844, gm_n1845, gm_n1846, gm_n1847, gm_n1848, gm_n1849, gm_n185, gm_n1850, gm_n1851, gm_n1852, gm_n1853, gm_n1854, gm_n1855, gm_n1856, gm_n1857, gm_n1858, gm_n1859, gm_n186, gm_n1860, gm_n1861, gm_n1862, gm_n1863, gm_n1864, gm_n1865, gm_n1866, gm_n1867, gm_n1868, gm_n1869, gm_n187, gm_n1870, gm_n1871, gm_n1872, gm_n1873, gm_n1874, gm_n1875, gm_n1876, gm_n1877, gm_n1878, gm_n1879, gm_n188, gm_n1880, gm_n1881, gm_n1882, gm_n1883, gm_n1884, gm_n1885, gm_n1886, gm_n1887, gm_n1888, gm_n1889, gm_n189, gm_n1890, gm_n1891, gm_n1892, gm_n1893, gm_n1894, gm_n1895, gm_n1896, gm_n1897, gm_n1898, gm_n1899, gm_n190, gm_n1900, gm_n1901, gm_n1902, gm_n1903, gm_n1904, gm_n1905, gm_n1906, gm_n1907, gm_n1908, gm_n1909, gm_n191, gm_n1910, gm_n1911, gm_n1912, gm_n1913, gm_n1914, gm_n1915, gm_n1916, gm_n1917, gm_n1918, gm_n1919, gm_n192, gm_n1920, gm_n1921, gm_n1922, gm_n1923, gm_n1924, gm_n1925, gm_n1926, gm_n1927, gm_n1928, gm_n1929, gm_n193, gm_n1930, gm_n1931, gm_n1932, gm_n1933, gm_n1934, gm_n1935, gm_n1936, gm_n1937, gm_n1938, gm_n1939, gm_n194, gm_n1940, gm_n1941, gm_n1942, gm_n1943, gm_n1944, gm_n1945, gm_n1946, gm_n1947, gm_n1948, gm_n1949, gm_n195, gm_n1950, gm_n1951, gm_n1952, gm_n1953, gm_n1954, gm_n1955, gm_n1956, gm_n1957, gm_n1958, gm_n1959, gm_n196, gm_n1960, gm_n1961, gm_n1962, gm_n1963, gm_n1964, gm_n1965, gm_n1966, gm_n1967, gm_n1968, gm_n1969, gm_n197, gm_n1970, gm_n1971, gm_n1972, gm_n1973, gm_n1974, gm_n1975, gm_n1976, gm_n1977, gm_n1978, gm_n1979, gm_n198, gm_n1980, gm_n1981, gm_n1982, gm_n1983, gm_n1984, gm_n1985, gm_n1986, gm_n1987, gm_n1988, gm_n1989, gm_n199, gm_n1990, gm_n1991, gm_n1992, gm_n1993, gm_n1994, gm_n1995, gm_n1996, gm_n1997, gm_n1998, gm_n1999, gm_n200, gm_n2000, gm_n2001, gm_n2002, gm_n2003, gm_n2004, gm_n2005, gm_n2006, gm_n2007, gm_n2008, gm_n2009, gm_n201, gm_n2010, gm_n2011, gm_n2012, gm_n2013, gm_n2014, gm_n2015, gm_n2016, gm_n2017, gm_n2018, gm_n2019, gm_n202, gm_n2020, gm_n2021, gm_n2022, gm_n2023, gm_n2024, gm_n2025, gm_n2026, gm_n2027, gm_n2028, gm_n2029, gm_n203, gm_n2030, gm_n2031, gm_n2032, gm_n2033, gm_n2034, gm_n2035, gm_n2036, gm_n2037, gm_n2038, gm_n2039, gm_n204, gm_n2040, gm_n2041, gm_n2042, gm_n2043, gm_n2044, gm_n2045, gm_n2046, gm_n2047, gm_n2048, gm_n2049, gm_n205, gm_n2050, gm_n2051, gm_n2052, gm_n2053, gm_n2054, gm_n2055, gm_n2056, gm_n2057, gm_n2058, gm_n2059, gm_n206, gm_n2060, gm_n2061, gm_n2062, gm_n2063, gm_n2064, gm_n2065, gm_n2066, gm_n2067, gm_n2068, gm_n2069, gm_n207, gm_n2070, gm_n2071, gm_n2072, gm_n2073, gm_n2074, gm_n2075, gm_n2076, gm_n2077, gm_n2078, gm_n2079, gm_n208, gm_n2080, gm_n2081, gm_n2082, gm_n2083, gm_n2084, gm_n2085, gm_n2086, gm_n2087, gm_n2088, gm_n2089, gm_n209, gm_n2090, gm_n2091, gm_n2092, gm_n2093, gm_n2094, gm_n2095, gm_n2096, gm_n2097, gm_n2098, gm_n2099, gm_n210, gm_n2100, gm_n2101, gm_n2102, gm_n2103, gm_n2104, gm_n2105, gm_n2106, gm_n2107, gm_n2108, gm_n2109, gm_n211, gm_n2110, gm_n2111, gm_n2112, gm_n2113, gm_n2114, gm_n2115, gm_n2116, gm_n2117, gm_n2118, gm_n2119, gm_n212, gm_n2120, gm_n2121, gm_n2122, gm_n2123, gm_n2124, gm_n2125, gm_n2126, gm_n2127, gm_n2128, gm_n2129, gm_n213, gm_n2130, gm_n2131, gm_n2132, gm_n2133, gm_n2134, gm_n2135, gm_n2136, gm_n2137, gm_n2138, gm_n2139, gm_n214, gm_n2140, gm_n2141, gm_n2142, gm_n2143, gm_n2144, gm_n2145, gm_n2146, gm_n2147, gm_n2148, gm_n2149, gm_n215, gm_n2150, gm_n2151, gm_n2152, gm_n2153, gm_n2154, gm_n2155, gm_n2156, gm_n2157, gm_n2158, gm_n2159, gm_n216, gm_n2160, gm_n2161, gm_n2162, gm_n2163, gm_n2164, gm_n2165, gm_n2166, gm_n2167, gm_n2168, gm_n2169, gm_n217, gm_n2170, gm_n2172, gm_n2173, gm_n2174, gm_n2175, gm_n2176, gm_n2177, gm_n2178, gm_n2179, gm_n218, gm_n2180, gm_n2181, gm_n2182, gm_n2183, gm_n2184, gm_n2185, gm_n2186, gm_n2187, gm_n2188, gm_n2189, gm_n219, gm_n2190, gm_n2191, gm_n2192, gm_n2193, gm_n2194, gm_n2195, gm_n2196, gm_n2197, gm_n2198, gm_n2199, gm_n220, gm_n2200, gm_n2201, gm_n2202, gm_n2203, gm_n2204, gm_n2205, gm_n2206, gm_n2207, gm_n2208, gm_n2209, gm_n221, gm_n2210, gm_n2211, gm_n2212, gm_n2213, gm_n2214, gm_n2215, gm_n2216, gm_n2217, gm_n2218, gm_n2219, gm_n222, gm_n2220, gm_n2221, gm_n2222, gm_n2223, gm_n2224, gm_n2225, gm_n2226, gm_n2227, gm_n2228, gm_n2229, gm_n223, gm_n2230, gm_n2231, gm_n2232, gm_n2233, gm_n2234, gm_n2235, gm_n2236, gm_n2237, gm_n2238, gm_n2239, gm_n224, gm_n2240, gm_n2241, gm_n2242, gm_n2243, gm_n2244, gm_n2245, gm_n2246, gm_n2247, gm_n2248, gm_n2249, gm_n225, gm_n2250, gm_n2251, gm_n2252, gm_n2253, gm_n2254, gm_n2255, gm_n2256, gm_n2257, gm_n2258, gm_n2259, gm_n226, gm_n2260, gm_n2261, gm_n2262, gm_n2263, gm_n2264, gm_n2265, gm_n2266, gm_n2267, gm_n2268, gm_n2269, gm_n227, gm_n2270, gm_n2271, gm_n2272, gm_n2273, gm_n2274, gm_n2275, gm_n2276, gm_n2277, gm_n2278, gm_n2279, gm_n228, gm_n2280, gm_n2281, gm_n2282, gm_n2283, gm_n2284, gm_n2285, gm_n2286, gm_n2287, gm_n2288, gm_n2289, gm_n229, gm_n2290, gm_n2291, gm_n2292, gm_n2293, gm_n2294, gm_n2295, gm_n2296, gm_n2297, gm_n2298, gm_n2299, gm_n230, gm_n2300, gm_n2301, gm_n2302, gm_n2303, gm_n2304, gm_n2305, gm_n2306, gm_n2307, gm_n2308, gm_n2309, gm_n231, gm_n2310, gm_n2311, gm_n2312, gm_n2313, gm_n2314, gm_n2315, gm_n2316, gm_n2317, gm_n2318, gm_n2319, gm_n232, gm_n2320, gm_n2321, gm_n2322, gm_n2323, gm_n2324, gm_n2325, gm_n2326, gm_n2327, gm_n2328, gm_n2329, gm_n233, gm_n2330, gm_n2331, gm_n2332, gm_n2333, gm_n2334, gm_n2335, gm_n2336, gm_n2337, gm_n2338, gm_n2339, gm_n234, gm_n2340, gm_n2341, gm_n2342, gm_n2343, gm_n2344, gm_n2345, gm_n2346, gm_n2347, gm_n2348, gm_n2349, gm_n235, gm_n2350, gm_n2351, gm_n2352, gm_n2353, gm_n2354, gm_n2355, gm_n2356, gm_n2357, gm_n2358, gm_n2359, gm_n236, gm_n2360, gm_n2361, gm_n2362, gm_n2363, gm_n2364, gm_n2365, gm_n2366, gm_n2367, gm_n2368, gm_n2369, gm_n237, gm_n2370, gm_n2371, gm_n2372, gm_n2373, gm_n2374, gm_n2375, gm_n2376, gm_n2377, gm_n2378, gm_n2379, gm_n238, gm_n2380, gm_n2381, gm_n2382, gm_n2383, gm_n2384, gm_n2385, gm_n2386, gm_n2387, gm_n2388, gm_n2389, gm_n239, gm_n2390, gm_n2391, gm_n2392, gm_n2393, gm_n2394, gm_n2395, gm_n2396, gm_n2397, gm_n2398, gm_n2399, gm_n240, gm_n2400, gm_n2401, gm_n2402, gm_n2403, gm_n2404, gm_n2405, gm_n2406, gm_n2407, gm_n2408, gm_n2409, gm_n241, gm_n2410, gm_n2411, gm_n2412, gm_n2413, gm_n2414, gm_n2415, gm_n2416, gm_n2417, gm_n2418, gm_n2419, gm_n242, gm_n2420, gm_n2421, gm_n2422, gm_n2423, gm_n2424, gm_n2425, gm_n2426, gm_n2427, gm_n2428, gm_n2429, gm_n243, gm_n2430, gm_n2431, gm_n2432, gm_n2433, gm_n2434, gm_n2435, gm_n2436, gm_n2437, gm_n2438, gm_n2439, gm_n244, gm_n2440, gm_n2441, gm_n2442, gm_n2443, gm_n2444, gm_n2445, gm_n2446, gm_n2447, gm_n2448, gm_n2449, gm_n245, gm_n2450, gm_n2451, gm_n2452, gm_n2453, gm_n2454, gm_n2455, gm_n2456, gm_n2457, gm_n2458, gm_n2459, gm_n246, gm_n2460, gm_n2461, gm_n2462, gm_n2463, gm_n2464, gm_n2465, gm_n2466, gm_n2467, gm_n2468, gm_n2469, gm_n247, gm_n2470, gm_n2471, gm_n2472, gm_n2473, gm_n2474, gm_n2475, gm_n2476, gm_n2477, gm_n2478, gm_n2479, gm_n248, gm_n2480, gm_n2481, gm_n2482, gm_n2483, gm_n2484, gm_n2485, gm_n2486, gm_n2487, gm_n2488, gm_n2489, gm_n249, gm_n2490, gm_n2491, gm_n2492, gm_n2493, gm_n2494, gm_n2495, gm_n2496, gm_n2497, gm_n2498, gm_n2499, gm_n250, gm_n2500, gm_n2501, gm_n2502, gm_n2503, gm_n2504, gm_n2505, gm_n2506, gm_n2507, gm_n2508, gm_n2509, gm_n251, gm_n2510, gm_n2511, gm_n2512, gm_n2513, gm_n2514, gm_n2515, gm_n2516, gm_n2517, gm_n2518, gm_n2519, gm_n252, gm_n2520, gm_n2521, gm_n2522, gm_n2523, gm_n2524, gm_n2525, gm_n2526, gm_n2527, gm_n2528, gm_n2529, gm_n253, gm_n2530, gm_n2531, gm_n2532, gm_n2533, gm_n2534, gm_n2535, gm_n2536, gm_n2537, gm_n2538, gm_n2539, gm_n254, gm_n2540, gm_n2541, gm_n2542, gm_n2543, gm_n2544, gm_n2545, gm_n2546, gm_n2547, gm_n2548, gm_n2549, gm_n255, gm_n2550, gm_n2551, gm_n2552, gm_n2553, gm_n2554, gm_n2555, gm_n2556, gm_n2557, gm_n2558, gm_n2559, gm_n256, gm_n2560, gm_n2561, gm_n2562, gm_n2563, gm_n2564, gm_n2565, gm_n2566, gm_n2567, gm_n2568, gm_n2569, gm_n257, gm_n2570, gm_n2571, gm_n2572, gm_n2573, gm_n2574, gm_n2575, gm_n2576, gm_n2577, gm_n2578, gm_n2579, gm_n258, gm_n2580, gm_n2581, gm_n2582, gm_n2583, gm_n2584, gm_n2585, gm_n2586, gm_n2587, gm_n2588, gm_n2589, gm_n259, gm_n2590, gm_n2591, gm_n2592, gm_n2593, gm_n2594, gm_n2595, gm_n2596, gm_n2597, gm_n2598, gm_n2599, gm_n260, gm_n2600, gm_n2601, gm_n2602, gm_n2603, gm_n2604, gm_n2605, gm_n2606, gm_n2607, gm_n2608, gm_n2609, gm_n261, gm_n2610, gm_n2611, gm_n2612, gm_n2613, gm_n2614, gm_n2615, gm_n2616, gm_n2617, gm_n2618, gm_n2619, gm_n262, gm_n2620, gm_n2621, gm_n2622, gm_n2623, gm_n2624, gm_n2625, gm_n2626, gm_n2627, gm_n2628, gm_n2629, gm_n263, gm_n2630, gm_n2631, gm_n2632, gm_n2633, gm_n2634, gm_n2635, gm_n2636, gm_n2637, gm_n2638, gm_n2639, gm_n264, gm_n2640, gm_n2641, gm_n2642, gm_n2643, gm_n2644, gm_n2645, gm_n2646, gm_n2647, gm_n2648, gm_n2649, gm_n265, gm_n2650, gm_n2651, gm_n2652, gm_n2653, gm_n2654, gm_n2655, gm_n2656, gm_n2657, gm_n2658, gm_n2659, gm_n266, gm_n2660, gm_n2661, gm_n2662, gm_n2663, gm_n2664, gm_n2665, gm_n2666, gm_n2667, gm_n2668, gm_n2669, gm_n267, gm_n2670, gm_n2671, gm_n2672, gm_n2673, gm_n2674, gm_n2675, gm_n2676, gm_n2677, gm_n2678, gm_n2679, gm_n268, gm_n2680, gm_n2681, gm_n2682, gm_n2683, gm_n2684, gm_n2685, gm_n2686, gm_n2687, gm_n2688, gm_n2689, gm_n269, gm_n2690, gm_n2691, gm_n2692, gm_n2693, gm_n2694, gm_n2695, gm_n2696, gm_n2697, gm_n2698, gm_n2699, gm_n270, gm_n2700, gm_n2701, gm_n2702, gm_n2703, gm_n2704, gm_n2705, gm_n2706, gm_n2707, gm_n2708, gm_n2709, gm_n271, gm_n2710, gm_n2711, gm_n2712, gm_n2713, gm_n2714, gm_n2715, gm_n2716, gm_n2717, gm_n2718, gm_n2719, gm_n272, gm_n2720, gm_n2721, gm_n2722, gm_n2723, gm_n2724, gm_n2725, gm_n2726, gm_n2727, gm_n2728, gm_n2729, gm_n273, gm_n2730, gm_n2731, gm_n2732, gm_n2733, gm_n2734, gm_n2735, gm_n2736, gm_n2737, gm_n2738, gm_n2739, gm_n274, gm_n2740, gm_n2741, gm_n2742, gm_n2743, gm_n2744, gm_n2745, gm_n2746, gm_n2747, gm_n2748, gm_n2749, gm_n275, gm_n2750, gm_n2751, gm_n2752, gm_n2753, gm_n2754, gm_n2755, gm_n2756, gm_n2757, gm_n2758, gm_n2759, gm_n276, gm_n2760, gm_n2761, gm_n2762, gm_n2763, gm_n2764, gm_n2765, gm_n2766, gm_n2767, gm_n2768, gm_n2769, gm_n277, gm_n2770, gm_n2771, gm_n2772, gm_n2773, gm_n2774, gm_n2775, gm_n2776, gm_n2777, gm_n2778, gm_n2779, gm_n278, gm_n2780, gm_n2781, gm_n2782, gm_n2783, gm_n2784, gm_n2785, gm_n2786, gm_n2787, gm_n2788, gm_n2789, gm_n279, gm_n2790, gm_n2791, gm_n2792, gm_n2793, gm_n2794, gm_n2795, gm_n2796, gm_n2797, gm_n2798, gm_n2799, gm_n280, gm_n2800, gm_n2802, gm_n2803, gm_n2804, gm_n2805, gm_n2806, gm_n2807, gm_n2808, gm_n2809, gm_n281, gm_n2810, gm_n2811, gm_n2812, gm_n2813, gm_n2814, gm_n2815, gm_n2816, gm_n2817, gm_n2818, gm_n2819, gm_n282, gm_n2820, gm_n2821, gm_n2822, gm_n2823, gm_n2824, gm_n2825, gm_n2826, gm_n2827, gm_n2828, gm_n2829, gm_n283, gm_n2830, gm_n2831, gm_n2832, gm_n2833, gm_n2834, gm_n2835, gm_n2836, gm_n2837, gm_n2838, gm_n2839, gm_n284, gm_n2840, gm_n2841, gm_n2842, gm_n2843, gm_n2844, gm_n2845, gm_n2846, gm_n2847, gm_n2848, gm_n2849, gm_n285, gm_n2850, gm_n2851, gm_n2852, gm_n2853, gm_n2854, gm_n2855, gm_n2856, gm_n2857, gm_n2858, gm_n2859, gm_n286, gm_n2860, gm_n2861, gm_n2862, gm_n2863, gm_n2864, gm_n2865, gm_n2866, gm_n2867, gm_n2868, gm_n2869, gm_n287, gm_n2870, gm_n2871, gm_n2872, gm_n2873, gm_n2874, gm_n2875, gm_n2876, gm_n2877, gm_n2878, gm_n2879, gm_n288, gm_n2880, gm_n2881, gm_n2882, gm_n2883, gm_n2884, gm_n2885, gm_n2886, gm_n2887, gm_n2888, gm_n2889, gm_n289, gm_n2890, gm_n2891, gm_n2892, gm_n2893, gm_n2894, gm_n2895, gm_n2896, gm_n2897, gm_n2898, gm_n2899, gm_n290, gm_n2900, gm_n2901, gm_n2902, gm_n2903, gm_n2904, gm_n2905, gm_n2906, gm_n2907, gm_n2908, gm_n2909, gm_n291, gm_n2910, gm_n2911, gm_n2912, gm_n2913, gm_n2914, gm_n2915, gm_n2916, gm_n2917, gm_n2918, gm_n2919, gm_n292, gm_n2920, gm_n2921, gm_n2922, gm_n2923, gm_n2924, gm_n2925, gm_n2926, gm_n2927, gm_n2928, gm_n2929, gm_n293, gm_n2930, gm_n2931, gm_n2932, gm_n2933, gm_n2934, gm_n2935, gm_n2936, gm_n2937, gm_n2938, gm_n2939, gm_n294, gm_n2940, gm_n2941, gm_n2942, gm_n2943, gm_n2944, gm_n2945, gm_n2946, gm_n2947, gm_n2948, gm_n2949, gm_n295, gm_n2950, gm_n2951, gm_n2952, gm_n2953, gm_n2954, gm_n2955, gm_n2956, gm_n2957, gm_n2958, gm_n2959, gm_n296, gm_n2960, gm_n2961, gm_n2962, gm_n2963, gm_n2964, gm_n2965, gm_n2966, gm_n2967, gm_n2968, gm_n2969, gm_n297, gm_n2970, gm_n2971, gm_n2972, gm_n2973, gm_n2974, gm_n2975, gm_n2976, gm_n2977, gm_n2978, gm_n2979, gm_n298, gm_n2980, gm_n2981, gm_n2982, gm_n2983, gm_n2984, gm_n2985, gm_n2986, gm_n2987, gm_n2988, gm_n2989, gm_n299, gm_n2990, gm_n2991, gm_n2992, gm_n2993, gm_n2994, gm_n2995, gm_n2996, gm_n2997, gm_n2998, gm_n2999, gm_n300, gm_n3000, gm_n3001, gm_n3002, gm_n3003, gm_n3004, gm_n3005, gm_n3006, gm_n3007, gm_n3008, gm_n3009, gm_n301, gm_n3010, gm_n3011, gm_n3012, gm_n3013, gm_n3014, gm_n3015, gm_n3016, gm_n3017, gm_n3018, gm_n3019, gm_n302, gm_n3020, gm_n3021, gm_n3022, gm_n3023, gm_n3024, gm_n3025, gm_n3026, gm_n3027, gm_n3028, gm_n3029, gm_n303, gm_n3030, gm_n3031, gm_n3032, gm_n3033, gm_n3034, gm_n3035, gm_n3036, gm_n3037, gm_n3038, gm_n3039, gm_n304, gm_n3040, gm_n3041, gm_n3042, gm_n3043, gm_n3044, gm_n3045, gm_n3046, gm_n3047, gm_n3048, gm_n3049, gm_n305, gm_n3050, gm_n3051, gm_n3052, gm_n3053, gm_n3054, gm_n3055, gm_n3056, gm_n3057, gm_n3058, gm_n3059, gm_n306, gm_n3060, gm_n3061, gm_n3062, gm_n3063, gm_n3064, gm_n3065, gm_n3066, gm_n3067, gm_n3068, gm_n3069, gm_n307, gm_n3070, gm_n3071, gm_n3072, gm_n3073, gm_n3074, gm_n3075, gm_n3076, gm_n3077, gm_n3078, gm_n3079, gm_n308, gm_n3080, gm_n3081, gm_n3082, gm_n3083, gm_n3084, gm_n3085, gm_n3086, gm_n3087, gm_n3088, gm_n3089, gm_n309, gm_n3090, gm_n3091, gm_n3092, gm_n3093, gm_n3094, gm_n3095, gm_n3096, gm_n3097, gm_n3098, gm_n3099, gm_n310, gm_n3100, gm_n3101, gm_n3102, gm_n3103, gm_n3104, gm_n3105, gm_n3106, gm_n3107, gm_n3108, gm_n3109, gm_n311, gm_n3110, gm_n3111, gm_n3112, gm_n3113, gm_n3114, gm_n3115, gm_n3116, gm_n3117, gm_n3118, gm_n3119, gm_n312, gm_n3120, gm_n3121, gm_n3122, gm_n3123, gm_n3124, gm_n3125, gm_n3126, gm_n3127, gm_n3128, gm_n3129, gm_n313, gm_n3130, gm_n3131, gm_n3132, gm_n3133, gm_n3134, gm_n3135, gm_n3136, gm_n3137, gm_n3138, gm_n3139, gm_n314, gm_n3140, gm_n3141, gm_n3142, gm_n3143, gm_n3144, gm_n3145, gm_n3146, gm_n3147, gm_n3148, gm_n3149, gm_n315, gm_n3150, gm_n3151, gm_n3152, gm_n3153, gm_n3154, gm_n3155, gm_n3156, gm_n3157, gm_n3158, gm_n3159, gm_n316, gm_n3160, gm_n3161, gm_n3162, gm_n3163, gm_n3164, gm_n3165, gm_n3166, gm_n3167, gm_n3168, gm_n3169, gm_n317, gm_n3170, gm_n3171, gm_n3172, gm_n3173, gm_n3174, gm_n3175, gm_n3176, gm_n3177, gm_n3178, gm_n3179, gm_n318, gm_n3180, gm_n3181, gm_n3182, gm_n3183, gm_n3184, gm_n3185, gm_n3186, gm_n3187, gm_n3188, gm_n3189, gm_n319, gm_n3190, gm_n3191, gm_n3192, gm_n3193, gm_n3194, gm_n3195, gm_n3196, gm_n3197, gm_n3198, gm_n3199, gm_n320, gm_n3200, gm_n3201, gm_n3202, gm_n3203, gm_n3204, gm_n3205, gm_n3206, gm_n3207, gm_n3208, gm_n3209, gm_n321, gm_n3210, gm_n3211, gm_n3212, gm_n3213, gm_n3214, gm_n3215, gm_n3216, gm_n3217, gm_n3218, gm_n3219, gm_n322, gm_n3220, gm_n3221, gm_n3222, gm_n3223, gm_n3224, gm_n3225, gm_n3226, gm_n3227, gm_n3228, gm_n3229, gm_n323, gm_n3230, gm_n3231, gm_n3232, gm_n3233, gm_n3234, gm_n3235, gm_n3236, gm_n3237, gm_n3238, gm_n3239, gm_n324, gm_n3240, gm_n3241, gm_n3242, gm_n3243, gm_n3244, gm_n3245, gm_n3246, gm_n3247, gm_n3248, gm_n3249, gm_n325, gm_n3250, gm_n3251, gm_n3252, gm_n3253, gm_n3254, gm_n3255, gm_n3256, gm_n3257, gm_n3258, gm_n3259, gm_n326, gm_n3260, gm_n3261, gm_n3262, gm_n3263, gm_n3264, gm_n3265, gm_n3266, gm_n3267, gm_n3268, gm_n3269, gm_n327, gm_n3270, gm_n3271, gm_n3272, gm_n3273, gm_n3274, gm_n3275, gm_n3276, gm_n3277, gm_n3278, gm_n3279, gm_n328, gm_n3280, gm_n3281, gm_n3282, gm_n3283, gm_n3284, gm_n3285, gm_n3286, gm_n3287, gm_n3288, gm_n3289, gm_n329, gm_n3290, gm_n3291, gm_n3292, gm_n3293, gm_n3294, gm_n3295, gm_n3296, gm_n3297, gm_n3298, gm_n3299, gm_n330, gm_n3300, gm_n3301, gm_n3302, gm_n3303, gm_n3304, gm_n3305, gm_n3306, gm_n3307, gm_n3308, gm_n3309, gm_n331, gm_n3310, gm_n3311, gm_n3312, gm_n3313, gm_n3314, gm_n3315, gm_n3316, gm_n3317, gm_n3318, gm_n3319, gm_n332, gm_n3320, gm_n3321, gm_n3322, gm_n3323, gm_n3324, gm_n3325, gm_n3326, gm_n3327, gm_n3328, gm_n3329, gm_n333, gm_n3330, gm_n3331, gm_n3332, gm_n3333, gm_n3334, gm_n3335, gm_n3336, gm_n3337, gm_n3338, gm_n3339, gm_n334, gm_n3340, gm_n3341, gm_n3342, gm_n3343, gm_n3344, gm_n3345, gm_n3346, gm_n3347, gm_n3348, gm_n3349, gm_n335, gm_n3350, gm_n3351, gm_n3352, gm_n3353, gm_n3354, gm_n3355, gm_n3356, gm_n3357, gm_n3358, gm_n3359, gm_n336, gm_n3360, gm_n3361, gm_n3362, gm_n3363, gm_n3364, gm_n3365, gm_n3366, gm_n3367, gm_n3368, gm_n3369, gm_n337, gm_n3370, gm_n3371, gm_n3372, gm_n3373, gm_n3374, gm_n3375, gm_n3376, gm_n3377, gm_n3378, gm_n3379, gm_n338, gm_n3380, gm_n3381, gm_n3382, gm_n3383, gm_n3384, gm_n3385, gm_n3386, gm_n3387, gm_n3388, gm_n3389, gm_n339, gm_n3390, gm_n3391, gm_n3392, gm_n3393, gm_n3394, gm_n3395, gm_n3396, gm_n3397, gm_n3398, gm_n3399, gm_n340, gm_n3400, gm_n3401, gm_n3402, gm_n3403, gm_n3404, gm_n3405, gm_n3406, gm_n3407, gm_n3408, gm_n3409, gm_n341, gm_n3410, gm_n3411, gm_n3413, gm_n3414, gm_n3415, gm_n3416, gm_n3417, gm_n3418, gm_n3419, gm_n342, gm_n3420, gm_n3421, gm_n3422, gm_n3423, gm_n3424, gm_n3425, gm_n3426, gm_n3427, gm_n3428, gm_n3429, gm_n343, gm_n3430, gm_n3431, gm_n3432, gm_n3433, gm_n3434, gm_n3435, gm_n3436, gm_n3437, gm_n3438, gm_n3439, gm_n344, gm_n3440, gm_n3441, gm_n3442, gm_n3443, gm_n3444, gm_n3445, gm_n3446, gm_n3447, gm_n3448, gm_n3449, gm_n345, gm_n3450, gm_n3451, gm_n3452, gm_n3453, gm_n3454, gm_n3455, gm_n3456, gm_n3457, gm_n3458, gm_n3459, gm_n346, gm_n3460, gm_n3461, gm_n3462, gm_n3463, gm_n3464, gm_n3465, gm_n3466, gm_n3467, gm_n3468, gm_n3469, gm_n347, gm_n3470, gm_n3471, gm_n3472, gm_n3473, gm_n3474, gm_n3475, gm_n3476, gm_n3477, gm_n3478, gm_n3479, gm_n348, gm_n3480, gm_n3481, gm_n3482, gm_n3483, gm_n3484, gm_n3485, gm_n3486, gm_n3487, gm_n3488, gm_n3489, gm_n349, gm_n3490, gm_n3491, gm_n3492, gm_n3493, gm_n3494, gm_n3495, gm_n3496, gm_n3497, gm_n3498, gm_n3499, gm_n350, gm_n3500, gm_n3501, gm_n3502, gm_n3503, gm_n3504, gm_n3505, gm_n3506, gm_n3507, gm_n3508, gm_n3509, gm_n351, gm_n3510, gm_n3511, gm_n3512, gm_n3513, gm_n3514, gm_n3515, gm_n3516, gm_n3517, gm_n3518, gm_n3519, gm_n352, gm_n3520, gm_n3521, gm_n3522, gm_n3523, gm_n3524, gm_n3525, gm_n3526, gm_n3527, gm_n3528, gm_n3529, gm_n353, gm_n3530, gm_n3531, gm_n3532, gm_n3533, gm_n3534, gm_n3535, gm_n3536, gm_n3537, gm_n3538, gm_n3539, gm_n354, gm_n3540, gm_n3541, gm_n3542, gm_n3543, gm_n3544, gm_n3545, gm_n3546, gm_n3547, gm_n3548, gm_n3549, gm_n355, gm_n3550, gm_n3551, gm_n3552, gm_n3553, gm_n3554, gm_n3555, gm_n3556, gm_n3557, gm_n3558, gm_n3559, gm_n356, gm_n3560, gm_n3561, gm_n3562, gm_n3563, gm_n3564, gm_n3565, gm_n3566, gm_n3567, gm_n3568, gm_n3569, gm_n357, gm_n3570, gm_n3571, gm_n3572, gm_n3573, gm_n3574, gm_n3575, gm_n3576, gm_n3577, gm_n3578, gm_n3579, gm_n358, gm_n3580, gm_n3581, gm_n3582, gm_n3583, gm_n3584, gm_n3585, gm_n3586, gm_n3587, gm_n3588, gm_n3589, gm_n359, gm_n3590, gm_n3591, gm_n3592, gm_n3593, gm_n3594, gm_n3595, gm_n3596, gm_n3597, gm_n3598, gm_n3599, gm_n360, gm_n3600, gm_n3601, gm_n3602, gm_n3603, gm_n3604, gm_n3605, gm_n3606, gm_n3607, gm_n3608, gm_n3609, gm_n361, gm_n3610, gm_n3611, gm_n3612, gm_n3613, gm_n3614, gm_n3615, gm_n3616, gm_n3617, gm_n3618, gm_n3619, gm_n362, gm_n3620, gm_n3621, gm_n3622, gm_n3623, gm_n3624, gm_n3625, gm_n3626, gm_n3627, gm_n3628, gm_n3629, gm_n363, gm_n3630, gm_n3631, gm_n3632, gm_n3633, gm_n3634, gm_n3635, gm_n3636, gm_n3637, gm_n3638, gm_n3639, gm_n364, gm_n3640, gm_n3641, gm_n3642, gm_n3643, gm_n3644, gm_n3645, gm_n3646, gm_n3647, gm_n3648, gm_n3649, gm_n365, gm_n3650, gm_n3651, gm_n3652, gm_n3653, gm_n3654, gm_n3655, gm_n3656, gm_n3657, gm_n3658, gm_n3659, gm_n366, gm_n3660, gm_n3661, gm_n3662, gm_n3663, gm_n3664, gm_n3665, gm_n3666, gm_n3667, gm_n3668, gm_n3669, gm_n367, gm_n3670, gm_n3671, gm_n3672, gm_n3673, gm_n3674, gm_n3675, gm_n3676, gm_n3677, gm_n3678, gm_n3679, gm_n368, gm_n3680, gm_n3681, gm_n3682, gm_n3683, gm_n3684, gm_n3685, gm_n3686, gm_n3687, gm_n3688, gm_n3689, gm_n369, gm_n3690, gm_n3691, gm_n3692, gm_n3693, gm_n3694, gm_n3695, gm_n3696, gm_n3697, gm_n3698, gm_n3699, gm_n370, gm_n3700, gm_n3701, gm_n3702, gm_n3703, gm_n3704, gm_n3705, gm_n3706, gm_n3707, gm_n3708, gm_n3709, gm_n371, gm_n3710, gm_n3711, gm_n3712, gm_n3713, gm_n3714, gm_n3715, gm_n3716, gm_n3717, gm_n3718, gm_n3719, gm_n372, gm_n3720, gm_n3721, gm_n3722, gm_n3723, gm_n3724, gm_n3725, gm_n3726, gm_n3727, gm_n3728, gm_n3729, gm_n373, gm_n3730, gm_n3731, gm_n3732, gm_n3733, gm_n3734, gm_n3735, gm_n3736, gm_n3737, gm_n3738, gm_n3739, gm_n374, gm_n3740, gm_n3741, gm_n3742, gm_n3743, gm_n3744, gm_n3745, gm_n3746, gm_n3747, gm_n3748, gm_n3749, gm_n375, gm_n3750, gm_n3751, gm_n3752, gm_n3753, gm_n3754, gm_n3755, gm_n3756, gm_n3757, gm_n3758, gm_n3759, gm_n376, gm_n3760, gm_n3761, gm_n3762, gm_n3763, gm_n3764, gm_n3765, gm_n3766, gm_n3767, gm_n3768, gm_n3769, gm_n377, gm_n3770, gm_n3771, gm_n3772, gm_n3773, gm_n3774, gm_n3775, gm_n3776, gm_n3777, gm_n3778, gm_n3779, gm_n378, gm_n3780, gm_n3781, gm_n3782, gm_n3783, gm_n3784, gm_n3785, gm_n3786, gm_n3787, gm_n3788, gm_n3789, gm_n379, gm_n3790, gm_n3791, gm_n3792, gm_n3793, gm_n3794, gm_n3795, gm_n3796, gm_n3797, gm_n3798, gm_n3799, gm_n380, gm_n3800, gm_n3801, gm_n3802, gm_n3803, gm_n3804, gm_n3805, gm_n3806, gm_n3807, gm_n3808, gm_n3809, gm_n381, gm_n3810, gm_n3811, gm_n3812, gm_n3813, gm_n3814, gm_n3815, gm_n3816, gm_n3817, gm_n3818, gm_n3819, gm_n382, gm_n3820, gm_n3821, gm_n3822, gm_n3823, gm_n3824, gm_n3825, gm_n3826, gm_n3827, gm_n3828, gm_n3829, gm_n383, gm_n3830, gm_n3831, gm_n3832, gm_n3833, gm_n3834, gm_n3835, gm_n3836, gm_n3837, gm_n3838, gm_n3839, gm_n384, gm_n3840, gm_n3841, gm_n3842, gm_n3843, gm_n3844, gm_n3845, gm_n3846, gm_n3847, gm_n3848, gm_n3849, gm_n385, gm_n3850, gm_n3851, gm_n3852, gm_n3853, gm_n3854, gm_n3855, gm_n3856, gm_n3857, gm_n3858, gm_n3859, gm_n386, gm_n3860, gm_n3861, gm_n3862, gm_n3863, gm_n3864, gm_n3865, gm_n3866, gm_n3867, gm_n3868, gm_n3869, gm_n387, gm_n3870, gm_n3871, gm_n3872, gm_n3873, gm_n3874, gm_n3875, gm_n3876, gm_n3877, gm_n3878, gm_n3879, gm_n388, gm_n3880, gm_n3881, gm_n3882, gm_n3883, gm_n3884, gm_n3885, gm_n3886, gm_n3887, gm_n3888, gm_n3889, gm_n389, gm_n3890, gm_n3891, gm_n3892, gm_n3893, gm_n3894, gm_n3895, gm_n3896, gm_n3897, gm_n3898, gm_n3899, gm_n390, gm_n3900, gm_n3901, gm_n3902, gm_n3903, gm_n3904, gm_n3905, gm_n3906, gm_n3907, gm_n3908, gm_n3909, gm_n391, gm_n3910, gm_n3911, gm_n3912, gm_n3913, gm_n3914, gm_n3915, gm_n3916, gm_n3917, gm_n3918, gm_n3919, gm_n392, gm_n3920, gm_n3921, gm_n3922, gm_n3923, gm_n3924, gm_n3925, gm_n3926, gm_n3927, gm_n3928, gm_n3929, gm_n393, gm_n3930, gm_n3931, gm_n3932, gm_n3933, gm_n3934, gm_n3935, gm_n3936, gm_n3937, gm_n3938, gm_n3939, gm_n394, gm_n3940, gm_n3941, gm_n3942, gm_n3943, gm_n3944, gm_n3945, gm_n3946, gm_n3947, gm_n3948, gm_n3949, gm_n395, gm_n3950, gm_n3951, gm_n3952, gm_n3953, gm_n3954, gm_n3955, gm_n3956, gm_n3957, gm_n3958, gm_n3959, gm_n396, gm_n3960, gm_n3961, gm_n3962, gm_n3963, gm_n3964, gm_n3965, gm_n3966, gm_n3967, gm_n3968, gm_n3969, gm_n397, gm_n3970, gm_n3971, gm_n3972, gm_n3973, gm_n3974, gm_n3975, gm_n3976, gm_n3977, gm_n3978, gm_n3979, gm_n398, gm_n3980, gm_n3981, gm_n3982, gm_n3983, gm_n3984, gm_n3985, gm_n3986, gm_n3987, gm_n3988, gm_n3989, gm_n399, gm_n3990, gm_n3991, gm_n3992, gm_n3993, gm_n3994, gm_n3995, gm_n3996, gm_n3997, gm_n3998, gm_n3999, gm_n400, gm_n4000, gm_n4001, gm_n4002, gm_n4003, gm_n4004, gm_n4005, gm_n4006, gm_n4007, gm_n4008, gm_n4009, gm_n401, gm_n4010, gm_n4011, gm_n4012, gm_n4013, gm_n4014, gm_n4015, gm_n4016, gm_n4017, gm_n4018, gm_n4019, gm_n402, gm_n4020, gm_n4021, gm_n4022, gm_n4023, gm_n4024, gm_n4026, gm_n4027, gm_n4028, gm_n4029, gm_n403, gm_n4030, gm_n4031, gm_n4032, gm_n4033, gm_n4034, gm_n4035, gm_n4036, gm_n4037, gm_n4038, gm_n4039, gm_n404, gm_n4040, gm_n4041, gm_n4042, gm_n4043, gm_n4044, gm_n4045, gm_n4046, gm_n4047, gm_n4048, gm_n4049, gm_n405, gm_n4050, gm_n4051, gm_n4052, gm_n4053, gm_n4054, gm_n4055, gm_n4056, gm_n4057, gm_n4058, gm_n4059, gm_n406, gm_n4060, gm_n4061, gm_n4062, gm_n4063, gm_n4064, gm_n4065, gm_n4066, gm_n4067, gm_n4068, gm_n4069, gm_n407, gm_n4070, gm_n4071, gm_n4072, gm_n4073, gm_n4074, gm_n4075, gm_n4076, gm_n4077, gm_n4078, gm_n4079, gm_n408, gm_n4080, gm_n4081, gm_n4082, gm_n4083, gm_n4084, gm_n4085, gm_n4086, gm_n4087, gm_n4088, gm_n4089, gm_n409, gm_n4090, gm_n4091, gm_n4092, gm_n4093, gm_n4094, gm_n4095, gm_n4096, gm_n4097, gm_n4098, gm_n4099, gm_n410, gm_n4100, gm_n4101, gm_n4102, gm_n4103, gm_n4104, gm_n4105, gm_n4106, gm_n4107, gm_n4108, gm_n4109, gm_n411, gm_n4110, gm_n4111, gm_n4112, gm_n4113, gm_n4114, gm_n4115, gm_n4116, gm_n4117, gm_n4118, gm_n4119, gm_n412, gm_n4120, gm_n4121, gm_n4122, gm_n4123, gm_n4124, gm_n4125, gm_n4126, gm_n4127, gm_n4128, gm_n4129, gm_n413, gm_n4130, gm_n4131, gm_n4132, gm_n4133, gm_n4134, gm_n4135, gm_n4136, gm_n4137, gm_n4138, gm_n4139, gm_n414, gm_n4140, gm_n4141, gm_n4142, gm_n4143, gm_n4144, gm_n4145, gm_n4146, gm_n4147, gm_n4148, gm_n4149, gm_n415, gm_n4150, gm_n4151, gm_n4152, gm_n4153, gm_n4154, gm_n4155, gm_n4156, gm_n4157, gm_n4158, gm_n4159, gm_n416, gm_n4160, gm_n4161, gm_n4162, gm_n4163, gm_n4164, gm_n4165, gm_n4166, gm_n4167, gm_n4168, gm_n4169, gm_n417, gm_n4170, gm_n4171, gm_n4172, gm_n4173, gm_n4174, gm_n4175, gm_n4176, gm_n4177, gm_n4178, gm_n4179, gm_n418, gm_n4180, gm_n4181, gm_n4182, gm_n4183, gm_n4184, gm_n4185, gm_n4186, gm_n4187, gm_n4188, gm_n4189, gm_n419, gm_n4190, gm_n4191, gm_n4192, gm_n4193, gm_n4194, gm_n4195, gm_n4196, gm_n4197, gm_n4198, gm_n4199, gm_n420, gm_n4200, gm_n4201, gm_n4202, gm_n4203, gm_n4204, gm_n4205, gm_n4206, gm_n4207, gm_n4208, gm_n4209, gm_n421, gm_n4210, gm_n4211, gm_n4212, gm_n4213, gm_n4214, gm_n4215, gm_n4216, gm_n4217, gm_n4218, gm_n4219, gm_n422, gm_n4220, gm_n4221, gm_n4222, gm_n4223, gm_n4224, gm_n4225, gm_n4226, gm_n4227, gm_n4228, gm_n4229, gm_n423, gm_n4230, gm_n4231, gm_n4232, gm_n4233, gm_n4234, gm_n4235, gm_n4236, gm_n4237, gm_n4238, gm_n4239, gm_n424, gm_n4240, gm_n4241, gm_n4242, gm_n4243, gm_n4244, gm_n4245, gm_n4246, gm_n4247, gm_n4248, gm_n4249, gm_n425, gm_n4250, gm_n4251, gm_n4252, gm_n4253, gm_n4254, gm_n4255, gm_n4256, gm_n4257, gm_n4258, gm_n4259, gm_n426, gm_n4260, gm_n4261, gm_n4262, gm_n4263, gm_n4264, gm_n4265, gm_n4266, gm_n4267, gm_n4268, gm_n4269, gm_n427, gm_n4270, gm_n4271, gm_n4272, gm_n4273, gm_n4274, gm_n4275, gm_n4276, gm_n4277, gm_n4278, gm_n4279, gm_n428, gm_n4280, gm_n4281, gm_n4282, gm_n4283, gm_n4284, gm_n4285, gm_n4286, gm_n4287, gm_n4288, gm_n4289, gm_n429, gm_n4290, gm_n4291, gm_n4292, gm_n4293, gm_n4294, gm_n4295, gm_n4296, gm_n4297, gm_n4298, gm_n4299, gm_n430, gm_n4300, gm_n4301, gm_n4302, gm_n4303, gm_n4304, gm_n4305, gm_n4306, gm_n4307, gm_n4308, gm_n4309, gm_n431, gm_n4310, gm_n4311, gm_n4312, gm_n4313, gm_n4314, gm_n4315, gm_n4316, gm_n4317, gm_n4318, gm_n4319, gm_n432, gm_n4320, gm_n4321, gm_n4322, gm_n4323, gm_n4324, gm_n4325, gm_n4326, gm_n4327, gm_n4328, gm_n4329, gm_n433, gm_n4330, gm_n4331, gm_n4332, gm_n4333, gm_n4334, gm_n4335, gm_n4336, gm_n4337, gm_n4338, gm_n4339, gm_n434, gm_n4340, gm_n4341, gm_n4342, gm_n4343, gm_n4344, gm_n4345, gm_n4346, gm_n4347, gm_n4348, gm_n4349, gm_n435, gm_n4350, gm_n4351, gm_n4352, gm_n4353, gm_n4354, gm_n4355, gm_n4356, gm_n4357, gm_n4358, gm_n4359, gm_n436, gm_n4360, gm_n4361, gm_n4362, gm_n4363, gm_n4364, gm_n4365, gm_n4366, gm_n4367, gm_n4368, gm_n4369, gm_n437, gm_n4370, gm_n4371, gm_n4372, gm_n4373, gm_n4374, gm_n4375, gm_n4376, gm_n4377, gm_n4378, gm_n4379, gm_n438, gm_n4380, gm_n4381, gm_n4382, gm_n4383, gm_n4384, gm_n4385, gm_n4386, gm_n4387, gm_n4388, gm_n4389, gm_n439, gm_n4390, gm_n4391, gm_n4392, gm_n4393, gm_n4394, gm_n4395, gm_n4396, gm_n4397, gm_n4398, gm_n4399, gm_n440, gm_n4400, gm_n4401, gm_n4402, gm_n4403, gm_n4404, gm_n4405, gm_n4406, gm_n4407, gm_n4408, gm_n4409, gm_n441, gm_n4410, gm_n4411, gm_n4412, gm_n4413, gm_n4414, gm_n4415, gm_n4416, gm_n4417, gm_n4418, gm_n4419, gm_n442, gm_n4420, gm_n4421, gm_n4422, gm_n4423, gm_n4424, gm_n4425, gm_n4426, gm_n4427, gm_n4428, gm_n4429, gm_n443, gm_n4430, gm_n4431, gm_n4432, gm_n4433, gm_n4434, gm_n4435, gm_n4436, gm_n4437, gm_n4438, gm_n4439, gm_n444, gm_n4440, gm_n4441, gm_n4442, gm_n4443, gm_n4444, gm_n4445, gm_n4446, gm_n4447, gm_n4448, gm_n4449, gm_n445, gm_n4450, gm_n4451, gm_n4452, gm_n4453, gm_n4454, gm_n4455, gm_n4456, gm_n4457, gm_n4458, gm_n4459, gm_n446, gm_n4460, gm_n4461, gm_n4462, gm_n4463, gm_n4464, gm_n4465, gm_n4466, gm_n4467, gm_n4468, gm_n4469, gm_n447, gm_n4470, gm_n4471, gm_n4472, gm_n4473, gm_n4474, gm_n4475, gm_n4476, gm_n4477, gm_n4478, gm_n4479, gm_n448, gm_n4480, gm_n4481, gm_n4482, gm_n4483, gm_n4484, gm_n4485, gm_n4486, gm_n4487, gm_n4488, gm_n4489, gm_n449, gm_n4490, gm_n4491, gm_n4492, gm_n4493, gm_n4494, gm_n4495, gm_n4496, gm_n4497, gm_n4498, gm_n4499, gm_n45, gm_n450, gm_n4500, gm_n4501, gm_n4502, gm_n4503, gm_n4504, gm_n4505, gm_n4506, gm_n4507, gm_n4508, gm_n4509, gm_n451, gm_n4510, gm_n4511, gm_n4512, gm_n4513, gm_n4514, gm_n4515, gm_n4516, gm_n4517, gm_n4518, gm_n4519, gm_n452, gm_n4520, gm_n4521, gm_n4522, gm_n4523, gm_n4524, gm_n4525, gm_n4526, gm_n4527, gm_n4528, gm_n4529, gm_n453, gm_n4530, gm_n4531, gm_n4532, gm_n4533, gm_n4534, gm_n4535, gm_n4536, gm_n4537, gm_n4538, gm_n4539, gm_n454, gm_n4540, gm_n4541, gm_n4542, gm_n4543, gm_n4544, gm_n4545, gm_n4546, gm_n4547, gm_n4548, gm_n4549, gm_n455, gm_n4550, gm_n4551, gm_n4552, gm_n4553, gm_n4554, gm_n4555, gm_n4556, gm_n4557, gm_n4558, gm_n4559, gm_n456, gm_n4560, gm_n4561, gm_n4562, gm_n4563, gm_n4564, gm_n4565, gm_n4566, gm_n4567, gm_n4568, gm_n4569, gm_n457, gm_n4570, gm_n4571, gm_n4572, gm_n4573, gm_n4574, gm_n4575, gm_n4576, gm_n4577, gm_n4578, gm_n4579, gm_n458, gm_n4580, gm_n4581, gm_n4582, gm_n4583, gm_n4584, gm_n4585, gm_n4586, gm_n4587, gm_n4588, gm_n4589, gm_n459, gm_n4590, gm_n4591, gm_n4592, gm_n4593, gm_n4594, gm_n4595, gm_n4596, gm_n4597, gm_n4598, gm_n4599, gm_n46, gm_n460, gm_n4600, gm_n4601, gm_n4602, gm_n4603, gm_n4604, gm_n4605, gm_n4606, gm_n4607, gm_n4608, gm_n4609, gm_n461, gm_n4610, gm_n4611, gm_n4612, gm_n4613, gm_n4614, gm_n4615, gm_n4616, gm_n4618, gm_n4619, gm_n462, gm_n4620, gm_n4621, gm_n4622, gm_n4623, gm_n4624, gm_n4625, gm_n4626, gm_n4627, gm_n4628, gm_n4629, gm_n463, gm_n4630, gm_n4631, gm_n4632, gm_n4633, gm_n4634, gm_n4635, gm_n4636, gm_n4637, gm_n4638, gm_n4639, gm_n464, gm_n4640, gm_n4641, gm_n4642, gm_n4643, gm_n4644, gm_n4645, gm_n4646, gm_n4647, gm_n4648, gm_n4649, gm_n465, gm_n4650, gm_n4651, gm_n4652, gm_n4653, gm_n4654, gm_n4655, gm_n4656, gm_n4657, gm_n4658, gm_n4659, gm_n466, gm_n4660, gm_n4661, gm_n4662, gm_n4663, gm_n4664, gm_n4665, gm_n4666, gm_n4667, gm_n4668, gm_n4669, gm_n467, gm_n4670, gm_n4671, gm_n4672, gm_n4673, gm_n4674, gm_n4675, gm_n4676, gm_n4677, gm_n4678, gm_n4679, gm_n468, gm_n4680, gm_n4681, gm_n4682, gm_n4683, gm_n4684, gm_n4685, gm_n4686, gm_n4687, gm_n4688, gm_n4689, gm_n469, gm_n4690, gm_n4691, gm_n4692, gm_n4693, gm_n4694, gm_n4695, gm_n4696, gm_n4697, gm_n4698, gm_n4699, gm_n47, gm_n470, gm_n4700, gm_n4701, gm_n4702, gm_n4703, gm_n4704, gm_n4705, gm_n4706, gm_n4707, gm_n4708, gm_n4709, gm_n471, gm_n4710, gm_n4711, gm_n4712, gm_n4713, gm_n4714, gm_n4715, gm_n4716, gm_n4717, gm_n4718, gm_n4719, gm_n472, gm_n4720, gm_n4721, gm_n4722, gm_n4723, gm_n4724, gm_n4725, gm_n4726, gm_n4727, gm_n4728, gm_n4729, gm_n473, gm_n4730, gm_n4731, gm_n4732, gm_n4733, gm_n4734, gm_n4735, gm_n4736, gm_n4737, gm_n4738, gm_n4739, gm_n474, gm_n4740, gm_n4741, gm_n4742, gm_n4743, gm_n4744, gm_n4745, gm_n4746, gm_n4747, gm_n4748, gm_n4749, gm_n475, gm_n4750, gm_n4751, gm_n4752, gm_n4753, gm_n4754, gm_n4755, gm_n4756, gm_n4757, gm_n4758, gm_n4759, gm_n476, gm_n4760, gm_n4761, gm_n4762, gm_n4763, gm_n4764, gm_n4765, gm_n4766, gm_n4767, gm_n4768, gm_n4769, gm_n477, gm_n4770, gm_n4771, gm_n4772, gm_n4773, gm_n4774, gm_n4775, gm_n4776, gm_n4777, gm_n4778, gm_n4779, gm_n478, gm_n4780, gm_n4781, gm_n4782, gm_n4783, gm_n4784, gm_n4785, gm_n4786, gm_n4787, gm_n4788, gm_n4789, gm_n479, gm_n4790, gm_n4791, gm_n4792, gm_n4793, gm_n4794, gm_n4795, gm_n4796, gm_n4797, gm_n4798, gm_n4799, gm_n48, gm_n480, gm_n4800, gm_n4801, gm_n4802, gm_n4803, gm_n4804, gm_n4805, gm_n4806, gm_n4807, gm_n4808, gm_n4809, gm_n481, gm_n4810, gm_n4811, gm_n4812, gm_n4813, gm_n4814, gm_n4815, gm_n4816, gm_n4817, gm_n4818, gm_n4819, gm_n482, gm_n4820, gm_n4821, gm_n4822, gm_n4823, gm_n4824, gm_n4825, gm_n4826, gm_n4827, gm_n4828, gm_n4829, gm_n483, gm_n4830, gm_n4831, gm_n4832, gm_n4833, gm_n4834, gm_n4835, gm_n4836, gm_n4837, gm_n4838, gm_n4839, gm_n484, gm_n4840, gm_n4841, gm_n4842, gm_n4843, gm_n4844, gm_n4845, gm_n4846, gm_n4847, gm_n4848, gm_n4849, gm_n485, gm_n4850, gm_n4851, gm_n4852, gm_n4853, gm_n4854, gm_n4855, gm_n4856, gm_n4857, gm_n4858, gm_n4859, gm_n486, gm_n4860, gm_n4861, gm_n4862, gm_n4863, gm_n4864, gm_n4865, gm_n4866, gm_n4867, gm_n4868, gm_n4869, gm_n487, gm_n4870, gm_n4871, gm_n4872, gm_n4873, gm_n4874, gm_n4875, gm_n4876, gm_n4877, gm_n4878, gm_n4879, gm_n488, gm_n4880, gm_n4881, gm_n4882, gm_n4883, gm_n4884, gm_n4885, gm_n4886, gm_n4887, gm_n4888, gm_n4889, gm_n489, gm_n4890, gm_n4891, gm_n4892, gm_n4893, gm_n4894, gm_n4895, gm_n4896, gm_n4897, gm_n4898, gm_n4899, gm_n49, gm_n490, gm_n4900, gm_n4901, gm_n4902, gm_n4903, gm_n4904, gm_n4905, gm_n4906, gm_n4907, gm_n4908, gm_n4909, gm_n491, gm_n4910, gm_n4911, gm_n4912, gm_n4913, gm_n4914, gm_n4915, gm_n4916, gm_n4917, gm_n4918, gm_n4919, gm_n492, gm_n4920, gm_n4921, gm_n4922, gm_n4923, gm_n4924, gm_n4925, gm_n4926, gm_n4927, gm_n4928, gm_n4929, gm_n493, gm_n4930, gm_n4931, gm_n4932, gm_n4933, gm_n4934, gm_n4935, gm_n4936, gm_n4937, gm_n4938, gm_n4939, gm_n494, gm_n4940, gm_n4941, gm_n4942, gm_n4943, gm_n4944, gm_n4945, gm_n4946, gm_n4947, gm_n4948, gm_n4949, gm_n495, gm_n4950, gm_n4951, gm_n4952, gm_n4953, gm_n4954, gm_n4955, gm_n4956, gm_n4957, gm_n4958, gm_n4959, gm_n496, gm_n4960, gm_n4961, gm_n4962, gm_n4963, gm_n4964, gm_n4965, gm_n4966, gm_n4967, gm_n4968, gm_n4969, gm_n497, gm_n4970, gm_n4971, gm_n4972, gm_n4973, gm_n4974, gm_n4975, gm_n4976, gm_n4977, gm_n4978, gm_n4979, gm_n498, gm_n4980, gm_n4981, gm_n4982, gm_n4983, gm_n4984, gm_n4985, gm_n4986, gm_n4987, gm_n4988, gm_n4989, gm_n499, gm_n4990, gm_n4991, gm_n4992, gm_n4993, gm_n4994, gm_n4995, gm_n4996, gm_n4997, gm_n4998, gm_n4999, gm_n50, gm_n500, gm_n5000, gm_n5001, gm_n5002, gm_n5003, gm_n5004, gm_n5005, gm_n5006, gm_n5007, gm_n5008, gm_n5009, gm_n501, gm_n5010, gm_n5011, gm_n5012, gm_n5013, gm_n5014, gm_n5015, gm_n5016, gm_n5017, gm_n5018, gm_n5019, gm_n502, gm_n5020, gm_n5021, gm_n5022, gm_n5023, gm_n5024, gm_n5025, gm_n5026, gm_n5027, gm_n5028, gm_n5029, gm_n503, gm_n5030, gm_n5031, gm_n5032, gm_n5033, gm_n5034, gm_n5035, gm_n5036, gm_n5037, gm_n5038, gm_n5039, gm_n504, gm_n5040, gm_n5041, gm_n5042, gm_n5043, gm_n5044, gm_n5045, gm_n5046, gm_n5047, gm_n5048, gm_n5049, gm_n505, gm_n5050, gm_n5051, gm_n5052, gm_n5053, gm_n5054, gm_n5055, gm_n5056, gm_n5057, gm_n5058, gm_n5059, gm_n506, gm_n5060, gm_n5061, gm_n5062, gm_n5063, gm_n5064, gm_n5065, gm_n5066, gm_n5067, gm_n5068, gm_n5069, gm_n507, gm_n5070, gm_n5071, gm_n5072, gm_n5073, gm_n5074, gm_n5075, gm_n5076, gm_n5077, gm_n5078, gm_n5079, gm_n508, gm_n5080, gm_n5081, gm_n5082, gm_n5083, gm_n5084, gm_n5085, gm_n5086, gm_n5087, gm_n5088, gm_n5089, gm_n509, gm_n5090, gm_n5091, gm_n5092, gm_n5093, gm_n5094, gm_n5095, gm_n5096, gm_n5097, gm_n5098, gm_n5099, gm_n51, gm_n510, gm_n5100, gm_n5101, gm_n5102, gm_n5103, gm_n5104, gm_n5105, gm_n5106, gm_n5107, gm_n5108, gm_n5109, gm_n511, gm_n5110, gm_n5111, gm_n5112, gm_n5113, gm_n5114, gm_n5115, gm_n5116, gm_n5117, gm_n5118, gm_n5119, gm_n512, gm_n5120, gm_n5121, gm_n5122, gm_n5123, gm_n5124, gm_n5125, gm_n5126, gm_n5127, gm_n5128, gm_n5129, gm_n513, gm_n5130, gm_n5131, gm_n5132, gm_n5133, gm_n5134, gm_n5135, gm_n5136, gm_n5137, gm_n5138, gm_n5139, gm_n514, gm_n5140, gm_n5141, gm_n5142, gm_n5143, gm_n5144, gm_n5145, gm_n5146, gm_n5147, gm_n5148, gm_n5149, gm_n515, gm_n5150, gm_n5151, gm_n5152, gm_n5153, gm_n5154, gm_n5155, gm_n5156, gm_n5157, gm_n5158, gm_n5159, gm_n516, gm_n5160, gm_n5161, gm_n5162, gm_n5163, gm_n5164, gm_n5165, gm_n5166, gm_n5167, gm_n5168, gm_n5169, gm_n517, gm_n5170, gm_n5171, gm_n5172, gm_n5173, gm_n5174, gm_n5175, gm_n5176, gm_n5177, gm_n5178, gm_n518, gm_n5180, gm_n5181, gm_n5182, gm_n5183, gm_n5184, gm_n5185, gm_n5186, gm_n5187, gm_n5188, gm_n5189, gm_n519, gm_n5190, gm_n5191, gm_n5192, gm_n5193, gm_n5194, gm_n5195, gm_n5196, gm_n5197, gm_n5198, gm_n5199, gm_n52, gm_n520, gm_n5200, gm_n5201, gm_n5202, gm_n5203, gm_n5204, gm_n5205, gm_n5206, gm_n5207, gm_n5208, gm_n5209, gm_n521, gm_n5210, gm_n5211, gm_n5212, gm_n5213, gm_n5214, gm_n5215, gm_n5216, gm_n5217, gm_n5218, gm_n5219, gm_n522, gm_n5220, gm_n5221, gm_n5222, gm_n5223, gm_n5224, gm_n5225, gm_n5226, gm_n5227, gm_n5228, gm_n5229, gm_n523, gm_n5230, gm_n5231, gm_n5232, gm_n5233, gm_n5234, gm_n5235, gm_n5236, gm_n5237, gm_n5238, gm_n5239, gm_n524, gm_n5240, gm_n5241, gm_n5242, gm_n5243, gm_n5244, gm_n5245, gm_n5246, gm_n5247, gm_n5248, gm_n5249, gm_n525, gm_n5250, gm_n5251, gm_n5252, gm_n5253, gm_n5254, gm_n5255, gm_n5256, gm_n5257, gm_n5258, gm_n5259, gm_n526, gm_n5260, gm_n5261, gm_n5262, gm_n5263, gm_n5264, gm_n5265, gm_n5266, gm_n5267, gm_n5268, gm_n5269, gm_n527, gm_n5270, gm_n5271, gm_n5272, gm_n5273, gm_n5274, gm_n5275, gm_n5276, gm_n5277, gm_n5278, gm_n5279, gm_n528, gm_n5280, gm_n5281, gm_n5282, gm_n5283, gm_n5284, gm_n5285, gm_n5286, gm_n5287, gm_n5288, gm_n5289, gm_n529, gm_n5290, gm_n5291, gm_n5292, gm_n5293, gm_n5294, gm_n5295, gm_n5296, gm_n5297, gm_n5298, gm_n5299, gm_n53, gm_n530, gm_n5300, gm_n5301, gm_n5302, gm_n5303, gm_n5304, gm_n5305, gm_n5306, gm_n5307, gm_n5308, gm_n5309, gm_n531, gm_n5310, gm_n5311, gm_n5312, gm_n5313, gm_n5314, gm_n5315, gm_n5316, gm_n5317, gm_n5318, gm_n5319, gm_n532, gm_n5320, gm_n5321, gm_n5322, gm_n5323, gm_n5324, gm_n5325, gm_n5326, gm_n5327, gm_n5328, gm_n5329, gm_n533, gm_n5330, gm_n5331, gm_n5332, gm_n5333, gm_n5334, gm_n5335, gm_n5336, gm_n5337, gm_n5338, gm_n5339, gm_n534, gm_n5340, gm_n5341, gm_n5342, gm_n5343, gm_n5344, gm_n5345, gm_n5346, gm_n5347, gm_n5348, gm_n5349, gm_n535, gm_n5350, gm_n5351, gm_n5352, gm_n5353, gm_n5354, gm_n5355, gm_n5356, gm_n5357, gm_n5358, gm_n5359, gm_n536, gm_n5360, gm_n5361, gm_n5362, gm_n5363, gm_n5364, gm_n5365, gm_n5366, gm_n5367, gm_n5368, gm_n5369, gm_n537, gm_n5370, gm_n5371, gm_n5372, gm_n5373, gm_n5374, gm_n5375, gm_n5376, gm_n5377, gm_n5378, gm_n5379, gm_n538, gm_n5380, gm_n5381, gm_n5382, gm_n5383, gm_n5384, gm_n5385, gm_n5386, gm_n5387, gm_n5388, gm_n5389, gm_n539, gm_n5390, gm_n5391, gm_n5392, gm_n5393, gm_n5394, gm_n5395, gm_n5396, gm_n5397, gm_n5398, gm_n5399, gm_n54, gm_n540, gm_n5400, gm_n5401, gm_n5402, gm_n5403, gm_n5404, gm_n5405, gm_n5406, gm_n5407, gm_n5408, gm_n5409, gm_n541, gm_n5410, gm_n5411, gm_n5412, gm_n5413, gm_n5414, gm_n5415, gm_n5416, gm_n5417, gm_n5418, gm_n5419, gm_n542, gm_n5420, gm_n5421, gm_n5422, gm_n5423, gm_n5424, gm_n5425, gm_n5426, gm_n5427, gm_n5428, gm_n5429, gm_n543, gm_n5430, gm_n5431, gm_n5432, gm_n5433, gm_n5434, gm_n5435, gm_n5436, gm_n5437, gm_n5438, gm_n5439, gm_n544, gm_n5440, gm_n5441, gm_n5442, gm_n5443, gm_n5444, gm_n5445, gm_n5446, gm_n5447, gm_n5448, gm_n5449, gm_n545, gm_n5450, gm_n5451, gm_n5452, gm_n5453, gm_n5454, gm_n5455, gm_n5456, gm_n5457, gm_n5458, gm_n5459, gm_n546, gm_n5460, gm_n5461, gm_n5462, gm_n5463, gm_n5464, gm_n5465, gm_n5466, gm_n5467, gm_n5468, gm_n5469, gm_n547, gm_n5470, gm_n5471, gm_n5472, gm_n5473, gm_n5474, gm_n5475, gm_n5476, gm_n5477, gm_n5478, gm_n5479, gm_n548, gm_n5480, gm_n5481, gm_n5482, gm_n5483, gm_n5484, gm_n5485, gm_n5486, gm_n5487, gm_n5488, gm_n5489, gm_n549, gm_n5490, gm_n5491, gm_n5492, gm_n5493, gm_n5494, gm_n5495, gm_n5496, gm_n5497, gm_n5498, gm_n5499, gm_n55, gm_n550, gm_n5500, gm_n5501, gm_n5502, gm_n5503, gm_n5504, gm_n5505, gm_n5506, gm_n5507, gm_n5508, gm_n5509, gm_n551, gm_n5510, gm_n5511, gm_n5512, gm_n5513, gm_n5514, gm_n5515, gm_n5516, gm_n5517, gm_n5518, gm_n5519, gm_n552, gm_n5520, gm_n5521, gm_n5522, gm_n5523, gm_n5524, gm_n5525, gm_n5526, gm_n5527, gm_n5528, gm_n5529, gm_n553, gm_n5530, gm_n5531, gm_n5532, gm_n5533, gm_n5534, gm_n5535, gm_n5536, gm_n5537, gm_n5538, gm_n5539, gm_n554, gm_n5540, gm_n5541, gm_n5542, gm_n5543, gm_n5544, gm_n5545, gm_n5546, gm_n5547, gm_n5548, gm_n5549, gm_n555, gm_n5550, gm_n5551, gm_n5552, gm_n5553, gm_n5554, gm_n5555, gm_n5556, gm_n5557, gm_n5558, gm_n5559, gm_n556, gm_n5560, gm_n5561, gm_n5562, gm_n5563, gm_n5564, gm_n5565, gm_n5566, gm_n5567, gm_n5568, gm_n5569, gm_n557, gm_n5570, gm_n5571, gm_n5572, gm_n5573, gm_n5574, gm_n5575, gm_n5576, gm_n5577, gm_n5578, gm_n5579, gm_n558, gm_n5580, gm_n5581, gm_n5582, gm_n5583, gm_n5584, gm_n5585, gm_n5586, gm_n5587, gm_n5588, gm_n5589, gm_n559, gm_n5590, gm_n5591, gm_n5592, gm_n5593, gm_n5594, gm_n5595, gm_n5596, gm_n5597, gm_n5598, gm_n5599, gm_n56, gm_n560, gm_n5600, gm_n5601, gm_n5602, gm_n5603, gm_n5604, gm_n5605, gm_n5606, gm_n5607, gm_n5608, gm_n5609, gm_n561, gm_n5610, gm_n5611, gm_n5612, gm_n5613, gm_n5614, gm_n5615, gm_n5616, gm_n5617, gm_n5618, gm_n5619, gm_n562, gm_n5620, gm_n5621, gm_n5622, gm_n5623, gm_n5624, gm_n5625, gm_n5626, gm_n5627, gm_n5628, gm_n5629, gm_n563, gm_n5630, gm_n5631, gm_n5632, gm_n5633, gm_n5634, gm_n5635, gm_n5636, gm_n5637, gm_n5638, gm_n5639, gm_n564, gm_n5640, gm_n5641, gm_n5642, gm_n5643, gm_n5644, gm_n5645, gm_n5646, gm_n5647, gm_n5648, gm_n5649, gm_n565, gm_n5650, gm_n5651, gm_n5652, gm_n5653, gm_n5654, gm_n5655, gm_n5656, gm_n5657, gm_n5658, gm_n5659, gm_n566, gm_n5660, gm_n5661, gm_n5662, gm_n5663, gm_n5664, gm_n5665, gm_n5666, gm_n5667, gm_n5668, gm_n5669, gm_n567, gm_n5670, gm_n5671, gm_n5672, gm_n5673, gm_n5674, gm_n5675, gm_n5676, gm_n5677, gm_n5678, gm_n5679, gm_n568, gm_n5680, gm_n5681, gm_n5682, gm_n5683, gm_n5684, gm_n5685, gm_n5686, gm_n5687, gm_n5688, gm_n5689, gm_n569, gm_n5690, gm_n5691, gm_n5692, gm_n5693, gm_n5694, gm_n5695, gm_n5696, gm_n5697, gm_n5698, gm_n5699, gm_n57, gm_n570, gm_n5700, gm_n5701, gm_n5702, gm_n5703, gm_n5704, gm_n5705, gm_n5706, gm_n5707, gm_n5708, gm_n5709, gm_n571, gm_n5710, gm_n5711, gm_n5712, gm_n5713, gm_n5714, gm_n5715, gm_n5716, gm_n5717, gm_n5718, gm_n5719, gm_n572, gm_n5720, gm_n5721, gm_n5722, gm_n5723, gm_n5724, gm_n5725, gm_n5726, gm_n5727, gm_n5728, gm_n5729, gm_n573, gm_n5730, gm_n5731, gm_n5732, gm_n5733, gm_n5734, gm_n5735, gm_n5736, gm_n5737, gm_n5738, gm_n5739, gm_n574, gm_n5741, gm_n5742, gm_n5743, gm_n5744, gm_n5745, gm_n5746, gm_n5747, gm_n5748, gm_n5749, gm_n575, gm_n5750, gm_n5751, gm_n5752, gm_n5753, gm_n5754, gm_n5755, gm_n5756, gm_n5757, gm_n5758, gm_n5759, gm_n576, gm_n5760, gm_n5761, gm_n5762, gm_n5763, gm_n5764, gm_n5765, gm_n5766, gm_n5767, gm_n5768, gm_n5769, gm_n577, gm_n5770, gm_n5771, gm_n5772, gm_n5773, gm_n5774, gm_n5775, gm_n5776, gm_n5777, gm_n5778, gm_n5779, gm_n578, gm_n5780, gm_n5781, gm_n5782, gm_n5783, gm_n5784, gm_n5785, gm_n5786, gm_n5787, gm_n5788, gm_n5789, gm_n579, gm_n5790, gm_n5791, gm_n5792, gm_n5793, gm_n5794, gm_n5795, gm_n5796, gm_n5797, gm_n5798, gm_n5799, gm_n58, gm_n580, gm_n5800, gm_n5801, gm_n5802, gm_n5803, gm_n5804, gm_n5805, gm_n5806, gm_n5807, gm_n5808, gm_n5809, gm_n581, gm_n5810, gm_n5811, gm_n5812, gm_n5813, gm_n5814, gm_n5815, gm_n5816, gm_n5817, gm_n5818, gm_n5819, gm_n582, gm_n5820, gm_n5821, gm_n5822, gm_n5823, gm_n5824, gm_n5825, gm_n5826, gm_n5827, gm_n5828, gm_n5829, gm_n583, gm_n5830, gm_n5831, gm_n5832, gm_n5833, gm_n5834, gm_n5835, gm_n5836, gm_n5837, gm_n5838, gm_n5839, gm_n584, gm_n5840, gm_n5841, gm_n5842, gm_n5843, gm_n5844, gm_n5845, gm_n5846, gm_n5847, gm_n5848, gm_n5849, gm_n585, gm_n5850, gm_n5851, gm_n5852, gm_n5853, gm_n5854, gm_n5855, gm_n5856, gm_n5857, gm_n5858, gm_n5859, gm_n586, gm_n5860, gm_n5861, gm_n5862, gm_n5863, gm_n5864, gm_n5865, gm_n5866, gm_n5867, gm_n5868, gm_n5869, gm_n587, gm_n5870, gm_n5871, gm_n5872, gm_n5873, gm_n5874, gm_n5875, gm_n5876, gm_n5877, gm_n5878, gm_n5879, gm_n588, gm_n5880, gm_n5881, gm_n5882, gm_n5883, gm_n5884, gm_n5885, gm_n5886, gm_n5887, gm_n5888, gm_n5889, gm_n589, gm_n5890, gm_n5891, gm_n5892, gm_n5893, gm_n5894, gm_n5895, gm_n5896, gm_n5897, gm_n5898, gm_n5899, gm_n59, gm_n590, gm_n5900, gm_n5901, gm_n5902, gm_n5903, gm_n5904, gm_n5905, gm_n5906, gm_n5907, gm_n5908, gm_n5909, gm_n591, gm_n5910, gm_n5911, gm_n5912, gm_n5913, gm_n5914, gm_n5915, gm_n5916, gm_n5917, gm_n5918, gm_n5919, gm_n592, gm_n5920, gm_n5921, gm_n5922, gm_n5923, gm_n5924, gm_n5925, gm_n5926, gm_n5927, gm_n5928, gm_n5929, gm_n593, gm_n5930, gm_n5931, gm_n5932, gm_n5933, gm_n5934, gm_n5935, gm_n5936, gm_n5937, gm_n5938, gm_n5939, gm_n594, gm_n5940, gm_n5941, gm_n5942, gm_n5943, gm_n5944, gm_n5945, gm_n5946, gm_n5947, gm_n5948, gm_n5949, gm_n595, gm_n5950, gm_n5951, gm_n5952, gm_n5953, gm_n5954, gm_n5955, gm_n5956, gm_n5957, gm_n5958, gm_n5959, gm_n596, gm_n5960, gm_n5961, gm_n5962, gm_n5963, gm_n5964, gm_n5965, gm_n5966, gm_n5967, gm_n5968, gm_n5969, gm_n597, gm_n5970, gm_n5971, gm_n5972, gm_n5973, gm_n5974, gm_n5975, gm_n5976, gm_n5977, gm_n5978, gm_n5979, gm_n598, gm_n5980, gm_n5981, gm_n5982, gm_n5983, gm_n5984, gm_n5985, gm_n5986, gm_n5987, gm_n5988, gm_n5989, gm_n599, gm_n5990, gm_n5991, gm_n5992, gm_n5993, gm_n5994, gm_n5995, gm_n5996, gm_n5997, gm_n5998, gm_n5999, gm_n60, gm_n600, gm_n6000, gm_n6001, gm_n6002, gm_n6003, gm_n6004, gm_n6005, gm_n6006, gm_n6007, gm_n6008, gm_n6009, gm_n601, gm_n6010, gm_n6011, gm_n6012, gm_n6013, gm_n6014, gm_n6015, gm_n6016, gm_n6017, gm_n6018, gm_n6019, gm_n602, gm_n6020, gm_n6021, gm_n6022, gm_n6023, gm_n6024, gm_n6025, gm_n6026, gm_n6027, gm_n6028, gm_n6029, gm_n603, gm_n6030, gm_n6031, gm_n6032, gm_n6033, gm_n6034, gm_n6035, gm_n6036, gm_n6037, gm_n6038, gm_n6039, gm_n604, gm_n6040, gm_n6041, gm_n6042, gm_n6043, gm_n6044, gm_n6045, gm_n6046, gm_n6047, gm_n6048, gm_n6049, gm_n605, gm_n6050, gm_n6051, gm_n6052, gm_n6053, gm_n6054, gm_n6055, gm_n6056, gm_n6057, gm_n6058, gm_n6059, gm_n606, gm_n6060, gm_n6061, gm_n6062, gm_n6063, gm_n6064, gm_n6065, gm_n6066, gm_n6067, gm_n6068, gm_n6069, gm_n607, gm_n6070, gm_n6071, gm_n6072, gm_n6073, gm_n6074, gm_n6075, gm_n6076, gm_n6077, gm_n6078, gm_n6079, gm_n608, gm_n6080, gm_n6081, gm_n6082, gm_n6083, gm_n6084, gm_n6085, gm_n6086, gm_n6087, gm_n6088, gm_n6089, gm_n609, gm_n6090, gm_n6091, gm_n6092, gm_n6093, gm_n6094, gm_n6095, gm_n6096, gm_n6097, gm_n6098, gm_n6099, gm_n61, gm_n610, gm_n6100, gm_n6101, gm_n6102, gm_n6103, gm_n6104, gm_n6105, gm_n6106, gm_n6107, gm_n6108, gm_n6109, gm_n611, gm_n6110, gm_n6111, gm_n6112, gm_n6113, gm_n6114, gm_n6115, gm_n6116, gm_n6117, gm_n6118, gm_n6119, gm_n612, gm_n6120, gm_n6121, gm_n6122, gm_n6123, gm_n6124, gm_n6125, gm_n6126, gm_n6127, gm_n6128, gm_n6129, gm_n613, gm_n6130, gm_n6131, gm_n6132, gm_n6133, gm_n6134, gm_n6135, gm_n6136, gm_n6137, gm_n6138, gm_n6139, gm_n614, gm_n6140, gm_n6141, gm_n6142, gm_n6143, gm_n6144, gm_n6145, gm_n6146, gm_n6147, gm_n6148, gm_n6149, gm_n615, gm_n6150, gm_n6151, gm_n6152, gm_n6153, gm_n6154, gm_n6155, gm_n6156, gm_n6157, gm_n6158, gm_n6159, gm_n616, gm_n6160, gm_n6161, gm_n6162, gm_n6163, gm_n6164, gm_n6165, gm_n6166, gm_n6167, gm_n6168, gm_n6169, gm_n617, gm_n6170, gm_n6171, gm_n6172, gm_n6173, gm_n6174, gm_n6175, gm_n6176, gm_n6177, gm_n6178, gm_n6179, gm_n618, gm_n6180, gm_n6181, gm_n6182, gm_n6183, gm_n6184, gm_n6185, gm_n6186, gm_n6187, gm_n6188, gm_n6189, gm_n619, gm_n6190, gm_n6191, gm_n6192, gm_n6193, gm_n6194, gm_n6195, gm_n6196, gm_n6197, gm_n6198, gm_n6199, gm_n62, gm_n620, gm_n6200, gm_n6201, gm_n6202, gm_n6203, gm_n6204, gm_n6205, gm_n6206, gm_n6207, gm_n6208, gm_n6209, gm_n621, gm_n6210, gm_n6211, gm_n6212, gm_n6213, gm_n6214, gm_n6215, gm_n6216, gm_n6217, gm_n6218, gm_n6219, gm_n622, gm_n6220, gm_n6221, gm_n6222, gm_n6223, gm_n6224, gm_n6225, gm_n6226, gm_n6227, gm_n6228, gm_n6229, gm_n623, gm_n6230, gm_n6231, gm_n6232, gm_n6233, gm_n6234, gm_n6235, gm_n6236, gm_n6237, gm_n6238, gm_n6239, gm_n624, gm_n6240, gm_n6241, gm_n6242, gm_n6243, gm_n6244, gm_n6245, gm_n6246, gm_n6247, gm_n6248, gm_n6249, gm_n625, gm_n6250, gm_n6251, gm_n6252, gm_n6253, gm_n6254, gm_n6255, gm_n6256, gm_n6257, gm_n6258, gm_n6259, gm_n626, gm_n6260, gm_n6261, gm_n6262, gm_n6263, gm_n6264, gm_n6265, gm_n6266, gm_n6267, gm_n6268, gm_n6269, gm_n627, gm_n6270, gm_n6271, gm_n6272, gm_n6273, gm_n6274, gm_n6275, gm_n6276, gm_n6277, gm_n6278, gm_n6279, gm_n628, gm_n6280, gm_n6281, gm_n6282, gm_n6283, gm_n6284, gm_n6285, gm_n6286, gm_n6288, gm_n6289, gm_n629, gm_n6290, gm_n6291, gm_n6292, gm_n6293, gm_n6294, gm_n6295, gm_n6296, gm_n6297, gm_n6298, gm_n6299, gm_n63, gm_n630, gm_n6300, gm_n6301, gm_n6302, gm_n6303, gm_n6304, gm_n6305, gm_n6306, gm_n6307, gm_n6308, gm_n6309, gm_n631, gm_n6310, gm_n6311, gm_n6312, gm_n6313, gm_n6314, gm_n6315, gm_n6316, gm_n6317, gm_n6318, gm_n6319, gm_n632, gm_n6320, gm_n6321, gm_n6322, gm_n6323, gm_n6324, gm_n6325, gm_n6326, gm_n6327, gm_n6328, gm_n6329, gm_n633, gm_n6330, gm_n6331, gm_n6332, gm_n6333, gm_n6334, gm_n6335, gm_n6336, gm_n6337, gm_n6338, gm_n6339, gm_n634, gm_n6340, gm_n6341, gm_n6342, gm_n6343, gm_n6344, gm_n6345, gm_n6346, gm_n6347, gm_n6348, gm_n6349, gm_n635, gm_n6350, gm_n6351, gm_n6352, gm_n6353, gm_n6354, gm_n6355, gm_n6356, gm_n6357, gm_n6358, gm_n6359, gm_n636, gm_n6360, gm_n6361, gm_n6362, gm_n6363, gm_n6364, gm_n6365, gm_n6366, gm_n6367, gm_n6368, gm_n6369, gm_n637, gm_n6370, gm_n6371, gm_n6372, gm_n6373, gm_n6374, gm_n6375, gm_n6376, gm_n6377, gm_n6378, gm_n6379, gm_n638, gm_n6380, gm_n6381, gm_n6382, gm_n6383, gm_n6384, gm_n6385, gm_n6386, gm_n6387, gm_n6388, gm_n6389, gm_n639, gm_n6390, gm_n6391, gm_n6392, gm_n6393, gm_n6394, gm_n6395, gm_n6396, gm_n6397, gm_n6398, gm_n6399, gm_n64, gm_n640, gm_n6400, gm_n6401, gm_n6402, gm_n6403, gm_n6404, gm_n6405, gm_n6406, gm_n6407, gm_n6408, gm_n6409, gm_n641, gm_n6410, gm_n6411, gm_n6412, gm_n6413, gm_n6414, gm_n6415, gm_n6416, gm_n6417, gm_n6418, gm_n6419, gm_n642, gm_n6420, gm_n6421, gm_n6422, gm_n6423, gm_n6424, gm_n6425, gm_n6426, gm_n6427, gm_n6428, gm_n6429, gm_n643, gm_n6430, gm_n6431, gm_n6432, gm_n6433, gm_n6434, gm_n6435, gm_n6436, gm_n6437, gm_n6438, gm_n6439, gm_n644, gm_n6440, gm_n6441, gm_n6442, gm_n6443, gm_n6444, gm_n6445, gm_n6446, gm_n6447, gm_n6448, gm_n6449, gm_n645, gm_n6450, gm_n6451, gm_n6452, gm_n6453, gm_n6454, gm_n6455, gm_n6456, gm_n6457, gm_n6458, gm_n6459, gm_n646, gm_n6460, gm_n6461, gm_n6462, gm_n6463, gm_n6464, gm_n6465, gm_n6466, gm_n6467, gm_n6468, gm_n6469, gm_n647, gm_n6470, gm_n6471, gm_n6472, gm_n6473, gm_n6474, gm_n6475, gm_n6476, gm_n6477, gm_n6478, gm_n6479, gm_n648, gm_n6480, gm_n6481, gm_n6482, gm_n6483, gm_n6484, gm_n6485, gm_n6486, gm_n6487, gm_n6488, gm_n6489, gm_n649, gm_n6490, gm_n6491, gm_n6492, gm_n6493, gm_n6494, gm_n6495, gm_n6496, gm_n6497, gm_n6498, gm_n6499, gm_n65, gm_n650, gm_n6500, gm_n6501, gm_n6502, gm_n6503, gm_n6504, gm_n6505, gm_n6506, gm_n6507, gm_n6508, gm_n6509, gm_n651, gm_n6510, gm_n6511, gm_n6512, gm_n6513, gm_n6514, gm_n6515, gm_n6516, gm_n6517, gm_n6518, gm_n6519, gm_n652, gm_n6520, gm_n6521, gm_n6522, gm_n6523, gm_n6524, gm_n6525, gm_n6526, gm_n6527, gm_n6528, gm_n6529, gm_n653, gm_n6530, gm_n6531, gm_n6532, gm_n6533, gm_n6534, gm_n6535, gm_n6536, gm_n6537, gm_n6538, gm_n6539, gm_n654, gm_n6540, gm_n6541, gm_n6542, gm_n6543, gm_n6544, gm_n6545, gm_n6546, gm_n6547, gm_n6548, gm_n6549, gm_n655, gm_n6550, gm_n6551, gm_n6552, gm_n6553, gm_n6554, gm_n6555, gm_n6556, gm_n6557, gm_n6558, gm_n6559, gm_n656, gm_n6560, gm_n6561, gm_n6562, gm_n6563, gm_n6564, gm_n6565, gm_n6566, gm_n6567, gm_n6568, gm_n6569, gm_n657, gm_n6570, gm_n6571, gm_n6572, gm_n6573, gm_n6574, gm_n6575, gm_n6576, gm_n6577, gm_n6578, gm_n6579, gm_n658, gm_n6580, gm_n6581, gm_n6582, gm_n6583, gm_n6584, gm_n6585, gm_n6586, gm_n6587, gm_n6588, gm_n6589, gm_n659, gm_n6590, gm_n6591, gm_n6592, gm_n6593, gm_n6594, gm_n6595, gm_n6596, gm_n6597, gm_n6598, gm_n6599, gm_n66, gm_n660, gm_n6600, gm_n6601, gm_n6602, gm_n6603, gm_n6604, gm_n6605, gm_n6606, gm_n6607, gm_n6608, gm_n6609, gm_n661, gm_n6610, gm_n6611, gm_n6612, gm_n6613, gm_n6614, gm_n6615, gm_n6616, gm_n6617, gm_n6618, gm_n6619, gm_n662, gm_n6620, gm_n6621, gm_n6622, gm_n6623, gm_n6624, gm_n6625, gm_n6626, gm_n6627, gm_n6628, gm_n6629, gm_n663, gm_n6630, gm_n6631, gm_n6632, gm_n6633, gm_n6634, gm_n6635, gm_n6636, gm_n6637, gm_n6638, gm_n6639, gm_n664, gm_n6640, gm_n6641, gm_n6642, gm_n6643, gm_n6644, gm_n6645, gm_n6646, gm_n6647, gm_n6648, gm_n6649, gm_n665, gm_n6650, gm_n6651, gm_n6652, gm_n6653, gm_n6654, gm_n6655, gm_n6656, gm_n6657, gm_n6658, gm_n6659, gm_n666, gm_n6660, gm_n6661, gm_n6662, gm_n6663, gm_n6664, gm_n6665, gm_n6666, gm_n6667, gm_n6668, gm_n6669, gm_n667, gm_n6670, gm_n6671, gm_n6672, gm_n6673, gm_n6674, gm_n6675, gm_n6676, gm_n6677, gm_n6678, gm_n6679, gm_n668, gm_n6680, gm_n6681, gm_n6682, gm_n6683, gm_n6684, gm_n6685, gm_n6686, gm_n6687, gm_n6688, gm_n6689, gm_n669, gm_n6690, gm_n6691, gm_n6692, gm_n6693, gm_n6694, gm_n6695, gm_n6696, gm_n6697, gm_n6698, gm_n6699, gm_n67, gm_n670, gm_n6700, gm_n6701, gm_n6702, gm_n6703, gm_n6704, gm_n6705, gm_n6706, gm_n6707, gm_n6708, gm_n6709, gm_n671, gm_n6710, gm_n6711, gm_n6712, gm_n6713, gm_n6714, gm_n6715, gm_n6716, gm_n6717, gm_n6718, gm_n6719, gm_n672, gm_n6720, gm_n6721, gm_n6722, gm_n6723, gm_n6724, gm_n6725, gm_n6726, gm_n6727, gm_n6728, gm_n6729, gm_n673, gm_n6730, gm_n6731, gm_n6732, gm_n6733, gm_n6734, gm_n6735, gm_n6736, gm_n6737, gm_n6738, gm_n6739, gm_n674, gm_n6740, gm_n6741, gm_n6742, gm_n6743, gm_n6744, gm_n6745, gm_n6746, gm_n6747, gm_n6748, gm_n6749, gm_n675, gm_n6750, gm_n6751, gm_n6752, gm_n6753, gm_n6754, gm_n6755, gm_n6756, gm_n6757, gm_n6758, gm_n6759, gm_n676, gm_n6760, gm_n6761, gm_n6762, gm_n6763, gm_n6764, gm_n6765, gm_n6766, gm_n6767, gm_n6768, gm_n6769, gm_n677, gm_n6770, gm_n6771, gm_n6772, gm_n6773, gm_n6774, gm_n6775, gm_n6776, gm_n6777, gm_n6778, gm_n6779, gm_n678, gm_n6780, gm_n6781, gm_n6782, gm_n6783, gm_n6784, gm_n6785, gm_n6786, gm_n6787, gm_n6788, gm_n6789, gm_n679, gm_n6790, gm_n6791, gm_n6792, gm_n6793, gm_n6794, gm_n6795, gm_n6796, gm_n6797, gm_n6798, gm_n6799, gm_n68, gm_n680, gm_n6800, gm_n6801, gm_n6802, gm_n6803, gm_n6804, gm_n6805, gm_n6806, gm_n6807, gm_n6808, gm_n6809, gm_n681, gm_n6810, gm_n6811, gm_n6812, gm_n6813, gm_n6814, gm_n6815, gm_n6816, gm_n6817, gm_n6818, gm_n6819, gm_n682, gm_n6820, gm_n6821, gm_n6822, gm_n6823, gm_n6824, gm_n6825, gm_n6826, gm_n6827, gm_n6828, gm_n6829, gm_n683, gm_n6830, gm_n6831, gm_n6832, gm_n6833, gm_n6834, gm_n6835, gm_n6836, gm_n6837, gm_n6838, gm_n6839, gm_n684, gm_n6840, gm_n6841, gm_n6842, gm_n6843, gm_n6844, gm_n6845, gm_n6846, gm_n6847, gm_n6848, gm_n6849, gm_n685, gm_n6850, gm_n6851, gm_n6853, gm_n6854, gm_n6855, gm_n6856, gm_n6857, gm_n6858, gm_n6859, gm_n686, gm_n6860, gm_n6861, gm_n6862, gm_n6863, gm_n6864, gm_n6865, gm_n6866, gm_n6867, gm_n6868, gm_n6869, gm_n687, gm_n6870, gm_n6871, gm_n6872, gm_n6873, gm_n6874, gm_n6875, gm_n6876, gm_n6877, gm_n6878, gm_n6879, gm_n688, gm_n6880, gm_n6881, gm_n6882, gm_n6883, gm_n6884, gm_n6885, gm_n6886, gm_n6887, gm_n6888, gm_n6889, gm_n689, gm_n6890, gm_n6891, gm_n6892, gm_n6893, gm_n6894, gm_n6895, gm_n6896, gm_n6897, gm_n6898, gm_n6899, gm_n69, gm_n690, gm_n6900, gm_n6901, gm_n6902, gm_n6903, gm_n6904, gm_n6905, gm_n6906, gm_n6907, gm_n6908, gm_n6909, gm_n691, gm_n6910, gm_n6911, gm_n6912, gm_n6913, gm_n6914, gm_n6915, gm_n6916, gm_n6917, gm_n6918, gm_n6919, gm_n692, gm_n6920, gm_n6921, gm_n6922, gm_n6923, gm_n6924, gm_n6925, gm_n6926, gm_n6927, gm_n6928, gm_n6929, gm_n693, gm_n6930, gm_n6931, gm_n6932, gm_n6933, gm_n6934, gm_n6935, gm_n6936, gm_n6937, gm_n6938, gm_n6939, gm_n694, gm_n6940, gm_n6941, gm_n6942, gm_n6943, gm_n6944, gm_n6945, gm_n6946, gm_n6947, gm_n6948, gm_n6949, gm_n695, gm_n6950, gm_n6951, gm_n6952, gm_n6953, gm_n6954, gm_n6955, gm_n6956, gm_n6957, gm_n6958, gm_n6959, gm_n696, gm_n6960, gm_n6961, gm_n6962, gm_n6963, gm_n6964, gm_n6965, gm_n6966, gm_n6967, gm_n6968, gm_n6969, gm_n697, gm_n6970, gm_n6971, gm_n6972, gm_n6973, gm_n6974, gm_n6975, gm_n6976, gm_n6977, gm_n6978, gm_n6979, gm_n698, gm_n6980, gm_n6981, gm_n6982, gm_n6983, gm_n6984, gm_n6985, gm_n6986, gm_n6987, gm_n6988, gm_n6989, gm_n699, gm_n6990, gm_n6991, gm_n6992, gm_n6993, gm_n6994, gm_n6995, gm_n6996, gm_n6997, gm_n6998, gm_n6999, gm_n70, gm_n700, gm_n7000, gm_n7001, gm_n7002, gm_n7003, gm_n7004, gm_n7005, gm_n7006, gm_n7007, gm_n7008, gm_n7009, gm_n701, gm_n7010, gm_n7011, gm_n7012, gm_n7013, gm_n7014, gm_n7015, gm_n7016, gm_n7017, gm_n7018, gm_n7019, gm_n702, gm_n7020, gm_n7021, gm_n7022, gm_n7023, gm_n7024, gm_n7025, gm_n7026, gm_n7027, gm_n7028, gm_n7029, gm_n703, gm_n7030, gm_n7031, gm_n7032, gm_n7033, gm_n7034, gm_n7035, gm_n7036, gm_n7037, gm_n7038, gm_n7039, gm_n704, gm_n7040, gm_n7041, gm_n7042, gm_n7043, gm_n7044, gm_n7045, gm_n7046, gm_n7047, gm_n7048, gm_n7049, gm_n705, gm_n7050, gm_n7051, gm_n7052, gm_n7053, gm_n7054, gm_n7055, gm_n7056, gm_n7057, gm_n7058, gm_n7059, gm_n706, gm_n7060, gm_n7061, gm_n7062, gm_n7063, gm_n7064, gm_n7065, gm_n7066, gm_n7067, gm_n7068, gm_n7069, gm_n707, gm_n7070, gm_n7071, gm_n7072, gm_n7073, gm_n7074, gm_n7075, gm_n7076, gm_n7077, gm_n7078, gm_n7079, gm_n708, gm_n7080, gm_n7081, gm_n7082, gm_n7083, gm_n7084, gm_n7085, gm_n7086, gm_n7087, gm_n7088, gm_n7089, gm_n709, gm_n7090, gm_n7091, gm_n7092, gm_n7093, gm_n7094, gm_n7095, gm_n7096, gm_n7097, gm_n7098, gm_n7099, gm_n71, gm_n710, gm_n7100, gm_n7101, gm_n7102, gm_n7103, gm_n7104, gm_n7105, gm_n7106, gm_n7107, gm_n7108, gm_n7109, gm_n711, gm_n7110, gm_n7111, gm_n7112, gm_n7113, gm_n7114, gm_n7115, gm_n7116, gm_n7117, gm_n7118, gm_n7119, gm_n712, gm_n7120, gm_n7121, gm_n7122, gm_n7123, gm_n7124, gm_n7125, gm_n7126, gm_n7127, gm_n7128, gm_n7129, gm_n713, gm_n7130, gm_n7131, gm_n7132, gm_n7133, gm_n7134, gm_n7135, gm_n7136, gm_n7137, gm_n7138, gm_n7139, gm_n714, gm_n7140, gm_n7141, gm_n7142, gm_n7143, gm_n7144, gm_n7145, gm_n7146, gm_n7147, gm_n7148, gm_n7149, gm_n715, gm_n7150, gm_n7151, gm_n7152, gm_n7153, gm_n7154, gm_n7155, gm_n7156, gm_n7157, gm_n7158, gm_n7159, gm_n716, gm_n7160, gm_n7161, gm_n7162, gm_n7163, gm_n7164, gm_n7165, gm_n7166, gm_n7167, gm_n7168, gm_n7169, gm_n717, gm_n7170, gm_n7171, gm_n7172, gm_n7173, gm_n7174, gm_n7175, gm_n7176, gm_n7177, gm_n7178, gm_n7179, gm_n718, gm_n7180, gm_n7181, gm_n7182, gm_n7183, gm_n7184, gm_n7185, gm_n7186, gm_n7187, gm_n7188, gm_n7189, gm_n719, gm_n7190, gm_n7191, gm_n7192, gm_n7193, gm_n7194, gm_n7195, gm_n7196, gm_n7197, gm_n7198, gm_n7199, gm_n72, gm_n720, gm_n7200, gm_n7201, gm_n7202, gm_n7203, gm_n7204, gm_n7205, gm_n7206, gm_n7207, gm_n7208, gm_n7209, gm_n721, gm_n7210, gm_n7211, gm_n7212, gm_n7213, gm_n7214, gm_n7215, gm_n7216, gm_n7217, gm_n7218, gm_n7219, gm_n722, gm_n7220, gm_n7221, gm_n7222, gm_n7223, gm_n7224, gm_n7225, gm_n7226, gm_n7227, gm_n7228, gm_n7229, gm_n723, gm_n7230, gm_n7231, gm_n7232, gm_n7233, gm_n7234, gm_n7235, gm_n7236, gm_n7237, gm_n7238, gm_n7239, gm_n724, gm_n7240, gm_n7241, gm_n7242, gm_n7243, gm_n7244, gm_n7245, gm_n7246, gm_n7247, gm_n7248, gm_n7249, gm_n725, gm_n7250, gm_n7251, gm_n7252, gm_n7253, gm_n7254, gm_n7255, gm_n7256, gm_n7257, gm_n7258, gm_n7259, gm_n726, gm_n7260, gm_n7261, gm_n7262, gm_n7263, gm_n7264, gm_n7265, gm_n7266, gm_n7267, gm_n7268, gm_n7269, gm_n727, gm_n7270, gm_n7271, gm_n7272, gm_n7273, gm_n7274, gm_n7275, gm_n7276, gm_n7277, gm_n7278, gm_n7279, gm_n728, gm_n7280, gm_n7281, gm_n7282, gm_n7283, gm_n7284, gm_n7285, gm_n7286, gm_n7287, gm_n7288, gm_n7289, gm_n729, gm_n7290, gm_n7291, gm_n7292, gm_n7293, gm_n7294, gm_n7295, gm_n7296, gm_n7297, gm_n7298, gm_n7299, gm_n73, gm_n730, gm_n7300, gm_n7301, gm_n7302, gm_n7303, gm_n7304, gm_n7305, gm_n7306, gm_n7307, gm_n7308, gm_n7309, gm_n731, gm_n7310, gm_n7311, gm_n7312, gm_n7313, gm_n7314, gm_n7315, gm_n7316, gm_n7317, gm_n7318, gm_n7319, gm_n732, gm_n7320, gm_n7321, gm_n7322, gm_n7323, gm_n7324, gm_n7325, gm_n7326, gm_n7327, gm_n7328, gm_n7329, gm_n733, gm_n7330, gm_n7331, gm_n7332, gm_n7333, gm_n7334, gm_n7335, gm_n7336, gm_n7337, gm_n7338, gm_n7339, gm_n734, gm_n7340, gm_n7341, gm_n7342, gm_n7343, gm_n7344, gm_n7345, gm_n7346, gm_n7347, gm_n7348, gm_n7349, gm_n735, gm_n7350, gm_n7351, gm_n7352, gm_n7353, gm_n7354, gm_n7355, gm_n7356, gm_n7357, gm_n7358, gm_n7359, gm_n736, gm_n7360, gm_n7361, gm_n7362, gm_n7363, gm_n7364, gm_n7365, gm_n7366, gm_n7367, gm_n7368, gm_n7369, gm_n737, gm_n7370, gm_n7371, gm_n7372, gm_n7373, gm_n7374, gm_n7375, gm_n7376, gm_n7377, gm_n7378, gm_n7379, gm_n738, gm_n7380, gm_n7381, gm_n7382, gm_n7383, gm_n7384, gm_n7385, gm_n7386, gm_n7387, gm_n7388, gm_n7389, gm_n739, gm_n7390, gm_n7391, gm_n7392, gm_n7393, gm_n7394, gm_n7395, gm_n7396, gm_n7397, gm_n7398, gm_n74, gm_n740, gm_n7400, gm_n7401, gm_n7402, gm_n7403, gm_n7404, gm_n7405, gm_n7406, gm_n7407, gm_n7408, gm_n7409, gm_n741, gm_n7410, gm_n7411, gm_n7412, gm_n7413, gm_n7414, gm_n7415, gm_n7416, gm_n7417, gm_n7418, gm_n7419, gm_n742, gm_n7420, gm_n7421, gm_n7422, gm_n7423, gm_n7424, gm_n7425, gm_n7426, gm_n7427, gm_n7428, gm_n7429, gm_n743, gm_n7430, gm_n7431, gm_n7432, gm_n7433, gm_n7434, gm_n7435, gm_n7436, gm_n7437, gm_n7438, gm_n7439, gm_n744, gm_n7440, gm_n7441, gm_n7442, gm_n7443, gm_n7444, gm_n7445, gm_n7446, gm_n7447, gm_n7448, gm_n7449, gm_n745, gm_n7450, gm_n7451, gm_n7452, gm_n7453, gm_n7454, gm_n7455, gm_n7456, gm_n7457, gm_n7458, gm_n7459, gm_n746, gm_n7460, gm_n7461, gm_n7462, gm_n7463, gm_n7464, gm_n7465, gm_n7466, gm_n7467, gm_n7468, gm_n7469, gm_n747, gm_n7470, gm_n7471, gm_n7472, gm_n7473, gm_n7474, gm_n7475, gm_n7476, gm_n7477, gm_n7478, gm_n7479, gm_n748, gm_n7480, gm_n7481, gm_n7482, gm_n7483, gm_n7484, gm_n7485, gm_n7486, gm_n7487, gm_n7488, gm_n7489, gm_n749, gm_n7490, gm_n7491, gm_n7492, gm_n7493, gm_n7494, gm_n7495, gm_n7496, gm_n7497, gm_n7498, gm_n7499, gm_n75, gm_n750, gm_n7500, gm_n7501, gm_n7502, gm_n7503, gm_n7504, gm_n7505, gm_n7506, gm_n7507, gm_n7508, gm_n7509, gm_n751, gm_n7510, gm_n7511, gm_n7512, gm_n7513, gm_n7514, gm_n7515, gm_n7516, gm_n7517, gm_n7518, gm_n7519, gm_n752, gm_n7520, gm_n7521, gm_n7522, gm_n7523, gm_n7524, gm_n7525, gm_n7526, gm_n7527, gm_n7528, gm_n7529, gm_n753, gm_n7530, gm_n7531, gm_n7532, gm_n7533, gm_n7534, gm_n7535, gm_n7536, gm_n7537, gm_n7538, gm_n7539, gm_n754, gm_n7540, gm_n7541, gm_n7542, gm_n7543, gm_n7544, gm_n7545, gm_n7546, gm_n7547, gm_n7548, gm_n7549, gm_n755, gm_n7550, gm_n7551, gm_n7552, gm_n7553, gm_n7554, gm_n7555, gm_n7556, gm_n7557, gm_n7558, gm_n7559, gm_n756, gm_n7560, gm_n7561, gm_n7562, gm_n7563, gm_n7564, gm_n7565, gm_n7566, gm_n7567, gm_n7568, gm_n7569, gm_n757, gm_n7570, gm_n7571, gm_n7572, gm_n7573, gm_n7574, gm_n7575, gm_n7576, gm_n7577, gm_n7578, gm_n7579, gm_n758, gm_n7580, gm_n7581, gm_n7582, gm_n7583, gm_n7584, gm_n7585, gm_n7586, gm_n7587, gm_n7588, gm_n7589, gm_n759, gm_n7590, gm_n7591, gm_n7592, gm_n7593, gm_n7594, gm_n7595, gm_n7596, gm_n7597, gm_n7598, gm_n7599, gm_n76, gm_n760, gm_n7600, gm_n7601, gm_n7602, gm_n7603, gm_n7604, gm_n7605, gm_n7606, gm_n7607, gm_n7608, gm_n7609, gm_n761, gm_n7610, gm_n7611, gm_n7612, gm_n7613, gm_n7614, gm_n7615, gm_n7616, gm_n7617, gm_n7618, gm_n7619, gm_n762, gm_n7620, gm_n7621, gm_n7622, gm_n7623, gm_n7624, gm_n7625, gm_n7626, gm_n7627, gm_n7628, gm_n7629, gm_n763, gm_n7630, gm_n7631, gm_n7632, gm_n7633, gm_n7634, gm_n7635, gm_n7636, gm_n7637, gm_n7638, gm_n7639, gm_n764, gm_n7640, gm_n7641, gm_n7642, gm_n7643, gm_n7644, gm_n7645, gm_n7646, gm_n7647, gm_n7648, gm_n7649, gm_n765, gm_n7650, gm_n7651, gm_n7652, gm_n7653, gm_n7654, gm_n7655, gm_n7656, gm_n7657, gm_n7658, gm_n7659, gm_n766, gm_n7660, gm_n7661, gm_n7662, gm_n7663, gm_n7664, gm_n7665, gm_n7666, gm_n7667, gm_n7668, gm_n7669, gm_n767, gm_n7670, gm_n7671, gm_n7672, gm_n7673, gm_n7674, gm_n7675, gm_n7676, gm_n7677, gm_n7678, gm_n7679, gm_n768, gm_n7680, gm_n7681, gm_n7682, gm_n7683, gm_n7684, gm_n7685, gm_n7686, gm_n7687, gm_n7688, gm_n7689, gm_n769, gm_n7690, gm_n7691, gm_n7692, gm_n7693, gm_n7694, gm_n7695, gm_n7696, gm_n7697, gm_n7698, gm_n7699, gm_n77, gm_n770, gm_n7700, gm_n7701, gm_n7702, gm_n7703, gm_n7704, gm_n7705, gm_n7706, gm_n7707, gm_n7708, gm_n7709, gm_n771, gm_n7710, gm_n7711, gm_n7712, gm_n7713, gm_n7714, gm_n7715, gm_n7716, gm_n7717, gm_n7718, gm_n7719, gm_n772, gm_n7720, gm_n7721, gm_n7722, gm_n7723, gm_n7724, gm_n7725, gm_n7726, gm_n7727, gm_n7728, gm_n7729, gm_n773, gm_n7730, gm_n7731, gm_n7732, gm_n7733, gm_n7734, gm_n7735, gm_n7736, gm_n7737, gm_n7738, gm_n7739, gm_n774, gm_n7740, gm_n7741, gm_n7742, gm_n7743, gm_n7744, gm_n7745, gm_n7746, gm_n7747, gm_n7748, gm_n7749, gm_n775, gm_n7750, gm_n7751, gm_n7752, gm_n7753, gm_n7754, gm_n7755, gm_n7756, gm_n7757, gm_n7758, gm_n7759, gm_n776, gm_n7760, gm_n7761, gm_n7762, gm_n7763, gm_n7764, gm_n7765, gm_n7766, gm_n7767, gm_n7768, gm_n7769, gm_n777, gm_n7770, gm_n7771, gm_n7772, gm_n7773, gm_n7774, gm_n7775, gm_n7776, gm_n7777, gm_n7778, gm_n7779, gm_n778, gm_n7780, gm_n7781, gm_n7782, gm_n7783, gm_n7784, gm_n7785, gm_n7786, gm_n7787, gm_n7788, gm_n7789, gm_n779, gm_n7790, gm_n7791, gm_n7792, gm_n7793, gm_n7794, gm_n7795, gm_n7796, gm_n7797, gm_n7798, gm_n7799, gm_n78, gm_n780, gm_n7800, gm_n7801, gm_n7802, gm_n7803, gm_n7804, gm_n7805, gm_n7806, gm_n7807, gm_n7808, gm_n7809, gm_n781, gm_n7810, gm_n7811, gm_n7812, gm_n7813, gm_n7814, gm_n7815, gm_n7816, gm_n7817, gm_n7818, gm_n7819, gm_n782, gm_n7820, gm_n7821, gm_n7822, gm_n7823, gm_n7824, gm_n7825, gm_n7826, gm_n7827, gm_n7828, gm_n7829, gm_n783, gm_n7830, gm_n7831, gm_n7832, gm_n7833, gm_n7834, gm_n7835, gm_n7836, gm_n7837, gm_n7838, gm_n7839, gm_n784, gm_n7840, gm_n7841, gm_n7842, gm_n7843, gm_n7844, gm_n7845, gm_n7846, gm_n7847, gm_n7848, gm_n7849, gm_n785, gm_n7850, gm_n7851, gm_n7852, gm_n7853, gm_n7854, gm_n7855, gm_n7856, gm_n7857, gm_n7858, gm_n7859, gm_n786, gm_n7860, gm_n7861, gm_n7862, gm_n7863, gm_n7864, gm_n7865, gm_n7866, gm_n7867, gm_n7868, gm_n7869, gm_n787, gm_n7870, gm_n7871, gm_n7872, gm_n7873, gm_n7874, gm_n7875, gm_n7876, gm_n7877, gm_n7878, gm_n7879, gm_n788, gm_n7880, gm_n7881, gm_n7882, gm_n7883, gm_n7884, gm_n7885, gm_n7886, gm_n7887, gm_n7888, gm_n7889, gm_n789, gm_n7890, gm_n7891, gm_n7892, gm_n7893, gm_n7894, gm_n7895, gm_n7896, gm_n7897, gm_n7898, gm_n7899, gm_n79, gm_n790, gm_n7900, gm_n7901, gm_n7902, gm_n7903, gm_n7904, gm_n7905, gm_n7906, gm_n7907, gm_n7908, gm_n7909, gm_n791, gm_n7910, gm_n7911, gm_n7912, gm_n7913, gm_n7914, gm_n7915, gm_n7916, gm_n7917, gm_n7918, gm_n7919, gm_n792, gm_n7920, gm_n7921, gm_n7922, gm_n7923, gm_n7925, gm_n7926, gm_n7927, gm_n7928, gm_n7929, gm_n793, gm_n7930, gm_n7931, gm_n7932, gm_n7933, gm_n7934, gm_n7935, gm_n7936, gm_n7937, gm_n7938, gm_n7939, gm_n794, gm_n7940, gm_n7941, gm_n7942, gm_n7943, gm_n7944, gm_n7945, gm_n7946, gm_n7947, gm_n7948, gm_n7949, gm_n795, gm_n7950, gm_n7951, gm_n7952, gm_n7953, gm_n7954, gm_n7955, gm_n7956, gm_n7957, gm_n7958, gm_n7959, gm_n796, gm_n7960, gm_n7961, gm_n7962, gm_n7963, gm_n7964, gm_n7965, gm_n7966, gm_n7967, gm_n7968, gm_n7969, gm_n797, gm_n7970, gm_n7971, gm_n7972, gm_n7973, gm_n7974, gm_n7975, gm_n7976, gm_n7977, gm_n7978, gm_n7979, gm_n798, gm_n7980, gm_n7981, gm_n7982, gm_n7983, gm_n7984, gm_n7985, gm_n7986, gm_n7987, gm_n7988, gm_n7989, gm_n799, gm_n7990, gm_n7991, gm_n7992, gm_n7993, gm_n7994, gm_n7995, gm_n7996, gm_n7997, gm_n7998, gm_n7999, gm_n80, gm_n800, gm_n8000, gm_n8001, gm_n8002, gm_n8003, gm_n8004, gm_n8005, gm_n8006, gm_n8007, gm_n8008, gm_n8009, gm_n801, gm_n8010, gm_n8011, gm_n8012, gm_n8013, gm_n8014, gm_n8015, gm_n8016, gm_n8017, gm_n8018, gm_n8019, gm_n802, gm_n8020, gm_n8021, gm_n8022, gm_n8023, gm_n8024, gm_n8025, gm_n8026, gm_n8027, gm_n8028, gm_n8029, gm_n803, gm_n8030, gm_n8031, gm_n8032, gm_n8033, gm_n8034, gm_n8035, gm_n8036, gm_n8037, gm_n8038, gm_n8039, gm_n804, gm_n8040, gm_n8041, gm_n8042, gm_n8043, gm_n8044, gm_n8045, gm_n8046, gm_n8047, gm_n8048, gm_n8049, gm_n805, gm_n8050, gm_n8051, gm_n8052, gm_n8053, gm_n8054, gm_n8055, gm_n8056, gm_n8057, gm_n8058, gm_n8059, gm_n806, gm_n8060, gm_n8061, gm_n8062, gm_n8063, gm_n8064, gm_n8065, gm_n8066, gm_n8067, gm_n8068, gm_n8069, gm_n807, gm_n8070, gm_n8071, gm_n8072, gm_n8073, gm_n8074, gm_n8075, gm_n8076, gm_n8077, gm_n8078, gm_n8079, gm_n808, gm_n8080, gm_n8081, gm_n8082, gm_n8083, gm_n8084, gm_n8085, gm_n8086, gm_n8087, gm_n8088, gm_n8089, gm_n809, gm_n8090, gm_n8091, gm_n8092, gm_n8093, gm_n8094, gm_n8095, gm_n8096, gm_n8097, gm_n8098, gm_n8099, gm_n81, gm_n810, gm_n8100, gm_n8101, gm_n8102, gm_n8103, gm_n8104, gm_n8105, gm_n8106, gm_n8107, gm_n8108, gm_n8109, gm_n811, gm_n8110, gm_n8111, gm_n8112, gm_n8113, gm_n8114, gm_n8115, gm_n8116, gm_n8117, gm_n8118, gm_n8119, gm_n812, gm_n8120, gm_n8121, gm_n8122, gm_n8123, gm_n8124, gm_n8125, gm_n8126, gm_n8127, gm_n8128, gm_n8129, gm_n813, gm_n8130, gm_n8131, gm_n8132, gm_n8133, gm_n8134, gm_n8135, gm_n8136, gm_n8137, gm_n8138, gm_n8139, gm_n814, gm_n8140, gm_n8141, gm_n8142, gm_n8143, gm_n8144, gm_n8145, gm_n8146, gm_n8147, gm_n8148, gm_n8149, gm_n815, gm_n8150, gm_n8151, gm_n8152, gm_n8153, gm_n8154, gm_n8155, gm_n8156, gm_n8157, gm_n8158, gm_n8159, gm_n816, gm_n8160, gm_n8161, gm_n8162, gm_n8163, gm_n8164, gm_n8165, gm_n8166, gm_n8167, gm_n8168, gm_n8169, gm_n817, gm_n8170, gm_n8171, gm_n8172, gm_n8173, gm_n8174, gm_n8175, gm_n8176, gm_n8177, gm_n8178, gm_n8179, gm_n818, gm_n8180, gm_n8181, gm_n8182, gm_n8183, gm_n8184, gm_n8185, gm_n8186, gm_n8187, gm_n8188, gm_n8189, gm_n819, gm_n8190, gm_n8191, gm_n8192, gm_n8193, gm_n8194, gm_n8195, gm_n8196, gm_n8197, gm_n8198, gm_n8199, gm_n82, gm_n820, gm_n8200, gm_n8201, gm_n8202, gm_n8203, gm_n8204, gm_n8205, gm_n8206, gm_n8207, gm_n8208, gm_n8209, gm_n821, gm_n8210, gm_n8211, gm_n8212, gm_n8213, gm_n8214, gm_n8215, gm_n8216, gm_n8217, gm_n8218, gm_n8219, gm_n822, gm_n8220, gm_n8221, gm_n8222, gm_n8223, gm_n8224, gm_n8225, gm_n8226, gm_n8227, gm_n8228, gm_n8229, gm_n823, gm_n8230, gm_n8231, gm_n8232, gm_n8233, gm_n8234, gm_n8235, gm_n8236, gm_n8237, gm_n8238, gm_n8239, gm_n824, gm_n8240, gm_n8241, gm_n8242, gm_n8243, gm_n8244, gm_n8245, gm_n8246, gm_n8247, gm_n8248, gm_n8249, gm_n825, gm_n8250, gm_n8251, gm_n8252, gm_n8253, gm_n8254, gm_n8255, gm_n8256, gm_n8257, gm_n8258, gm_n8259, gm_n826, gm_n8260, gm_n8261, gm_n8262, gm_n8263, gm_n8264, gm_n8265, gm_n8266, gm_n8267, gm_n8268, gm_n8269, gm_n827, gm_n8270, gm_n8271, gm_n8272, gm_n8273, gm_n8274, gm_n8275, gm_n8276, gm_n8277, gm_n8278, gm_n8279, gm_n828, gm_n8280, gm_n8281, gm_n8282, gm_n8283, gm_n8284, gm_n8285, gm_n8286, gm_n8287, gm_n8288, gm_n8289, gm_n829, gm_n8290, gm_n8291, gm_n8292, gm_n8293, gm_n8294, gm_n8295, gm_n8296, gm_n8297, gm_n8298, gm_n8299, gm_n83, gm_n830, gm_n8300, gm_n8301, gm_n8302, gm_n8303, gm_n8304, gm_n8305, gm_n8306, gm_n8307, gm_n8308, gm_n8309, gm_n831, gm_n8310, gm_n8311, gm_n8312, gm_n8313, gm_n8314, gm_n8315, gm_n8316, gm_n8317, gm_n8318, gm_n8319, gm_n832, gm_n8320, gm_n8321, gm_n8322, gm_n8323, gm_n8324, gm_n8325, gm_n8326, gm_n8327, gm_n8328, gm_n8329, gm_n833, gm_n8330, gm_n8331, gm_n8332, gm_n8333, gm_n8334, gm_n8335, gm_n8336, gm_n8337, gm_n8338, gm_n8339, gm_n8340, gm_n8341, gm_n8342, gm_n8343, gm_n8344, gm_n8345, gm_n8346, gm_n8347, gm_n8348, gm_n8349, gm_n835, gm_n8350, gm_n8351, gm_n8352, gm_n8353, gm_n8354, gm_n8355, gm_n8356, gm_n8357, gm_n8358, gm_n8359, gm_n836, gm_n8360, gm_n8361, gm_n8362, gm_n8363, gm_n8364, gm_n8365, gm_n8366, gm_n8367, gm_n8368, gm_n8369, gm_n837, gm_n8370, gm_n8371, gm_n8372, gm_n8373, gm_n8374, gm_n8375, gm_n8376, gm_n8377, gm_n8378, gm_n8379, gm_n838, gm_n8380, gm_n8381, gm_n8382, gm_n8383, gm_n8384, gm_n8385, gm_n8386, gm_n8387, gm_n8388, gm_n8389, gm_n839, gm_n8390, gm_n8391, gm_n8392, gm_n8393, gm_n8394, gm_n8395, gm_n8396, gm_n8397, gm_n8398, gm_n8399, gm_n84, gm_n840, gm_n8400, gm_n8401, gm_n8402, gm_n8403, gm_n8404, gm_n8405, gm_n8406, gm_n8407, gm_n8408, gm_n8409, gm_n841, gm_n8410, gm_n8411, gm_n8412, gm_n8413, gm_n8414, gm_n8415, gm_n8416, gm_n8417, gm_n8418, gm_n8419, gm_n842, gm_n8420, gm_n8421, gm_n8422, gm_n8423, gm_n8424, gm_n8425, gm_n8426, gm_n8427, gm_n8428, gm_n8429, gm_n843, gm_n8430, gm_n8431, gm_n8432, gm_n8433, gm_n8434, gm_n8435, gm_n8436, gm_n8437, gm_n8438, gm_n8439, gm_n844, gm_n8440, gm_n8441, gm_n8442, gm_n8443, gm_n8444, gm_n8445, gm_n8446, gm_n8447, gm_n8448, gm_n8449, gm_n845, gm_n8450, gm_n8451, gm_n8452, gm_n8454, gm_n8455, gm_n8456, gm_n8457, gm_n8458, gm_n8459, gm_n846, gm_n8460, gm_n8461, gm_n8462, gm_n8463, gm_n8464, gm_n8465, gm_n8466, gm_n8467, gm_n8468, gm_n8469, gm_n847, gm_n8470, gm_n8471, gm_n8472, gm_n8473, gm_n8474, gm_n8475, gm_n8476, gm_n8477, gm_n8478, gm_n8479, gm_n848, gm_n8480, gm_n8481, gm_n8482, gm_n8483, gm_n8484, gm_n8485, gm_n8486, gm_n8487, gm_n8488, gm_n8489, gm_n849, gm_n8490, gm_n8491, gm_n8492, gm_n8493, gm_n8494, gm_n8495, gm_n8496, gm_n8497, gm_n8498, gm_n8499, gm_n85, gm_n850, gm_n8500, gm_n8501, gm_n8502, gm_n8503, gm_n8504, gm_n8505, gm_n8506, gm_n8507, gm_n8508, gm_n8509, gm_n851, gm_n8510, gm_n8511, gm_n8512, gm_n8513, gm_n8514, gm_n8515, gm_n8516, gm_n8517, gm_n8518, gm_n8519, gm_n852, gm_n8520, gm_n8521, gm_n8522, gm_n8523, gm_n8524, gm_n8525, gm_n8526, gm_n8527, gm_n8528, gm_n8529, gm_n853, gm_n8530, gm_n8531, gm_n8532, gm_n8533, gm_n8534, gm_n8535, gm_n8536, gm_n8537, gm_n8538, gm_n8539, gm_n854, gm_n8540, gm_n8541, gm_n8542, gm_n8543, gm_n8544, gm_n8545, gm_n8546, gm_n8547, gm_n8548, gm_n8549, gm_n855, gm_n8550, gm_n8551, gm_n8552, gm_n8553, gm_n8554, gm_n8555, gm_n8556, gm_n8557, gm_n8558, gm_n8559, gm_n856, gm_n8560, gm_n8561, gm_n8562, gm_n8563, gm_n8564, gm_n8565, gm_n8566, gm_n8567, gm_n8568, gm_n8569, gm_n857, gm_n8570, gm_n8571, gm_n8572, gm_n8573, gm_n8574, gm_n8575, gm_n8576, gm_n8577, gm_n8578, gm_n8579, gm_n858, gm_n8580, gm_n8581, gm_n8582, gm_n8583, gm_n8584, gm_n8585, gm_n8586, gm_n8587, gm_n8588, gm_n8589, gm_n859, gm_n8590, gm_n8591, gm_n8592, gm_n8593, gm_n8594, gm_n8595, gm_n8596, gm_n8597, gm_n8598, gm_n8599, gm_n86, gm_n860, gm_n8600, gm_n8601, gm_n8602, gm_n8603, gm_n8604, gm_n8605, gm_n8606, gm_n8607, gm_n8608, gm_n8609, gm_n861, gm_n8610, gm_n8611, gm_n8612, gm_n8613, gm_n8614, gm_n8615, gm_n8616, gm_n8617, gm_n8618, gm_n8619, gm_n862, gm_n8620, gm_n8621, gm_n8622, gm_n8623, gm_n8624, gm_n8625, gm_n8626, gm_n8627, gm_n8628, gm_n8629, gm_n863, gm_n8630, gm_n8631, gm_n8632, gm_n8633, gm_n8634, gm_n8635, gm_n8636, gm_n8637, gm_n8638, gm_n8639, gm_n864, gm_n8640, gm_n8641, gm_n8642, gm_n8643, gm_n8644, gm_n8645, gm_n8646, gm_n8647, gm_n8648, gm_n8649, gm_n865, gm_n8650, gm_n8651, gm_n8652, gm_n8653, gm_n8654, gm_n8655, gm_n8656, gm_n8657, gm_n8658, gm_n8659, gm_n866, gm_n8660, gm_n8661, gm_n8662, gm_n8663, gm_n8664, gm_n8665, gm_n8666, gm_n8667, gm_n8668, gm_n8669, gm_n867, gm_n8670, gm_n8671, gm_n8672, gm_n8673, gm_n8674, gm_n8675, gm_n8676, gm_n8677, gm_n8678, gm_n8679, gm_n868, gm_n8680, gm_n8681, gm_n8682, gm_n8683, gm_n8684, gm_n8685, gm_n8686, gm_n8687, gm_n8688, gm_n8689, gm_n869, gm_n8690, gm_n8691, gm_n8692, gm_n8693, gm_n8694, gm_n8695, gm_n8696, gm_n8697, gm_n8698, gm_n8699, gm_n87, gm_n870, gm_n8700, gm_n8701, gm_n8702, gm_n8703, gm_n8704, gm_n8705, gm_n8706, gm_n8707, gm_n8708, gm_n8709, gm_n871, gm_n8710, gm_n8711, gm_n8712, gm_n8713, gm_n8714, gm_n8715, gm_n8716, gm_n8717, gm_n8718, gm_n8719, gm_n872, gm_n8720, gm_n8721, gm_n8722, gm_n8723, gm_n8724, gm_n8725, gm_n8726, gm_n8727, gm_n8728, gm_n8729, gm_n873, gm_n8730, gm_n8731, gm_n8732, gm_n8733, gm_n8734, gm_n8735, gm_n8736, gm_n8737, gm_n8738, gm_n8739, gm_n874, gm_n8740, gm_n8741, gm_n8742, gm_n8743, gm_n8744, gm_n8745, gm_n8746, gm_n8747, gm_n8748, gm_n8749, gm_n875, gm_n8750, gm_n8751, gm_n8752, gm_n8753, gm_n8754, gm_n8755, gm_n8756, gm_n8757, gm_n8758, gm_n8759, gm_n876, gm_n8760, gm_n8761, gm_n8762, gm_n8763, gm_n8764, gm_n8765, gm_n8766, gm_n8767, gm_n8768, gm_n8769, gm_n877, gm_n8770, gm_n8771, gm_n8772, gm_n8773, gm_n8774, gm_n8775, gm_n8776, gm_n8777, gm_n8778, gm_n8779, gm_n878, gm_n8780, gm_n8781, gm_n8782, gm_n8783, gm_n8784, gm_n8785, gm_n8786, gm_n8787, gm_n8788, gm_n8789, gm_n879, gm_n8790, gm_n8791, gm_n8792, gm_n8793, gm_n8794, gm_n8795, gm_n8796, gm_n8797, gm_n8798, gm_n8799, gm_n88, gm_n880, gm_n8800, gm_n8801, gm_n8802, gm_n8803, gm_n8804, gm_n8805, gm_n8806, gm_n8807, gm_n8808, gm_n8809, gm_n881, gm_n8810, gm_n8811, gm_n8812, gm_n8813, gm_n8814, gm_n8815, gm_n8816, gm_n8817, gm_n8818, gm_n8819, gm_n882, gm_n8820, gm_n8821, gm_n8822, gm_n8823, gm_n8824, gm_n8825, gm_n8826, gm_n8827, gm_n8828, gm_n8829, gm_n883, gm_n8830, gm_n8831, gm_n8832, gm_n8833, gm_n8834, gm_n8835, gm_n8836, gm_n8837, gm_n8838, gm_n8839, gm_n884, gm_n8840, gm_n8841, gm_n8842, gm_n8843, gm_n8844, gm_n8845, gm_n8846, gm_n8847, gm_n8848, gm_n8849, gm_n885, gm_n8850, gm_n8851, gm_n8852, gm_n8853, gm_n8854, gm_n8855, gm_n8856, gm_n8857, gm_n8858, gm_n8859, gm_n886, gm_n8860, gm_n8861, gm_n8862, gm_n8863, gm_n8864, gm_n8865, gm_n8866, gm_n8867, gm_n8868, gm_n8869, gm_n887, gm_n8870, gm_n8871, gm_n8872, gm_n8873, gm_n8874, gm_n8875, gm_n8876, gm_n8877, gm_n8878, gm_n8879, gm_n888, gm_n8880, gm_n8881, gm_n8882, gm_n8883, gm_n8884, gm_n8885, gm_n8886, gm_n8887, gm_n8888, gm_n8889, gm_n889, gm_n8890, gm_n8891, gm_n8892, gm_n8893, gm_n8894, gm_n8895, gm_n8896, gm_n8897, gm_n8898, gm_n8899, gm_n89, gm_n890, gm_n8900, gm_n8901, gm_n8902, gm_n8903, gm_n8904, gm_n8905, gm_n8906, gm_n8907, gm_n8908, gm_n8909, gm_n891, gm_n8910, gm_n8911, gm_n8912, gm_n8913, gm_n8914, gm_n8915, gm_n8916, gm_n8917, gm_n8918, gm_n8919, gm_n892, gm_n8920, gm_n8921, gm_n8922, gm_n8923, gm_n8924, gm_n8925, gm_n8926, gm_n8927, gm_n8928, gm_n8929, gm_n893, gm_n8930, gm_n8931, gm_n8932, gm_n8933, gm_n8934, gm_n8935, gm_n8936, gm_n8937, gm_n8938, gm_n8939, gm_n894, gm_n8940, gm_n8941, gm_n8942, gm_n8943, gm_n8944, gm_n8945, gm_n8946, gm_n8947, gm_n8948, gm_n8949, gm_n895, gm_n8950, gm_n8951, gm_n8952, gm_n8953, gm_n8954, gm_n8955, gm_n8956, gm_n8957, gm_n8958, gm_n8959, gm_n896, gm_n8960, gm_n8961, gm_n8962, gm_n8963, gm_n8964, gm_n8965, gm_n8966, gm_n8967, gm_n8968, gm_n897, gm_n8970, gm_n8971, gm_n8972, gm_n8973, gm_n8974, gm_n8975, gm_n8976, gm_n8977, gm_n8978, gm_n8979, gm_n898, gm_n8980, gm_n8981, gm_n8982, gm_n8983, gm_n8984, gm_n8985, gm_n8986, gm_n8987, gm_n8988, gm_n8989, gm_n899, gm_n8990, gm_n8991, gm_n8992, gm_n8993, gm_n8994, gm_n8995, gm_n8996, gm_n8997, gm_n8998, gm_n8999, gm_n90, gm_n900, gm_n9000, gm_n9001, gm_n9002, gm_n9003, gm_n9004, gm_n9005, gm_n9006, gm_n9007, gm_n9008, gm_n9009, gm_n901, gm_n9010, gm_n9011, gm_n9012, gm_n9013, gm_n9014, gm_n9015, gm_n9016, gm_n9017, gm_n9018, gm_n9019, gm_n902, gm_n9020, gm_n9021, gm_n9022, gm_n9023, gm_n9024, gm_n9025, gm_n9026, gm_n9027, gm_n9028, gm_n9029, gm_n903, gm_n9030, gm_n9031, gm_n9032, gm_n9033, gm_n9034, gm_n9035, gm_n9036, gm_n9037, gm_n9038, gm_n9039, gm_n904, gm_n9040, gm_n9041, gm_n9042, gm_n9043, gm_n9044, gm_n9045, gm_n9046, gm_n9047, gm_n9048, gm_n9049, gm_n905, gm_n9050, gm_n9051, gm_n9052, gm_n9053, gm_n9054, gm_n9055, gm_n9056, gm_n9057, gm_n9058, gm_n9059, gm_n906, gm_n9060, gm_n9061, gm_n9062, gm_n9063, gm_n9064, gm_n9065, gm_n9066, gm_n9067, gm_n9068, gm_n9069, gm_n907, gm_n9070, gm_n9071, gm_n9072, gm_n9073, gm_n9074, gm_n9075, gm_n9076, gm_n9077, gm_n9078, gm_n9079, gm_n908, gm_n9080, gm_n9081, gm_n9082, gm_n9083, gm_n9084, gm_n9085, gm_n9086, gm_n9087, gm_n9088, gm_n9089, gm_n909, gm_n9090, gm_n9091, gm_n9092, gm_n9093, gm_n9094, gm_n9095, gm_n9096, gm_n9097, gm_n9098, gm_n9099, gm_n91, gm_n910, gm_n9100, gm_n9101, gm_n9102, gm_n9103, gm_n9104, gm_n9105, gm_n9106, gm_n9107, gm_n9108, gm_n9109, gm_n911, gm_n9110, gm_n9111, gm_n9112, gm_n9113, gm_n9114, gm_n9115, gm_n9116, gm_n9117, gm_n9118, gm_n9119, gm_n912, gm_n9120, gm_n9121, gm_n9122, gm_n9123, gm_n9124, gm_n9125, gm_n9126, gm_n9127, gm_n9128, gm_n9129, gm_n913, gm_n9130, gm_n9131, gm_n9132, gm_n9133, gm_n9134, gm_n9135, gm_n9136, gm_n9137, gm_n9138, gm_n9139, gm_n914, gm_n9140, gm_n9141, gm_n9142, gm_n9143, gm_n9144, gm_n9145, gm_n9146, gm_n9147, gm_n9148, gm_n9149, gm_n915, gm_n9150, gm_n9151, gm_n9152, gm_n9153, gm_n9154, gm_n9155, gm_n9156, gm_n9157, gm_n9158, gm_n9159, gm_n916, gm_n9160, gm_n9161, gm_n9162, gm_n9163, gm_n9164, gm_n9165, gm_n9166, gm_n9167, gm_n9168, gm_n9169, gm_n917, gm_n9170, gm_n9171, gm_n9172, gm_n9173, gm_n9174, gm_n9175, gm_n9176, gm_n9177, gm_n9178, gm_n9179, gm_n918, gm_n9180, gm_n9181, gm_n9182, gm_n9183, gm_n9184, gm_n9185, gm_n9186, gm_n9187, gm_n9188, gm_n9189, gm_n919, gm_n9190, gm_n9191, gm_n9192, gm_n9193, gm_n9194, gm_n9195, gm_n9196, gm_n9197, gm_n9198, gm_n9199, gm_n92, gm_n920, gm_n9200, gm_n9201, gm_n9202, gm_n9203, gm_n9204, gm_n9205, gm_n9206, gm_n9207, gm_n9208, gm_n9209, gm_n921, gm_n9210, gm_n9211, gm_n9212, gm_n9213, gm_n9214, gm_n9215, gm_n9216, gm_n9217, gm_n9218, gm_n9219, gm_n922, gm_n9220, gm_n9221, gm_n9222, gm_n9223, gm_n9224, gm_n9225, gm_n9226, gm_n9227, gm_n9228, gm_n9229, gm_n923, gm_n9230, gm_n9231, gm_n9232, gm_n9233, gm_n9234, gm_n9235, gm_n9236, gm_n9237, gm_n9238, gm_n9239, gm_n924, gm_n9240, gm_n9241, gm_n9242, gm_n9243, gm_n9244, gm_n9245, gm_n9246, gm_n9247, gm_n9248, gm_n9249, gm_n925, gm_n9250, gm_n9251, gm_n9252, gm_n9253, gm_n9254, gm_n9255, gm_n9256, gm_n9257, gm_n9258, gm_n9259, gm_n926, gm_n9260, gm_n9261, gm_n9262, gm_n9263, gm_n9264, gm_n9265, gm_n9266, gm_n9267, gm_n9268, gm_n9269, gm_n927, gm_n9270, gm_n9271, gm_n9272, gm_n9273, gm_n9274, gm_n9275, gm_n9276, gm_n9277, gm_n9278, gm_n9279, gm_n928, gm_n9280, gm_n9281, gm_n9282, gm_n9283, gm_n9284, gm_n9285, gm_n9286, gm_n9287, gm_n9288, gm_n9289, gm_n929, gm_n9290, gm_n9291, gm_n9292, gm_n9293, gm_n9294, gm_n9295, gm_n9296, gm_n9297, gm_n9298, gm_n9299, gm_n93, gm_n930, gm_n9300, gm_n9301, gm_n9302, gm_n9303, gm_n9304, gm_n9305, gm_n9306, gm_n9307, gm_n9308, gm_n9309, gm_n931, gm_n9310, gm_n9311, gm_n9312, gm_n9313, gm_n9314, gm_n9315, gm_n9316, gm_n9317, gm_n9318, gm_n9319, gm_n932, gm_n9320, gm_n9321, gm_n9322, gm_n9323, gm_n9324, gm_n9325, gm_n9326, gm_n9327, gm_n9328, gm_n9329, gm_n933, gm_n9330, gm_n9331, gm_n9332, gm_n9333, gm_n9334, gm_n9335, gm_n9336, gm_n9337, gm_n9338, gm_n9339, gm_n934, gm_n9340, gm_n9341, gm_n9342, gm_n9343, gm_n9344, gm_n9345, gm_n9346, gm_n9347, gm_n9348, gm_n9349, gm_n935, gm_n9350, gm_n9351, gm_n9352, gm_n9353, gm_n9354, gm_n9355, gm_n9356, gm_n9357, gm_n9358, gm_n9359, gm_n936, gm_n9360, gm_n9361, gm_n9362, gm_n9363, gm_n9364, gm_n9365, gm_n9366, gm_n9367, gm_n9368, gm_n9369, gm_n937, gm_n9370, gm_n9371, gm_n9372, gm_n9373, gm_n9374, gm_n9375, gm_n9376, gm_n9377, gm_n9378, gm_n9379, gm_n938, gm_n9380, gm_n9381, gm_n9382, gm_n9383, gm_n9384, gm_n9385, gm_n9386, gm_n9387, gm_n9388, gm_n9389, gm_n939, gm_n9390, gm_n9391, gm_n9392, gm_n9393, gm_n9394, gm_n9395, gm_n9396, gm_n9397, gm_n9398, gm_n9399, gm_n94, gm_n940, gm_n9400, gm_n9401, gm_n9402, gm_n9403, gm_n9404, gm_n9405, gm_n9406, gm_n9407, gm_n9408, gm_n9409, gm_n941, gm_n9410, gm_n9411, gm_n9412, gm_n9413, gm_n9414, gm_n9415, gm_n9416, gm_n9417, gm_n9418, gm_n9419, gm_n942, gm_n9420, gm_n9421, gm_n9422, gm_n9423, gm_n9424, gm_n9425, gm_n9426, gm_n9427, gm_n9428, gm_n9429, gm_n943, gm_n9430, gm_n9431, gm_n9432, gm_n9433, gm_n9434, gm_n9435, gm_n9436, gm_n9437, gm_n9438, gm_n9439, gm_n944, gm_n9440, gm_n9441, gm_n9442, gm_n9443, gm_n9444, gm_n9445, gm_n9446, gm_n9447, gm_n9448, gm_n9449, gm_n945, gm_n9450, gm_n9451, gm_n9452, gm_n9453, gm_n9454, gm_n9455, gm_n9456, gm_n9457, gm_n9458, gm_n9459, gm_n946, gm_n9460, gm_n9461, gm_n9462, gm_n9463, gm_n9464, gm_n9465, gm_n9466, gm_n9467, gm_n9468, gm_n9469, gm_n947, gm_n9470, gm_n9471, gm_n9472, gm_n9473, gm_n9474, gm_n9475, gm_n9476, gm_n9477, gm_n9478, gm_n9479, gm_n948, gm_n9481, gm_n9482, gm_n9483, gm_n9484, gm_n9485, gm_n9486, gm_n9487, gm_n9488, gm_n9489, gm_n949, gm_n9490, gm_n9491, gm_n9492, gm_n9493, gm_n9494, gm_n9495, gm_n9496, gm_n9497, gm_n9498, gm_n9499, gm_n95, gm_n950, gm_n9500, gm_n9501, gm_n9502, gm_n9503, gm_n9504, gm_n9505, gm_n9506, gm_n9507, gm_n9508, gm_n9509, gm_n951, gm_n9510, gm_n9511, gm_n9512, gm_n9513, gm_n9514, gm_n9515, gm_n9516, gm_n9517, gm_n9518, gm_n9519, gm_n952, gm_n9520, gm_n9521, gm_n9522, gm_n9523, gm_n9524, gm_n9525, gm_n9526, gm_n9527, gm_n9528, gm_n9529, gm_n953, gm_n9530, gm_n9531, gm_n9532, gm_n9533, gm_n9534, gm_n9535, gm_n9536, gm_n9537, gm_n9538, gm_n9539, gm_n954, gm_n9540, gm_n9541, gm_n9542, gm_n9543, gm_n9544, gm_n9545, gm_n9546, gm_n9547, gm_n9548, gm_n9549, gm_n955, gm_n9550, gm_n9551, gm_n9552, gm_n9553, gm_n9554, gm_n9555, gm_n9556, gm_n9557, gm_n9558, gm_n9559, gm_n956, gm_n9560, gm_n9561, gm_n9562, gm_n9563, gm_n9564, gm_n9565, gm_n9566, gm_n9567, gm_n9568, gm_n9569, gm_n957, gm_n9570, gm_n9571, gm_n9572, gm_n9573, gm_n9574, gm_n9575, gm_n9576, gm_n9577, gm_n9578, gm_n9579, gm_n958, gm_n9580, gm_n9581, gm_n9582, gm_n9583, gm_n9584, gm_n9585, gm_n9586, gm_n9587, gm_n9588, gm_n9589, gm_n959, gm_n9590, gm_n9591, gm_n9592, gm_n9593, gm_n9594, gm_n9595, gm_n9596, gm_n9597, gm_n9598, gm_n9599, gm_n96, gm_n960, gm_n9600, gm_n9601, gm_n9602, gm_n9603, gm_n9604, gm_n9605, gm_n9606, gm_n9607, gm_n9608, gm_n9609, gm_n961, gm_n9610, gm_n9611, gm_n9612, gm_n9613, gm_n9614, gm_n9615, gm_n9616, gm_n9617, gm_n9618, gm_n9619, gm_n962, gm_n9620, gm_n9621, gm_n9622, gm_n9623, gm_n9624, gm_n9625, gm_n9626, gm_n9627, gm_n9628, gm_n9629, gm_n963, gm_n9630, gm_n9631, gm_n9632, gm_n9633, gm_n9634, gm_n9635, gm_n9636, gm_n9637, gm_n9638, gm_n9639, gm_n964, gm_n9640, gm_n9641, gm_n9642, gm_n9643, gm_n9644, gm_n9645, gm_n9646, gm_n9647, gm_n9648, gm_n9649, gm_n965, gm_n9650, gm_n9651, gm_n9652, gm_n9653, gm_n9654, gm_n9655, gm_n9656, gm_n9657, gm_n9658, gm_n9659, gm_n966, gm_n9660, gm_n9661, gm_n9662, gm_n9663, gm_n9664, gm_n9665, gm_n9666, gm_n9667, gm_n9668, gm_n9669, gm_n967, gm_n9670, gm_n9671, gm_n9672, gm_n9673, gm_n9674, gm_n9675, gm_n9676, gm_n9677, gm_n9678, gm_n9679, gm_n968, gm_n9680, gm_n9681, gm_n9682, gm_n9683, gm_n9684, gm_n9685, gm_n9686, gm_n9687, gm_n9688, gm_n9689, gm_n969, gm_n9690, gm_n9691, gm_n9692, gm_n9693, gm_n9694, gm_n9695, gm_n9696, gm_n9697, gm_n9698, gm_n9699, gm_n97, gm_n970, gm_n9700, gm_n9701, gm_n9702, gm_n9703, gm_n9704, gm_n9705, gm_n9706, gm_n9707, gm_n9708, gm_n9709, gm_n971, gm_n9710, gm_n9711, gm_n9712, gm_n9713, gm_n9714, gm_n9715, gm_n9716, gm_n9717, gm_n9718, gm_n9719, gm_n972, gm_n9720, gm_n9721, gm_n9722, gm_n9723, gm_n9724, gm_n9725, gm_n9726, gm_n9727, gm_n9728, gm_n9729, gm_n973, gm_n9730, gm_n9731, gm_n9732, gm_n9733, gm_n9734, gm_n9735, gm_n9736, gm_n9737, gm_n9738, gm_n9739, gm_n974, gm_n9740, gm_n9741, gm_n9742, gm_n9743, gm_n9744, gm_n9745, gm_n9746, gm_n9747, gm_n9748, gm_n9749, gm_n975, gm_n9750, gm_n9751, gm_n9752, gm_n9753, gm_n9754, gm_n9755, gm_n9756, gm_n9757, gm_n9758, gm_n9759, gm_n976, gm_n9760, gm_n9761, gm_n9762, gm_n9763, gm_n9764, gm_n9765, gm_n9766, gm_n9767, gm_n9768, gm_n9769, gm_n977, gm_n9770, gm_n9771, gm_n9772, gm_n9773, gm_n9774, gm_n9775, gm_n9776, gm_n9777, gm_n9778, gm_n9779, gm_n978, gm_n9780, gm_n9781, gm_n9782, gm_n9783, gm_n9784, gm_n9785, gm_n9786, gm_n9787, gm_n9788, gm_n9789, gm_n979, gm_n9790, gm_n9791, gm_n9792, gm_n9793, gm_n9794, gm_n9795, gm_n9796, gm_n9797, gm_n9798, gm_n9799, gm_n98, gm_n980, gm_n9800, gm_n9801, gm_n9802, gm_n9803, gm_n9804, gm_n9805, gm_n9806, gm_n9807, gm_n9808, gm_n9809, gm_n981, gm_n9810, gm_n9811, gm_n9812, gm_n9813, gm_n9814, gm_n9815, gm_n9816, gm_n9817, gm_n9818, gm_n9819, gm_n982, gm_n9820, gm_n9821, gm_n9822, gm_n9823, gm_n9824, gm_n9825, gm_n9826, gm_n9827, gm_n9828, gm_n9829, gm_n983, gm_n9830, gm_n9831, gm_n9832, gm_n9833, gm_n9834, gm_n9835, gm_n9836, gm_n9837, gm_n9838, gm_n9839, gm_n984, gm_n9840, gm_n9841, gm_n9842, gm_n9843, gm_n9844, gm_n9845, gm_n9846, gm_n9847, gm_n9848, gm_n9849, gm_n985, gm_n9850, gm_n9851, gm_n9852, gm_n9853, gm_n9854, gm_n9855, gm_n9856, gm_n9857, gm_n9858, gm_n9859, gm_n986, gm_n9860, gm_n9861, gm_n9862, gm_n9863, gm_n9864, gm_n9865, gm_n9866, gm_n9867, gm_n9868, gm_n9869, gm_n987, gm_n9870, gm_n9871, gm_n9872, gm_n9873, gm_n9874, gm_n9875, gm_n9876, gm_n9877, gm_n9878, gm_n9879, gm_n988, gm_n9880, gm_n9881, gm_n9882, gm_n9883, gm_n9884, gm_n9885, gm_n9886, gm_n9887, gm_n9888, gm_n9889, gm_n989, gm_n9890, gm_n9891, gm_n9892, gm_n9893, gm_n9894, gm_n9895, gm_n9896, gm_n9897, gm_n9898, gm_n9899, gm_n99, gm_n990, gm_n9900, gm_n9901, gm_n9902, gm_n9903, gm_n9904, gm_n9905, gm_n9906, gm_n9907, gm_n9908, gm_n9909, gm_n991, gm_n9910, gm_n9911, gm_n9912, gm_n9913, gm_n9914, gm_n9915, gm_n9916, gm_n9917, gm_n9918, gm_n9919, gm_n992, gm_n9920, gm_n9921, gm_n9922, gm_n9923, gm_n9924, gm_n9925, gm_n9926, gm_n9927, gm_n9928, gm_n9929, gm_n993, gm_n9930, gm_n9931, gm_n9932, gm_n9933, gm_n9934, gm_n9935, gm_n9936, gm_n9937, gm_n9938, gm_n9939, gm_n994, gm_n9940, gm_n9941, gm_n9942, gm_n9943, gm_n9944, gm_n9945, gm_n9946, gm_n9947, gm_n9948, gm_n9949, gm_n995, gm_n9950, gm_n9951, gm_n9952, gm_n9953, gm_n9954, gm_n9955, gm_n9956, gm_n9957, gm_n9958, gm_n9959, gm_n996, gm_n9960, gm_n9961, gm_n9962, gm_n9963, gm_n9964, gm_n9965, gm_n9966, gm_n9967, gm_n9968, gm_n9969, gm_n997, gm_n9970, gm_n9971, gm_n9972, gm_n9973, gm_n9974, gm_n9975, gm_n9976, gm_n9977, gm_n9978, gm_n9979, gm_n998, gm_n9980, gm_n9981, gm_n9982, gm_n9983, gm_n9984, gm_n9985, gm_n9986, gm_n9987, gm_n9988, gm_n9989, gm_n999, gm_n9990, gm_n9991, gm_n9992, gm_n9993, gm_n9995, gm_n9996, gm_n9997, gm_n9998, gm_n9999;
	not (gm_n45, in_20);
	not (gm_n46, in_16);
	not (gm_n47, in_18);
	not (gm_n48, in_12);
	not (gm_n49, in_13);
	not (gm_n50, in_14);
	not (gm_n51, in_9);
	not (gm_n52, in_10);
	not (gm_n53, in_11);
	not (gm_n54, in_4);
	not (gm_n55, in_7);
	or (gm_n56, in_2, in_1, in_0, in_3);
	nor (gm_n57, in_6, in_5, gm_n54, gm_n56, gm_n55);
	and (gm_n58, gm_n52, gm_n51, in_8, gm_n57, gm_n53);
	and (gm_n59, gm_n50, gm_n49, gm_n48, gm_n58, in_15);
	nand (gm_n60, gm_n47, in_17, gm_n46, gm_n59, in_19);
	nor (gm_n61, gm_n60, in_21, gm_n45);
	not (gm_n62, in_19);
	not (gm_n63, in_15);
	not (gm_n64, in_8);
	nand (gm_n65, in_2, in_1, in_0);
	nor (gm_n66, in_5, in_4, in_3, gm_n65, in_6);
	and (gm_n67, gm_n51, gm_n64, in_7, gm_n66, gm_n52);
	nand (gm_n68, in_13, gm_n48, gm_n53, gm_n67, gm_n50);
	nor (gm_n69, in_17, gm_n46, gm_n63, gm_n68, in_18);
	nand (gm_n70, in_21, gm_n45, gm_n62, gm_n69);
	not (gm_n71, in_21);
	not (gm_n72, in_5);
	not (gm_n73, in_0);
	not (gm_n74, in_3);
	nand (gm_n75, in_2, in_1, gm_n73, gm_n54, gm_n74);
	nor (gm_n76, gm_n55, in_6, gm_n72, gm_n75, gm_n64);
	and (gm_n77, gm_n53, gm_n52, in_9, gm_n76, in_12);
	nand (gm_n78, gm_n63, in_14, gm_n49, gm_n77, in_16);
	nor (gm_n79, gm_n62, in_18, in_17, gm_n78, in_20);
	nand (gm_n80, gm_n79, gm_n71);
	not (gm_n81, in_17);
	not (gm_n82, in_6);
	nor (gm_n83, in_2, in_1, in_0);
	nand (gm_n84, in_5, in_4, in_3, gm_n83, gm_n82);
	nor (gm_n85, gm_n51, gm_n64, gm_n55, gm_n84, gm_n52);
	nand (gm_n86, in_13, gm_n48, gm_n53, gm_n85, gm_n50);
	nor (gm_n87, gm_n81, gm_n46, in_15, gm_n86, in_18);
	nand (gm_n88, in_21, in_20, in_19, gm_n87);
	nor (gm_n89, in_2, in_1, gm_n73, gm_n54, gm_n74);
	nand (gm_n90, in_7, in_6, in_5, gm_n89, in_8);
	nor (gm_n91, gm_n53, in_10, gm_n51, gm_n90, in_12);
	nand (gm_n92, in_15, gm_n50, gm_n49, gm_n91, gm_n46);
	nor (gm_n93, gm_n62, in_18, gm_n81, gm_n92, in_20);
	nand (gm_n94, gm_n93, gm_n71);
	nor (gm_n95, in_1, in_0);
	nand (gm_n96, in_4, in_3, in_2, gm_n95, in_5);
	or (gm_n97, gm_n64, in_7, in_6, gm_n96, gm_n51);
	nor (gm_n98, gm_n48, in_11, gm_n52, gm_n97, gm_n49);
	nand (gm_n99, in_16, gm_n63, gm_n50, gm_n98, in_17);
	nor (gm_n100, gm_n45, gm_n62, in_18, gm_n99, gm_n71);
	not (gm_n101, in_2);
	and (gm_n102, in_1, in_0);
	nand (gm_n103, in_4, gm_n74, gm_n101, gm_n102, in_5);
	or (gm_n104, gm_n64, in_7, in_6, gm_n103, in_9);
	nor (gm_n105, gm_n48, in_11, gm_n52, gm_n104, in_13);
	nand (gm_n106, gm_n46, gm_n63, gm_n50, gm_n105, in_17);
	nor (gm_n107, gm_n45, in_19, in_18, gm_n106, in_21);
	nand (gm_n108, in_2, in_1, in_0, in_4, in_3);
	nor (gm_n109, gm_n55, in_6, gm_n72, gm_n108, in_8);
	nand (gm_n110, gm_n53, gm_n52, in_9, gm_n109, in_12);
	nor (gm_n111, gm_n63, in_14, gm_n49, gm_n110, in_16);
	nand (gm_n112, in_19, gm_n47, in_17, gm_n111, gm_n45);
	nor (gm_n113, gm_n112, gm_n71);
	nor (gm_n114, in_7, in_6, in_5, gm_n108, gm_n64);
	nand (gm_n115, in_11, in_10, gm_n51, gm_n114, gm_n48);
	nor (gm_n116, gm_n63, in_14, gm_n49, gm_n115);
	nand (gm_n117, in_18, in_17, gm_n46, gm_n116, in_19);
	nor (gm_n118, gm_n117, in_21, gm_n45);
	nand (gm_n119, in_4, in_3, gm_n101, gm_n102, gm_n72);
	nor (gm_n120, in_8, in_7, gm_n82, gm_n119, gm_n51);
	nand (gm_n121, in_12, gm_n53, gm_n52, gm_n120, in_13);
	nor (gm_n122, gm_n46, in_15, in_14, gm_n121, gm_n81);
	nand (gm_n123, in_20, in_19, gm_n47, gm_n122, gm_n71);
	nand (gm_n124, gm_n101, in_1, gm_n73, in_4, in_3);
	nor (gm_n125, gm_n55, gm_n82, in_5, gm_n124, gm_n64);
	nand (gm_n126, gm_n53, in_10, in_9, gm_n125, gm_n48);
	nor (gm_n127, in_15, in_14, gm_n49, gm_n126);
	and (gm_n128, in_18, gm_n81, gm_n46, gm_n127, gm_n62);
	nand (gm_n129, gm_n128, gm_n71, gm_n45);
	or (gm_n130, in_2, in_1, in_0, in_4, in_3);
	or (gm_n131, gm_n55, in_6, in_5, gm_n130, in_8);
	nor (gm_n132, in_11, gm_n52, in_9, gm_n131, in_12);
	nand (gm_n133, gm_n63, gm_n50, gm_n49, gm_n132, gm_n46);
	nor (gm_n134, gm_n62, gm_n47, in_17, gm_n133, in_20);
	nand (gm_n135, gm_n134, gm_n71);
	nor (gm_n136, in_5, gm_n54, in_3, gm_n65, gm_n82);
	and (gm_n137, in_9, gm_n64, gm_n55, gm_n136, in_10);
	nand (gm_n138, in_13, in_12, in_11, gm_n137, in_14);
	nor (gm_n139, in_17, in_16, gm_n63, gm_n138, in_18);
	nand (gm_n140, in_21, in_20, gm_n62, gm_n139);
	nand (gm_n141, gm_n54, gm_n74, in_2, gm_n95, in_5);
	nor (gm_n142, in_8, gm_n55, in_6, gm_n141, in_9);
	and (gm_n143, gm_n48, in_11, in_10, gm_n142, in_13);
	nand (gm_n144, in_16, in_15, in_14, gm_n143, in_17);
	nor (gm_n145, gm_n45, gm_n62, in_18, gm_n144, gm_n71);
	nor (gm_n146, gm_n64, in_7, in_6, gm_n141, gm_n51);
	and (gm_n147, gm_n48, gm_n53, gm_n52, gm_n146, gm_n49);
	nand (gm_n148, gm_n46, in_15, gm_n50, gm_n147, in_17);
	nor (gm_n149, gm_n45, in_19, in_18, gm_n148, gm_n71);
	or (gm_n150, in_2, in_1, in_0);
	nor (gm_n151, in_5, in_4, gm_n74, gm_n150, gm_n82);
	nand (gm_n152, gm_n51, gm_n64, in_7, gm_n151, gm_n52);
	nor (gm_n153, in_13, gm_n48, in_11, gm_n152, gm_n50);
	nand (gm_n154, gm_n81, gm_n46, in_15, gm_n153, gm_n47);
	nor (gm_n155, gm_n71, in_20, in_19, gm_n154);
	nand (gm_n156, gm_n54, in_3, gm_n101, gm_n102, gm_n72);
	nor (gm_n157, gm_n64, in_7, in_6, gm_n156, gm_n51);
	and (gm_n158, in_12, gm_n53, gm_n52, gm_n157, in_13);
	nand (gm_n159, gm_n46, in_15, gm_n50, gm_n158, in_17);
	nor (gm_n160, gm_n45, in_19, in_18, gm_n159, in_21);
	nand (gm_n161, in_4, gm_n74, in_2, gm_n95, in_5);
	or (gm_n162, in_8, in_7, gm_n82, gm_n161, in_9);
	or (gm_n163, in_12, gm_n53, gm_n52, gm_n162, gm_n49);
	nor (gm_n164, in_16, in_15, gm_n50, gm_n163, in_17);
	nand (gm_n165, gm_n45, in_19, gm_n47, gm_n164, in_21);
	not (gm_n166, in_1);
	nand (gm_n167, in_2, gm_n166, in_0, in_4, gm_n74);
	nor (gm_n168, in_7, gm_n82, gm_n72, gm_n167, gm_n64);
	nand (gm_n169, gm_n168, in_10, in_9);
	or (gm_n170, in_13, in_12, gm_n53, gm_n169, in_14);
	nor (gm_n171, gm_n81, in_16, gm_n63, gm_n170, gm_n47);
	nand (gm_n172, gm_n71, gm_n45, in_19, gm_n171);
	and (gm_n173, gm_n55, in_6, in_5, gm_n89, gm_n64);
	and (gm_n174, gm_n173, in_9);
	nand (gm_n175, gm_n48, gm_n53, gm_n52, gm_n174, in_13);
	nor (gm_n176, gm_n46, in_15, in_14, gm_n175, in_17);
	nand (gm_n177, in_20, gm_n62, in_18, gm_n176, in_21);
	nand (gm_n178, in_7, gm_n82, in_5, gm_n89, in_8);
	nor (gm_n179, in_11, in_10, gm_n51, gm_n178, gm_n48);
	nand (gm_n180, in_15, gm_n50, gm_n49, gm_n179, in_16);
	nor (gm_n181, gm_n62, gm_n47, gm_n81, gm_n180, gm_n45);
	nand (gm_n182, gm_n181, in_21);
	or (gm_n183, in_7, gm_n82, in_5, gm_n167, gm_n64);
	or (gm_n184, in_11, in_10, gm_n51, gm_n183, in_12);
	nor (gm_n185, in_15, gm_n50, in_13, gm_n184, in_16);
	nand (gm_n186, in_19, in_18, gm_n81, gm_n185, gm_n45);
	nor (gm_n187, gm_n186, in_21);
	nand (gm_n188, gm_n101, in_1, gm_n73, gm_n54, gm_n74);
	nor (gm_n189, gm_n55, gm_n82, in_5, gm_n188, gm_n64);
	nand (gm_n190, gm_n53, in_10, in_9, gm_n189, gm_n48);
	nor (gm_n191, gm_n63, in_14, gm_n49, gm_n190, gm_n46);
	nand (gm_n192, in_19, in_18, in_17, gm_n191, gm_n45);
	nor (gm_n193, gm_n192, gm_n71);
	nor (gm_n194, gm_n55, in_6, in_5, gm_n124, gm_n64);
	nand (gm_n195, in_11, gm_n52, in_9, gm_n194, gm_n48);
	nor (gm_n196, in_15, gm_n50, in_13, gm_n195, gm_n46);
	nand (gm_n197, in_19, in_18, gm_n81, gm_n196, gm_n45);
	nor (gm_n198, gm_n197, in_21);
	nand (gm_n199, in_4, gm_n74, gm_n101, gm_n102, gm_n72);
	nor (gm_n200, in_8, gm_n55, gm_n82, gm_n199, in_9);
	and (gm_n201, gm_n48, gm_n53, gm_n52, gm_n200, in_13);
	nand (gm_n202, gm_n46, gm_n63, in_14, gm_n201, gm_n81);
	nor (gm_n203, gm_n45, in_19, gm_n47, gm_n202, in_21);
	nand (gm_n204, gm_n54, gm_n74, in_2, gm_n95, gm_n72);
	nor (gm_n205, gm_n64, in_7, in_6, gm_n204, in_9);
	nand (gm_n206, in_12, in_11, gm_n52, gm_n205, gm_n49);
	nor (gm_n207, in_16, gm_n63, gm_n50, gm_n206, in_17);
	nand (gm_n208, in_20, in_19, gm_n47, gm_n207, in_21);
	nor (gm_n209, gm_n101, gm_n166, in_0, gm_n54, in_3);
	and (gm_n210, gm_n55, in_6, gm_n72, gm_n209, in_8);
	and (gm_n211, in_11, gm_n52, in_9, gm_n210, in_12);
	nand (gm_n212, in_15, in_14, in_13, gm_n211, gm_n46);
	nor (gm_n213, in_19, in_18, gm_n81, gm_n212, in_20);
	nand (gm_n214, gm_n213, gm_n71);
	and (gm_n215, gm_n48, gm_n53, gm_n52, gm_n120, in_13);
	and (gm_n216, gm_n46, in_15, gm_n50, gm_n215, in_17);
	nand (gm_n217, in_20, gm_n62, gm_n47, gm_n216, gm_n71);
	or (gm_n218, in_7, in_6, gm_n72, gm_n130, in_8);
	nor (gm_n219, gm_n218, gm_n52, gm_n51);
	nand (gm_n220, in_13, in_12, gm_n53, gm_n219, gm_n50);
	nor (gm_n221, gm_n81, gm_n46, in_15, gm_n220, gm_n47);
	nand (gm_n222, in_21, in_20, in_19, gm_n221);
	nand (gm_n223, gm_n72, in_4, in_3, gm_n83, in_6);
	nor (gm_n224, gm_n51, in_8, in_7, gm_n223, in_10);
	and (gm_n225, gm_n49, in_12, gm_n53, gm_n224, gm_n50);
	nand (gm_n226, gm_n81, in_16, in_15, gm_n225, in_18);
	nor (gm_n227, gm_n71, gm_n45, in_19, gm_n226);
	or (gm_n228, in_8, in_7, in_6, gm_n96, in_9);
	nor (gm_n229, gm_n48, gm_n53, gm_n52, gm_n228, in_13);
	nand (gm_n230, in_16, in_15, in_14, gm_n229, gm_n81);
	nor (gm_n231, in_20, gm_n62, in_18, gm_n230, gm_n71);
	nor (gm_n232, gm_n55, in_6, gm_n72, gm_n108, gm_n64);
	nand (gm_n233, gm_n232, in_9);
	nor (gm_n234, in_12, gm_n53, gm_n52, gm_n233, in_13);
	nand (gm_n235, gm_n46, gm_n63, in_14, gm_n234, gm_n81);
	nor (gm_n236, gm_n45, gm_n62, gm_n47, gm_n235, gm_n71);
	nand (gm_n237, in_11, gm_n52, gm_n51, gm_n194, in_12);
	nor (gm_n238, gm_n63, in_14, in_13, gm_n237, gm_n46);
	nand (gm_n239, in_19, gm_n47, gm_n81, gm_n238, gm_n45);
	nor (gm_n240, gm_n239, gm_n71);
	nor (gm_n241, in_2, in_1, gm_n73, in_4, gm_n74);
	and (gm_n242, in_7, gm_n82, in_5, gm_n241, gm_n64);
	and (gm_n243, gm_n53, gm_n52, in_9, gm_n242, gm_n48);
	nand (gm_n244, gm_n63, in_14, gm_n49, gm_n243, gm_n46);
	nor (gm_n245, gm_n62, gm_n47, in_17, gm_n244, gm_n45);
	nand (gm_n246, gm_n245, in_21);
	nand (gm_n247, gm_n55, in_6, in_5, gm_n241, in_8);
	nor (gm_n248, in_11, in_10, gm_n51, gm_n247, gm_n48);
	nand (gm_n249, in_15, in_14, in_13, gm_n248, in_16);
	nor (gm_n250, gm_n62, gm_n47, in_17, gm_n249, gm_n45);
	nand (gm_n251, gm_n250, gm_n71);
	nor (gm_n252, gm_n101, in_1, gm_n73, in_4, in_3);
	nand (gm_n253, in_7, gm_n82, in_5, gm_n252, gm_n64);
	nor (gm_n254, in_11, in_10, gm_n51, gm_n253, gm_n48);
	nand (gm_n255, gm_n254, in_13);
	nor (gm_n256, in_16, gm_n63, gm_n50, gm_n255, gm_n81);
	nand (gm_n257, in_20, gm_n62, gm_n47, gm_n256, in_21);
	and (gm_n258, in_2, in_1, in_0);
	nand (gm_n259, gm_n72, in_4, gm_n74, gm_n258, gm_n82);
	nor (gm_n260, in_9, in_8, in_7, gm_n259, gm_n52);
	nand (gm_n261, gm_n49, in_12, in_11, gm_n260, in_14);
	nor (gm_n262, gm_n81, gm_n46, in_15, gm_n261, gm_n47);
	nand (gm_n263, gm_n71, gm_n45, in_19, gm_n262);
	or (gm_n264, in_8, in_7, in_6, gm_n156, gm_n51);
	nor (gm_n265, gm_n48, gm_n53, gm_n52, gm_n264, gm_n49);
	nand (gm_n266, gm_n46, gm_n63, gm_n50, gm_n265, in_17);
	nor (gm_n267, gm_n45, gm_n62, gm_n47, gm_n266, in_21);
	nor (gm_n268, in_8, gm_n55, gm_n82, gm_n119, gm_n51);
	and (gm_n269, in_12, in_11, in_10, gm_n268, gm_n49);
	nand (gm_n270, in_16, gm_n63, gm_n50, gm_n269, in_17);
	nor (gm_n271, gm_n45, gm_n62, gm_n47, gm_n270, gm_n71);
	nor (gm_n272, in_12, in_11, gm_n52, gm_n162, in_13);
	nand (gm_n273, in_16, gm_n63, gm_n50, gm_n272, in_17);
	nor (gm_n274, gm_n45, in_19, gm_n47, gm_n273, gm_n71);
	nand (gm_n275, gm_n53, gm_n52, gm_n51, gm_n109, in_12);
	nor (gm_n276, in_15, in_14, gm_n49, gm_n275, gm_n46);
	nand (gm_n277, in_19, in_18, in_17, gm_n276, in_20);
	nor (gm_n278, gm_n277, in_21);
	nand (gm_n279, in_5, in_4, gm_n74, gm_n258, gm_n82);
	nor (gm_n280, gm_n51, gm_n64, gm_n55, gm_n279);
	nand (gm_n281, gm_n48, in_11, gm_n52, gm_n280, gm_n49);
	nor (gm_n282, gm_n46, in_15, gm_n50, gm_n281, in_17);
	nand (gm_n283, in_20, gm_n62, gm_n47, gm_n282, in_21);
	nor (gm_n284, gm_n101, in_1, gm_n73, gm_n54, gm_n74);
	nand (gm_n285, gm_n55, in_6, gm_n72, gm_n284, in_8);
	nor (gm_n286, gm_n53, gm_n52, in_9, gm_n285);
	nand (gm_n287, in_14, in_13, in_12, gm_n286, gm_n63);
	nor (gm_n288, in_18, gm_n81, in_16, gm_n287, in_19);
	nand (gm_n289, gm_n288, in_21, in_20);
	nand (gm_n290, gm_n101, gm_n166, in_0, gm_n54, gm_n74);
	nor (gm_n291, in_7, in_6, in_5, gm_n290, gm_n64);
	nand (gm_n292, in_11, in_10, gm_n51, gm_n291, in_12);
	nor (gm_n293, gm_n292, in_14, in_13);
	and (gm_n294, in_17, in_16, in_15, gm_n293, gm_n47);
	nand (gm_n295, in_21, gm_n45, gm_n62, gm_n294);
	nor (gm_n296, in_2, in_1, gm_n73, gm_n54, in_3);
	and (gm_n297, gm_n55, gm_n82, gm_n72, gm_n296, in_8);
	and (gm_n298, in_11, in_10, gm_n51, gm_n297);
	nand (gm_n299, in_14, gm_n49, in_12, gm_n298, gm_n63);
	nor (gm_n300, gm_n47, gm_n81, in_16, gm_n299, gm_n62);
	nand (gm_n301, gm_n300, gm_n71, in_20);
	and (gm_n302, gm_n55, in_6, in_5, gm_n209);
	and (gm_n303, gm_n52, gm_n51, in_8, gm_n302, in_11);
	and (gm_n304, gm_n50, gm_n49, gm_n48, gm_n303, in_15);
	nand (gm_n305, in_18, in_17, in_16, gm_n304, in_19);
	nor (gm_n306, gm_n305, gm_n71, in_20);
	or (gm_n307, gm_n53, in_10, in_9, gm_n183, in_12);
	nor (gm_n308, in_15, in_14, gm_n49, gm_n307, gm_n46);
	nand (gm_n309, gm_n62, in_18, in_17, gm_n308, in_20);
	nor (gm_n310, gm_n309, in_21);
	nor (gm_n311, gm_n64, in_7, gm_n82, gm_n141, gm_n51);
	and (gm_n312, in_12, in_11, in_10, gm_n311, in_13);
	nand (gm_n313, in_16, gm_n63, in_14, gm_n312, gm_n81);
	nor (gm_n314, in_20, gm_n62, gm_n47, gm_n313, gm_n71);
	nand (gm_n315, in_2, in_1, in_0, in_3);
	nor (gm_n316, in_6, gm_n72, in_4, gm_n315, in_7);
	nand (gm_n317, gm_n52, gm_n51, gm_n64, gm_n316, in_11);
	nor (gm_n318, in_14, in_13, gm_n48, gm_n317);
	nand (gm_n319, gm_n81, gm_n46, gm_n63, gm_n318, gm_n47);
	nor (gm_n320, in_21, gm_n45, gm_n62, gm_n319);
	nand (gm_n321, gm_n101, in_1, gm_n73, gm_n54, in_3);
	or (gm_n322, gm_n55, in_6, gm_n72, gm_n321, in_8);
	nor (gm_n323, gm_n53, gm_n52, gm_n51, gm_n322);
	nand (gm_n324, in_14, gm_n49, gm_n48, gm_n323, gm_n63);
	nor (gm_n325, gm_n47, in_17, gm_n46, gm_n324, in_19);
	nand (gm_n326, gm_n325, gm_n71, gm_n45);
	nor (gm_n327, gm_n101, in_1, gm_n73, in_4, gm_n74);
	nand (gm_n328, gm_n55, gm_n82, in_5, gm_n327, in_8);
	nor (gm_n329, gm_n328, in_10, in_9);
	nand (gm_n330, gm_n49, gm_n48, gm_n53, gm_n329, gm_n50);
	nor (gm_n331, gm_n81, gm_n46, in_15, gm_n330, gm_n47);
	nand (gm_n332, gm_n71, in_20, gm_n62, gm_n331);
	nand (gm_n333, in_7, in_6, in_5, gm_n327, gm_n64);
	or (gm_n334, in_11, gm_n52, in_9, gm_n333, gm_n48);
	or (gm_n335, in_15, in_14, in_13, gm_n334, gm_n46);
	nor (gm_n336, gm_n62, in_18, gm_n81, gm_n335, gm_n45);
	nand (gm_n337, gm_n336, gm_n71);
	nor (gm_n338, gm_n82, gm_n72, gm_n54, gm_n56, gm_n55);
	and (gm_n339, gm_n338, gm_n51, in_8);
	nand (gm_n340, in_12, gm_n53, gm_n52, gm_n339, in_13);
	nor (gm_n341, in_16, in_15, gm_n50, gm_n340, in_17);
	nand (gm_n342, gm_n45, in_19, gm_n47, gm_n341, in_21);
	nor (gm_n343, in_8, in_7, gm_n82, gm_n96, gm_n51);
	and (gm_n344, gm_n48, gm_n53, in_10, gm_n343, in_13);
	nand (gm_n345, in_16, gm_n63, in_14, gm_n344, in_17);
	nor (gm_n346, gm_n45, gm_n62, in_18, gm_n345, in_21);
	or (gm_n347, in_9, in_8, in_7, gm_n84);
	nor (gm_n348, gm_n48, gm_n53, in_10, gm_n347, gm_n49);
	nand (gm_n349, in_16, in_15, in_14, gm_n348, in_17);
	nor (gm_n350, in_20, gm_n62, gm_n47, gm_n349, gm_n71);
	nor (gm_n351, gm_n328, gm_n52, gm_n51);
	and (gm_n352, in_13, in_12, gm_n53, gm_n351, gm_n50);
	nand (gm_n353, gm_n81, in_16, gm_n63, gm_n352, in_18);
	nor (gm_n354, gm_n71, in_20, gm_n62, gm_n353);
	nor (gm_n355, gm_n55, in_6, in_5, gm_n108, in_8);
	and (gm_n356, in_11, in_10, gm_n51, gm_n355, gm_n48);
	and (gm_n357, in_15, gm_n50, gm_n49, gm_n356, gm_n46);
	nand (gm_n358, in_19, in_18, gm_n81, gm_n357, gm_n45);
	nor (gm_n359, gm_n358, gm_n71);
	and (gm_n360, gm_n48, in_11, gm_n52, gm_n146, gm_n49);
	and (gm_n361, gm_n46, gm_n63, in_14, gm_n360, gm_n81);
	nand (gm_n362, gm_n45, gm_n62, in_18, gm_n361, gm_n71);
	or (gm_n363, gm_n55, in_6, in_5, gm_n75, in_8);
	nor (gm_n364, in_11, in_10, in_9, gm_n363, in_12);
	nand (gm_n365, in_15, gm_n50, in_13, gm_n364, gm_n46);
	nor (gm_n366, gm_n62, in_18, gm_n81, gm_n365, in_20);
	nand (gm_n367, gm_n366, in_21);
	or (gm_n368, in_7, in_6, gm_n72, gm_n130, gm_n64);
	or (gm_n369, gm_n53, in_10, in_9, gm_n368);
	nor (gm_n370, in_14, gm_n49, in_12, gm_n369, in_15);
	and (gm_n371, in_18, gm_n81, gm_n46, gm_n370, in_19);
	nand (gm_n372, gm_n371, gm_n71, in_20);
	nand (gm_n373, in_1, in_0);
	nor (gm_n374, in_4, in_3, in_2, gm_n373, in_5);
	and (gm_n375, gm_n64, gm_n55, gm_n82, gm_n374, gm_n51);
	nand (gm_n376, gm_n48, gm_n53, in_10, gm_n375, gm_n49);
	nor (gm_n377, in_16, gm_n63, gm_n50, gm_n376, in_17);
	nand (gm_n378, in_20, gm_n62, in_18, gm_n377, in_21);
	nor (gm_n379, gm_n54, gm_n74, in_2, gm_n373, gm_n72);
	and (gm_n380, in_8, in_7, in_6, gm_n379, gm_n51);
	and (gm_n381, gm_n48, gm_n53, in_10, gm_n380, in_13);
	nand (gm_n382, in_16, gm_n63, in_14, gm_n381, gm_n81);
	nor (gm_n383, gm_n45, gm_n62, in_18, gm_n382, in_21);
	nor (gm_n384, in_7, in_6, gm_n72, gm_n124);
	nand (gm_n385, in_10, gm_n51, in_8, gm_n384);
	nor (gm_n386, in_13, gm_n48, gm_n53, gm_n385);
	nand (gm_n387, gm_n46, in_15, gm_n50, gm_n386, gm_n81);
	nor (gm_n388, gm_n45, in_19, gm_n47, gm_n387, in_21);
	and (gm_n389, in_2, in_1, in_0, in_3);
	nand (gm_n390, gm_n82, in_5, gm_n54, gm_n389, in_7);
	or (gm_n391, in_10, gm_n51, gm_n64, gm_n390);
	nor (gm_n392, in_13, gm_n48, in_11, gm_n391, in_14);
	nand (gm_n393, in_17, in_16, gm_n63, gm_n392, in_18);
	nor (gm_n394, in_21, in_20, in_19, gm_n393);
	nand (gm_n395, gm_n55, gm_n82, in_5, gm_n296, in_8);
	nor (gm_n396, gm_n53, in_10, gm_n51, gm_n395);
	and (gm_n397, in_14, in_13, in_12, gm_n396, gm_n63);
	nand (gm_n398, gm_n47, in_17, gm_n46, gm_n397, gm_n62);
	nor (gm_n399, gm_n398, gm_n71, gm_n45);
	nor (gm_n400, in_8, gm_n55, gm_n82, gm_n199, gm_n51);
	and (gm_n401, gm_n48, in_11, in_10, gm_n400, gm_n49);
	and (gm_n402, in_16, gm_n63, in_14, gm_n401, in_17);
	nand (gm_n403, gm_n45, in_19, in_18, gm_n402, gm_n71);
	nor (gm_n404, gm_n72, gm_n54, in_3, gm_n65, gm_n82);
	nand (gm_n405, in_9, in_8, gm_n55, gm_n404, gm_n52);
	nor (gm_n406, gm_n405, in_11);
	nand (gm_n407, in_14, in_13, in_12, gm_n406, in_15);
	nor (gm_n408, in_18, in_17, in_16, gm_n407, in_19);
	nand (gm_n409, gm_n408, gm_n71, in_20);
	or (gm_n410, gm_n55, in_6, in_5, gm_n321, in_8);
	or (gm_n411, gm_n410, gm_n51);
	or (gm_n412, gm_n48, in_11, in_10, gm_n411, in_13);
	nor (gm_n413, in_16, in_15, gm_n50, gm_n412, in_17);
	nand (gm_n414, in_20, gm_n62, in_18, gm_n413, gm_n71);
	or (gm_n415, gm_n55, gm_n82, in_5, gm_n75, gm_n64);
	nor (gm_n416, gm_n415, in_10, gm_n51);
	nand (gm_n417, gm_n49, in_12, in_11, gm_n416, in_14);
	nor (gm_n418, gm_n81, gm_n46, gm_n63, gm_n417, gm_n47);
	nand (gm_n419, gm_n71, gm_n45, gm_n62, gm_n418);
	nor (gm_n420, gm_n101, gm_n166, in_0, gm_n54, gm_n74);
	and (gm_n421, gm_n55, in_6, gm_n72, gm_n420, gm_n64);
	nand (gm_n422, in_11, in_10, in_9, gm_n421, gm_n48);
	nor (gm_n423, in_15, gm_n50, in_13, gm_n422, gm_n46);
	nand (gm_n424, gm_n423, gm_n47, gm_n81);
	nor (gm_n425, gm_n71, in_20, in_19, gm_n424);
	nand (gm_n426, in_7, gm_n82, in_5, gm_n284, in_8);
	nor (gm_n427, gm_n426, in_9);
	and (gm_n428, in_12, in_11, gm_n52, gm_n427, in_13);
	nand (gm_n429, gm_n46, in_15, in_14, gm_n428, gm_n81);
	nor (gm_n430, gm_n45, in_19, gm_n47, gm_n429, gm_n71);
	nor (gm_n431, in_6, in_5, in_4, gm_n315, in_7);
	nand (gm_n432, gm_n431, gm_n51, in_8);
	nor (gm_n433, gm_n48, gm_n53, gm_n52, gm_n432, gm_n49);
	nand (gm_n434, in_16, in_15, gm_n50, gm_n433, gm_n81);
	nor (gm_n435, gm_n45, in_19, in_18, gm_n434, gm_n71);
	nor (gm_n436, in_9, in_8, in_7, gm_n279, in_10);
	and (gm_n437, gm_n49, in_12, gm_n53, gm_n436);
	nand (gm_n438, gm_n46, gm_n63, in_14, gm_n437, gm_n81);
	nor (gm_n439, in_20, in_19, gm_n47, gm_n438, in_21);
	or (gm_n440, in_7, in_6, in_5, gm_n167, in_8);
	nor (gm_n441, gm_n53, gm_n52, in_9, gm_n440, in_12);
	nand (gm_n442, gm_n63, gm_n50, in_13, gm_n441, in_16);
	nor (gm_n443, gm_n62, in_18, in_17, gm_n442, in_20);
	nand (gm_n444, gm_n443, gm_n71);
	or (gm_n445, gm_n51, gm_n64, in_7, gm_n259, gm_n52);
	or (gm_n446, gm_n49, in_12, gm_n53, gm_n445);
	nor (gm_n447, gm_n46, gm_n63, gm_n50, gm_n446, gm_n81);
	nand (gm_n448, in_20, in_19, gm_n47, gm_n447, in_21);
	nor (gm_n449, gm_n51, in_8, in_7, gm_n259);
	nand (gm_n450, gm_n48, gm_n53, in_10, gm_n449, in_13);
	nor (gm_n451, gm_n46, in_15, in_14, gm_n450, in_17);
	nand (gm_n452, in_20, in_19, in_18, gm_n451, gm_n71);
	or (gm_n453, in_7, in_6, in_5, gm_n167, gm_n64);
	nor (gm_n454, in_11, gm_n52, gm_n51, gm_n453, gm_n48);
	nand (gm_n455, gm_n454, in_14, in_13);
	nor (gm_n456, in_17, gm_n46, in_15, gm_n455, gm_n47);
	nand (gm_n457, gm_n71, gm_n45, in_19, gm_n456);
	and (gm_n458, in_7, gm_n82, gm_n72, gm_n296, gm_n64);
	and (gm_n459, in_11, in_10, gm_n51, gm_n458, gm_n48);
	and (gm_n460, gm_n63, in_14, gm_n49, gm_n459, in_16);
	nand (gm_n461, in_19, gm_n47, gm_n81, gm_n460, gm_n45);
	nor (gm_n462, gm_n461, gm_n71);
	nand (gm_n463, in_5, gm_n54, in_3, gm_n83, in_6);
	or (gm_n464, in_9, in_8, in_7, gm_n463, gm_n52);
	nor (gm_n465, gm_n49, gm_n48, gm_n53, gm_n464, in_14);
	nand (gm_n466, in_17, gm_n46, in_15, gm_n465, in_18);
	nor (gm_n467, in_21, in_20, gm_n62, gm_n466);
	or (gm_n468, gm_n82, in_5, gm_n54, gm_n56, gm_n55);
	nor (gm_n469, gm_n52, gm_n51, gm_n64, gm_n468, in_11);
	and (gm_n470, gm_n50, in_13, in_12, gm_n469, gm_n63);
	nand (gm_n471, gm_n47, gm_n81, gm_n46, gm_n470, gm_n62);
	nor (gm_n472, gm_n471, in_21, gm_n45);
	nor (gm_n473, in_7, in_6, gm_n72, gm_n321, gm_n64);
	nand (gm_n474, in_11, in_10, in_9, gm_n473, in_12);
	nor (gm_n475, in_15, gm_n50, gm_n49, gm_n474, gm_n46);
	nand (gm_n476, in_19, in_18, in_17, gm_n475, in_20);
	nor (gm_n477, gm_n476, in_21);
	nand (gm_n478, in_6, in_5, gm_n54, gm_n389, in_7);
	nor (gm_n479, gm_n52, gm_n51, gm_n64, gm_n478, in_11);
	nand (gm_n480, in_14, gm_n49, in_12, gm_n479, in_15);
	nor (gm_n481, in_18, gm_n81, gm_n46, gm_n480, gm_n62);
	nand (gm_n482, gm_n481, gm_n71, gm_n45);
	nand (gm_n483, in_2, gm_n166, in_0, gm_n54, gm_n74);
	nor (gm_n484, in_7, in_6, in_5, gm_n483, in_8);
	and (gm_n485, gm_n53, gm_n52, in_9, gm_n484);
	nand (gm_n486, gm_n50, in_13, gm_n48, gm_n485, in_15);
	nor (gm_n487, gm_n47, gm_n81, in_16, gm_n486, in_19);
	nand (gm_n488, gm_n487, in_21, in_20);
	nor (gm_n489, gm_n53, in_10, in_9, gm_n453, in_12);
	nand (gm_n490, in_15, in_14, gm_n49, gm_n489, in_16);
	nor (gm_n491, gm_n62, gm_n47, gm_n81, gm_n490, gm_n45);
	nand (gm_n492, gm_n491, gm_n71);
	nor (gm_n493, gm_n101, gm_n166, in_0, in_4, gm_n74);
	and (gm_n494, gm_n55, in_6, in_5, gm_n493, gm_n64);
	and (gm_n495, in_11, gm_n52, in_9, gm_n494, gm_n48);
	nand (gm_n496, in_15, gm_n50, in_13, gm_n495, gm_n46);
	nor (gm_n497, gm_n62, gm_n47, in_17, gm_n496, in_20);
	nand (gm_n498, gm_n497, gm_n71);
	or (gm_n499, gm_n64, in_7, in_6, gm_n199, gm_n51);
	nor (gm_n500, gm_n499, in_10);
	and (gm_n501, gm_n49, in_12, in_11, gm_n500, gm_n50);
	nand (gm_n502, gm_n81, gm_n46, in_15, gm_n501, in_18);
	nor (gm_n503, in_21, gm_n45, in_19, gm_n502);
	nor (gm_n504, in_5, in_4, in_3, gm_n65, gm_n82);
	and (gm_n505, gm_n51, gm_n64, in_7, gm_n504, gm_n52);
	and (gm_n506, in_13, in_12, in_11, gm_n505, gm_n50);
	nand (gm_n507, in_17, gm_n46, gm_n63, gm_n506, gm_n47);
	nor (gm_n508, in_21, gm_n45, gm_n62, gm_n507);
	nor (gm_n509, gm_n55, gm_n82, in_5, gm_n290, gm_n64);
	nand (gm_n510, gm_n509, gm_n51);
	nor (gm_n511, in_12, gm_n53, in_10, gm_n510, gm_n49);
	nand (gm_n512, gm_n46, gm_n63, gm_n50, gm_n511, gm_n81);
	nor (gm_n513, in_20, in_19, in_18, gm_n512, gm_n71);
	nand (gm_n514, in_7, in_6, in_5, gm_n420, in_8);
	or (gm_n515, in_11, in_10, gm_n51, gm_n514, in_12);
	nor (gm_n516, gm_n515, gm_n50, in_13);
	nand (gm_n517, gm_n81, gm_n46, gm_n63, gm_n516, gm_n47);
	nor (gm_n518, in_21, gm_n45, gm_n62, gm_n517);
	nor (gm_n519, in_2, gm_n166, in_0, in_4, in_3);
	nand (gm_n520, in_7, in_6, in_5, gm_n519, gm_n64);
	nor (gm_n521, in_11, in_10, in_9, gm_n520, in_12);
	nand (gm_n522, gm_n63, in_14, in_13, gm_n521, in_16);
	nor (gm_n523, in_19, in_18, in_17, gm_n522, gm_n45);
	nand (gm_n524, gm_n523, in_21);
	nand (gm_n525, in_5, in_4, in_3, gm_n83, in_6);
	nor (gm_n526, gm_n51, gm_n64, in_7, gm_n525, gm_n52);
	nand (gm_n527, gm_n49, in_12, gm_n53, gm_n526, gm_n50);
	nor (gm_n528, gm_n81, gm_n46, in_15, gm_n527, gm_n47);
	nand (gm_n529, in_21, in_20, gm_n62, gm_n528);
	nand (gm_n530, in_4, gm_n74, in_2, gm_n95, gm_n72);
	or (gm_n531, gm_n64, in_7, gm_n82, gm_n530, gm_n51);
	or (gm_n532, gm_n48, gm_n53, in_10, gm_n531, in_13);
	nor (gm_n533, in_16, gm_n63, gm_n50, gm_n532, in_17);
	nand (gm_n534, gm_n45, gm_n62, in_18, gm_n533, gm_n71);
	nand (gm_n535, in_14, in_13, in_12, gm_n303, in_15);
	nor (gm_n536, gm_n47, gm_n81, in_16, gm_n535, gm_n62);
	nand (gm_n537, gm_n536, in_21, in_20);
	nor (gm_n538, gm_n55, gm_n82, gm_n72, gm_n75, in_8);
	and (gm_n539, gm_n538, in_10, in_9);
	and (gm_n540, in_13, in_12, in_11, gm_n539, gm_n50);
	nand (gm_n541, in_17, in_16, gm_n63, gm_n540, gm_n47);
	nor (gm_n542, gm_n71, in_20, gm_n62, gm_n541);
	and (gm_n543, gm_n55, gm_n82, in_5, gm_n296, gm_n64);
	and (gm_n544, gm_n543, in_9);
	and (gm_n545, in_12, gm_n53, gm_n52, gm_n544, gm_n49);
	nand (gm_n546, in_16, in_15, gm_n50, gm_n545, gm_n81);
	nor (gm_n547, gm_n45, gm_n62, gm_n47, gm_n546, in_21);
	nor (gm_n548, gm_n55, gm_n82, in_5, gm_n321, in_8);
	and (gm_n549, gm_n53, gm_n52, in_9, gm_n548);
	and (gm_n550, in_14, in_13, in_12, gm_n549, gm_n63);
	nand (gm_n551, in_18, in_17, gm_n46, gm_n550, in_19);
	nor (gm_n552, gm_n551, in_21, gm_n45);
	nand (gm_n553, in_5, gm_n54, gm_n74, gm_n258, in_6);
	or (gm_n554, gm_n51, gm_n64, in_7, gm_n553, gm_n52);
	nor (gm_n555, in_13, gm_n48, in_11, gm_n554, gm_n50);
	nand (gm_n556, in_17, gm_n46, in_15, gm_n555, gm_n47);
	nor (gm_n557, gm_n71, in_20, in_19, gm_n556);
	nor (gm_n558, in_11, gm_n52, in_9, gm_n178, gm_n48);
	nand (gm_n559, gm_n63, gm_n50, gm_n49, gm_n558, gm_n46);
	nor (gm_n560, in_19, in_18, in_17, gm_n559, gm_n45);
	nand (gm_n561, gm_n560, in_21);
	nor (gm_n562, in_8, gm_n55, in_6, gm_n161, gm_n51);
	nand (gm_n563, in_12, gm_n53, in_10, gm_n562, gm_n49);
	nor (gm_n564, gm_n46, gm_n63, gm_n50, gm_n563, gm_n81);
	nand (gm_n565, gm_n45, gm_n62, gm_n47, gm_n564, in_21);
	and (gm_n566, in_7, gm_n82, gm_n72, gm_n493, in_8);
	and (gm_n567, in_11, gm_n52, in_9, gm_n566);
	nand (gm_n568, in_14, gm_n49, in_12, gm_n567, gm_n63);
	nor (gm_n569, gm_n47, in_17, gm_n46, gm_n568, gm_n62);
	nand (gm_n570, gm_n569, gm_n71, gm_n45);
	nand (gm_n571, in_7, in_6, in_5, gm_n493, in_8);
	nor (gm_n572, in_11, gm_n52, gm_n51, gm_n571);
	nand (gm_n573, in_14, gm_n49, in_12, gm_n572, gm_n63);
	nor (gm_n574, in_18, gm_n81, in_16, gm_n573, in_19);
	nand (gm_n575, gm_n574, gm_n71, gm_n45);
	and (gm_n576, gm_n48, in_11, in_10, gm_n120, gm_n49);
	nand (gm_n577, gm_n46, in_15, in_14, gm_n576, gm_n81);
	nor (gm_n578, in_20, in_19, gm_n47, gm_n577, gm_n71);
	nor (gm_n579, gm_n51, gm_n64, gm_n55, gm_n553, gm_n52);
	and (gm_n580, in_13, in_12, in_11, gm_n579, in_14);
	nand (gm_n581, gm_n81, gm_n46, gm_n63, gm_n580, in_18);
	nor (gm_n582, gm_n71, gm_n45, in_19, gm_n581);
	or (gm_n583, gm_n55, gm_n82, in_5, gm_n167, in_8);
	nor (gm_n584, in_11, in_10, in_9, gm_n583);
	and (gm_n585, gm_n50, gm_n49, in_12, gm_n584, gm_n63);
	nand (gm_n586, in_18, gm_n81, gm_n46, gm_n585, in_19);
	nor (gm_n587, gm_n586, in_21, gm_n45);
	nand (gm_n588, in_5, gm_n54, in_3, gm_n83, gm_n82);
	nor (gm_n589, gm_n51, gm_n64, in_7, gm_n588);
	and (gm_n590, in_12, in_11, gm_n52, gm_n589, gm_n49);
	nand (gm_n591, in_16, in_15, in_14, gm_n590, in_17);
	nor (gm_n592, in_20, gm_n62, gm_n47, gm_n591, gm_n71);
	nor (gm_n593, gm_n55, in_6, in_5, gm_n290, in_8);
	and (gm_n594, gm_n593, in_10, in_9);
	nand (gm_n595, in_13, gm_n48, gm_n53, gm_n594, gm_n50);
	nor (gm_n596, in_17, in_16, in_15, gm_n595, gm_n47);
	nand (gm_n597, in_21, in_20, gm_n62, gm_n596);
	and (gm_n598, in_2, in_1, in_0, in_4, in_3);
	nand (gm_n599, gm_n55, gm_n82, in_5, gm_n598, gm_n64);
	nor (gm_n600, in_11, in_10, gm_n51, gm_n599, in_12);
	nand (gm_n601, in_15, in_14, gm_n49, gm_n600, gm_n46);
	nor (gm_n602, in_19, gm_n47, in_17, gm_n601, in_20);
	nand (gm_n603, gm_n602, gm_n71);
	nand (gm_n604, gm_n48, in_11, in_10, gm_n174, in_13);
	nor (gm_n605, in_16, in_15, in_14, gm_n604, in_17);
	nand (gm_n606, in_20, gm_n62, gm_n47, gm_n605, gm_n71);
	or (gm_n607, in_7, gm_n82, gm_n72, gm_n321, gm_n64);
	nor (gm_n608, in_11, gm_n52, in_9, gm_n607, gm_n48);
	nand (gm_n609, in_15, gm_n50, in_13, gm_n608, in_16);
	nor (gm_n610, gm_n62, gm_n47, in_17, gm_n609, gm_n45);
	nand (gm_n611, gm_n610, gm_n71);
	nor (gm_n612, gm_n55, gm_n82, gm_n72, gm_n290, gm_n64);
	nand (gm_n613, in_11, in_10, in_9, gm_n612);
	nor (gm_n614, gm_n50, in_13, gm_n48, gm_n613, in_15);
	nand (gm_n615, in_18, in_17, gm_n46, gm_n614, gm_n62);
	nor (gm_n616, gm_n615, gm_n71, gm_n45);
	nor (gm_n617, gm_n64, gm_n55, in_6, gm_n204, in_9);
	and (gm_n618, gm_n48, gm_n53, in_10, gm_n617, gm_n49);
	nand (gm_n619, gm_n46, in_15, gm_n50, gm_n618, in_17);
	nor (gm_n620, gm_n45, gm_n62, gm_n47, gm_n619, in_21);
	and (gm_n621, gm_n55, gm_n82, in_5, gm_n493, gm_n64);
	nand (gm_n622, gm_n621, in_10, in_9);
	nor (gm_n623, in_13, in_12, gm_n53, gm_n622, gm_n50);
	nand (gm_n624, gm_n81, in_16, in_15, gm_n623, in_18);
	nor (gm_n625, gm_n71, gm_n45, gm_n62, gm_n624);
	or (gm_n626, gm_n52, gm_n51, in_8, gm_n478, gm_n53);
	nor (gm_n627, in_14, in_13, gm_n48, gm_n626, in_15);
	nand (gm_n628, gm_n47, gm_n81, gm_n46, gm_n627, gm_n62);
	nor (gm_n629, gm_n628, in_21, in_20);
	or (gm_n630, in_9, in_8, gm_n55, gm_n279, gm_n52);
	nor (gm_n631, gm_n49, gm_n48, gm_n53, gm_n630, in_14);
	and (gm_n632, in_17, gm_n46, gm_n63, gm_n631, in_18);
	nand (gm_n633, gm_n71, in_20, in_19, gm_n632);
	nor (gm_n634, in_11, gm_n52, in_9, gm_n571);
	nand (gm_n635, gm_n50, gm_n49, gm_n48, gm_n634, gm_n63);
	nor (gm_n636, gm_n47, in_17, gm_n46, gm_n635, in_19);
	nand (gm_n637, gm_n636, gm_n71, gm_n45);
	nor (gm_n638, in_4, gm_n74, in_2, gm_n373, gm_n72);
	nand (gm_n639, gm_n64, gm_n55, in_6, gm_n638, gm_n51);
	or (gm_n640, gm_n48, in_11, gm_n52, gm_n639, in_13);
	nor (gm_n641, in_16, gm_n63, gm_n50, gm_n640, gm_n81);
	nand (gm_n642, gm_n45, in_19, gm_n47, gm_n641, gm_n71);
	nand (gm_n643, gm_n101, in_1, gm_n73, in_4, gm_n74);
	nor (gm_n644, in_7, in_6, gm_n72, gm_n643, gm_n64);
	and (gm_n645, in_11, in_10, in_9, gm_n644, gm_n48);
	nand (gm_n646, in_15, in_14, in_13, gm_n645, gm_n46);
	nor (gm_n647, gm_n62, in_18, in_17, gm_n646, gm_n45);
	nand (gm_n648, gm_n647, gm_n71);
	or (gm_n649, in_7, in_6, in_5, gm_n130, in_8);
	or (gm_n650, in_11, in_10, gm_n51, gm_n649);
	nor (gm_n651, in_14, gm_n49, gm_n48, gm_n650, gm_n63);
	nand (gm_n652, gm_n47, gm_n81, gm_n46, gm_n651, gm_n62);
	nor (gm_n653, gm_n652, in_21, in_20);
	nor (gm_n654, in_8, in_7, in_6, gm_n141, gm_n51);
	and (gm_n655, in_12, in_11, in_10, gm_n654, gm_n49);
	nand (gm_n656, in_16, gm_n63, gm_n50, gm_n655, gm_n81);
	nor (gm_n657, in_20, gm_n62, gm_n47, gm_n656, gm_n71);
	and (gm_n658, in_7, in_6, gm_n72, gm_n284, gm_n64);
	nand (gm_n659, in_11, in_10, in_9, gm_n658, gm_n48);
	nor (gm_n660, gm_n63, gm_n50, gm_n49, gm_n659, gm_n46);
	nand (gm_n661, in_19, in_18, gm_n81, gm_n660, gm_n45);
	nor (gm_n662, gm_n661, in_21);
	nor (gm_n663, in_7, gm_n82, in_5, gm_n130);
	and (gm_n664, gm_n52, in_9, gm_n64, gm_n663, in_11);
	and (gm_n665, in_14, in_13, in_12, gm_n664, gm_n63);
	nand (gm_n666, in_18, in_17, in_16, gm_n665, gm_n62);
	nor (gm_n667, gm_n666, in_21, gm_n45);
	nor (gm_n668, gm_n55, gm_n82, in_5, gm_n321, gm_n64);
	nand (gm_n669, gm_n53, in_10, in_9, gm_n668, in_12);
	nor (gm_n670, gm_n669, in_13);
	and (gm_n671, in_16, in_15, in_14, gm_n670, gm_n81);
	nand (gm_n672, gm_n45, in_19, gm_n47, gm_n671, gm_n71);
	and (gm_n673, in_7, in_6, in_5, gm_n296, gm_n64);
	and (gm_n674, in_11, gm_n52, gm_n51, gm_n673, gm_n48);
	nand (gm_n675, gm_n63, in_14, in_13, gm_n674, gm_n46);
	nor (gm_n676, gm_n62, in_18, in_17, gm_n675, gm_n45);
	nand (gm_n677, gm_n676, gm_n71);
	and (gm_n678, in_9, gm_n64, in_7, gm_n504);
	nand (gm_n679, gm_n48, gm_n53, gm_n52, gm_n678, gm_n49);
	nor (gm_n680, in_16, gm_n63, in_14, gm_n679, in_17);
	nand (gm_n681, gm_n45, gm_n62, gm_n47, gm_n680, in_21);
	nor (gm_n682, gm_n51, in_8, gm_n55, gm_n84, gm_n52);
	nand (gm_n683, in_13, in_12, gm_n53, gm_n682, in_14);
	nor (gm_n684, gm_n81, in_16, gm_n63, gm_n683, in_18);
	nand (gm_n685, in_21, in_20, in_19, gm_n684);
	or (gm_n686, in_7, gm_n82, gm_n72, gm_n124, in_8);
	nor (gm_n687, gm_n686, in_10, in_9);
	and (gm_n688, gm_n49, gm_n48, in_11, gm_n687, gm_n50);
	nand (gm_n689, in_17, gm_n46, in_15, gm_n688, in_18);
	nor (gm_n690, gm_n71, in_20, in_19, gm_n689);
	nor (gm_n691, gm_n82, in_5, gm_n54, gm_n56, in_7);
	and (gm_n692, gm_n691, gm_n51, gm_n64);
	and (gm_n693, gm_n48, in_11, gm_n52, gm_n692, in_13);
	nand (gm_n694, in_16, gm_n63, gm_n50, gm_n693, gm_n81);
	nor (gm_n695, gm_n45, in_19, in_18, gm_n694, in_21);
	nor (gm_n696, in_8, in_7, in_6, gm_n199, gm_n51);
	and (gm_n697, gm_n48, in_11, in_10, gm_n696, in_13);
	nand (gm_n698, in_16, in_15, in_14, gm_n697, in_17);
	nor (gm_n699, gm_n45, gm_n62, gm_n47, gm_n698, in_21);
	and (gm_n700, in_7, gm_n82, in_5, gm_n296, in_8);
	nand (gm_n701, gm_n53, in_10, in_9, gm_n700);
	nor (gm_n702, in_14, gm_n49, gm_n48, gm_n701, in_15);
	nand (gm_n703, gm_n47, gm_n81, in_16, gm_n702, gm_n62);
	nor (gm_n704, gm_n703, in_21, in_20);
	nor (gm_n705, gm_n53, gm_n52, in_9, gm_n415, gm_n48);
	nand (gm_n706, gm_n63, gm_n50, gm_n49, gm_n705, gm_n46);
	nor (gm_n707, in_19, gm_n47, gm_n81, gm_n706, gm_n45);
	nand (gm_n708, gm_n707, in_21);
	nor (gm_n709, gm_n53, gm_n52, gm_n51, gm_n607);
	nand (gm_n710, in_14, gm_n49, in_12, gm_n709, gm_n63);
	nor (gm_n711, in_18, gm_n81, gm_n46, gm_n710, gm_n62);
	nand (gm_n712, gm_n711, gm_n71, gm_n45);
	nor (gm_n713, in_9, gm_n64, gm_n55, gm_n223, in_10);
	nand (gm_n714, in_13, in_12, in_11, gm_n713);
	nor (gm_n715, in_16, gm_n63, gm_n50, gm_n714, in_17);
	nand (gm_n716, gm_n45, in_19, in_18, gm_n715, in_21);
	nor (gm_n717, in_7, in_6, in_5, gm_n321, gm_n64);
	and (gm_n718, in_11, gm_n52, gm_n51, gm_n717, gm_n48);
	nand (gm_n719, in_15, gm_n50, gm_n49, gm_n718, gm_n46);
	nor (gm_n720, in_19, gm_n47, in_17, gm_n719, gm_n45);
	nand (gm_n721, gm_n720, gm_n71);
	nand (gm_n722, gm_n51, in_8, in_7, gm_n136, gm_n52);
	nor (gm_n723, gm_n49, in_12, gm_n53, gm_n722, gm_n50);
	nand (gm_n724, in_17, in_16, gm_n63, gm_n723, gm_n47);
	nor (gm_n725, gm_n71, in_20, gm_n62, gm_n724);
	or (gm_n726, in_11, in_10, in_9, gm_n607);
	nor (gm_n727, gm_n50, gm_n49, gm_n48, gm_n726, in_15);
	nand (gm_n728, gm_n47, in_17, gm_n46, gm_n727, gm_n62);
	nor (gm_n729, gm_n728, in_21, gm_n45);
	nand (gm_n730, in_9, gm_n64, gm_n55, gm_n66);
	nor (gm_n731, in_12, in_11, in_10, gm_n730, in_13);
	nand (gm_n732, in_16, in_15, gm_n50, gm_n731, in_17);
	nor (gm_n733, gm_n45, gm_n62, gm_n47, gm_n732, gm_n71);
	nand (gm_n734, in_11, gm_n52, gm_n51, gm_n473, gm_n48);
	nor (gm_n735, gm_n63, in_14, in_13, gm_n734, in_16);
	nand (gm_n736, gm_n62, in_18, gm_n81, gm_n735, gm_n45);
	nor (gm_n737, gm_n736, in_21);
	or (gm_n738, gm_n55, gm_n82, gm_n72, gm_n124, gm_n64);
	nor (gm_n739, in_11, in_10, in_9, gm_n738, gm_n48);
	nand (gm_n740, gm_n63, in_14, gm_n49, gm_n739, in_16);
	nor (gm_n741, gm_n62, in_18, in_17, gm_n740, gm_n45);
	nand (gm_n742, gm_n741, in_21);
	nor (gm_n743, gm_n738, gm_n52, in_9);
	nand (gm_n744, gm_n49, gm_n48, in_11, gm_n743, gm_n50);
	nor (gm_n745, in_17, in_16, gm_n63, gm_n744, in_18);
	nand (gm_n746, in_21, in_20, in_19, gm_n745);
	and (gm_n747, in_8, gm_n55, in_6, gm_n638, in_9);
	nand (gm_n748, gm_n48, gm_n53, gm_n52, gm_n747, gm_n49);
	nor (gm_n749, in_16, in_15, in_14, gm_n748, gm_n81);
	nand (gm_n750, in_20, gm_n62, gm_n47, gm_n749, in_21);
	or (gm_n751, gm_n55, in_6, in_5, gm_n643, in_8);
	nor (gm_n752, in_11, gm_n52, gm_n51, gm_n751, gm_n48);
	nand (gm_n753, gm_n63, gm_n50, gm_n49, gm_n752, gm_n46);
	nor (gm_n754, gm_n62, in_18, in_17, gm_n753, in_20);
	nand (gm_n755, gm_n754, gm_n71);
	or (gm_n756, in_1, in_0);
	nor (gm_n757, in_4, gm_n74, gm_n101, gm_n756, in_5);
	nand (gm_n758, in_8, in_7, in_6, gm_n757, gm_n51);
	nor (gm_n759, in_12, gm_n53, in_10, gm_n758, in_13);
	nand (gm_n760, gm_n46, gm_n63, gm_n50, gm_n759, in_17);
	nor (gm_n761, gm_n45, in_19, in_18, gm_n760, in_21);
	or (gm_n762, in_9, gm_n64, in_7, gm_n463, gm_n52);
	nor (gm_n763, gm_n49, gm_n48, gm_n53, gm_n762, gm_n50);
	nand (gm_n764, in_17, in_16, in_15, gm_n763, in_18);
	nor (gm_n765, in_21, gm_n45, in_19, gm_n764);
	or (gm_n766, gm_n64, in_7, gm_n82, gm_n530, in_9);
	nor (gm_n767, gm_n48, gm_n53, in_10, gm_n766, in_13);
	nand (gm_n768, gm_n46, gm_n63, in_14, gm_n767, in_17);
	nor (gm_n769, gm_n45, gm_n62, in_18, gm_n768, in_21);
	nand (gm_n770, in_11, in_10, in_9, gm_n114);
	nor (gm_n771, gm_n50, in_13, gm_n48, gm_n770);
	nand (gm_n772, in_17, in_16, gm_n63, gm_n771, in_18);
	nor (gm_n773, in_21, gm_n45, gm_n62, gm_n772);
	nand (gm_n774, in_7, in_6, gm_n72, gm_n420, gm_n64);
	nor (gm_n775, gm_n53, gm_n52, gm_n51, gm_n774, gm_n48);
	nand (gm_n776, gm_n775, gm_n50, in_13);
	nor (gm_n777, in_17, gm_n46, gm_n63, gm_n776, gm_n47);
	nand (gm_n778, in_21, gm_n45, gm_n62, gm_n777);
	nor (gm_n779, in_9, gm_n64, in_7, gm_n84, in_10);
	nand (gm_n780, gm_n49, gm_n48, gm_n53, gm_n779);
	nor (gm_n781, gm_n46, gm_n63, gm_n50, gm_n780, in_17);
	nand (gm_n782, in_20, in_19, gm_n47, gm_n781, in_21);
	or (gm_n783, gm_n55, in_6, in_5, gm_n167, gm_n64);
	nor (gm_n784, gm_n783, in_9);
	nand (gm_n785, in_12, in_11, gm_n52, gm_n784, gm_n49);
	nor (gm_n786, gm_n46, in_15, gm_n50, gm_n785, in_17);
	nand (gm_n787, in_20, in_19, gm_n47, gm_n786, in_21);
	nand (gm_n788, gm_n64, in_7, in_6, gm_n757, gm_n51);
	nor (gm_n789, gm_n48, gm_n53, gm_n52, gm_n788, in_13);
	and (gm_n790, in_16, gm_n63, gm_n50, gm_n789, gm_n81);
	nand (gm_n791, gm_n45, gm_n62, gm_n47, gm_n790, in_21);
	and (gm_n792, gm_n55, in_6, in_5, gm_n420, in_8);
	and (gm_n793, gm_n53, gm_n52, gm_n51, gm_n792, in_12);
	nand (gm_n794, in_15, in_14, gm_n49, gm_n793, in_16);
	nor (gm_n795, gm_n62, gm_n47, gm_n81, gm_n794, gm_n45);
	nand (gm_n796, gm_n795, gm_n71);
	nand (gm_n797, gm_n787, gm_n782, gm_n778, gm_n796, gm_n791);
	nor (gm_n798, gm_n769, gm_n765, gm_n761, gm_n797, gm_n773);
	nand (gm_n799, gm_n750, gm_n746, gm_n742, gm_n798, gm_n755);
	nor (gm_n800, gm_n733, gm_n729, gm_n725, gm_n799, gm_n737);
	nand (gm_n801, gm_n716, gm_n712, gm_n708, gm_n800, gm_n721);
	nor (gm_n802, gm_n699, gm_n695, gm_n690, gm_n801, gm_n704);
	nand (gm_n803, gm_n681, gm_n677, gm_n672, gm_n802, gm_n685);
	nor (gm_n804, gm_n662, gm_n657, gm_n653, gm_n803, gm_n667);
	nand (gm_n805, gm_n642, gm_n637, gm_n633, gm_n804, gm_n648);
	nor (gm_n806, gm_n625, gm_n620, gm_n616, gm_n805, gm_n629);
	nand (gm_n807, gm_n606, gm_n603, gm_n597, gm_n806, gm_n611);
	nor (gm_n808, gm_n587, gm_n582, gm_n578, gm_n807, gm_n592);
	nand (gm_n809, gm_n570, gm_n565, gm_n561, gm_n808, gm_n575);
	nor (gm_n810, gm_n552, gm_n547, gm_n542, gm_n809, gm_n557);
	nand (gm_n811, gm_n534, gm_n529, gm_n524, gm_n810, gm_n537);
	nor (gm_n812, gm_n513, gm_n508, gm_n503, gm_n811, gm_n518);
	nand (gm_n813, gm_n492, gm_n488, gm_n482, gm_n812, gm_n498);
	nor (gm_n814, gm_n472, gm_n467, gm_n462, gm_n813, gm_n477);
	nand (gm_n815, gm_n452, gm_n448, gm_n444, gm_n814, gm_n457);
	nor (gm_n816, gm_n435, gm_n430, gm_n425, gm_n815, gm_n439);
	nand (gm_n817, gm_n414, gm_n409, gm_n403, gm_n816, gm_n419);
	nor (gm_n818, gm_n394, gm_n388, gm_n383, gm_n817, gm_n399);
	nand (gm_n819, gm_n372, gm_n367, gm_n362, gm_n818, gm_n378);
	nor (gm_n820, gm_n354, gm_n350, gm_n346, gm_n819, gm_n359);
	nand (gm_n821, gm_n337, gm_n332, gm_n326, gm_n820, gm_n342);
	nor (gm_n822, gm_n314, gm_n310, gm_n306, gm_n821, gm_n320);
	nand (gm_n823, gm_n295, gm_n289, gm_n283, gm_n822, gm_n301);
	nor (gm_n824, gm_n274, gm_n271, gm_n267, gm_n823, gm_n278);
	nand (gm_n825, gm_n257, gm_n251, gm_n246, gm_n824, gm_n263);
	nor (gm_n826, gm_n236, gm_n231, gm_n227, gm_n825, gm_n240);
	nand (gm_n827, gm_n217, gm_n214, gm_n208, gm_n826, gm_n222);
	nor (gm_n828, gm_n198, gm_n193, gm_n187, gm_n827, gm_n203);
	nand (gm_n829, gm_n177, gm_n172, gm_n165, gm_n828, gm_n182);
	nor (gm_n830, gm_n155, gm_n149, gm_n145, gm_n829, gm_n160);
	nand (gm_n831, gm_n135, gm_n129, gm_n123, gm_n830, gm_n140);
	nor (gm_n832, gm_n113, gm_n107, gm_n100, gm_n831, gm_n118);
	nand (gm_n833, gm_n88, gm_n80, gm_n70, gm_n832, gm_n94);
	nor (out_0, gm_n833, gm_n61);
	and (gm_n835, gm_n48, in_11, gm_n52, gm_n562, gm_n49);
	nand (gm_n836, in_16, in_15, in_14, gm_n835, in_17);
	nor (gm_n837, in_20, in_19, in_18, gm_n836, in_21);
	nor (gm_n838, gm_n82, gm_n72, gm_n54, gm_n56, in_7);
	and (gm_n839, gm_n52, in_9, in_8, gm_n838, gm_n53);
	nand (gm_n840, gm_n50, gm_n49, gm_n48, gm_n839, gm_n63);
	nor (gm_n841, in_18, in_17, gm_n46, gm_n840, gm_n62);
	nand (gm_n842, gm_n841, gm_n71, in_20);
	nand (gm_n843, gm_n72, in_4, in_3, gm_n83, gm_n82);
	nor (gm_n844, gm_n51, gm_n64, in_7, gm_n843, gm_n52);
	nand (gm_n845, gm_n49, in_12, gm_n53, gm_n844, gm_n50);
	nor (gm_n846, in_17, in_16, gm_n63, gm_n845, in_18);
	nand (gm_n847, in_21, in_20, gm_n62, gm_n846);
	and (gm_n848, in_7, in_6, in_5, gm_n209, in_8);
	and (gm_n849, gm_n53, gm_n52, in_9, gm_n848, gm_n48);
	nand (gm_n850, gm_n63, in_14, gm_n49, gm_n849, gm_n46);
	nor (gm_n851, gm_n62, gm_n47, in_17, gm_n850, gm_n45);
	nand (gm_n852, gm_n851, gm_n71);
	or (gm_n853, in_6, in_5, gm_n54, gm_n56, in_7);
	or (gm_n854, in_10, gm_n51, in_8, gm_n853, in_11);
	or (gm_n855, gm_n50, gm_n49, in_12, gm_n854, gm_n63);
	nor (gm_n856, in_18, in_17, gm_n46, gm_n855, in_19);
	nand (gm_n857, gm_n856, gm_n71, in_20);
	nor (gm_n858, gm_n55, gm_n82, gm_n72, gm_n108, in_8);
	nand (gm_n859, gm_n858, gm_n52, in_9);
	nor (gm_n860, gm_n49, in_12, gm_n53, gm_n859, gm_n50);
	nand (gm_n861, in_17, in_16, in_15, gm_n860, gm_n47);
	nor (gm_n862, in_21, gm_n45, in_19, gm_n861);
	nand (gm_n863, gm_n64, in_7, gm_n82, gm_n379, in_9);
	nor (gm_n864, in_12, gm_n53, in_10, gm_n863, gm_n49);
	nand (gm_n865, in_16, gm_n63, in_14, gm_n864, gm_n81);
	nor (gm_n866, gm_n45, gm_n62, in_18, gm_n865, gm_n71);
	nand (gm_n867, in_2, gm_n166, in_0, gm_n54, in_3);
	nor (gm_n868, in_7, gm_n82, gm_n72, gm_n867, gm_n64);
	nand (gm_n869, in_11, gm_n52, in_9, gm_n868);
	nor (gm_n870, in_14, in_13, in_12, gm_n869, gm_n63);
	nand (gm_n871, in_18, in_17, in_16, gm_n870, in_19);
	nor (gm_n872, gm_n871, in_21, gm_n45);
	or (gm_n873, gm_n55, gm_n82, in_5, gm_n167, gm_n64);
	nor (gm_n874, gm_n53, gm_n52, in_9, gm_n873);
	and (gm_n875, gm_n50, in_13, gm_n48, gm_n874, gm_n63);
	nand (gm_n876, gm_n47, gm_n81, gm_n46, gm_n875, gm_n62);
	nor (gm_n877, gm_n876, gm_n71, in_20);
	nand (gm_n878, gm_n48, gm_n53, in_10, gm_n120, gm_n49);
	nor (gm_n879, in_16, in_15, in_14, gm_n878, gm_n81);
	nand (gm_n880, in_20, gm_n62, in_18, gm_n879, gm_n71);
	nor (gm_n881, gm_n52, in_9, in_8, gm_n478);
	nand (gm_n882, in_13, gm_n48, gm_n53, gm_n881, in_14);
	nor (gm_n883, gm_n81, in_16, in_15, gm_n882, in_18);
	nand (gm_n884, gm_n71, gm_n45, gm_n62, gm_n883);
	nor (gm_n885, gm_n751, in_9);
	nand (gm_n886, in_12, gm_n53, gm_n52, gm_n885, in_13);
	nor (gm_n887, in_16, gm_n63, in_14, gm_n886, in_17);
	nand (gm_n888, gm_n45, in_19, in_18, gm_n887, gm_n71);
	nor (gm_n889, in_8, in_7, gm_n82, gm_n119, in_9);
	nand (gm_n890, in_12, gm_n53, gm_n52, gm_n889, in_13);
	nor (gm_n891, gm_n46, in_15, in_14, gm_n890, gm_n81);
	nand (gm_n892, gm_n45, in_19, gm_n47, gm_n891, gm_n71);
	nand (gm_n893, gm_n64, gm_n55, gm_n82, gm_n757, gm_n51);
	nor (gm_n894, gm_n48, in_11, in_10, gm_n893, in_13);
	nand (gm_n895, in_16, in_15, gm_n50, gm_n894, in_17);
	nor (gm_n896, in_20, gm_n62, gm_n47, gm_n895, in_21);
	nand (gm_n897, in_5, gm_n54, gm_n74, gm_n258, gm_n82);
	or (gm_n898, in_9, gm_n64, gm_n55, gm_n897);
	nor (gm_n899, in_12, gm_n53, in_10, gm_n898, in_13);
	nand (gm_n900, in_16, gm_n63, in_14, gm_n899, in_17);
	nor (gm_n901, gm_n45, in_19, gm_n47, gm_n900, gm_n71);
	nor (gm_n902, in_7, in_6, gm_n72, gm_n75, in_8);
	and (gm_n903, gm_n902, in_10, gm_n51);
	nand (gm_n904, in_13, in_12, gm_n53, gm_n903);
	or (gm_n905, in_16, gm_n63, gm_n50, gm_n904, gm_n81);
	nor (gm_n906, gm_n45, gm_n62, in_18, gm_n905, gm_n71);
	or (gm_n907, in_6, gm_n72, gm_n54, gm_n56, in_7);
	nor (gm_n908, gm_n52, in_9, gm_n64, gm_n907, gm_n53);
	and (gm_n909, gm_n50, gm_n49, gm_n48, gm_n908, in_15);
	nand (gm_n910, gm_n47, gm_n81, gm_n46, gm_n909, gm_n62);
	nor (gm_n911, gm_n910, gm_n71, gm_n45);
	nor (gm_n912, gm_n64, in_7, gm_n82, gm_n204, in_9);
	nand (gm_n913, in_12, gm_n53, gm_n52, gm_n912, in_13);
	nor (gm_n914, gm_n46, gm_n63, gm_n50, gm_n913, gm_n81);
	nand (gm_n915, gm_n45, gm_n62, gm_n47, gm_n914, gm_n71);
	nand (gm_n916, in_7, in_6, in_5, gm_n252, in_8);
	nor (gm_n917, in_11, in_10, in_9, gm_n916, gm_n48);
	nand (gm_n918, gm_n63, in_14, in_13, gm_n917, in_16);
	nor (gm_n919, gm_n62, gm_n47, in_17, gm_n918, in_20);
	nand (gm_n920, gm_n919, in_21);
	nor (gm_n921, gm_n55, in_6, in_5, gm_n867);
	nand (gm_n922, gm_n52, gm_n51, gm_n64, gm_n921, gm_n53);
	nor (gm_n923, gm_n922, gm_n49, gm_n48);
	and (gm_n924, gm_n46, in_15, in_14, gm_n923, in_17);
	nand (gm_n925, gm_n45, in_19, gm_n47, gm_n924, in_21);
	nand (gm_n926, gm_n48, in_11, in_10, gm_n157, gm_n49);
	nor (gm_n927, gm_n46, gm_n63, gm_n50, gm_n926, in_17);
	nand (gm_n928, in_20, in_19, in_18, gm_n927, gm_n71);
	and (gm_n929, in_7, gm_n82, gm_n72, gm_n89, in_8);
	nand (gm_n930, gm_n929, in_9);
	nor (gm_n931, gm_n48, in_11, in_10, gm_n930, gm_n49);
	nand (gm_n932, gm_n46, in_15, gm_n50, gm_n931, gm_n81);
	nor (gm_n933, gm_n45, in_19, in_18, gm_n932, gm_n71);
	nor (gm_n934, in_8, in_7, gm_n82, gm_n156, gm_n51);
	and (gm_n935, in_12, in_11, gm_n52, gm_n934, in_13);
	nand (gm_n936, in_16, in_15, in_14, gm_n935, gm_n81);
	nor (gm_n937, gm_n45, gm_n62, gm_n47, gm_n936, in_21);
	or (gm_n938, gm_n51, gm_n64, gm_n55, gm_n897, in_10);
	nor (gm_n939, in_13, gm_n48, in_11, gm_n938, in_14);
	nand (gm_n940, in_17, gm_n46, gm_n63, gm_n939, in_18);
	nor (gm_n941, gm_n71, in_20, in_19, gm_n940);
	or (gm_n942, gm_n51, in_8, gm_n55, gm_n897, in_10);
	nor (gm_n943, in_13, gm_n48, in_11, gm_n942, in_14);
	nand (gm_n944, in_17, in_16, in_15, gm_n943, in_18);
	nor (gm_n945, gm_n71, gm_n45, in_19, gm_n944);
	and (gm_n946, gm_n64, gm_n55, in_6, gm_n757, gm_n51);
	nand (gm_n947, gm_n48, gm_n53, in_10, gm_n946, in_13);
	nor (gm_n948, gm_n46, in_15, in_14, gm_n947, gm_n81);
	nand (gm_n949, in_20, gm_n62, gm_n47, gm_n948, in_21);
	or (gm_n950, gm_n55, gm_n82, gm_n72, gm_n167, gm_n64);
	nor (gm_n951, gm_n53, gm_n52, in_9, gm_n950, in_12);
	nand (gm_n952, gm_n951, gm_n50, in_13);
	nor (gm_n953, gm_n81, gm_n46, in_15, gm_n952, in_18);
	nand (gm_n954, gm_n71, in_20, in_19, gm_n953);
	or (gm_n955, gm_n55, gm_n82, gm_n72, gm_n643, gm_n64);
	nor (gm_n956, in_11, gm_n52, gm_n51, gm_n955);
	nand (gm_n957, gm_n50, in_13, in_12, gm_n956, in_15);
	nor (gm_n958, in_18, in_17, gm_n46, gm_n957, gm_n62);
	nand (gm_n959, gm_n958, gm_n71, in_20);
	nand (gm_n960, gm_n55, in_6, gm_n72, gm_n296, gm_n64);
	nor (gm_n961, gm_n53, in_10, in_9, gm_n960);
	nand (gm_n962, gm_n50, in_13, in_12, gm_n961, in_15);
	nor (gm_n963, in_18, in_17, in_16, gm_n962, in_19);
	nand (gm_n964, gm_n963, in_21, in_20);
	nor (gm_n965, in_12, gm_n53, gm_n52, gm_n510, gm_n49);
	nand (gm_n966, in_16, gm_n63, in_14, gm_n965, in_17);
	nor (gm_n967, gm_n45, in_19, gm_n47, gm_n966, gm_n71);
	nor (gm_n968, gm_n64, in_7, in_6, gm_n141, in_9);
	and (gm_n969, in_12, gm_n53, gm_n52, gm_n968, gm_n49);
	nand (gm_n970, gm_n46, in_15, in_14, gm_n969, in_17);
	nor (gm_n971, gm_n45, gm_n62, gm_n47, gm_n970, in_21);
	nor (gm_n972, in_8, in_7, gm_n82, gm_n141, in_9);
	and (gm_n973, gm_n48, in_11, in_10, gm_n972, gm_n49);
	nand (gm_n974, in_16, in_15, in_14, gm_n973, in_17);
	nor (gm_n975, gm_n45, gm_n62, gm_n47, gm_n974, in_21);
	nor (gm_n976, in_11, gm_n52, in_9, gm_n960, in_12);
	and (gm_n977, in_15, gm_n50, gm_n49, gm_n976, in_16);
	nand (gm_n978, gm_n62, in_18, gm_n81, gm_n977, gm_n45);
	nor (gm_n979, gm_n978, gm_n71);
	nor (gm_n980, in_8, in_7, in_6, gm_n161, in_9);
	and (gm_n981, in_12, in_11, gm_n52, gm_n980, gm_n49);
	and (gm_n982, in_16, gm_n63, gm_n50, gm_n981, in_17);
	nand (gm_n983, gm_n45, in_19, gm_n47, gm_n982, in_21);
	nor (gm_n984, gm_n53, gm_n52, gm_n51, gm_n686, gm_n48);
	nand (gm_n985, gm_n63, gm_n50, gm_n49, gm_n984, gm_n46);
	nor (gm_n986, gm_n62, in_18, in_17, gm_n985, in_20);
	nand (gm_n987, gm_n986, in_21);
	nor (gm_n988, gm_n64, gm_n55, in_6, gm_n161, in_9);
	nand (gm_n989, gm_n988, gm_n52);
	or (gm_n990, gm_n49, gm_n48, gm_n53, gm_n989, in_14);
	nor (gm_n991, in_17, in_16, gm_n63, gm_n990, gm_n47);
	nand (gm_n992, in_21, gm_n45, gm_n62, gm_n991);
	nor (gm_n993, gm_n53, in_10, gm_n51, gm_n328, gm_n48);
	nand (gm_n994, gm_n993, in_14, gm_n49);
	nor (gm_n995, gm_n81, gm_n46, in_15, gm_n994, in_18);
	nand (gm_n996, in_21, in_20, in_19, gm_n995);
	nor (gm_n997, gm_n55, in_6, in_5, gm_n321, gm_n64);
	and (gm_n998, gm_n997, gm_n52, gm_n51);
	and (gm_n999, in_13, gm_n48, in_11, gm_n998, gm_n50);
	nand (gm_n1000, in_17, in_16, gm_n63, gm_n999, in_18);
	nor (gm_n1001, in_21, in_20, in_19, gm_n1000);
	nor (gm_n1002, gm_n55, gm_n82, in_5, gm_n643, in_8);
	nand (gm_n1003, gm_n1002, gm_n52, in_9);
	nor (gm_n1004, in_13, gm_n48, gm_n53, gm_n1003, gm_n50);
	nand (gm_n1005, gm_n81, in_16, gm_n63, gm_n1004, in_18);
	nor (gm_n1006, gm_n71, in_20, in_19, gm_n1005);
	nor (gm_n1007, in_5, gm_n54, gm_n74, gm_n150, gm_n82);
	nand (gm_n1008, gm_n51, in_8, gm_n55, gm_n1007, in_10);
	nor (gm_n1009, gm_n49, gm_n48, in_11, gm_n1008, in_14);
	nand (gm_n1010, in_17, gm_n46, gm_n63, gm_n1009, in_18);
	nor (gm_n1011, gm_n71, gm_n45, gm_n62, gm_n1010);
	nand (gm_n1012, in_11, in_10, in_9, gm_n355, in_12);
	nor (gm_n1013, gm_n63, in_14, in_13, gm_n1012, gm_n46);
	nand (gm_n1014, in_19, in_18, in_17, gm_n1013, gm_n45);
	nor (gm_n1015, gm_n1014, gm_n71);
	and (gm_n1016, gm_n53, in_10, gm_n51, gm_n858);
	nand (gm_n1017, gm_n50, gm_n49, in_12, gm_n1016, in_15);
	nor (gm_n1018, gm_n47, in_17, gm_n46, gm_n1017, in_19);
	nand (gm_n1019, gm_n1018, gm_n71, in_20);
	nand (gm_n1020, gm_n48, in_11, in_10, gm_n912, gm_n49);
	nor (gm_n1021, gm_n46, in_15, gm_n50, gm_n1020, in_17);
	nand (gm_n1022, gm_n45, gm_n62, gm_n47, gm_n1021, gm_n71);
	nand (gm_n1023, gm_n55, gm_n82, gm_n72, gm_n296, gm_n64);
	or (gm_n1024, gm_n1023, gm_n52, gm_n51);
	nor (gm_n1025, gm_n49, in_12, gm_n53, gm_n1024, gm_n50);
	and (gm_n1026, gm_n81, gm_n46, in_15, gm_n1025, gm_n47);
	nand (gm_n1027, in_21, gm_n45, in_19, gm_n1026);
	nand (gm_n1028, in_12, gm_n53, in_10, gm_n339, gm_n49);
	nor (gm_n1029, in_16, gm_n63, in_14, gm_n1028, gm_n81);
	nand (gm_n1030, gm_n45, in_19, in_18, gm_n1029, gm_n71);
	nand (gm_n1031, gm_n242, in_10, in_9);
	nor (gm_n1032, gm_n49, in_12, gm_n53, gm_n1031, gm_n50);
	nand (gm_n1033, in_17, in_16, in_15, gm_n1032, in_18);
	nor (gm_n1034, gm_n71, in_20, in_19, gm_n1033);
	nand (gm_n1035, gm_n55, in_6, gm_n72, gm_n209, gm_n64);
	nor (gm_n1036, gm_n1035, in_10, in_9);
	and (gm_n1037, in_13, gm_n48, in_11, gm_n1036, gm_n50);
	nand (gm_n1038, gm_n81, in_16, in_15, gm_n1037, gm_n47);
	nor (gm_n1039, in_21, gm_n45, gm_n62, gm_n1038);
	nand (gm_n1040, in_11, in_10, gm_n51, gm_n232, gm_n48);
	nor (gm_n1041, gm_n63, in_14, in_13, gm_n1040, gm_n46);
	nand (gm_n1042, in_19, gm_n47, in_17, gm_n1041, gm_n45);
	nor (gm_n1043, gm_n1042, gm_n71);
	and (gm_n1044, in_7, in_6, in_5, gm_n493, in_8);
	nand (gm_n1045, in_11, in_10, gm_n51, gm_n1044, in_12);
	nor (gm_n1046, in_15, gm_n50, gm_n49, gm_n1045, gm_n46);
	nand (gm_n1047, gm_n62, in_18, in_17, gm_n1046, gm_n45);
	nor (gm_n1048, gm_n1047, in_21);
	nand (gm_n1049, in_13, in_12, in_11, gm_n844, gm_n50);
	nor (gm_n1050, in_17, in_16, in_15, gm_n1049, gm_n47);
	nand (gm_n1051, gm_n71, in_20, gm_n62, gm_n1050);
	nand (gm_n1052, in_7, in_6, in_5, gm_n420, gm_n64);
	nor (gm_n1053, gm_n1052, gm_n52, gm_n51);
	nand (gm_n1054, in_13, in_12, gm_n53, gm_n1053, gm_n50);
	nor (gm_n1055, gm_n81, in_16, gm_n63, gm_n1054, gm_n47);
	nand (gm_n1056, gm_n71, gm_n45, gm_n62, gm_n1055);
	and (gm_n1057, in_7, gm_n82, in_5, gm_n420, in_8);
	and (gm_n1058, gm_n1057, in_10, in_9);
	nand (gm_n1059, in_13, in_12, in_11, gm_n1058, in_14);
	nor (gm_n1060, gm_n81, in_16, gm_n63, gm_n1059, gm_n47);
	nand (gm_n1061, gm_n71, in_20, gm_n62, gm_n1060);
	nor (gm_n1062, in_9, in_8, gm_n55, gm_n843, in_10);
	nand (gm_n1063, gm_n49, gm_n48, in_11, gm_n1062, in_14);
	nor (gm_n1064, gm_n81, gm_n46, gm_n63, gm_n1063, in_18);
	nand (gm_n1065, in_21, gm_n45, in_19, gm_n1064);
	nand (gm_n1066, gm_n53, gm_n52, gm_n51, gm_n210);
	nor (gm_n1067, gm_n1066, gm_n49, in_12);
	nand (gm_n1068, gm_n46, in_15, in_14, gm_n1067, in_17);
	nor (gm_n1069, gm_n45, in_19, gm_n47, gm_n1068, in_21);
	nor (gm_n1070, gm_n55, gm_n82, in_5, gm_n130, gm_n64);
	nand (gm_n1071, in_11, in_10, gm_n51, gm_n1070);
	nor (gm_n1072, gm_n50, in_13, gm_n48, gm_n1071, gm_n63);
	nand (gm_n1073, in_18, gm_n81, in_16, gm_n1072, in_19);
	nor (gm_n1074, gm_n1073, in_21, gm_n45);
	nor (gm_n1075, in_4, gm_n74, gm_n101, gm_n756, gm_n72);
	nand (gm_n1076, in_8, gm_n55, in_6, gm_n1075, in_9);
	nor (gm_n1077, in_12, gm_n53, in_10, gm_n1076, in_13);
	nand (gm_n1078, gm_n46, gm_n63, in_14, gm_n1077, gm_n81);
	nor (gm_n1079, gm_n45, in_19, gm_n47, gm_n1078, in_21);
	and (gm_n1080, in_8, gm_n55, in_6, gm_n374, gm_n51);
	and (gm_n1081, gm_n48, in_11, in_10, gm_n1080, in_13);
	nand (gm_n1082, in_16, gm_n63, gm_n50, gm_n1081, gm_n81);
	nor (gm_n1083, in_20, gm_n62, in_18, gm_n1082, gm_n71);
	nor (gm_n1084, in_11, gm_n52, gm_n51, gm_n183, gm_n48);
	nand (gm_n1085, in_15, in_14, in_13, gm_n1084, in_16);
	nor (gm_n1086, gm_n62, gm_n47, in_17, gm_n1085, in_20);
	nand (gm_n1087, gm_n1086, gm_n71);
	nor (gm_n1088, gm_n82, gm_n72, in_4, gm_n315, in_7);
	and (gm_n1089, gm_n52, in_9, in_8, gm_n1088, gm_n53);
	nand (gm_n1090, in_14, gm_n49, gm_n48, gm_n1089, in_15);
	nor (gm_n1091, in_18, gm_n81, in_16, gm_n1090, gm_n62);
	nand (gm_n1092, gm_n1091, in_21, gm_n45);
	nor (gm_n1093, in_7, gm_n82, in_5, gm_n167);
	and (gm_n1094, gm_n52, gm_n51, gm_n64, gm_n1093);
	nand (gm_n1095, in_13, in_12, gm_n53, gm_n1094, in_14);
	nor (gm_n1096, in_17, gm_n46, gm_n63, gm_n1095, in_18);
	nand (gm_n1097, in_21, gm_n45, in_19, gm_n1096);
	nand (gm_n1098, in_7, in_6, gm_n72, gm_n241, in_8);
	nor (gm_n1099, gm_n1098, in_10, in_9);
	nand (gm_n1100, in_13, in_12, in_11, gm_n1099, gm_n50);
	nor (gm_n1101, gm_n81, in_16, in_15, gm_n1100, in_18);
	nand (gm_n1102, gm_n71, in_20, in_19, gm_n1101);
	or (gm_n1103, gm_n52, in_9, gm_n64, gm_n853, gm_n53);
	nor (gm_n1104, gm_n50, in_13, in_12, gm_n1103, in_15);
	nand (gm_n1105, in_18, gm_n81, in_16, gm_n1104, in_19);
	nor (gm_n1106, gm_n1105, gm_n71, gm_n45);
	and (gm_n1107, gm_n792, in_10, in_9);
	and (gm_n1108, gm_n49, gm_n48, gm_n53, gm_n1107, in_14);
	nand (gm_n1109, in_17, in_16, gm_n63, gm_n1108, in_18);
	nor (gm_n1110, in_21, in_20, gm_n62, gm_n1109);
	nor (gm_n1111, in_7, gm_n82, in_5, gm_n290, gm_n64);
	nand (gm_n1112, in_11, gm_n52, in_9, gm_n1111, in_12);
	nor (gm_n1113, gm_n1112, in_13);
	nand (gm_n1114, gm_n46, gm_n63, gm_n50, gm_n1113, gm_n81);
	nor (gm_n1115, in_20, gm_n62, gm_n47, gm_n1114, gm_n71);
	and (gm_n1116, in_7, gm_n82, gm_n72, gm_n420, gm_n64);
	nand (gm_n1117, gm_n1116, in_9);
	nor (gm_n1118, gm_n48, in_11, in_10, gm_n1117, in_13);
	nand (gm_n1119, gm_n46, gm_n63, gm_n50, gm_n1118, gm_n81);
	nor (gm_n1120, in_20, in_19, in_18, gm_n1119, in_21);
	nand (gm_n1121, in_7, gm_n82, gm_n72, gm_n296, in_8);
	nor (gm_n1122, gm_n53, gm_n52, in_9, gm_n1121);
	nand (gm_n1123, gm_n50, in_13, in_12, gm_n1122, gm_n63);
	nor (gm_n1124, gm_n47, in_17, gm_n46, gm_n1123, gm_n62);
	nand (gm_n1125, gm_n1124, gm_n71, gm_n45);
	nor (gm_n1126, in_2, in_1, gm_n73, in_4, in_3);
	nand (gm_n1127, in_7, in_6, gm_n72, gm_n1126, gm_n64);
	nor (gm_n1128, gm_n1127, in_9);
	nand (gm_n1129, in_12, in_11, in_10, gm_n1128, gm_n49);
	nor (gm_n1130, gm_n46, gm_n63, gm_n50, gm_n1129, gm_n81);
	nand (gm_n1131, gm_n45, in_19, in_18, gm_n1130, in_21);
	nor (gm_n1132, gm_n46, gm_n63, gm_n50, gm_n913, in_17);
	nand (gm_n1133, in_20, gm_n62, gm_n47, gm_n1132, in_21);
	and (gm_n1134, gm_n55, gm_n82, in_5, gm_n420, gm_n64);
	and (gm_n1135, gm_n1134, in_10, gm_n51);
	nand (gm_n1136, gm_n49, gm_n48, gm_n53, gm_n1135, gm_n50);
	nor (gm_n1137, in_17, gm_n46, in_15, gm_n1136, gm_n47);
	nand (gm_n1138, gm_n71, in_20, in_19, gm_n1137);
	nor (gm_n1139, in_12, in_11, gm_n52, gm_n930, in_13);
	nand (gm_n1140, gm_n46, gm_n63, gm_n50, gm_n1139, gm_n81);
	nor (gm_n1141, in_20, in_19, in_18, gm_n1140, gm_n71);
	nor (gm_n1142, in_7, gm_n82, in_5, gm_n75, gm_n64);
	nand (gm_n1143, gm_n53, in_10, gm_n51, gm_n1142, gm_n48);
	nor (gm_n1144, in_15, gm_n50, in_13, gm_n1143, gm_n46);
	nand (gm_n1145, gm_n62, gm_n47, gm_n81, gm_n1144, in_20);
	nor (gm_n1146, gm_n1145, gm_n71);
	nor (gm_n1147, in_7, in_6, gm_n72, gm_n483, in_8);
	and (gm_n1148, in_11, in_10, gm_n51, gm_n1147, in_12);
	and (gm_n1149, in_15, in_14, gm_n49, gm_n1148);
	nand (gm_n1150, gm_n47, in_17, in_16, gm_n1149, in_19);
	nor (gm_n1151, gm_n1150, in_21, in_20);
	nand (gm_n1152, gm_n431, gm_n51, gm_n64);
	nor (gm_n1153, gm_n48, gm_n53, gm_n52, gm_n1152, gm_n49);
	nand (gm_n1154, in_16, in_15, in_14, gm_n1153, in_17);
	nor (gm_n1155, gm_n45, gm_n62, gm_n47, gm_n1154, in_21);
	and (gm_n1156, in_7, in_6, gm_n72, gm_n493, gm_n64);
	and (gm_n1157, in_11, in_10, in_9, gm_n1156, gm_n48);
	nand (gm_n1158, in_15, gm_n50, gm_n49, gm_n1157, in_16);
	nor (gm_n1159, in_19, in_18, gm_n81, gm_n1158, gm_n45);
	nand (gm_n1160, gm_n1159, in_21);
	nor (gm_n1161, gm_n51, gm_n64, gm_n55, gm_n259, in_10);
	nand (gm_n1162, gm_n49, gm_n48, gm_n53, gm_n1161, in_14);
	nor (gm_n1163, in_17, in_16, gm_n63, gm_n1162, gm_n47);
	nand (gm_n1164, in_21, gm_n45, gm_n62, gm_n1163);
	and (gm_n1165, in_7, in_6, in_5, gm_n209, gm_n64);
	and (gm_n1166, gm_n53, in_10, gm_n51, gm_n1165, in_12);
	nand (gm_n1167, in_15, gm_n50, in_13, gm_n1166, in_16);
	nor (gm_n1168, gm_n62, in_18, gm_n81, gm_n1167, in_20);
	nand (gm_n1169, gm_n1168, gm_n71);
	nor (gm_n1170, in_9, gm_n64, gm_n55, gm_n463);
	nand (gm_n1171, in_12, in_11, in_10, gm_n1170, in_13);
	nor (gm_n1172, in_16, gm_n63, gm_n50, gm_n1171, gm_n81);
	nand (gm_n1173, gm_n45, in_19, in_18, gm_n1172, in_21);
	or (gm_n1174, gm_n64, in_7, gm_n82, gm_n161, in_9);
	nor (gm_n1175, in_12, in_11, gm_n52, gm_n1174, in_13);
	nand (gm_n1176, in_16, gm_n63, gm_n50, gm_n1175, in_17);
	nor (gm_n1177, gm_n45, in_19, in_18, gm_n1176, in_21);
	nor (gm_n1178, in_7, gm_n82, in_5, gm_n321, gm_n64);
	nand (gm_n1179, gm_n1178, in_10, in_9);
	nor (gm_n1180, in_13, gm_n48, in_11, gm_n1179, in_14);
	nand (gm_n1181, in_17, in_16, in_15, gm_n1180, gm_n47);
	nor (gm_n1182, in_21, gm_n45, gm_n62, gm_n1181);
	and (gm_n1183, gm_n55, gm_n82, gm_n72, gm_n241, gm_n64);
	nand (gm_n1184, in_11, gm_n52, gm_n51, gm_n1183, in_12);
	nor (gm_n1185, gm_n63, in_14, gm_n49, gm_n1184, in_16);
	nand (gm_n1186, gm_n62, gm_n47, in_17, gm_n1185, gm_n45);
	nor (gm_n1187, gm_n1186, in_21);
	and (gm_n1188, in_11, in_10, in_9, gm_n997);
	and (gm_n1189, gm_n50, gm_n49, in_12, gm_n1188, in_15);
	nand (gm_n1190, gm_n47, gm_n81, in_16, gm_n1189, gm_n62);
	nor (gm_n1191, gm_n1190, in_21, in_20);
	nor (gm_n1192, in_7, gm_n82, gm_n72, gm_n130, in_8);
	nand (gm_n1193, in_11, in_10, in_9, gm_n1192);
	or (gm_n1194, in_14, gm_n49, gm_n48, gm_n1193, in_15);
	nor (gm_n1195, in_18, gm_n81, in_16, gm_n1194, gm_n62);
	nand (gm_n1196, gm_n1195, in_21, in_20);
	nor (gm_n1197, gm_n53, in_10, in_9, gm_n520, gm_n48);
	nand (gm_n1198, gm_n63, gm_n50, in_13, gm_n1197, gm_n46);
	nor (gm_n1199, in_19, gm_n47, gm_n81, gm_n1198, in_20);
	nand (gm_n1200, gm_n1199, gm_n71);
	nor (gm_n1201, in_8, gm_n55, in_6, gm_n161, in_9);
	nand (gm_n1202, in_12, gm_n53, gm_n52, gm_n1201, in_13);
	nor (gm_n1203, gm_n46, gm_n63, gm_n50, gm_n1202, gm_n81);
	nand (gm_n1204, gm_n45, in_19, in_18, gm_n1203, in_21);
	or (gm_n1205, in_12, in_11, gm_n52, gm_n264, gm_n49);
	nor (gm_n1206, in_16, gm_n63, in_14, gm_n1205, gm_n81);
	nand (gm_n1207, gm_n45, gm_n62, in_18, gm_n1206, gm_n71);
	nand (gm_n1208, in_10, gm_n51, in_8, gm_n316);
	nor (gm_n1209, gm_n49, gm_n48, gm_n53, gm_n1208, gm_n50);
	nand (gm_n1210, in_17, gm_n46, in_15, gm_n1209, gm_n47);
	nor (gm_n1211, gm_n71, gm_n45, in_19, gm_n1210);
	nor (gm_n1212, in_7, gm_n82, gm_n72, gm_n108, gm_n64);
	and (gm_n1213, in_11, gm_n52, gm_n51, gm_n1212);
	and (gm_n1214, in_14, in_13, gm_n48, gm_n1213, gm_n63);
	and (gm_n1215, in_18, gm_n81, in_16, gm_n1214, in_19);
	and (gm_n1216, gm_n1215, gm_n71, in_20);
	or (gm_n1217, in_7, in_6, gm_n72, gm_n124, in_8);
	or (gm_n1218, in_11, in_10, in_9, gm_n1217, in_12);
	nor (gm_n1219, in_15, in_14, in_13, gm_n1218, in_16);
	nand (gm_n1220, gm_n62, gm_n47, in_17, gm_n1219, gm_n45);
	nor (gm_n1221, gm_n1220, in_21);
	and (gm_n1222, in_7, in_6, in_5, gm_n241, gm_n64);
	and (gm_n1223, in_11, in_10, gm_n51, gm_n1222);
	and (gm_n1224, gm_n50, gm_n49, in_12, gm_n1223, gm_n63);
	nand (gm_n1225, in_18, gm_n81, gm_n46, gm_n1224, in_19);
	nor (gm_n1226, gm_n1225, in_21, in_20);
	nor (gm_n1227, in_8, gm_n55, gm_n82, gm_n156, gm_n51);
	nand (gm_n1228, in_12, gm_n53, in_10, gm_n1227, gm_n49);
	nor (gm_n1229, in_16, in_15, in_14, gm_n1228, gm_n81);
	nand (gm_n1230, in_20, in_19, in_18, gm_n1229, gm_n71);
	nor (gm_n1231, gm_n64, gm_n55, in_6, gm_n103, gm_n51);
	nand (gm_n1232, gm_n48, gm_n53, in_10, gm_n1231, in_13);
	nor (gm_n1233, gm_n46, in_15, in_14, gm_n1232, in_17);
	nand (gm_n1234, gm_n45, in_19, in_18, gm_n1233, gm_n71);
	and (gm_n1235, gm_n51, in_8, in_7, gm_n504, in_10);
	nand (gm_n1236, gm_n49, in_12, in_11, gm_n1235, in_14);
	nor (gm_n1237, in_17, gm_n46, in_15, gm_n1236, gm_n47);
	nand (gm_n1238, gm_n71, in_20, in_19, gm_n1237);
	nand (gm_n1239, in_7, gm_n82, gm_n72, gm_n89, gm_n64);
	nor (gm_n1240, gm_n1239, in_10, gm_n51);
	nand (gm_n1241, in_13, in_12, gm_n53, gm_n1240, in_14);
	nor (gm_n1242, in_17, in_16, in_15, gm_n1241, gm_n47);
	nand (gm_n1243, gm_n71, gm_n45, gm_n62, gm_n1242);
	nor (gm_n1244, gm_n49, in_12, in_11, gm_n464, gm_n50);
	nand (gm_n1245, in_17, gm_n46, gm_n63, gm_n1244, in_18);
	nor (gm_n1246, gm_n71, gm_n45, in_19, gm_n1245);
	nand (gm_n1247, in_7, in_6, in_5, gm_n89, gm_n64);
	nor (gm_n1248, in_11, gm_n52, in_9, gm_n1247, gm_n48);
	and (gm_n1249, gm_n1248, in_13);
	nand (gm_n1250, gm_n46, gm_n63, in_14, gm_n1249, in_17);
	nor (gm_n1251, in_20, in_19, gm_n47, gm_n1250, gm_n71);
	nand (gm_n1252, gm_n593, gm_n51);
	nor (gm_n1253, in_12, in_11, gm_n52, gm_n1252, in_13);
	nand (gm_n1254, gm_n46, in_15, gm_n50, gm_n1253, in_17);
	nor (gm_n1255, in_20, gm_n62, in_18, gm_n1254, gm_n71);
	nand (gm_n1256, gm_n72, gm_n54, in_3, gm_n83, gm_n82);
	nor (gm_n1257, gm_n51, in_8, in_7, gm_n1256, in_10);
	and (gm_n1258, gm_n49, in_12, in_11, gm_n1257, gm_n50);
	nand (gm_n1259, in_17, in_16, gm_n63, gm_n1258, in_18);
	nor (gm_n1260, gm_n71, gm_n45, gm_n62, gm_n1259);
	nand (gm_n1261, gm_n55, gm_n82, in_5, gm_n598, in_8);
	nor (gm_n1262, gm_n1261, gm_n51);
	nand (gm_n1263, in_12, in_11, gm_n52, gm_n1262, gm_n49);
	nor (gm_n1264, gm_n46, gm_n63, in_14, gm_n1263, in_17);
	nand (gm_n1265, in_20, gm_n62, gm_n47, gm_n1264, gm_n71);
	nor (gm_n1266, in_11, in_10, gm_n51, gm_n395, gm_n48);
	nand (gm_n1267, in_15, gm_n50, in_13, gm_n1266, in_16);
	nor (gm_n1268, gm_n62, in_18, gm_n81, gm_n1267, in_20);
	nand (gm_n1269, gm_n1268, gm_n71);
	and (gm_n1270, gm_n53, in_10, in_9, gm_n1212, gm_n48);
	nand (gm_n1271, gm_n63, in_14, gm_n49, gm_n1270, in_16);
	nor (gm_n1272, in_19, gm_n47, gm_n81, gm_n1271, in_20);
	nand (gm_n1273, gm_n1272, gm_n71);
	nor (gm_n1274, gm_n55, in_6, gm_n72, gm_n483, gm_n64);
	and (gm_n1275, gm_n53, in_10, gm_n51, gm_n1274, in_12);
	nand (gm_n1276, in_15, in_14, gm_n49, gm_n1275, gm_n46);
	nor (gm_n1277, gm_n62, in_18, gm_n81, gm_n1276, gm_n45);
	nand (gm_n1278, gm_n1277, in_21);
	nor (gm_n1279, gm_n55, in_6, gm_n72, gm_n188, gm_n64);
	nand (gm_n1280, gm_n1279, gm_n51);
	nor (gm_n1281, in_12, in_11, in_10, gm_n1280, gm_n49);
	nand (gm_n1282, in_16, gm_n63, in_14, gm_n1281, in_17);
	nor (gm_n1283, gm_n45, in_19, gm_n47, gm_n1282, gm_n71);
	nor (gm_n1284, in_7, in_6, gm_n72, gm_n75, gm_n64);
	nand (gm_n1285, in_11, gm_n52, in_9, gm_n1284, in_12);
	nor (gm_n1286, in_15, in_14, in_13, gm_n1285, gm_n46);
	nand (gm_n1287, in_19, in_18, gm_n81, gm_n1286, in_20);
	nor (gm_n1288, gm_n1287, gm_n71);
	or (gm_n1289, gm_n453, in_10, gm_n51);
	nor (gm_n1290, in_13, in_12, in_11, gm_n1289, gm_n50);
	nand (gm_n1291, in_17, in_16, in_15, gm_n1290, in_18);
	nor (gm_n1292, in_21, in_20, in_19, gm_n1291);
	nor (gm_n1293, in_7, gm_n82, gm_n72, gm_n130, gm_n64);
	nand (gm_n1294, gm_n53, in_10, in_9, gm_n1293, gm_n48);
	nor (gm_n1295, in_15, gm_n50, in_13, gm_n1294, gm_n46);
	nand (gm_n1296, gm_n62, gm_n47, gm_n81, gm_n1295, in_20);
	nor (gm_n1297, gm_n1296, gm_n71);
	and (gm_n1298, gm_n51, gm_n64, in_7, gm_n66, in_10);
	nand (gm_n1299, in_13, gm_n48, gm_n53, gm_n1298, gm_n50);
	nor (gm_n1300, in_17, gm_n46, in_15, gm_n1299, gm_n47);
	nand (gm_n1301, in_21, gm_n45, gm_n62, gm_n1300);
	nor (gm_n1302, in_7, gm_n82, in_5, gm_n643, in_8);
	and (gm_n1303, in_11, gm_n52, in_9, gm_n1302);
	nand (gm_n1304, in_14, in_13, gm_n48, gm_n1303, in_15);
	nor (gm_n1305, in_18, gm_n81, gm_n46, gm_n1304, gm_n62);
	nand (gm_n1306, gm_n1305, in_21, in_20);
	and (gm_n1307, gm_n64, in_7, in_6, gm_n757, in_9);
	nand (gm_n1308, in_12, gm_n53, in_10, gm_n1307, gm_n49);
	nor (gm_n1309, gm_n46, in_15, in_14, gm_n1308, gm_n81);
	nand (gm_n1310, gm_n45, in_19, in_18, gm_n1309, in_21);
	nor (gm_n1311, gm_n950, in_10, in_9);
	nand (gm_n1312, gm_n49, gm_n48, in_11, gm_n1311);
	nor (gm_n1313, gm_n46, in_15, in_14, gm_n1312, gm_n81);
	nand (gm_n1314, gm_n45, in_19, gm_n47, gm_n1313, gm_n71);
	nor (gm_n1315, in_7, in_6, in_5, gm_n108, in_8);
	nand (gm_n1316, gm_n53, in_10, gm_n51, gm_n1315, in_12);
	nor (gm_n1317, gm_n63, in_14, gm_n49, gm_n1316, in_16);
	nand (gm_n1318, in_19, gm_n47, in_17, gm_n1317, in_20);
	nor (gm_n1319, gm_n1318, in_21);
	nand (gm_n1320, gm_n53, gm_n52, gm_n51, gm_n1183);
	nor (gm_n1321, gm_n50, gm_n49, in_12, gm_n1320, gm_n63);
	nand (gm_n1322, gm_n47, gm_n81, in_16, gm_n1321, in_19);
	nor (gm_n1323, gm_n1322, gm_n71, gm_n45);
	or (gm_n1324, in_9, in_8, in_7, gm_n553, in_10);
	nor (gm_n1325, gm_n49, in_12, gm_n53, gm_n1324, gm_n50);
	nand (gm_n1326, in_17, gm_n46, in_15, gm_n1325, in_18);
	nor (gm_n1327, gm_n71, in_20, in_19, gm_n1326);
	and (gm_n1328, gm_n52, gm_n51, in_8, gm_n838);
	and (gm_n1329, gm_n49, in_12, gm_n53, gm_n1328, in_14);
	nand (gm_n1330, in_17, in_16, in_15, gm_n1329, gm_n47);
	nor (gm_n1331, gm_n71, gm_n45, in_19, gm_n1330);
	nor (gm_n1332, in_8, in_7, in_6, gm_n103, in_9);
	nand (gm_n1333, in_12, in_11, in_10, gm_n1332, in_13);
	nor (gm_n1334, gm_n46, in_15, gm_n50, gm_n1333, in_17);
	nand (gm_n1335, in_20, in_19, gm_n47, gm_n1334, in_21);
	and (gm_n1336, gm_n48, in_11, in_10, gm_n784, in_13);
	and (gm_n1337, gm_n46, in_15, gm_n50, gm_n1336, in_17);
	nand (gm_n1338, gm_n45, in_19, gm_n47, gm_n1337, gm_n71);
	and (gm_n1339, in_7, in_6, gm_n72, gm_n420, in_8);
	and (gm_n1340, in_11, in_10, in_9, gm_n1339);
	nand (gm_n1341, in_14, in_13, gm_n48, gm_n1340, gm_n63);
	nor (gm_n1342, gm_n47, gm_n81, in_16, gm_n1341, in_19);
	nand (gm_n1343, gm_n1342, in_21, in_20);
	nor (gm_n1344, gm_n51, in_8, in_7, gm_n525, gm_n52);
	nand (gm_n1345, gm_n49, gm_n48, in_11, gm_n1344, gm_n50);
	nor (gm_n1346, in_17, in_16, gm_n63, gm_n1345, in_18);
	nand (gm_n1347, gm_n71, gm_n45, gm_n62, gm_n1346);
	or (gm_n1348, gm_n53, gm_n52, in_9, gm_n178);
	nor (gm_n1349, in_14, in_13, gm_n48, gm_n1348, in_15);
	nand (gm_n1350, in_18, gm_n81, in_16, gm_n1349, in_19);
	nor (gm_n1351, gm_n1350, gm_n71, in_20);
	nand (gm_n1352, gm_n53, in_10, gm_n51, gm_n1274, gm_n48);
	nor (gm_n1353, in_15, in_14, gm_n49, gm_n1352, gm_n46);
	nand (gm_n1354, gm_n62, gm_n47, gm_n81, gm_n1353, gm_n45);
	nor (gm_n1355, gm_n1354, in_21);
	nand (gm_n1356, gm_n64, in_7, in_6, gm_n1075, in_9);
	nor (gm_n1357, in_12, gm_n53, in_10, gm_n1356, in_13);
	nand (gm_n1358, gm_n46, in_15, in_14, gm_n1357, gm_n81);
	nor (gm_n1359, in_20, in_19, gm_n47, gm_n1358, gm_n71);
	nor (gm_n1360, gm_n55, gm_n82, gm_n72, gm_n321, in_8);
	nand (gm_n1361, gm_n53, in_10, gm_n51, gm_n1360, in_12);
	nor (gm_n1362, in_15, gm_n50, gm_n49, gm_n1361, in_16);
	nand (gm_n1363, in_19, gm_n47, in_17, gm_n1362, gm_n45);
	nor (gm_n1364, gm_n1363, gm_n71);
	nor (gm_n1365, gm_n64, gm_n55, gm_n82, gm_n96, in_9);
	nand (gm_n1366, in_12, in_11, gm_n52, gm_n1365, in_13);
	nor (gm_n1367, gm_n46, gm_n63, in_14, gm_n1366, in_17);
	nand (gm_n1368, in_20, in_19, in_18, gm_n1367, gm_n71);
	nand (gm_n1369, in_12, gm_n53, in_10, gm_n1201, in_13);
	nor (gm_n1370, gm_n46, in_15, gm_n50, gm_n1369, gm_n81);
	nand (gm_n1371, gm_n45, in_19, gm_n47, gm_n1370, in_21);
	nand (gm_n1372, gm_n64, gm_n55, gm_n82, gm_n1075, in_9);
	or (gm_n1373, in_12, gm_n53, in_10, gm_n1372, gm_n49);
	nor (gm_n1374, in_16, gm_n63, in_14, gm_n1373, in_17);
	nand (gm_n1375, gm_n45, in_19, gm_n47, gm_n1374, in_21);
	and (gm_n1376, gm_n51, in_8, gm_n55, gm_n504);
	nand (gm_n1377, gm_n48, gm_n53, in_10, gm_n1376, gm_n49);
	nor (gm_n1378, in_16, gm_n63, in_14, gm_n1377, gm_n81);
	nand (gm_n1379, gm_n45, in_19, in_18, gm_n1378, gm_n71);
	nor (gm_n1380, in_7, in_6, in_5, gm_n867, gm_n64);
	nand (gm_n1381, gm_n1380, in_10, in_9);
	nor (gm_n1382, in_13, gm_n48, in_11, gm_n1381, gm_n50);
	nand (gm_n1383, in_17, gm_n46, gm_n63, gm_n1382, in_18);
	nor (gm_n1384, gm_n71, gm_n45, gm_n62, gm_n1383);
	nor (gm_n1385, gm_n64, in_7, in_6, gm_n530, in_9);
	and (gm_n1386, gm_n48, gm_n53, in_10, gm_n1385, in_13);
	nand (gm_n1387, gm_n46, gm_n63, gm_n50, gm_n1386, in_17);
	nor (gm_n1388, in_20, gm_n62, gm_n47, gm_n1387, in_21);
	nand (gm_n1389, in_11, in_10, in_9, gm_n1293, gm_n48);
	nor (gm_n1390, gm_n1389, gm_n49);
	nand (gm_n1391, in_16, gm_n63, gm_n50, gm_n1390, gm_n81);
	nor (gm_n1392, in_20, in_19, in_18, gm_n1391, gm_n71);
	nand (gm_n1393, in_7, gm_n82, gm_n72, gm_n284, in_8);
	nor (gm_n1394, gm_n1393, in_9);
	and (gm_n1395, gm_n48, in_11, gm_n52, gm_n1394, gm_n49);
	nand (gm_n1396, in_16, in_15, in_14, gm_n1395, gm_n81);
	nor (gm_n1397, gm_n45, gm_n62, in_18, gm_n1396, in_21);
	or (gm_n1398, gm_n64, in_7, in_6, gm_n119, in_9);
	or (gm_n1399, in_12, gm_n53, gm_n52, gm_n1398, gm_n49);
	nor (gm_n1400, in_16, gm_n63, gm_n50, gm_n1399, in_17);
	nand (gm_n1401, gm_n45, gm_n62, gm_n47, gm_n1400, in_21);
	nor (gm_n1402, in_11, gm_n52, gm_n51, gm_n960, in_12);
	nand (gm_n1403, in_15, gm_n50, in_13, gm_n1402, in_16);
	nor (gm_n1404, in_19, gm_n47, in_17, gm_n1403, gm_n45);
	nand (gm_n1405, gm_n1404, gm_n71);
	nor (gm_n1406, in_8, gm_n55, gm_n82, gm_n161, gm_n51);
	nand (gm_n1407, gm_n48, gm_n53, in_10, gm_n1406, in_13);
	nor (gm_n1408, gm_n46, gm_n63, in_14, gm_n1407, gm_n81);
	nand (gm_n1409, gm_n45, gm_n62, gm_n47, gm_n1408, gm_n71);
	nand (gm_n1410, in_12, gm_n53, gm_n52, gm_n142, in_13);
	nor (gm_n1411, gm_n46, gm_n63, gm_n50, gm_n1410, gm_n81);
	nand (gm_n1412, in_20, in_19, in_18, gm_n1411, gm_n71);
	nor (gm_n1413, gm_n64, in_7, in_6, gm_n119, gm_n51);
	and (gm_n1414, gm_n48, in_11, in_10, gm_n1413, gm_n49);
	nand (gm_n1415, gm_n46, in_15, gm_n50, gm_n1414, in_17);
	nor (gm_n1416, gm_n45, gm_n62, in_18, gm_n1415, in_21);
	nand (gm_n1417, gm_n53, gm_n52, gm_n51, gm_n297, in_12);
	nor (gm_n1418, gm_n63, in_14, in_13, gm_n1417, in_16);
	nand (gm_n1419, in_19, gm_n47, gm_n81, gm_n1418, in_20);
	nor (gm_n1420, gm_n1419, in_21);
	nor (gm_n1421, gm_n55, in_6, gm_n72, gm_n167, in_8);
	nand (gm_n1422, in_11, gm_n52, gm_n51, gm_n1421, gm_n48);
	nor (gm_n1423, gm_n63, in_14, gm_n49, gm_n1422, gm_n46);
	nand (gm_n1424, gm_n62, in_18, in_17, gm_n1423, in_20);
	nor (gm_n1425, gm_n1424, in_21);
	and (gm_n1426, gm_n49, in_12, in_11, gm_n137, gm_n50);
	nand (gm_n1427, in_17, gm_n46, in_15, gm_n1426, in_18);
	nor (gm_n1428, in_21, in_20, gm_n62, gm_n1427);
	nand (gm_n1429, in_4, in_3, in_2, gm_n95, gm_n72);
	or (gm_n1430, gm_n64, in_7, in_6, gm_n1429, gm_n51);
	or (gm_n1431, gm_n48, gm_n53, gm_n52, gm_n1430, in_13);
	nor (gm_n1432, in_16, gm_n63, in_14, gm_n1431, in_17);
	nand (gm_n1433, gm_n45, in_19, in_18, gm_n1432, in_21);
	nand (gm_n1434, in_7, in_6, gm_n72, gm_n89, in_8);
	nor (gm_n1435, gm_n1434, in_10, in_9);
	nand (gm_n1436, gm_n49, in_12, gm_n53, gm_n1435, in_14);
	nor (gm_n1437, in_17, in_16, gm_n63, gm_n1436, gm_n47);
	nand (gm_n1438, gm_n71, gm_n45, in_19, gm_n1437);
	nand (gm_n1439, gm_n55, in_6, gm_n72, gm_n284, gm_n64);
	nor (gm_n1440, gm_n1439, gm_n51);
	nand (gm_n1441, gm_n48, gm_n53, in_10, gm_n1440, in_13);
	nor (gm_n1442, gm_n46, gm_n63, gm_n50, gm_n1441, in_17);
	nand (gm_n1443, in_20, gm_n62, gm_n47, gm_n1442, in_21);
	and (gm_n1444, gm_n53, gm_n52, in_9, gm_n355);
	nand (gm_n1445, in_14, gm_n49, gm_n48, gm_n1444, gm_n63);
	nor (gm_n1446, gm_n47, gm_n81, in_16, gm_n1445, in_19);
	nand (gm_n1447, gm_n1446, gm_n71, in_20);
	nand (gm_n1448, gm_n53, gm_n52, in_9, gm_n1156, in_12);
	nor (gm_n1449, in_15, gm_n50, in_13, gm_n1448, gm_n46);
	nand (gm_n1450, in_19, in_18, in_17, gm_n1449, in_20);
	nor (gm_n1451, gm_n1450, gm_n71);
	or (gm_n1452, gm_n64, gm_n55, in_6, gm_n96, gm_n51);
	nor (gm_n1453, gm_n48, in_11, in_10, gm_n1452, in_13);
	nand (gm_n1454, in_16, gm_n63, in_14, gm_n1453, in_17);
	nor (gm_n1455, gm_n45, gm_n62, gm_n47, gm_n1454, gm_n71);
	nor (gm_n1456, gm_n50, in_13, in_12, gm_n922, gm_n63);
	nand (gm_n1457, in_18, in_17, gm_n46, gm_n1456, gm_n62);
	nor (gm_n1458, gm_n1457, gm_n71, gm_n45);
	and (gm_n1459, gm_n55, gm_n82, in_5, gm_n241, gm_n64);
	nand (gm_n1460, gm_n53, gm_n52, in_9, gm_n1459);
	nor (gm_n1461, gm_n50, gm_n49, gm_n48, gm_n1460, gm_n63);
	nand (gm_n1462, gm_n47, gm_n81, in_16, gm_n1461, gm_n62);
	nor (gm_n1463, gm_n1462, gm_n71, in_20);
	nand (gm_n1464, in_7, gm_n82, in_5, gm_n493, gm_n64);
	nor (gm_n1465, in_11, gm_n52, gm_n51, gm_n1464, gm_n48);
	nand (gm_n1466, gm_n1465, in_13);
	nor (gm_n1467, in_16, gm_n63, in_14, gm_n1466, in_17);
	nand (gm_n1468, gm_n45, in_19, in_18, gm_n1467, gm_n71);
	nor (gm_n1469, gm_n55, gm_n82, gm_n72, gm_n124, in_8);
	and (gm_n1470, gm_n53, in_10, in_9, gm_n1469);
	nand (gm_n1471, gm_n50, gm_n49, gm_n48, gm_n1470);
	nor (gm_n1472, in_17, gm_n46, gm_n63, gm_n1471, in_18);
	nand (gm_n1473, in_21, in_20, in_19, gm_n1472);
	nand (gm_n1474, gm_n55, in_6, gm_n72, gm_n493, gm_n64);
	nor (gm_n1475, gm_n53, gm_n52, in_9, gm_n1474, gm_n48);
	nand (gm_n1476, gm_n63, gm_n50, in_13, gm_n1475, gm_n46);
	nor (gm_n1477, gm_n1476, in_18, in_17);
	nand (gm_n1478, gm_n71, in_20, gm_n62, gm_n1477);
	nor (gm_n1479, gm_n46, gm_n63, in_14, gm_n255, gm_n81);
	nand (gm_n1480, gm_n45, in_19, in_18, gm_n1479, gm_n71);
	or (gm_n1481, in_7, in_6, in_5, gm_n643, in_8);
	nor (gm_n1482, in_11, gm_n52, in_9, gm_n1481, in_12);
	nand (gm_n1483, in_15, in_14, gm_n49, gm_n1482, gm_n46);
	nor (gm_n1484, gm_n62, gm_n47, gm_n81, gm_n1483, gm_n45);
	nand (gm_n1485, gm_n1484, in_21);
	nand (gm_n1486, gm_n1478, gm_n1473, gm_n1468, gm_n1485, gm_n1480);
	nor (gm_n1487, gm_n1458, gm_n1455, gm_n1451, gm_n1486, gm_n1463);
	nand (gm_n1488, gm_n1443, gm_n1438, gm_n1433, gm_n1487, gm_n1447);
	nor (gm_n1489, gm_n1425, gm_n1420, gm_n1416, gm_n1488, gm_n1428);
	nand (gm_n1490, gm_n1409, gm_n1405, gm_n1401, gm_n1489, gm_n1412);
	nor (gm_n1491, gm_n1392, gm_n1388, gm_n1384, gm_n1490, gm_n1397);
	nand (gm_n1492, gm_n1375, gm_n1371, gm_n1368, gm_n1491, gm_n1379);
	nor (gm_n1493, gm_n1359, gm_n1355, gm_n1351, gm_n1492, gm_n1364);
	nand (gm_n1494, gm_n1343, gm_n1338, gm_n1335, gm_n1493, gm_n1347);
	nor (gm_n1495, gm_n1327, gm_n1323, gm_n1319, gm_n1494, gm_n1331);
	nand (gm_n1496, gm_n1310, gm_n1306, gm_n1301, gm_n1495, gm_n1314);
	nor (gm_n1497, gm_n1292, gm_n1288, gm_n1283, gm_n1496, gm_n1297);
	nand (gm_n1498, gm_n1273, gm_n1269, gm_n1265, gm_n1497, gm_n1278);
	nor (gm_n1499, gm_n1255, gm_n1251, gm_n1246, gm_n1498, gm_n1260);
	nand (gm_n1500, gm_n1238, gm_n1234, gm_n1230, gm_n1499, gm_n1243);
	nor (gm_n1501, gm_n1221, gm_n1216, gm_n1211, gm_n1500, gm_n1226);
	nand (gm_n1502, gm_n1204, gm_n1200, gm_n1196, gm_n1501, gm_n1207);
	nor (gm_n1503, gm_n1187, gm_n1182, gm_n1177, gm_n1502, gm_n1191);
	nand (gm_n1504, gm_n1169, gm_n1164, gm_n1160, gm_n1503, gm_n1173);
	nor (gm_n1505, gm_n1151, gm_n1146, gm_n1141, gm_n1504, gm_n1155);
	nand (gm_n1506, gm_n1133, gm_n1131, gm_n1125, gm_n1505, gm_n1138);
	nor (gm_n1507, gm_n1115, gm_n1110, gm_n1106, gm_n1506, gm_n1120);
	nand (gm_n1508, gm_n1097, gm_n1092, gm_n1087, gm_n1507, gm_n1102);
	nor (gm_n1509, gm_n1079, gm_n1074, gm_n1069, gm_n1508, gm_n1083);
	nand (gm_n1510, gm_n1061, gm_n1056, gm_n1051, gm_n1509, gm_n1065);
	nor (gm_n1511, gm_n1043, gm_n1039, gm_n1034, gm_n1510, gm_n1048);
	nand (gm_n1512, gm_n1027, gm_n1022, gm_n1019, gm_n1511, gm_n1030);
	nor (gm_n1513, gm_n1011, gm_n1006, gm_n1001, gm_n1512, gm_n1015);
	nand (gm_n1514, gm_n992, gm_n987, gm_n983, gm_n1513, gm_n996);
	nor (gm_n1515, gm_n975, gm_n971, gm_n967, gm_n1514, gm_n979);
	nand (gm_n1516, gm_n959, gm_n954, gm_n949, gm_n1515, gm_n964);
	nor (gm_n1517, gm_n941, gm_n937, gm_n933, gm_n1516, gm_n945);
	nand (gm_n1518, gm_n925, gm_n920, gm_n915, gm_n1517, gm_n928);
	nor (gm_n1519, gm_n906, gm_n901, gm_n896, gm_n1518, gm_n911);
	nand (gm_n1520, gm_n888, gm_n884, gm_n880, gm_n1519, gm_n892);
	nor (gm_n1521, gm_n872, gm_n866, gm_n862, gm_n1520, gm_n877);
	nand (gm_n1522, gm_n852, gm_n847, gm_n842, gm_n1521, gm_n857);
	nor (out_1, gm_n1522, gm_n837);
	nand (gm_n1524, in_8, in_7, gm_n82, gm_n374, gm_n51);
	nor (gm_n1525, gm_n48, gm_n53, in_10, gm_n1524, gm_n49);
	nand (gm_n1526, gm_n46, gm_n63, gm_n50, gm_n1525, in_17);
	nor (gm_n1527, gm_n45, gm_n62, in_18, gm_n1526, gm_n71);
	nor (gm_n1528, in_7, in_6, in_5, gm_n75, in_8);
	and (gm_n1529, gm_n53, in_10, gm_n51, gm_n1528, gm_n48);
	and (gm_n1530, gm_n1529, gm_n49);
	and (gm_n1531, gm_n46, gm_n63, in_14, gm_n1530, in_17);
	nand (gm_n1532, gm_n45, gm_n62, in_18, gm_n1531, gm_n71);
	nand (gm_n1533, gm_n55, in_6, in_5, gm_n296, gm_n64);
	nor (gm_n1534, gm_n53, in_10, gm_n51, gm_n1533, in_12);
	nand (gm_n1535, in_15, gm_n50, in_13, gm_n1534, in_16);
	nor (gm_n1536, in_19, gm_n47, in_17, gm_n1535, in_20);
	nand (gm_n1537, gm_n1536, gm_n71);
	nor (gm_n1538, in_10, in_9, gm_n64, gm_n478);
	nand (gm_n1539, gm_n49, in_12, gm_n53, gm_n1538, in_14);
	nor (gm_n1540, in_17, in_16, in_15, gm_n1539, in_18);
	nand (gm_n1541, gm_n71, in_20, in_19, gm_n1540);
	and (gm_n1542, in_10, in_9, gm_n64, gm_n1088);
	nand (gm_n1543, gm_n49, in_12, in_11, gm_n1542, gm_n50);
	nor (gm_n1544, gm_n81, gm_n46, gm_n63, gm_n1543, in_18);
	nand (gm_n1545, in_21, in_20, gm_n62, gm_n1544);
	nand (gm_n1546, in_11, gm_n52, in_9, gm_n644);
	nor (gm_n1547, in_14, gm_n49, gm_n48, gm_n1546, in_15);
	nand (gm_n1548, in_18, gm_n81, in_16, gm_n1547, in_19);
	nor (gm_n1549, gm_n1548, gm_n71, in_20);
	and (gm_n1550, in_7, in_6, in_5, gm_n296, in_8);
	and (gm_n1551, gm_n1550, in_10, gm_n51);
	and (gm_n1552, gm_n49, gm_n48, in_11, gm_n1551, gm_n50);
	nand (gm_n1553, gm_n81, in_16, in_15, gm_n1552, gm_n47);
	nor (gm_n1554, in_21, in_20, in_19, gm_n1553);
	nor (gm_n1555, in_7, gm_n82, gm_n72, gm_n483, in_8);
	and (gm_n1556, in_11, in_10, in_9, gm_n1555, in_12);
	and (gm_n1557, in_15, in_14, gm_n49, gm_n1556, gm_n46);
	nand (gm_n1558, in_19, in_18, in_17, gm_n1557, gm_n45);
	nor (gm_n1559, gm_n1558, gm_n71);
	nor (gm_n1560, in_13, in_12, in_11, gm_n445, in_14);
	nand (gm_n1561, in_17, gm_n46, in_15, gm_n1560, gm_n47);
	nor (gm_n1562, in_21, gm_n45, in_19, gm_n1561);
	nor (gm_n1563, gm_n55, gm_n82, gm_n72, gm_n290, in_8);
	and (gm_n1564, in_11, in_10, gm_n51, gm_n1563, gm_n48);
	nand (gm_n1565, in_15, in_14, in_13, gm_n1564, in_16);
	nor (gm_n1566, in_19, gm_n47, gm_n81, gm_n1565, in_20);
	nand (gm_n1567, gm_n1566, in_21);
	nor (gm_n1568, in_11, gm_n52, gm_n51, gm_n583, gm_n48);
	nand (gm_n1569, gm_n1568, in_13);
	nor (gm_n1570, gm_n46, in_15, in_14, gm_n1569, gm_n81);
	nand (gm_n1571, gm_n45, in_19, in_18, gm_n1570, gm_n71);
	and (gm_n1572, in_7, in_6, in_5, gm_n284, gm_n64);
	and (gm_n1573, in_11, gm_n52, in_9, gm_n1572, gm_n48);
	and (gm_n1574, gm_n1573, gm_n49);
	and (gm_n1575, gm_n46, gm_n63, in_14, gm_n1574, gm_n81);
	nand (gm_n1576, gm_n45, gm_n62, in_18, gm_n1575, gm_n71);
	nand (gm_n1577, in_11, gm_n52, in_9, gm_n1293, gm_n48);
	or (gm_n1578, gm_n63, gm_n50, gm_n49, gm_n1577, gm_n46);
	nor (gm_n1579, in_19, gm_n47, in_17, gm_n1578, in_20);
	nand (gm_n1580, gm_n1579, gm_n71);
	nand (gm_n1581, gm_n46, gm_n63, gm_n50, gm_n923, gm_n81);
	nor (gm_n1582, in_20, in_19, in_18, gm_n1581, gm_n71);
	nor (gm_n1583, in_7, gm_n82, gm_n72, gm_n643, in_8);
	and (gm_n1584, gm_n1583, in_10, gm_n51);
	and (gm_n1585, gm_n49, gm_n48, gm_n53, gm_n1584, in_14);
	nand (gm_n1586, in_17, gm_n46, in_15, gm_n1585, in_18);
	nor (gm_n1587, gm_n71, gm_n45, in_19, gm_n1586);
	nand (gm_n1588, gm_n51, gm_n64, in_7, gm_n404, gm_n52);
	nor (gm_n1589, in_13, in_12, in_11, gm_n1588, in_14);
	nand (gm_n1590, gm_n81, gm_n46, in_15, gm_n1589, gm_n47);
	nor (gm_n1591, gm_n71, in_20, in_19, gm_n1590);
	and (gm_n1592, gm_n49, in_12, in_11, gm_n1240, gm_n50);
	nand (gm_n1593, gm_n81, gm_n46, in_15, gm_n1592, in_18);
	nor (gm_n1594, gm_n71, gm_n45, in_19, gm_n1593);
	nand (gm_n1595, in_11, in_10, in_9, gm_n902, gm_n48);
	or (gm_n1596, gm_n63, in_14, gm_n49, gm_n1595, in_16);
	nor (gm_n1597, in_19, gm_n47, gm_n81, gm_n1596, gm_n45);
	nand (gm_n1598, gm_n1597, gm_n71);
	or (gm_n1599, gm_n64, in_7, gm_n82, gm_n199, gm_n51);
	or (gm_n1600, gm_n48, in_11, gm_n52, gm_n1599, gm_n49);
	nor (gm_n1601, in_16, in_15, gm_n50, gm_n1600, in_17);
	nand (gm_n1602, in_20, gm_n62, in_18, gm_n1601, in_21);
	nor (gm_n1603, gm_n55, gm_n82, in_5, gm_n130, in_8);
	and (gm_n1604, gm_n53, gm_n52, gm_n51, gm_n1603);
	nand (gm_n1605, in_14, gm_n49, gm_n48, gm_n1604, in_15);
	nor (gm_n1606, gm_n47, gm_n81, in_16, gm_n1605, in_19);
	nand (gm_n1607, gm_n1606, in_21, in_20);
	nor (gm_n1608, gm_n82, in_5, in_4, gm_n315, gm_n55);
	and (gm_n1609, gm_n52, gm_n51, in_8, gm_n1608);
	nand (gm_n1610, gm_n49, gm_n48, gm_n53, gm_n1609, gm_n50);
	nor (gm_n1611, gm_n81, in_16, gm_n63, gm_n1610, in_18);
	nand (gm_n1612, gm_n71, in_20, in_19, gm_n1611);
	nand (gm_n1613, gm_n53, gm_n52, in_9, gm_n1555, in_12);
	nor (gm_n1614, in_15, in_14, in_13, gm_n1613, in_16);
	nand (gm_n1615, gm_n62, in_18, in_17, gm_n1614, in_20);
	nor (gm_n1616, gm_n1615, gm_n71);
	nand (gm_n1617, gm_n57, in_9, gm_n64);
	nor (gm_n1618, in_12, gm_n53, gm_n52, gm_n1617, in_13);
	nand (gm_n1619, in_16, gm_n63, gm_n50, gm_n1618, gm_n81);
	nor (gm_n1620, gm_n45, gm_n62, in_18, gm_n1619, in_21);
	nand (gm_n1621, in_9, in_8, in_7, gm_n504);
	nor (gm_n1622, in_12, in_11, gm_n52, gm_n1621, in_13);
	nand (gm_n1623, in_16, in_15, gm_n50, gm_n1622, in_17);
	nor (gm_n1624, gm_n45, gm_n62, in_18, gm_n1623, in_21);
	nand (gm_n1625, in_11, gm_n52, in_9, gm_n109);
	nor (gm_n1626, gm_n50, gm_n49, gm_n48, gm_n1625, gm_n63);
	nand (gm_n1627, in_18, gm_n81, gm_n46, gm_n1626, in_19);
	nor (gm_n1628, gm_n1627, in_21, gm_n45);
	nand (gm_n1629, in_7, in_6, gm_n72, gm_n209, in_8);
	nor (gm_n1630, in_11, in_10, in_9, gm_n1629, gm_n48);
	nand (gm_n1631, gm_n63, in_14, in_13, gm_n1630, in_16);
	nor (gm_n1632, gm_n62, gm_n47, gm_n81, gm_n1631, gm_n45);
	nand (gm_n1633, gm_n1632, gm_n71);
	nor (gm_n1634, in_7, gm_n82, in_5, gm_n867, in_8);
	and (gm_n1635, gm_n53, gm_n52, in_9, gm_n1634, in_12);
	nand (gm_n1636, in_15, in_14, gm_n49, gm_n1635, gm_n46);
	nor (gm_n1637, in_19, gm_n47, in_17, gm_n1636, in_20);
	nand (gm_n1638, gm_n1637, gm_n71);
	nor (gm_n1639, in_11, in_10, gm_n51, gm_n285, in_12);
	and (gm_n1640, gm_n63, gm_n50, gm_n49, gm_n1639, gm_n46);
	and (gm_n1641, gm_n1640, gm_n47, in_17);
	nand (gm_n1642, in_21, gm_n45, gm_n62, gm_n1641);
	and (gm_n1643, gm_n55, gm_n82, in_5, gm_n493, in_8);
	and (gm_n1644, gm_n1643, in_10, gm_n51);
	nand (gm_n1645, in_13, gm_n48, gm_n53, gm_n1644, in_14);
	nor (gm_n1646, gm_n81, in_16, in_15, gm_n1645, in_18);
	nand (gm_n1647, gm_n71, gm_n45, in_19, gm_n1646);
	or (gm_n1648, gm_n51, in_8, in_7, gm_n1256, gm_n52);
	nor (gm_n1649, in_13, gm_n48, in_11, gm_n1648, gm_n50);
	nand (gm_n1650, gm_n81, in_16, in_15, gm_n1649, gm_n47);
	nor (gm_n1651, in_21, in_20, in_19, gm_n1650);
	nor (gm_n1652, gm_n51, gm_n64, gm_n55, gm_n84, in_10);
	and (gm_n1653, gm_n49, in_12, in_11, gm_n1652);
	nand (gm_n1654, gm_n46, in_15, gm_n50, gm_n1653, gm_n81);
	nor (gm_n1655, in_20, in_19, in_18, gm_n1654, gm_n71);
	nand (gm_n1656, in_11, in_10, gm_n51, gm_n668, gm_n48);
	nor (gm_n1657, in_15, gm_n50, in_13, gm_n1656, gm_n46);
	nand (gm_n1658, in_19, in_18, in_17, gm_n1657, in_20);
	nor (gm_n1659, gm_n1658, gm_n71);
	nand (gm_n1660, gm_n53, gm_n52, gm_n51, gm_n1315, in_12);
	nor (gm_n1661, gm_n63, gm_n50, gm_n49, gm_n1660, in_16);
	nand (gm_n1662, gm_n62, gm_n47, gm_n81, gm_n1661, gm_n45);
	nor (gm_n1663, gm_n1662, in_21);
	nand (gm_n1664, gm_n49, gm_n48, gm_n53, gm_n881, in_14);
	nor (gm_n1665, in_17, gm_n46, in_15, gm_n1664, gm_n47);
	nand (gm_n1666, gm_n71, in_20, in_19, gm_n1665);
	and (gm_n1667, in_11, gm_n52, gm_n51, gm_n1603, in_12);
	nand (gm_n1668, gm_n63, in_14, in_13, gm_n1667, gm_n46);
	nor (gm_n1669, in_19, in_18, gm_n81, gm_n1668, gm_n45);
	nand (gm_n1670, gm_n1669, gm_n71);
	nor (gm_n1671, in_8, in_7, in_6, gm_n119, in_9);
	nand (gm_n1672, in_12, in_11, gm_n52, gm_n1671, in_13);
	nor (gm_n1673, in_16, gm_n63, in_14, gm_n1672, gm_n81);
	nand (gm_n1674, in_20, gm_n62, gm_n47, gm_n1673, in_21);
	nor (gm_n1675, gm_n64, in_7, gm_n82, gm_n141, in_9);
	nand (gm_n1676, in_12, in_11, in_10, gm_n1675, gm_n49);
	nor (gm_n1677, gm_n46, gm_n63, in_14, gm_n1676, gm_n81);
	nand (gm_n1678, gm_n45, in_19, gm_n47, gm_n1677, gm_n71);
	or (gm_n1679, in_8, gm_n55, in_6, gm_n1429, gm_n51);
	nor (gm_n1680, gm_n48, gm_n53, gm_n52, gm_n1679, in_13);
	nand (gm_n1681, in_16, in_15, gm_n50, gm_n1680, gm_n81);
	nor (gm_n1682, gm_n45, in_19, gm_n47, gm_n1681, in_21);
	nor (gm_n1683, gm_n55, in_6, gm_n72, gm_n130, in_8);
	nand (gm_n1684, gm_n1683, in_9);
	nor (gm_n1685, in_12, in_11, gm_n52, gm_n1684, gm_n49);
	nand (gm_n1686, gm_n46, in_15, in_14, gm_n1685, gm_n81);
	nor (gm_n1687, in_20, gm_n62, in_18, gm_n1686, gm_n71);
	nor (gm_n1688, gm_n64, gm_n55, gm_n82, gm_n161, in_9);
	and (gm_n1689, in_12, in_11, gm_n52, gm_n1688, in_13);
	nand (gm_n1690, in_16, gm_n63, gm_n50, gm_n1689, gm_n81);
	nor (gm_n1691, in_20, gm_n62, gm_n47, gm_n1690, in_21);
	nor (gm_n1692, gm_n64, in_7, in_6, gm_n1429, in_9);
	and (gm_n1693, in_12, gm_n53, gm_n52, gm_n1692, gm_n49);
	nand (gm_n1694, in_16, gm_n63, gm_n50, gm_n1693, in_17);
	nor (gm_n1695, gm_n45, gm_n62, in_18, gm_n1694, in_21);
	nor (gm_n1696, in_10, in_9, in_8, gm_n853);
	nand (gm_n1697, in_13, gm_n48, in_11, gm_n1696, in_14);
	nor (gm_n1698, in_17, gm_n46, in_15, gm_n1697, gm_n47);
	nand (gm_n1699, gm_n71, in_20, gm_n62, gm_n1698);
	nor (gm_n1700, gm_n64, gm_n55, gm_n82, gm_n156, in_9);
	nand (gm_n1701, in_12, gm_n53, gm_n52, gm_n1700, in_13);
	nor (gm_n1702, gm_n46, gm_n63, in_14, gm_n1701, in_17);
	nand (gm_n1703, gm_n45, gm_n62, gm_n47, gm_n1702, gm_n71);
	and (gm_n1704, gm_n55, gm_n82, gm_n72, gm_n284, in_8);
	and (gm_n1705, in_11, in_10, in_9, gm_n1704, in_12);
	nand (gm_n1706, gm_n63, gm_n50, in_13, gm_n1705, gm_n46);
	nor (gm_n1707, gm_n62, gm_n47, gm_n81, gm_n1706, gm_n45);
	nand (gm_n1708, gm_n1707, in_21);
	nand (gm_n1709, gm_n55, gm_n82, gm_n72, gm_n420, gm_n64);
	nor (gm_n1710, gm_n53, in_10, gm_n51, gm_n1709, in_12);
	nand (gm_n1711, gm_n63, gm_n50, gm_n49, gm_n1710, gm_n46);
	nor (gm_n1712, gm_n62, in_18, gm_n81, gm_n1711, in_20);
	nand (gm_n1713, gm_n1712, in_21);
	and (gm_n1714, gm_n55, gm_n82, in_5, gm_n284, in_8);
	nand (gm_n1715, gm_n53, in_10, in_9, gm_n1714, in_12);
	nor (gm_n1716, gm_n63, in_14, in_13, gm_n1715, gm_n46);
	nand (gm_n1717, in_19, gm_n47, gm_n81, gm_n1716, gm_n45);
	nor (gm_n1718, gm_n1717, gm_n71);
	and (gm_n1719, gm_n64, gm_n55, gm_n82, gm_n638, in_9);
	and (gm_n1720, in_12, gm_n53, gm_n52, gm_n1719, gm_n49);
	nand (gm_n1721, gm_n46, gm_n63, in_14, gm_n1720, gm_n81);
	nor (gm_n1722, in_20, gm_n62, in_18, gm_n1721, gm_n71);
	nand (gm_n1723, in_8, in_7, in_6, gm_n1075, in_9);
	nor (gm_n1724, gm_n48, in_11, in_10, gm_n1723, gm_n49);
	nand (gm_n1725, in_16, gm_n63, in_14, gm_n1724, gm_n81);
	nor (gm_n1726, gm_n45, gm_n62, in_18, gm_n1725, in_21);
	and (gm_n1727, gm_n53, in_10, gm_n51, gm_n1315, gm_n48);
	and (gm_n1728, gm_n63, gm_n50, gm_n49, gm_n1727, gm_n46);
	nand (gm_n1729, gm_n62, in_18, gm_n81, gm_n1728, gm_n45);
	nor (gm_n1730, gm_n1729, gm_n71);
	nor (gm_n1731, gm_n64, gm_n55, gm_n82, gm_n1429, in_9);
	nand (gm_n1732, gm_n48, gm_n53, in_10, gm_n1731, in_13);
	nor (gm_n1733, in_16, gm_n63, in_14, gm_n1732, gm_n81);
	nand (gm_n1734, in_20, in_19, gm_n47, gm_n1733, in_21);
	or (gm_n1735, gm_n55, in_6, gm_n72, gm_n130, gm_n64);
	nor (gm_n1736, in_11, gm_n52, in_9, gm_n1735, in_12);
	nand (gm_n1737, gm_n63, in_14, gm_n49, gm_n1736);
	nor (gm_n1738, in_18, gm_n81, gm_n46, gm_n1737, in_19);
	nand (gm_n1739, gm_n1738, gm_n71, in_20);
	nor (gm_n1740, in_11, gm_n52, in_9, gm_n363);
	nand (gm_n1741, in_14, gm_n49, gm_n48, gm_n1740, gm_n63);
	nor (gm_n1742, gm_n47, gm_n81, in_16, gm_n1741, in_19);
	nand (gm_n1743, gm_n1742, gm_n71, gm_n45);
	or (gm_n1744, gm_n64, in_7, in_6, gm_n530, gm_n51);
	or (gm_n1745, gm_n48, gm_n53, gm_n52, gm_n1744, gm_n49);
	nor (gm_n1746, in_16, gm_n63, gm_n50, gm_n1745, gm_n81);
	nand (gm_n1747, in_20, in_19, in_18, gm_n1746, gm_n71);
	nand (gm_n1748, gm_n62, gm_n47, gm_n81, gm_n191, in_20);
	nor (gm_n1749, gm_n1748, gm_n71);
	nand (gm_n1750, in_7, gm_n82, gm_n72, gm_n252, in_8);
	nor (gm_n1751, gm_n53, in_10, gm_n51, gm_n1750);
	and (gm_n1752, gm_n50, in_13, in_12, gm_n1751, in_15);
	nand (gm_n1753, gm_n47, gm_n81, gm_n46, gm_n1752, in_19);
	nor (gm_n1754, gm_n1753, gm_n71, in_20);
	nor (gm_n1755, in_8, gm_n55, gm_n82, gm_n530, gm_n51);
	and (gm_n1756, in_12, in_11, in_10, gm_n1755, gm_n49);
	nand (gm_n1757, in_16, gm_n63, in_14, gm_n1756, gm_n81);
	nor (gm_n1758, gm_n45, in_19, in_18, gm_n1757, gm_n71);
	nor (gm_n1759, gm_n64, in_7, gm_n82, gm_n103, gm_n51);
	and (gm_n1760, gm_n48, in_11, in_10, gm_n1759, in_13);
	nand (gm_n1761, gm_n46, gm_n63, gm_n50, gm_n1760, in_17);
	nor (gm_n1762, in_20, gm_n62, in_18, gm_n1761, in_21);
	nand (gm_n1763, in_7, in_6, in_5, gm_n493, gm_n64);
	nor (gm_n1764, gm_n53, in_10, gm_n51, gm_n1763, gm_n48);
	nand (gm_n1765, in_15, in_14, gm_n49, gm_n1764, in_16);
	nor (gm_n1766, gm_n62, in_18, gm_n81, gm_n1765, in_20);
	nand (gm_n1767, gm_n1766, in_21);
	nand (gm_n1768, gm_n49, gm_n48, gm_n53, gm_n505, in_14);
	nor (gm_n1769, in_17, in_16, in_15, gm_n1768, gm_n47);
	nand (gm_n1770, gm_n71, in_20, gm_n62, gm_n1769);
	nand (gm_n1771, gm_n71, gm_n45, in_19, gm_n1477);
	nor (gm_n1772, in_10, gm_n51, in_8, gm_n390, gm_n53);
	nand (gm_n1773, gm_n50, gm_n49, in_12, gm_n1772, in_15);
	nor (gm_n1774, gm_n47, in_17, in_16, gm_n1773, gm_n62);
	nand (gm_n1775, gm_n1774, gm_n71, in_20);
	nor (gm_n1776, gm_n285, gm_n52, gm_n51);
	and (gm_n1777, gm_n49, in_12, in_11, gm_n1776, gm_n50);
	nand (gm_n1778, gm_n81, gm_n46, gm_n63, gm_n1777, gm_n47);
	nor (gm_n1779, in_21, gm_n45, gm_n62, gm_n1778);
	nor (gm_n1780, gm_n64, gm_n55, gm_n82, gm_n119, gm_n51);
	and (gm_n1781, in_12, in_11, in_10, gm_n1780, in_13);
	nand (gm_n1782, in_16, in_15, gm_n50, gm_n1781, in_17);
	nor (gm_n1783, gm_n45, gm_n62, in_18, gm_n1782, gm_n71);
	nand (gm_n1784, in_8, gm_n55, in_6, gm_n379, gm_n51);
	nor (gm_n1785, gm_n48, in_11, in_10, gm_n1784, in_13);
	nand (gm_n1786, in_16, gm_n63, in_14, gm_n1785, in_17);
	nor (gm_n1787, in_20, gm_n62, in_18, gm_n1786, in_21);
	nor (gm_n1788, in_7, in_6, gm_n72, gm_n867, in_8);
	and (gm_n1789, in_11, in_10, in_9, gm_n1788);
	and (gm_n1790, in_14, in_13, in_12, gm_n1789, in_15);
	nand (gm_n1791, gm_n47, in_17, in_16, gm_n1790, gm_n62);
	nor (gm_n1792, gm_n1791, in_21, gm_n45);
	nor (gm_n1793, gm_n46, in_15, in_14, gm_n412, in_17);
	nand (gm_n1794, in_20, gm_n62, gm_n47, gm_n1793, gm_n71);
	nand (gm_n1795, gm_n48, in_11, gm_n52, gm_n1365, in_13);
	nor (gm_n1796, in_16, in_15, gm_n50, gm_n1795, in_17);
	nand (gm_n1797, gm_n45, in_19, gm_n47, gm_n1796, gm_n71);
	nand (gm_n1798, gm_n64, in_7, gm_n82, gm_n757, in_9);
	nor (gm_n1799, gm_n1798, gm_n52);
	nand (gm_n1800, in_13, gm_n48, gm_n53, gm_n1799, gm_n50);
	nor (gm_n1801, gm_n81, in_16, gm_n63, gm_n1800, gm_n47);
	nand (gm_n1802, in_21, gm_n45, gm_n62, gm_n1801);
	nand (gm_n1803, in_7, in_6, in_5, gm_n327, in_8);
	nor (gm_n1804, gm_n1803, in_9);
	nand (gm_n1805, gm_n48, in_11, gm_n52, gm_n1804, gm_n49);
	nor (gm_n1806, in_16, gm_n63, gm_n50, gm_n1805, gm_n81);
	nand (gm_n1807, gm_n45, in_19, gm_n47, gm_n1806, in_21);
	and (gm_n1808, gm_n431, in_9, gm_n64);
	and (gm_n1809, in_12, in_11, gm_n52, gm_n1808, in_13);
	nand (gm_n1810, gm_n46, in_15, gm_n50, gm_n1809, gm_n81);
	nor (gm_n1811, gm_n45, in_19, gm_n47, gm_n1810, gm_n71);
	nand (gm_n1812, gm_n566, in_10, gm_n51);
	nor (gm_n1813, in_13, in_12, gm_n53, gm_n1812, gm_n50);
	nand (gm_n1814, gm_n81, gm_n46, in_15, gm_n1813, in_18);
	nor (gm_n1815, gm_n71, in_20, in_19, gm_n1814);
	nand (gm_n1816, gm_n53, in_10, gm_n51, gm_n1603, in_12);
	nor (gm_n1817, gm_n1816, in_14, in_13);
	nand (gm_n1818, in_17, in_16, gm_n63, gm_n1817, gm_n47);
	nor (gm_n1819, gm_n71, gm_n45, gm_n62, gm_n1818);
	and (gm_n1820, in_11, in_10, in_9, gm_n458);
	and (gm_n1821, gm_n50, in_13, gm_n48, gm_n1820, gm_n63);
	nand (gm_n1822, in_18, gm_n81, gm_n46, gm_n1821, in_19);
	nor (gm_n1823, gm_n1822, in_21, in_20);
	or (gm_n1824, in_8, gm_n55, gm_n82, gm_n103, in_9);
	or (gm_n1825, gm_n48, in_11, gm_n52, gm_n1824, in_13);
	nor (gm_n1826, gm_n46, in_15, in_14, gm_n1825, gm_n81);
	nand (gm_n1827, gm_n45, gm_n62, in_18, gm_n1826, gm_n71);
	or (gm_n1828, in_12, in_11, in_10, gm_n1398, in_13);
	nor (gm_n1829, in_16, in_15, in_14, gm_n1828, gm_n81);
	nand (gm_n1830, in_20, in_19, gm_n47, gm_n1829, in_21);
	or (gm_n1831, gm_n55, gm_n82, gm_n72, gm_n75, gm_n64);
	nor (gm_n1832, in_11, in_10, gm_n51, gm_n1831, in_12);
	nand (gm_n1833, gm_n63, gm_n50, in_13, gm_n1832, in_16);
	nor (gm_n1834, gm_n62, in_18, in_17, gm_n1833, in_20);
	nand (gm_n1835, gm_n1834, in_21);
	or (gm_n1836, in_8, in_7, gm_n82, gm_n103, gm_n51);
	nor (gm_n1837, in_12, in_11, gm_n52, gm_n1836, in_13);
	and (gm_n1838, in_16, in_15, in_14, gm_n1837, in_17);
	nand (gm_n1839, gm_n45, gm_n62, gm_n47, gm_n1838, in_21);
	and (gm_n1840, gm_n64, gm_n55, gm_n82, gm_n379, gm_n51);
	nand (gm_n1841, gm_n48, gm_n53, gm_n52, gm_n1840, gm_n49);
	or (gm_n1842, in_16, in_15, in_14, gm_n1841, gm_n81);
	nor (gm_n1843, in_20, gm_n62, in_18, gm_n1842, in_21);
	or (gm_n1844, in_9, gm_n64, gm_n55, gm_n843, gm_n52);
	nor (gm_n1845, in_13, gm_n48, gm_n53, gm_n1844, gm_n50);
	nand (gm_n1846, gm_n81, in_16, in_15, gm_n1845, in_18);
	nor (gm_n1847, in_21, gm_n45, gm_n62, gm_n1846);
	nand (gm_n1848, in_9, in_8, in_7, gm_n404, gm_n52);
	nor (gm_n1849, in_13, gm_n48, in_11, gm_n1848, in_14);
	nand (gm_n1850, gm_n81, gm_n46, in_15, gm_n1849, gm_n47);
	nor (gm_n1851, in_21, gm_n45, in_19, gm_n1850);
	or (gm_n1852, in_9, in_8, in_7, gm_n1256, in_10);
	nor (gm_n1853, gm_n49, in_12, in_11, gm_n1852, gm_n50);
	nand (gm_n1854, in_17, in_16, in_15, gm_n1853, gm_n47);
	nor (gm_n1855, in_21, in_20, in_19, gm_n1854);
	nor (gm_n1856, in_7, in_6, in_5, gm_n130, gm_n64);
	and (gm_n1857, gm_n53, in_10, in_9, gm_n1856);
	nand (gm_n1858, in_14, in_13, in_12, gm_n1857, in_15);
	nor (gm_n1859, gm_n47, gm_n81, gm_n46, gm_n1858, gm_n62);
	nand (gm_n1860, gm_n1859, in_21, gm_n45);
	nor (gm_n1861, in_8, in_7, gm_n82, gm_n199, gm_n51);
	nand (gm_n1862, in_12, in_11, in_10, gm_n1861, gm_n49);
	nor (gm_n1863, in_16, in_15, in_14, gm_n1862, gm_n81);
	nand (gm_n1864, in_20, gm_n62, in_18, gm_n1863, gm_n71);
	nor (gm_n1865, gm_n51, gm_n64, in_7, gm_n897, in_10);
	nand (gm_n1866, in_13, in_12, gm_n53, gm_n1865, in_14);
	nor (gm_n1867, gm_n81, in_16, in_15, gm_n1866, gm_n47);
	nand (gm_n1868, gm_n71, gm_n45, gm_n62, gm_n1867);
	or (gm_n1869, in_7, in_6, gm_n72, gm_n167, in_8);
	nor (gm_n1870, gm_n53, in_10, in_9, gm_n1869);
	nand (gm_n1871, in_14, in_13, in_12, gm_n1870, gm_n63);
	nor (gm_n1872, gm_n47, in_17, in_16, gm_n1871, gm_n62);
	nand (gm_n1873, gm_n1872, in_21, gm_n45);
	and (gm_n1874, gm_n55, gm_n82, gm_n72, gm_n89, gm_n64);
	nand (gm_n1875, in_11, in_10, in_9, gm_n1874);
	nor (gm_n1876, gm_n50, in_13, in_12, gm_n1875, in_15);
	nand (gm_n1877, in_18, in_17, gm_n46, gm_n1876, in_19);
	nor (gm_n1878, gm_n1877, in_21, gm_n45);
	nand (gm_n1879, gm_n55, in_6, in_5, gm_n519, in_8);
	or (gm_n1880, in_11, in_10, gm_n51, gm_n1879, gm_n48);
	nor (gm_n1881, in_15, in_14, gm_n49, gm_n1880);
	nand (gm_n1882, in_18, in_17, in_16, gm_n1881, gm_n62);
	nor (gm_n1883, gm_n1882, gm_n71, gm_n45);
	or (gm_n1884, gm_n328, gm_n52, in_9);
	nor (gm_n1885, gm_n49, in_12, gm_n53, gm_n1884, gm_n50);
	nand (gm_n1886, gm_n81, gm_n46, in_15, gm_n1885, gm_n47);
	nor (gm_n1887, in_21, gm_n45, in_19, gm_n1886);
	or (gm_n1888, gm_n64, in_7, in_6, gm_n161, in_9);
	nor (gm_n1889, gm_n1888, in_10);
	and (gm_n1890, gm_n49, gm_n48, in_11, gm_n1889, in_14);
	nand (gm_n1891, gm_n81, in_16, gm_n63, gm_n1890, gm_n47);
	nor (gm_n1892, in_21, in_20, gm_n62, gm_n1891);
	and (gm_n1893, in_16, in_15, in_14, gm_n835, gm_n81);
	nand (gm_n1894, in_20, gm_n62, gm_n47, gm_n1893, in_21);
	and (gm_n1895, gm_n55, in_6, in_5, gm_n89, in_8);
	and (gm_n1896, in_11, in_10, in_9, gm_n1895, in_12);
	nand (gm_n1897, gm_n63, gm_n50, in_13, gm_n1896, gm_n46);
	nor (gm_n1898, gm_n62, gm_n47, gm_n81, gm_n1897, in_20);
	nand (gm_n1899, gm_n1898, in_21);
	nand (gm_n1900, gm_n64, in_7, gm_n82, gm_n1075, in_9);
	or (gm_n1901, gm_n48, in_11, gm_n52, gm_n1900, in_13);
	nor (gm_n1902, in_16, gm_n63, in_14, gm_n1901, in_17);
	nand (gm_n1903, in_20, gm_n62, gm_n47, gm_n1902, gm_n71);
	nor (gm_n1904, gm_n53, in_10, gm_n51, gm_n1098, in_12);
	nand (gm_n1905, gm_n63, gm_n50, in_13, gm_n1904, in_16);
	nor (gm_n1906, gm_n62, gm_n47, gm_n81, gm_n1905, gm_n45);
	nand (gm_n1907, gm_n1906, in_21);
	or (gm_n1908, in_9, gm_n64, gm_n55, gm_n279, in_10);
	nor (gm_n1909, in_13, in_12, gm_n53, gm_n1908, gm_n50);
	nand (gm_n1910, gm_n81, gm_n46, gm_n63, gm_n1909, in_18);
	nor (gm_n1911, in_21, gm_n45, in_19, gm_n1910);
	or (gm_n1912, gm_n53, gm_n52, in_9, gm_n520, in_12);
	nor (gm_n1913, gm_n1912, gm_n49);
	nand (gm_n1914, gm_n46, in_15, in_14, gm_n1913, in_17);
	nor (gm_n1915, in_20, in_19, gm_n47, gm_n1914, in_21);
	nand (gm_n1916, gm_n1116, gm_n52, gm_n51);
	nor (gm_n1917, in_13, gm_n48, gm_n53, gm_n1916, gm_n50);
	nand (gm_n1918, in_17, in_16, in_15, gm_n1917, in_18);
	nor (gm_n1919, gm_n71, in_20, gm_n62, gm_n1918);
	nand (gm_n1920, gm_n51, in_8, gm_n55, gm_n1007, gm_n52);
	nor (gm_n1921, gm_n49, in_12, in_11, gm_n1920, gm_n50);
	nand (gm_n1922, gm_n81, in_16, gm_n63, gm_n1921, gm_n47);
	nor (gm_n1923, in_21, in_20, in_19, gm_n1922);
	and (gm_n1924, in_11, gm_n52, in_9, gm_n1315);
	nand (gm_n1925, gm_n50, in_13, in_12, gm_n1924, in_15);
	nor (gm_n1926, in_18, gm_n81, in_16, gm_n1925, in_19);
	nand (gm_n1927, gm_n1926, gm_n71, in_20);
	nor (gm_n1928, gm_n53, in_10, gm_n51, gm_n178, in_12);
	nand (gm_n1929, in_15, in_14, gm_n49, gm_n1928, in_16);
	nor (gm_n1930, in_19, gm_n47, in_17, gm_n1929, in_20);
	nand (gm_n1931, gm_n1930, in_21);
	nor (gm_n1932, in_8, in_7, gm_n82, gm_n96, in_9);
	nand (gm_n1933, in_12, in_11, gm_n52, gm_n1932, in_13);
	nor (gm_n1934, gm_n46, in_15, in_14, gm_n1933, in_17);
	nand (gm_n1935, in_20, in_19, gm_n47, gm_n1934, gm_n71);
	nor (gm_n1936, gm_n55, gm_n82, gm_n72, gm_n188, gm_n64);
	and (gm_n1937, gm_n53, in_10, in_9, gm_n1936);
	and (gm_n1938, gm_n1937, in_13, gm_n48);
	and (gm_n1939, in_16, in_15, gm_n50, gm_n1938, gm_n81);
	nand (gm_n1940, in_20, gm_n62, in_18, gm_n1939, in_21);
	nor (gm_n1941, gm_n64, gm_n55, gm_n82, gm_n119, in_9);
	and (gm_n1942, gm_n48, gm_n53, gm_n52, gm_n1941, in_13);
	nand (gm_n1943, in_16, in_15, gm_n50, gm_n1942, in_17);
	nor (gm_n1944, gm_n45, in_19, gm_n47, gm_n1943, gm_n71);
	and (gm_n1945, in_8, gm_n55, in_6, gm_n757, in_9);
	and (gm_n1946, in_12, in_11, in_10, gm_n1945, gm_n49);
	nand (gm_n1947, in_16, in_15, in_14, gm_n1946, gm_n81);
	nor (gm_n1948, gm_n45, gm_n62, in_18, gm_n1947, in_21);
	nor (gm_n1949, in_12, gm_n53, in_10, gm_n1599, gm_n49);
	nand (gm_n1950, in_16, in_15, gm_n50, gm_n1949, in_17);
	nor (gm_n1951, in_20, gm_n62, in_18, gm_n1950, gm_n71);
	nor (gm_n1952, in_7, gm_n82, in_5, gm_n483, in_8);
	nand (gm_n1953, gm_n1952, in_10, gm_n51);
	nor (gm_n1954, gm_n49, in_12, gm_n53, gm_n1953, in_14);
	nand (gm_n1955, gm_n81, in_16, in_15, gm_n1954, in_18);
	nor (gm_n1956, in_21, in_20, in_19, gm_n1955);
	nand (gm_n1957, in_7, gm_n82, gm_n72, gm_n284, gm_n64);
	nor (gm_n1958, gm_n1957, gm_n52, in_9);
	nand (gm_n1959, in_13, gm_n48, gm_n53, gm_n1958, gm_n50);
	nor (gm_n1960, gm_n81, gm_n46, gm_n63, gm_n1959, in_18);
	nand (gm_n1961, in_21, gm_n45, gm_n62, gm_n1960);
	nor (gm_n1962, in_8, gm_n55, gm_n82, gm_n161, in_9);
	nand (gm_n1963, gm_n48, gm_n53, gm_n52, gm_n1962, in_13);
	nor (gm_n1964, in_16, gm_n63, in_14, gm_n1963, gm_n81);
	nand (gm_n1965, gm_n45, in_19, gm_n47, gm_n1964, in_21);
	nor (gm_n1966, gm_n64, gm_n55, in_6, gm_n119, in_9);
	nand (gm_n1967, gm_n48, in_11, in_10, gm_n1966, in_13);
	nor (gm_n1968, gm_n46, gm_n63, gm_n50, gm_n1967, gm_n81);
	nand (gm_n1969, in_20, in_19, in_18, gm_n1968, in_21);
	or (gm_n1970, in_7, gm_n82, in_5, gm_n643, gm_n64);
	nor (gm_n1971, in_11, gm_n52, gm_n51, gm_n1970, in_12);
	nand (gm_n1972, in_15, gm_n50, in_13, gm_n1971, gm_n46);
	nor (gm_n1973, gm_n62, gm_n47, gm_n81, gm_n1972, gm_n45);
	nand (gm_n1974, gm_n1973, in_21);
	and (gm_n1975, gm_n64, gm_n55, in_6, gm_n757, in_9);
	and (gm_n1976, in_12, in_11, gm_n52, gm_n1975, gm_n49);
	nand (gm_n1977, gm_n46, in_15, gm_n50, gm_n1976, gm_n81);
	nor (gm_n1978, gm_n45, gm_n62, gm_n47, gm_n1977, in_21);
	nor (gm_n1979, gm_n49, gm_n48, gm_n53, gm_n1008, in_14);
	nand (gm_n1980, gm_n81, gm_n46, gm_n63, gm_n1979, gm_n47);
	nor (gm_n1981, gm_n71, in_20, gm_n62, gm_n1980);
	and (gm_n1982, in_8, gm_n55, gm_n82, gm_n374, in_9);
	nand (gm_n1983, in_12, gm_n53, gm_n52, gm_n1982, in_13);
	or (gm_n1984, in_16, gm_n63, gm_n50, gm_n1983, in_17);
	nor (gm_n1985, in_20, gm_n62, gm_n47, gm_n1984, in_21);
	nor (gm_n1986, gm_n55, in_6, gm_n72, gm_n643, gm_n64);
	and (gm_n1987, in_11, in_10, gm_n51, gm_n1986);
	and (gm_n1988, gm_n50, gm_n49, gm_n48, gm_n1987, gm_n63);
	nand (gm_n1989, in_18, in_17, in_16, gm_n1988, gm_n62);
	nor (gm_n1990, gm_n1989, gm_n71, gm_n45);
	nand (gm_n1991, in_14, gm_n49, in_12, gm_n1820, gm_n63);
	nor (gm_n1992, in_18, gm_n81, in_16, gm_n1991, in_19);
	nand (gm_n1993, gm_n1992, gm_n71, in_20);
	nand (gm_n1994, gm_n48, in_11, in_10, gm_n1932, gm_n49);
	nor (gm_n1995, gm_n46, in_15, in_14, gm_n1994, in_17);
	nand (gm_n1996, in_20, gm_n62, gm_n47, gm_n1995, in_21);
	and (gm_n1997, in_11, in_10, gm_n51, gm_n1315, gm_n48);
	nand (gm_n1998, gm_n1997, in_14, gm_n49);
	nor (gm_n1999, in_17, gm_n46, in_15, gm_n1998, gm_n47);
	nand (gm_n2000, gm_n71, in_20, gm_n62, gm_n1999);
	nor (gm_n2001, in_9, gm_n64, gm_n55, gm_n84);
	nand (gm_n2002, gm_n48, gm_n53, in_10, gm_n2001, gm_n49);
	nor (gm_n2003, gm_n46, gm_n63, in_14, gm_n2002, gm_n81);
	nand (gm_n2004, in_20, gm_n62, in_18, gm_n2003, in_21);
	nand (gm_n2005, gm_n55, in_6, gm_n72, gm_n420, in_8);
	or (gm_n2006, gm_n2005, in_10, gm_n51);
	nor (gm_n2007, in_13, gm_n48, gm_n53, gm_n2006);
	nand (gm_n2008, gm_n46, gm_n63, in_14, gm_n2007, gm_n81);
	nor (gm_n2009, in_20, in_19, in_18, gm_n2008, in_21);
	nand (gm_n2010, gm_n53, gm_n52, in_9, gm_n593, in_12);
	nor (gm_n2011, gm_n63, gm_n50, in_13, gm_n2010, gm_n46);
	nand (gm_n2012, gm_n62, in_18, in_17, gm_n2011, in_20);
	nor (gm_n2013, gm_n2012, in_21);
	and (gm_n2014, gm_n55, gm_n82, gm_n72, gm_n493, in_8);
	nand (gm_n2015, gm_n2014, gm_n52, in_9);
	nor (gm_n2016, gm_n49, in_12, in_11, gm_n2015, in_14);
	nand (gm_n2017, in_17, gm_n46, in_15, gm_n2016, in_18);
	nor (gm_n2018, in_21, in_20, in_19, gm_n2017);
	and (gm_n2019, in_11, in_10, gm_n51, gm_n868);
	and (gm_n2020, gm_n50, gm_n49, gm_n48, gm_n2019, in_15);
	nand (gm_n2021, in_18, gm_n81, gm_n46, gm_n2020, gm_n62);
	nor (gm_n2022, gm_n2021, in_21, gm_n45);
	and (gm_n2023, in_11, gm_n52, gm_n51, gm_n1315);
	nand (gm_n2024, in_14, in_13, gm_n48, gm_n2023, gm_n63);
	nor (gm_n2025, in_18, in_17, gm_n46, gm_n2024, gm_n62);
	nand (gm_n2026, gm_n2025, in_21, gm_n45);
	nand (gm_n2027, in_11, gm_n52, in_9, gm_n242, gm_n48);
	or (gm_n2028, gm_n63, gm_n50, in_13, gm_n2027, in_16);
	nor (gm_n2029, gm_n62, in_18, gm_n81, gm_n2028, in_20);
	nand (gm_n2030, gm_n2029, in_21);
	or (gm_n2031, in_12, in_11, in_10, gm_n228, gm_n49);
	nor (gm_n2032, in_16, gm_n63, gm_n50, gm_n2031, in_17);
	nand (gm_n2033, in_20, gm_n62, gm_n47, gm_n2032, in_21);
	nor (gm_n2034, in_7, gm_n82, in_5, gm_n188, gm_n64);
	and (gm_n2035, in_11, gm_n52, gm_n51, gm_n2034);
	nand (gm_n2036, in_14, in_13, in_12, gm_n2035, in_15);
	nor (gm_n2037, in_18, gm_n81, in_16, gm_n2036, gm_n62);
	nand (gm_n2038, gm_n2037, in_21, gm_n45);
	and (gm_n2039, in_11, in_10, gm_n51, gm_n858);
	and (gm_n2040, gm_n50, in_13, in_12, gm_n2039, gm_n63);
	nand (gm_n2041, gm_n47, gm_n81, in_16, gm_n2040, in_19);
	nor (gm_n2042, gm_n2041, in_21, gm_n45);
	nand (gm_n2043, gm_n64, gm_n55, gm_n82, gm_n638, gm_n51);
	or (gm_n2044, gm_n48, gm_n53, gm_n52, gm_n2043, gm_n49);
	or (gm_n2045, in_16, in_15, gm_n50, gm_n2044, gm_n81);
	nor (gm_n2046, in_20, in_19, gm_n47, gm_n2045, gm_n71);
	and (gm_n2047, in_7, in_6, gm_n72, gm_n493, in_8);
	nand (gm_n2048, gm_n53, in_10, in_9, gm_n2047);
	nor (gm_n2049, gm_n50, gm_n49, gm_n48, gm_n2048, gm_n63);
	nand (gm_n2050, gm_n47, in_17, gm_n46, gm_n2049, in_19);
	nor (gm_n2051, gm_n2050, gm_n71, in_20);
	nand (gm_n2052, gm_n64, gm_n55, in_6, gm_n374, gm_n51);
	nor (gm_n2053, in_12, gm_n53, gm_n52, gm_n2052, in_13);
	nand (gm_n2054, gm_n46, in_15, gm_n50, gm_n2053, in_17);
	nor (gm_n2055, gm_n45, gm_n62, gm_n47, gm_n2054, gm_n71);
	and (gm_n2056, gm_n64, gm_n55, in_6, gm_n1075, in_9);
	nand (gm_n2057, gm_n48, gm_n53, gm_n52, gm_n2056, in_13);
	nor (gm_n2058, gm_n46, gm_n63, gm_n50, gm_n2057, gm_n81);
	nand (gm_n2059, in_20, gm_n62, in_18, gm_n2058, in_21);
	nand (gm_n2060, gm_n55, gm_n82, gm_n72, gm_n89, in_8);
	nor (gm_n2061, gm_n53, in_10, gm_n51, gm_n2060, in_12);
	nand (gm_n2062, gm_n63, in_14, gm_n49, gm_n2061, in_16);
	nor (gm_n2063, gm_n62, in_18, in_17, gm_n2062, in_20);
	nand (gm_n2064, gm_n2063, in_21);
	nor (gm_n2065, in_16, gm_n63, in_14, gm_n714, gm_n81);
	nand (gm_n2066, in_20, in_19, in_18, gm_n2065, in_21);
	nor (gm_n2067, gm_n51, in_8, gm_n55, gm_n279);
	nand (gm_n2068, gm_n48, gm_n53, in_10, gm_n2067, gm_n49);
	nor (gm_n2069, gm_n46, in_15, in_14, gm_n2068, in_17);
	nand (gm_n2070, in_20, gm_n62, gm_n47, gm_n2069, gm_n71);
	and (gm_n2071, in_12, gm_n53, in_10, gm_n1365, gm_n49);
	nand (gm_n2072, in_16, in_15, in_14, gm_n2071, gm_n81);
	nor (gm_n2073, gm_n45, gm_n62, gm_n47, gm_n2072, gm_n71);
	nor (gm_n2074, in_12, in_11, gm_n52, gm_n863, gm_n49);
	nand (gm_n2075, gm_n46, gm_n63, gm_n50, gm_n2074, in_17);
	nor (gm_n2076, gm_n45, gm_n62, in_18, gm_n2075, in_21);
	or (gm_n2077, in_7, gm_n82, gm_n72, gm_n75, gm_n64);
	nor (gm_n2078, gm_n2077, in_10, gm_n51);
	and (gm_n2079, in_13, gm_n48, gm_n53, gm_n2078);
	nand (gm_n2080, gm_n46, gm_n63, gm_n50, gm_n2079, gm_n81);
	nor (gm_n2081, gm_n45, gm_n62, gm_n47, gm_n2080, in_21);
	nand (gm_n2082, gm_n47, gm_n81, gm_n46, gm_n1881, in_19);
	nor (gm_n2083, gm_n2082, in_21, in_20);
	nor (gm_n2084, gm_n53, gm_n52, in_9, gm_n607, in_12);
	nand (gm_n2085, gm_n63, gm_n50, in_13, gm_n2084, gm_n46);
	nor (gm_n2086, gm_n62, in_18, in_17, gm_n2085, gm_n45);
	nand (gm_n2087, gm_n2086, in_21);
	nor (gm_n2088, in_7, gm_n82, in_5, gm_n130, gm_n64);
	and (gm_n2089, gm_n53, gm_n52, gm_n51, gm_n2088, gm_n48);
	nand (gm_n2090, gm_n2089, in_13);
	nor (gm_n2091, in_16, gm_n63, gm_n50, gm_n2090, gm_n81);
	nand (gm_n2092, gm_n45, gm_n62, in_18, gm_n2091, gm_n71);
	nor (gm_n2093, gm_n64, in_7, in_6, gm_n96, in_9);
	nand (gm_n2094, in_12, in_11, in_10, gm_n2093, gm_n49);
	nor (gm_n2095, gm_n46, gm_n63, in_14, gm_n2094, in_17);
	nand (gm_n2096, gm_n45, in_19, gm_n47, gm_n2095, in_21);
	nor (gm_n2097, gm_n64, in_7, gm_n82, gm_n1429, gm_n51);
	nand (gm_n2098, in_12, gm_n53, in_10, gm_n2097, gm_n49);
	nor (gm_n2099, in_16, in_15, gm_n50, gm_n2098, in_17);
	nand (gm_n2100, in_20, in_19, in_18, gm_n2099, gm_n71);
	nor (gm_n2101, in_15, gm_n50, in_13, gm_n1352, gm_n46);
	nand (gm_n2102, in_19, gm_n47, in_17, gm_n2101, gm_n45);
	nor (gm_n2103, gm_n2102, gm_n71);
	or (gm_n2104, in_11, gm_n52, in_9, gm_n218, in_12);
	nor (gm_n2105, gm_n63, gm_n50, gm_n49, gm_n2104, in_16);
	nand (gm_n2106, gm_n62, in_18, gm_n81, gm_n2105, in_20);
	nor (gm_n2107, gm_n2106, gm_n71);
	nor (gm_n2108, gm_n50, gm_n49, gm_n48, gm_n854, in_15);
	nand (gm_n2109, in_18, in_17, gm_n46, gm_n2108, gm_n62);
	nor (gm_n2110, gm_n2109, in_21, in_20);
	nor (gm_n2111, in_15, in_14, in_13, gm_n1595, gm_n46);
	nand (gm_n2112, gm_n62, in_18, in_17, gm_n2111, in_20);
	nor (gm_n2113, gm_n2112, in_21);
	nand (gm_n2114, gm_n55, in_6, in_5, gm_n420, gm_n64);
	nor (gm_n2115, gm_n53, gm_n52, in_9, gm_n2114, gm_n48);
	nand (gm_n2116, gm_n63, in_14, gm_n49, gm_n2115, in_16);
	nor (gm_n2117, gm_n62, gm_n47, gm_n81, gm_n2116, in_20);
	nand (gm_n2118, gm_n2117, in_21);
	nand (gm_n2119, gm_n55, in_6, gm_n72, gm_n296, in_8);
	nor (gm_n2120, gm_n2119, in_10, gm_n51);
	nand (gm_n2121, in_13, in_12, in_11, gm_n2120);
	nor (gm_n2122, in_16, in_15, gm_n50, gm_n2121, gm_n81);
	nand (gm_n2123, gm_n45, in_19, gm_n47, gm_n2122, in_21);
	nand (gm_n2124, in_13, in_12, in_11, gm_n682, gm_n50);
	nor (gm_n2125, gm_n81, in_16, in_15, gm_n2124, in_18);
	nand (gm_n2126, gm_n71, gm_n45, gm_n62, gm_n2125);
	nor (gm_n2127, gm_n2114, in_10, in_9);
	nand (gm_n2128, gm_n49, in_12, in_11, gm_n2127);
	nor (gm_n2129, in_16, in_15, in_14, gm_n2128, gm_n81);
	nand (gm_n2130, gm_n45, gm_n62, gm_n47, gm_n2129, gm_n71);
	nand (gm_n2131, in_14, gm_n49, in_12, gm_n634, in_15);
	nor (gm_n2132, gm_n47, gm_n81, in_16, gm_n2131, in_19);
	nand (gm_n2133, gm_n2132, in_21, in_20);
	nand (gm_n2134, gm_n2126, gm_n2123, gm_n2118, gm_n2133, gm_n2130);
	nor (gm_n2135, gm_n2110, gm_n2107, gm_n2103, gm_n2134, gm_n2113);
	nand (gm_n2136, gm_n2096, gm_n2092, gm_n2087, gm_n2135, gm_n2100);
	nor (gm_n2137, gm_n2081, gm_n2076, gm_n2073, gm_n2136, gm_n2083);
	nand (gm_n2138, gm_n2066, gm_n2064, gm_n2059, gm_n2137, gm_n2070);
	nor (gm_n2139, gm_n2051, gm_n2046, gm_n2042, gm_n2138, gm_n2055);
	nand (gm_n2140, gm_n2033, gm_n2030, gm_n2026, gm_n2139, gm_n2038);
	nor (gm_n2141, gm_n2018, gm_n2013, gm_n2009, gm_n2140, gm_n2022);
	nand (gm_n2142, gm_n2000, gm_n1996, gm_n1993, gm_n2141, gm_n2004);
	nor (gm_n2143, gm_n1985, gm_n1981, gm_n1978, gm_n2142, gm_n1990);
	nand (gm_n2144, gm_n1969, gm_n1965, gm_n1961, gm_n2143, gm_n1974);
	nor (gm_n2145, gm_n1951, gm_n1948, gm_n1944, gm_n2144, gm_n1956);
	nand (gm_n2146, gm_n1935, gm_n1931, gm_n1927, gm_n2145, gm_n1940);
	nor (gm_n2147, gm_n1919, gm_n1915, gm_n1911, gm_n2146, gm_n1923);
	nand (gm_n2148, gm_n1903, gm_n1899, gm_n1894, gm_n2147, gm_n1907);
	nor (gm_n2149, gm_n1887, gm_n1883, gm_n1878, gm_n2148, gm_n1892);
	nand (gm_n2150, gm_n1868, gm_n1864, gm_n1860, gm_n2149, gm_n1873);
	nor (gm_n2151, gm_n1851, gm_n1847, gm_n1843, gm_n2150, gm_n1855);
	nand (gm_n2152, gm_n1835, gm_n1830, gm_n1827, gm_n2151, gm_n1839);
	nor (gm_n2153, gm_n1819, gm_n1815, gm_n1811, gm_n2152, gm_n1823);
	nand (gm_n2154, gm_n1802, gm_n1797, gm_n1794, gm_n2153, gm_n1807);
	nor (gm_n2155, gm_n1787, gm_n1783, gm_n1779, gm_n2154, gm_n1792);
	nand (gm_n2156, gm_n1771, gm_n1770, gm_n1767, gm_n2155, gm_n1775);
	nor (gm_n2157, gm_n1758, gm_n1754, gm_n1749, gm_n2156, gm_n1762);
	nand (gm_n2158, gm_n1743, gm_n1739, gm_n1734, gm_n2157, gm_n1747);
	nor (gm_n2159, gm_n1726, gm_n1722, gm_n1718, gm_n2158, gm_n1730);
	nand (gm_n2160, gm_n1708, gm_n1703, gm_n1699, gm_n2159, gm_n1713);
	nor (gm_n2161, gm_n1691, gm_n1687, gm_n1682, gm_n2160, gm_n1695);
	nand (gm_n2162, gm_n1674, gm_n1670, gm_n1666, gm_n2161, gm_n1678);
	nor (gm_n2163, gm_n1659, gm_n1655, gm_n1651, gm_n2162, gm_n1663);
	nand (gm_n2164, gm_n1642, gm_n1638, gm_n1633, gm_n2163, gm_n1647);
	nor (gm_n2165, gm_n1624, gm_n1620, gm_n1616, gm_n2164, gm_n1628);
	nand (gm_n2166, gm_n1607, gm_n1602, gm_n1598, gm_n2165, gm_n1612);
	nor (gm_n2167, gm_n1591, gm_n1587, gm_n1582, gm_n2166, gm_n1594);
	nand (gm_n2168, gm_n1576, gm_n1571, gm_n1567, gm_n2167, gm_n1580);
	nor (gm_n2169, gm_n1559, gm_n1554, gm_n1549, gm_n2168, gm_n1562);
	nand (gm_n2170, gm_n1541, gm_n1537, gm_n1532, gm_n2169, gm_n1545);
	nor (out_2, gm_n2170, gm_n1527);
	nor (gm_n2172, in_12, in_11, in_10, gm_n1900, in_13);
	nand (gm_n2173, in_16, in_15, in_14, gm_n2172, in_17);
	nor (gm_n2174, gm_n45, in_19, in_18, gm_n2173, in_21);
	nand (gm_n2175, gm_n48, in_11, gm_n52, gm_n343, in_13);
	nor (gm_n2176, gm_n46, gm_n63, in_14, gm_n2175, gm_n81);
	nand (gm_n2177, gm_n45, gm_n62, in_18, gm_n2176, gm_n71);
	nand (gm_n2178, gm_n50, in_13, gm_n48, gm_n664, in_15);
	nor (gm_n2179, in_18, in_17, in_16, gm_n2178, gm_n62);
	nand (gm_n2180, gm_n2179, in_21, in_20);
	nor (gm_n2181, gm_n55, in_6, in_5, gm_n130, gm_n64);
	and (gm_n2182, gm_n2181, in_9);
	nand (gm_n2183, in_12, gm_n53, gm_n52, gm_n2182, in_13);
	nor (gm_n2184, gm_n46, in_15, in_14, gm_n2183, in_17);
	nand (gm_n2185, in_20, gm_n62, in_18, gm_n2184, gm_n71);
	and (gm_n2186, gm_n1274, gm_n52, gm_n51);
	nand (gm_n2187, gm_n49, in_12, in_11, gm_n2186, gm_n50);
	nor (gm_n2188, gm_n81, gm_n46, gm_n63, gm_n2187, in_18);
	nand (gm_n2189, in_21, gm_n45, in_19, gm_n2188);
	and (gm_n2190, in_11, gm_n52, in_9, gm_n509, gm_n48);
	and (gm_n2191, gm_n63, in_14, gm_n49, gm_n2190, gm_n46);
	nand (gm_n2192, in_19, in_18, in_17, gm_n2191, gm_n45);
	nor (gm_n2193, gm_n2192, gm_n71);
	nor (gm_n2194, in_7, gm_n82, in_5, gm_n108, gm_n64);
	nand (gm_n2195, gm_n53, gm_n52, in_9, gm_n2194, gm_n48);
	nor (gm_n2196, in_15, gm_n50, in_13, gm_n2195, in_16);
	nand (gm_n2197, gm_n62, gm_n47, gm_n81, gm_n2196, in_20);
	nor (gm_n2198, gm_n2197, in_21);
	nand (gm_n2199, in_11, gm_n52, gm_n51, gm_n242, in_12);
	nor (gm_n2200, gm_n63, in_14, in_13, gm_n2199, gm_n46);
	nand (gm_n2201, in_19, gm_n47, in_17, gm_n2200, in_20);
	nor (gm_n2202, gm_n2201, gm_n71);
	nor (gm_n2203, in_9, in_8, gm_n55, gm_n897, in_10);
	and (gm_n2204, gm_n49, in_12, in_11, gm_n2203, gm_n50);
	nand (gm_n2205, gm_n81, in_16, in_15, gm_n2204, in_18);
	nor (gm_n2206, gm_n71, gm_n45, gm_n62, gm_n2205);
	nand (gm_n2207, gm_n50, in_13, gm_n48, gm_n584, in_15);
	nor (gm_n2208, in_18, in_17, gm_n46, gm_n2207, gm_n62);
	nand (gm_n2209, gm_n2208, in_21, gm_n45);
	nor (gm_n2210, gm_n53, gm_n52, in_9, gm_n2114, in_12);
	nand (gm_n2211, in_15, in_14, gm_n49, gm_n2210, gm_n46);
	nor (gm_n2212, gm_n62, gm_n47, gm_n81, gm_n2211, in_20);
	nand (gm_n2213, gm_n2212, in_21);
	nor (gm_n2214, gm_n1750, gm_n52, gm_n51);
	nand (gm_n2215, in_13, in_12, in_11, gm_n2214, gm_n50);
	nor (gm_n2216, gm_n81, in_16, in_15, gm_n2215, in_18);
	nand (gm_n2217, gm_n71, gm_n45, gm_n62, gm_n2216);
	and (gm_n2218, in_9, in_8, in_7, gm_n151, in_10);
	nand (gm_n2219, in_13, in_12, gm_n53, gm_n2218, in_14);
	nor (gm_n2220, gm_n81, in_16, gm_n63, gm_n2219, in_18);
	nand (gm_n2221, in_21, gm_n45, in_19, gm_n2220);
	nor (gm_n2222, in_12, gm_n53, gm_n52, gm_n104, gm_n49);
	nand (gm_n2223, gm_n46, gm_n63, in_14, gm_n2222, gm_n81);
	nor (gm_n2224, in_20, gm_n62, in_18, gm_n2223, in_21);
	or (gm_n2225, gm_n51, in_8, in_7, gm_n279, gm_n52);
	nor (gm_n2226, in_13, gm_n48, gm_n53, gm_n2225, gm_n50);
	nand (gm_n2227, gm_n81, in_16, gm_n63, gm_n2226, gm_n47);
	nor (gm_n2228, in_21, gm_n45, gm_n62, gm_n2227);
	nor (gm_n2229, in_7, gm_n82, gm_n72, gm_n290, in_8);
	nand (gm_n2230, gm_n53, in_10, gm_n51, gm_n2229, gm_n48);
	nor (gm_n2231, gm_n2230, gm_n50, in_13);
	nand (gm_n2232, gm_n81, in_16, gm_n63, gm_n2231, in_18);
	nor (gm_n2233, gm_n71, gm_n45, gm_n62, gm_n2232);
	nor (gm_n2234, gm_n55, gm_n82, in_5, gm_n867, in_8);
	and (gm_n2235, gm_n2234, in_9);
	and (gm_n2236, in_12, in_11, gm_n52, gm_n2235, gm_n49);
	nand (gm_n2237, in_16, gm_n63, in_14, gm_n2236, gm_n81);
	nor (gm_n2238, gm_n45, in_19, gm_n47, gm_n2237, gm_n71);
	nand (gm_n2239, in_7, gm_n82, in_5, gm_n284);
	nor (gm_n2240, in_10, gm_n51, in_8, gm_n2239, in_11);
	nand (gm_n2241, gm_n50, in_13, in_12, gm_n2240, gm_n63);
	nor (gm_n2242, gm_n47, gm_n81, gm_n46, gm_n2241, in_19);
	nand (gm_n2243, gm_n2242, gm_n71, in_20);
	nor (gm_n2244, gm_n1957, in_10, gm_n51);
	nand (gm_n2245, in_13, in_12, in_11, gm_n2244, gm_n50);
	nor (gm_n2246, gm_n81, gm_n46, in_15, gm_n2245, in_18);
	nand (gm_n2247, gm_n71, gm_n45, in_19, gm_n2246);
	nand (gm_n2248, in_12, in_11, gm_n52, gm_n1755, in_13);
	nor (gm_n2249, in_16, in_15, gm_n50, gm_n2248, in_17);
	nand (gm_n2250, in_20, gm_n62, in_18, gm_n2249, gm_n71);
	nand (gm_n2251, in_14, in_13, in_12, gm_n874, gm_n63);
	nor (gm_n2252, gm_n47, gm_n81, gm_n46, gm_n2251, gm_n62);
	nand (gm_n2253, gm_n2252, gm_n71, gm_n45);
	nor (gm_n2254, gm_n55, gm_n82, gm_n72, gm_n643, in_8);
	nand (gm_n2255, in_11, in_10, gm_n51, gm_n2254, in_12);
	nor (gm_n2256, gm_n63, gm_n50, gm_n49, gm_n2255, in_16);
	nand (gm_n2257, gm_n62, in_18, gm_n81, gm_n2256, gm_n45);
	nor (gm_n2258, gm_n2257, gm_n71);
	nor (gm_n2259, gm_n49, gm_n48, in_11, gm_n630, in_14);
	nand (gm_n2260, in_17, gm_n46, gm_n63, gm_n2259, in_18);
	nor (gm_n2261, gm_n71, in_20, in_19, gm_n2260);
	nor (gm_n2262, in_9, in_8, in_7, gm_n525, gm_n52);
	and (gm_n2263, gm_n49, gm_n48, in_11, gm_n2262, in_14);
	nand (gm_n2264, gm_n81, gm_n46, in_15, gm_n2263, in_18);
	nor (gm_n2265, in_21, in_20, gm_n62, gm_n2264);
	or (gm_n2266, gm_n55, gm_n82, in_5, gm_n75, in_8);
	nor (gm_n2267, gm_n53, gm_n52, gm_n51, gm_n2266);
	and (gm_n2268, in_14, gm_n49, in_12, gm_n2267, gm_n63);
	nand (gm_n2269, in_18, in_17, gm_n46, gm_n2268, in_19);
	nor (gm_n2270, gm_n2269, in_21, in_20);
	nor (gm_n2271, in_11, gm_n52, gm_n51, gm_n2119, in_12);
	and (gm_n2272, gm_n2271, in_14, in_13);
	and (gm_n2273, gm_n81, gm_n46, in_15, gm_n2272, in_18);
	nand (gm_n2274, gm_n71, gm_n45, in_19, gm_n2273);
	nand (gm_n2275, gm_n55, gm_n82, gm_n72, gm_n519, gm_n64);
	nor (gm_n2276, gm_n2275, in_10, gm_n51);
	nand (gm_n2277, in_13, gm_n48, in_11, gm_n2276, in_14);
	nor (gm_n2278, gm_n81, gm_n46, gm_n63, gm_n2277, gm_n47);
	nand (gm_n2279, in_21, gm_n45, in_19, gm_n2278);
	or (gm_n2280, gm_n64, in_7, gm_n82, gm_n161, gm_n51);
	or (gm_n2281, in_12, in_11, gm_n52, gm_n2280, gm_n49);
	nor (gm_n2282, in_16, gm_n63, in_14, gm_n2281, gm_n81);
	nand (gm_n2283, in_20, in_19, in_18, gm_n2282, gm_n71);
	nor (gm_n2284, in_8, in_7, gm_n82, gm_n156, in_9);
	nand (gm_n2285, in_12, gm_n53, gm_n52, gm_n2284, in_13);
	nor (gm_n2286, in_16, in_15, in_14, gm_n2285, in_17);
	nand (gm_n2287, in_20, in_19, gm_n47, gm_n2286, gm_n71);
	nand (gm_n2288, gm_n1421, gm_n52, in_9);
	nor (gm_n2289, in_13, gm_n48, gm_n53, gm_n2288, gm_n50);
	nand (gm_n2290, gm_n81, in_16, gm_n63, gm_n2289, gm_n47);
	nor (gm_n2291, gm_n71, gm_n45, gm_n62, gm_n2290);
	nand (gm_n2292, in_10, in_9, in_8, gm_n1608, gm_n53);
	nor (gm_n2293, in_14, in_13, in_12, gm_n2292, gm_n63);
	nand (gm_n2294, in_18, in_17, in_16, gm_n2293, gm_n62);
	nor (gm_n2295, gm_n2294, gm_n71, in_20);
	or (gm_n2296, gm_n686, gm_n52, in_9);
	nor (gm_n2297, in_13, in_12, gm_n53, gm_n2296, in_14);
	nand (gm_n2298, gm_n81, gm_n46, gm_n63, gm_n2297, in_18);
	nor (gm_n2299, gm_n71, gm_n45, in_19, gm_n2298);
	nand (gm_n2300, in_7, in_6, in_5, gm_n598, in_8);
	or (gm_n2301, gm_n53, in_10, gm_n51, gm_n2300, gm_n48);
	nor (gm_n2302, in_15, in_14, gm_n49, gm_n2301);
	nand (gm_n2303, gm_n47, gm_n81, in_16, gm_n2302, in_19);
	nor (gm_n2304, gm_n2303, in_21, gm_n45);
	nor (gm_n2305, gm_n51, gm_n64, gm_n55, gm_n588, in_10);
	nand (gm_n2306, in_13, gm_n48, gm_n53, gm_n2305, in_14);
	nor (gm_n2307, gm_n81, gm_n46, in_15, gm_n2306, in_18);
	nand (gm_n2308, in_21, gm_n45, in_19, gm_n2307);
	or (gm_n2309, in_12, in_11, in_10, gm_n264, in_13);
	nor (gm_n2310, gm_n46, gm_n63, gm_n50, gm_n2309, in_17);
	nand (gm_n2311, gm_n45, in_19, in_18, gm_n2310, in_21);
	nor (gm_n2312, in_9, gm_n64, in_7, gm_n279, in_10);
	nand (gm_n2313, in_13, in_12, gm_n53, gm_n2312, gm_n50);
	nor (gm_n2314, in_17, in_16, gm_n63, gm_n2313, gm_n47);
	nand (gm_n2315, in_21, in_20, gm_n62, gm_n2314);
	nor (gm_n2316, gm_n52, in_9, gm_n64, gm_n478, gm_n53);
	nand (gm_n2317, in_14, gm_n49, in_12, gm_n2316, gm_n63);
	nor (gm_n2318, gm_n47, in_17, in_16, gm_n2317, gm_n62);
	nand (gm_n2319, gm_n2318, gm_n71, gm_n45);
	nor (gm_n2320, gm_n53, in_10, gm_n51, gm_n410, gm_n48);
	and (gm_n2321, in_15, gm_n50, in_13, gm_n2320, gm_n46);
	nand (gm_n2322, in_19, in_18, in_17, gm_n2321, in_20);
	nor (gm_n2323, gm_n2322, gm_n71);
	nor (gm_n2324, in_13, gm_n48, gm_n53, gm_n1920, gm_n50);
	nand (gm_n2325, in_17, gm_n46, in_15, gm_n2324, gm_n47);
	nor (gm_n2326, gm_n71, in_20, in_19, gm_n2325);
	nand (gm_n2327, gm_n64, in_7, gm_n82, gm_n638, in_9);
	nor (gm_n2328, gm_n48, in_11, gm_n52, gm_n2327, in_13);
	nand (gm_n2329, in_16, in_15, in_14, gm_n2328, gm_n81);
	nor (gm_n2330, gm_n45, in_19, gm_n47, gm_n2329, in_21);
	nor (gm_n2331, in_13, gm_n48, gm_n53, gm_n1289, in_14);
	nand (gm_n2332, gm_n81, in_16, in_15, gm_n2331, in_18);
	nor (gm_n2333, in_21, in_20, in_19, gm_n2332);
	and (gm_n2334, gm_n64, in_7, gm_n82, gm_n757, gm_n51);
	nand (gm_n2335, in_12, in_11, gm_n52, gm_n2334, gm_n49);
	nor (gm_n2336, gm_n46, gm_n63, in_14, gm_n2335, gm_n81);
	nand (gm_n2337, in_20, in_19, in_18, gm_n2336, in_21);
	or (gm_n2338, gm_n48, in_11, gm_n52, gm_n228, gm_n49);
	nor (gm_n2339, gm_n46, in_15, gm_n50, gm_n2338, gm_n81);
	nand (gm_n2340, gm_n45, in_19, in_18, gm_n2339, gm_n71);
	and (gm_n2341, gm_n53, in_10, in_9, gm_n1643, in_12);
	nand (gm_n2342, gm_n63, in_14, in_13, gm_n2341, gm_n46);
	nor (gm_n2343, gm_n62, gm_n47, in_17, gm_n2342, gm_n45);
	nand (gm_n2344, gm_n2343, gm_n71);
	nand (gm_n2345, in_7, gm_n82, gm_n72, gm_n209, gm_n64);
	nor (gm_n2346, gm_n53, gm_n52, in_9, gm_n2345, gm_n48);
	nand (gm_n2347, gm_n63, in_14, gm_n49, gm_n2346, gm_n46);
	nor (gm_n2348, gm_n2347, gm_n81);
	nand (gm_n2349, in_20, in_19, in_18, gm_n2348, gm_n71);
	nand (gm_n2350, in_17, in_16, gm_n63, gm_n1025, gm_n47);
	nor (gm_n2351, gm_n71, gm_n45, in_19, gm_n2350);
	nor (gm_n2352, in_12, gm_n53, in_10, gm_n162, in_13);
	nand (gm_n2353, in_16, in_15, in_14, gm_n2352, gm_n81);
	nor (gm_n2354, gm_n45, gm_n62, gm_n47, gm_n2353, in_21);
	or (gm_n2355, gm_n64, gm_n55, in_6, gm_n156, in_9);
	nor (gm_n2356, gm_n48, in_11, gm_n52, gm_n2355, gm_n49);
	nand (gm_n2357, gm_n46, in_15, gm_n50, gm_n2356, gm_n81);
	nor (gm_n2358, gm_n45, gm_n62, in_18, gm_n2357, gm_n71);
	nand (gm_n2359, gm_n612, in_10, gm_n51);
	nor (gm_n2360, gm_n49, in_12, in_11, gm_n2359, gm_n50);
	nand (gm_n2361, in_17, in_16, gm_n63, gm_n2360, in_18);
	nor (gm_n2362, in_21, gm_n45, gm_n62, gm_n2361);
	or (gm_n2363, in_12, in_11, gm_n52, gm_n898, gm_n49);
	nor (gm_n2364, in_16, in_15, gm_n50, gm_n2363, gm_n81);
	nand (gm_n2365, gm_n45, gm_n62, gm_n47, gm_n2364, in_21);
	nor (gm_n2366, in_11, in_10, in_9, gm_n322);
	nand (gm_n2367, gm_n50, gm_n49, in_12, gm_n2366, in_15);
	nor (gm_n2368, gm_n47, in_17, gm_n46, gm_n2367, in_19);
	nand (gm_n2369, gm_n2368, in_21, in_20);
	or (gm_n2370, gm_n64, gm_n55, in_6, gm_n199, gm_n51);
	nor (gm_n2371, gm_n2370, gm_n53, gm_n52);
	nand (gm_n2372, gm_n50, in_13, gm_n48, gm_n2371, gm_n63);
	nor (gm_n2373, in_18, gm_n81, gm_n46, gm_n2372, in_19);
	nand (gm_n2374, gm_n2373, gm_n71, in_20);
	nor (gm_n2375, gm_n53, gm_n52, gm_n51, gm_n426, gm_n48);
	nand (gm_n2376, gm_n63, gm_n50, gm_n49, gm_n2375, gm_n46);
	nor (gm_n2377, gm_n62, gm_n47, gm_n81, gm_n2376, gm_n45);
	nand (gm_n2378, gm_n2377, in_21);
	nor (gm_n2379, in_15, gm_n50, gm_n49, gm_n184, gm_n46);
	nand (gm_n2380, gm_n62, in_18, in_17, gm_n2379, in_20);
	nor (gm_n2381, gm_n2380, gm_n71);
	nand (gm_n2382, gm_n53, gm_n52, gm_n51, gm_n1643);
	nor (gm_n2383, in_14, gm_n49, gm_n48, gm_n2382, in_15);
	nand (gm_n2384, in_18, in_17, gm_n46, gm_n2383, in_19);
	nor (gm_n2385, gm_n2384, gm_n71, gm_n45);
	and (gm_n2386, in_13, in_12, in_11, gm_n85, gm_n50);
	nand (gm_n2387, in_17, gm_n46, gm_n63, gm_n2386, in_18);
	nor (gm_n2388, in_21, in_20, in_19, gm_n2387);
	nand (gm_n2389, gm_n621, gm_n52, in_9);
	nor (gm_n2390, in_13, in_12, gm_n53, gm_n2389, in_14);
	nand (gm_n2391, in_17, in_16, gm_n63, gm_n2390, in_18);
	nor (gm_n2392, in_21, gm_n45, gm_n62, gm_n2391);
	nor (gm_n2393, in_9, in_8, gm_n55, gm_n588, gm_n52);
	nand (gm_n2394, gm_n49, gm_n48, gm_n53, gm_n2393, gm_n50);
	nor (gm_n2395, gm_n81, gm_n46, gm_n63, gm_n2394, in_18);
	nand (gm_n2396, in_21, gm_n45, gm_n62, gm_n2395);
	nand (gm_n2397, in_7, gm_n82, in_5, gm_n209, in_8);
	nor (gm_n2398, in_11, in_10, in_9, gm_n2397, in_12);
	nand (gm_n2399, in_15, in_14, gm_n49, gm_n2398, in_16);
	nor (gm_n2400, gm_n62, in_18, in_17, gm_n2399, gm_n45);
	nand (gm_n2401, gm_n2400, gm_n71);
	nand (gm_n2402, gm_n48, gm_n53, gm_n52, gm_n968, gm_n49);
	nor (gm_n2403, in_16, gm_n63, gm_n50, gm_n2402, in_17);
	nand (gm_n2404, in_20, in_19, in_18, gm_n2403, in_21);
	and (gm_n2405, gm_n53, gm_n52, gm_n51, gm_n1142, in_12);
	nand (gm_n2406, gm_n2405, in_13);
	nor (gm_n2407, gm_n46, gm_n63, in_14, gm_n2406, in_17);
	nand (gm_n2408, in_20, in_19, gm_n47, gm_n2407, gm_n71);
	nor (gm_n2409, in_12, in_11, in_10, gm_n1836, in_13);
	nand (gm_n2410, in_16, gm_n63, in_14, gm_n2409, gm_n81);
	nor (gm_n2411, in_20, in_19, in_18, gm_n2410, in_21);
	nor (gm_n2412, in_12, gm_n53, gm_n52, gm_n1524, gm_n49);
	nand (gm_n2413, in_16, in_15, in_14, gm_n2412, gm_n81);
	nor (gm_n2414, gm_n45, gm_n62, in_18, gm_n2413, gm_n71);
	and (gm_n2415, gm_n51, gm_n64, gm_n55, gm_n136);
	and (gm_n2416, in_12, gm_n53, in_10, gm_n2415, in_13);
	nand (gm_n2417, in_16, in_15, gm_n50, gm_n2416, in_17);
	nor (gm_n2418, in_20, in_19, gm_n47, gm_n2417, in_21);
	nand (gm_n2419, gm_n55, gm_n82, in_5, gm_n252, in_8);
	nor (gm_n2420, gm_n53, gm_n52, gm_n51, gm_n2419);
	and (gm_n2421, gm_n50, in_13, in_12, gm_n2420, gm_n63);
	nand (gm_n2422, gm_n47, in_17, in_16, gm_n2421, in_19);
	nor (gm_n2423, gm_n2422, gm_n71, in_20);
	and (gm_n2424, in_11, gm_n52, in_9, gm_n612, in_12);
	nand (gm_n2425, gm_n63, gm_n50, in_13, gm_n2424, in_16);
	nor (gm_n2426, in_19, in_18, gm_n81, gm_n2425, gm_n45);
	nand (gm_n2427, gm_n2426, in_21);
	nand (gm_n2428, gm_n1528, gm_n52, in_9);
	or (gm_n2429, gm_n49, in_12, in_11, gm_n2428, gm_n50);
	nor (gm_n2430, gm_n81, in_16, in_15, gm_n2429, in_18);
	nand (gm_n2431, in_21, gm_n45, in_19, gm_n2430);
	and (gm_n2432, gm_n55, gm_n82, in_5, gm_n209, in_8);
	and (gm_n2433, gm_n53, gm_n52, in_9, gm_n2432);
	nand (gm_n2434, in_14, in_13, gm_n48, gm_n2433, gm_n63);
	nor (gm_n2435, gm_n47, gm_n81, in_16, gm_n2434, gm_n62);
	nand (gm_n2436, gm_n2435, in_21, in_20);
	nor (gm_n2437, gm_n52, in_9, gm_n64, gm_n853, in_11);
	nand (gm_n2438, gm_n50, gm_n49, gm_n48, gm_n2437, in_15);
	nor (gm_n2439, gm_n47, in_17, gm_n46, gm_n2438, gm_n62);
	nand (gm_n2440, gm_n2439, gm_n71, in_20);
	nor (gm_n2441, in_9, in_8, gm_n55, gm_n279);
	and (gm_n2442, gm_n48, in_11, gm_n52, gm_n2441, gm_n49);
	nand (gm_n2443, in_16, gm_n63, gm_n50, gm_n2442, gm_n81);
	nor (gm_n2444, in_20, in_19, in_18, gm_n2443, in_21);
	nand (gm_n2445, in_7, in_6, gm_n72, gm_n296, in_8);
	nor (gm_n2446, in_11, in_10, in_9, gm_n2445, in_12);
	and (gm_n2447, gm_n63, in_14, in_13, gm_n2446);
	nand (gm_n2448, gm_n47, gm_n81, gm_n46, gm_n2447, in_19);
	nor (gm_n2449, gm_n2448, gm_n71, in_20);
	nand (gm_n2450, in_11, gm_n52, gm_n51, gm_n673, in_12);
	nor (gm_n2451, gm_n63, gm_n50, in_13, gm_n2450, gm_n46);
	nand (gm_n2452, gm_n62, gm_n47, gm_n81, gm_n2451, gm_n45);
	nor (gm_n2453, gm_n2452, gm_n71);
	nor (gm_n2454, gm_n48, in_11, gm_n52, gm_n1836, in_13);
	nand (gm_n2455, in_16, gm_n63, in_14, gm_n2454, gm_n81);
	nor (gm_n2456, gm_n45, in_19, gm_n47, gm_n2455, gm_n71);
	nand (gm_n2457, in_14, in_13, gm_n48, gm_n1870, gm_n63);
	nor (gm_n2458, gm_n47, gm_n81, gm_n46, gm_n2457, gm_n62);
	nand (gm_n2459, gm_n2458, gm_n71, gm_n45);
	and (gm_n2460, in_11, gm_n52, gm_n51, gm_n1302, gm_n48);
	nand (gm_n2461, in_15, gm_n50, in_13, gm_n2460, gm_n46);
	nor (gm_n2462, in_19, in_18, gm_n81, gm_n2461, gm_n45);
	nand (gm_n2463, gm_n2462, gm_n71);
	nor (gm_n2464, gm_n1261, in_10, in_9);
	nand (gm_n2465, gm_n49, gm_n48, in_11, gm_n2464, gm_n50);
	nor (gm_n2466, gm_n81, gm_n46, gm_n63, gm_n2465, in_18);
	nand (gm_n2467, in_21, gm_n45, gm_n62, gm_n2466);
	nor (gm_n2468, in_11, in_10, in_9, gm_n649, in_12);
	nand (gm_n2469, in_15, in_14, in_13, gm_n2468, in_16);
	nor (gm_n2470, in_19, gm_n47, in_17, gm_n2469, gm_n45);
	nand (gm_n2471, gm_n2470, in_21);
	nor (gm_n2472, in_7, gm_n82, in_5, gm_n867, gm_n64);
	nand (gm_n2473, gm_n2472, in_10, in_9);
	nor (gm_n2474, gm_n49, in_12, gm_n53, gm_n2473, in_14);
	nand (gm_n2475, in_17, gm_n46, in_15, gm_n2474, gm_n47);
	nor (gm_n2476, in_21, gm_n45, gm_n62, gm_n2475);
	nand (gm_n2477, in_9, gm_n64, gm_n55, gm_n504, in_10);
	nor (gm_n2478, gm_n49, gm_n48, gm_n53, gm_n2477, in_14);
	nand (gm_n2479, in_17, in_16, in_15, gm_n2478, in_18);
	nor (gm_n2480, in_21, in_20, gm_n62, gm_n2479);
	and (gm_n2481, gm_n55, gm_n82, gm_n72, gm_n493, gm_n64);
	and (gm_n2482, gm_n2481, in_9);
	and (gm_n2483, in_12, gm_n53, in_10, gm_n2482, gm_n49);
	nand (gm_n2484, in_16, in_15, gm_n50, gm_n2483, in_17);
	nor (gm_n2485, in_20, in_19, gm_n47, gm_n2484, gm_n71);
	and (gm_n2486, in_12, in_11, gm_n52, gm_n1376, in_13);
	nand (gm_n2487, in_16, gm_n63, gm_n50, gm_n2486, gm_n81);
	nor (gm_n2488, in_20, gm_n62, in_18, gm_n2487, in_21);
	nand (gm_n2489, gm_n48, gm_n53, gm_n52, gm_n1945, gm_n49);
	nor (gm_n2490, gm_n46, in_15, gm_n50, gm_n2489, gm_n81);
	nand (gm_n2491, in_20, gm_n62, gm_n47, gm_n2490, in_21);
	nand (gm_n2492, gm_n48, in_11, gm_n52, gm_n889, gm_n49);
	nor (gm_n2493, in_16, gm_n63, gm_n50, gm_n2492, in_17);
	nand (gm_n2494, gm_n45, gm_n62, in_18, gm_n2493, gm_n71);
	nor (gm_n2495, in_9, gm_n64, in_7, gm_n843, gm_n52);
	nand (gm_n2496, in_13, gm_n48, gm_n53, gm_n2495, in_14);
	nor (gm_n2497, gm_n81, gm_n46, in_15, gm_n2496, in_18);
	nand (gm_n2498, in_21, in_20, in_19, gm_n2497);
	and (gm_n2499, gm_n1070, in_10, in_9);
	nand (gm_n2500, gm_n49, in_12, in_11, gm_n2499, in_14);
	nor (gm_n2501, gm_n81, in_16, in_15, gm_n2500, in_18);
	nand (gm_n2502, gm_n71, gm_n45, in_19, gm_n2501);
	nand (gm_n2503, in_7, in_6, gm_n72, gm_n598, gm_n64);
	or (gm_n2504, gm_n53, gm_n52, in_9, gm_n2503);
	nor (gm_n2505, in_14, gm_n49, in_12, gm_n2504);
	nand (gm_n2506, gm_n81, in_16, gm_n63, gm_n2505, gm_n47);
	nor (gm_n2507, in_21, gm_n45, gm_n62, gm_n2506);
	nor (gm_n2508, gm_n55, gm_n82, in_5, gm_n483, gm_n64);
	nand (gm_n2509, in_11, gm_n52, gm_n51, gm_n2508, in_12);
	nor (gm_n2510, gm_n63, in_14, in_13, gm_n2509, in_16);
	nand (gm_n2511, gm_n62, gm_n47, gm_n81, gm_n2510, in_20);
	nor (gm_n2512, gm_n2511, gm_n71);
	nor (gm_n2513, gm_n55, gm_n82, gm_n72, gm_n321, gm_n64);
	nand (gm_n2514, gm_n2513, gm_n52, gm_n51);
	nor (gm_n2515, gm_n49, in_12, in_11, gm_n2514, gm_n50);
	nand (gm_n2516, in_17, in_16, in_15, gm_n2515, in_18);
	nor (gm_n2517, in_21, gm_n45, gm_n62, gm_n2516);
	or (gm_n2518, gm_n51, in_8, in_7, gm_n463, gm_n52);
	nor (gm_n2519, in_13, gm_n48, in_11, gm_n2518, in_14);
	nand (gm_n2520, in_17, gm_n46, in_15, gm_n2519, in_18);
	nor (gm_n2521, in_21, in_20, in_19, gm_n2520);
	nor (gm_n2522, in_8, gm_n55, in_6, gm_n156, in_9);
	nand (gm_n2523, gm_n48, gm_n53, gm_n52, gm_n2522, in_13);
	nor (gm_n2524, gm_n46, in_15, gm_n50, gm_n2523, in_17);
	nand (gm_n2525, in_20, gm_n62, gm_n47, gm_n2524, gm_n71);
	nor (gm_n2526, in_7, gm_n82, gm_n72, gm_n867, in_8);
	and (gm_n2527, in_11, gm_n52, in_9, gm_n2526, in_12);
	nand (gm_n2528, in_15, in_14, gm_n49, gm_n2527, gm_n46);
	nor (gm_n2529, in_19, in_18, in_17, gm_n2528, gm_n45);
	nand (gm_n2530, gm_n2529, gm_n71);
	or (gm_n2531, gm_n48, gm_n53, gm_n52, gm_n162, gm_n49);
	nor (gm_n2532, gm_n46, gm_n63, gm_n50, gm_n2531, gm_n81);
	nand (gm_n2533, gm_n45, gm_n62, in_18, gm_n2532, in_21);
	nor (gm_n2534, in_9, gm_n64, gm_n55, gm_n553, in_10);
	nand (gm_n2535, in_13, in_12, in_11, gm_n2534, in_14);
	nor (gm_n2536, in_17, gm_n46, in_15, gm_n2535, gm_n47);
	nand (gm_n2537, in_21, in_20, in_19, gm_n2536);
	and (gm_n2538, in_10, in_9, gm_n64, gm_n1608, gm_n53);
	and (gm_n2539, in_14, gm_n49, gm_n48, gm_n2538, gm_n63);
	nand (gm_n2540, gm_n47, in_17, in_16, gm_n2539, gm_n62);
	nor (gm_n2541, gm_n2540, in_21, in_20);
	nand (gm_n2542, in_10, in_9, gm_n64, gm_n663, gm_n53);
	nor (gm_n2543, in_14, in_13, in_12, gm_n2542, gm_n63);
	nand (gm_n2544, in_18, gm_n81, in_16, gm_n2543, gm_n62);
	nor (gm_n2545, gm_n2544, gm_n71, in_20);
	nand (gm_n2546, gm_n55, gm_n82, in_5, gm_n420, in_8);
	or (gm_n2547, gm_n53, in_10, gm_n51, gm_n2546, gm_n48);
	nor (gm_n2548, gm_n2547, in_14, gm_n49);
	nand (gm_n2549, gm_n81, gm_n46, in_15, gm_n2548, gm_n47);
	nor (gm_n2550, gm_n71, gm_n45, gm_n62, gm_n2549);
	nor (gm_n2551, in_8, in_7, in_6, gm_n161, gm_n51);
	and (gm_n2552, gm_n48, gm_n53, gm_n52, gm_n2551, gm_n49);
	nand (gm_n2553, in_16, in_15, in_14, gm_n2552, gm_n81);
	nor (gm_n2554, in_20, gm_n62, in_18, gm_n2553, gm_n71);
	nor (gm_n2555, in_8, in_7, in_6, gm_n103, gm_n51);
	nand (gm_n2556, in_12, in_11, in_10, gm_n2555, gm_n49);
	nor (gm_n2557, in_16, in_15, in_14, gm_n2556, gm_n81);
	nand (gm_n2558, in_20, in_19, in_18, gm_n2557, gm_n71);
	nand (gm_n2559, gm_n55, gm_n82, gm_n72, gm_n1126, gm_n64);
	nor (gm_n2560, in_11, gm_n52, in_9, gm_n2559, gm_n48);
	nand (gm_n2561, gm_n63, gm_n50, in_13, gm_n2560, in_16);
	nor (gm_n2562, gm_n62, gm_n47, in_17, gm_n2561, gm_n45);
	nand (gm_n2563, gm_n2562, gm_n71);
	nand (gm_n2564, gm_n55, in_6, gm_n72, gm_n598, gm_n64);
	nor (gm_n2565, in_11, in_10, gm_n51, gm_n2564, in_12);
	nand (gm_n2566, gm_n63, gm_n50, gm_n49, gm_n2565, gm_n46);
	nor (gm_n2567, gm_n62, in_18, in_17, gm_n2566, gm_n45);
	nand (gm_n2568, gm_n2567, in_21);
	nand (gm_n2569, in_12, in_11, gm_n52, gm_n146, in_13);
	nor (gm_n2570, gm_n46, in_15, gm_n50, gm_n2569, gm_n81);
	nand (gm_n2571, gm_n45, in_19, in_18, gm_n2570, in_21);
	and (gm_n2572, gm_n49, in_12, in_11, gm_n1644);
	nand (gm_n2573, gm_n46, in_15, gm_n50, gm_n2572, in_17);
	nor (gm_n2574, gm_n45, gm_n62, in_18, gm_n2573, gm_n71);
	nand (gm_n2575, in_9, gm_n64, in_7, gm_n1007, in_10);
	nor (gm_n2576, gm_n49, gm_n48, in_11, gm_n2575, gm_n50);
	nand (gm_n2577, in_17, gm_n46, gm_n63, gm_n2576, gm_n47);
	nor (gm_n2578, gm_n71, in_20, in_19, gm_n2577);
	nor (gm_n2579, gm_n49, gm_n48, gm_n53, gm_n2225, in_14);
	nand (gm_n2580, gm_n81, in_16, gm_n63, gm_n2579, gm_n47);
	nor (gm_n2581, gm_n71, in_20, in_19, gm_n2580);
	nand (gm_n2582, in_9, gm_n64, in_7, gm_n404, gm_n52);
	nor (gm_n2583, in_13, in_12, in_11, gm_n2582, gm_n50);
	nand (gm_n2584, gm_n81, gm_n46, gm_n63, gm_n2583, gm_n47);
	nor (gm_n2585, gm_n71, in_20, in_19, gm_n2584);
	nand (gm_n2586, in_13, in_12, in_11, gm_n1435, gm_n50);
	nor (gm_n2587, in_17, in_16, in_15, gm_n2586, in_18);
	nand (gm_n2588, in_21, gm_n45, in_19, gm_n2587);
	nand (gm_n2589, gm_n2047, in_10, gm_n51);
	nor (gm_n2590, in_13, in_12, in_11, gm_n2589, gm_n50);
	and (gm_n2591, gm_n81, gm_n46, gm_n63, gm_n2590, in_18);
	nand (gm_n2592, in_21, in_20, in_19, gm_n2591);
	nor (gm_n2593, gm_n2419, in_9);
	nand (gm_n2594, gm_n48, in_11, in_10, gm_n2593, in_13);
	nor (gm_n2595, gm_n46, gm_n63, in_14, gm_n2594, gm_n81);
	nand (gm_n2596, gm_n45, in_19, in_18, gm_n2595, gm_n71);
	nand (gm_n2597, gm_n51, in_8, gm_n55, gm_n404);
	nor (gm_n2598, gm_n48, gm_n53, in_10, gm_n2597, gm_n49);
	and (gm_n2599, in_16, gm_n63, in_14, gm_n2598, gm_n81);
	nand (gm_n2600, gm_n45, gm_n62, gm_n47, gm_n2599, in_21);
	and (gm_n2601, gm_n55, in_6, in_5, gm_n296, in_8);
	nand (gm_n2602, gm_n2601, gm_n52, in_9);
	nor (gm_n2603, gm_n49, in_12, gm_n53, gm_n2602, gm_n50);
	nand (gm_n2604, gm_n81, in_16, in_15, gm_n2603, in_18);
	nor (gm_n2605, in_21, gm_n45, gm_n62, gm_n2604);
	nand (gm_n2606, gm_n53, gm_n52, gm_n51, gm_n2601, gm_n48);
	nor (gm_n2607, gm_n63, gm_n50, gm_n49, gm_n2606, in_16);
	nand (gm_n2608, in_19, gm_n47, in_17, gm_n2607, in_20);
	nor (gm_n2609, gm_n2608, gm_n71);
	nand (gm_n2610, gm_n55, gm_n82, in_5, gm_n89, in_8);
	nor (gm_n2611, gm_n2610, in_10, gm_n51);
	and (gm_n2612, in_13, gm_n48, in_11, gm_n2611, gm_n50);
	nand (gm_n2613, in_17, in_16, gm_n63, gm_n2612, in_18);
	nor (gm_n2614, in_21, gm_n45, gm_n62, gm_n2613);
	or (gm_n2615, gm_n53, gm_n52, in_9, gm_n1098, gm_n48);
	nor (gm_n2616, in_15, gm_n50, in_13, gm_n2615, gm_n46);
	nand (gm_n2617, gm_n62, in_18, in_17, gm_n2616, gm_n45);
	nor (gm_n2618, gm_n2617, in_21);
	nor (gm_n2619, in_8, gm_n55, gm_n82, gm_n119, in_9);
	nand (gm_n2620, in_12, gm_n53, in_10, gm_n2619, in_13);
	nor (gm_n2621, in_16, gm_n63, in_14, gm_n2620, in_17);
	nand (gm_n2622, in_20, in_19, in_18, gm_n2621, gm_n71);
	nand (gm_n2623, gm_n1165, in_9);
	or (gm_n2624, gm_n48, gm_n53, gm_n52, gm_n2623, in_13);
	nor (gm_n2625, gm_n46, in_15, gm_n50, gm_n2624, gm_n81);
	nand (gm_n2626, gm_n45, in_19, gm_n47, gm_n2625, in_21);
	and (gm_n2627, gm_n53, in_10, gm_n51, gm_n2088);
	nand (gm_n2628, in_14, gm_n49, gm_n48, gm_n2627, gm_n63);
	nor (gm_n2629, gm_n47, gm_n81, in_16, gm_n2628, in_19);
	nand (gm_n2630, gm_n2629, gm_n71, gm_n45);
	and (gm_n2631, in_7, in_6, gm_n72, gm_n296, gm_n64);
	and (gm_n2632, gm_n53, gm_n52, gm_n51, gm_n2631, in_12);
	nand (gm_n2633, gm_n63, in_14, gm_n49, gm_n2632, gm_n46);
	nor (gm_n2634, gm_n62, in_18, gm_n81, gm_n2633, in_20);
	nand (gm_n2635, gm_n2634, gm_n71);
	nand (gm_n2636, in_11, in_10, gm_n51, gm_n1156, in_12);
	nor (gm_n2637, in_15, gm_n50, gm_n49, gm_n2636, in_16);
	nand (gm_n2638, in_19, in_18, in_17, gm_n2637, gm_n45);
	nor (gm_n2639, gm_n2638, in_21);
	nor (gm_n2640, in_4, in_3, in_2, gm_n373, gm_n72);
	and (gm_n2641, gm_n64, gm_n55, gm_n82, gm_n2640, in_9);
	and (gm_n2642, gm_n48, in_11, in_10, gm_n2641, gm_n49);
	nand (gm_n2643, in_16, gm_n63, gm_n50, gm_n2642, in_17);
	nor (gm_n2644, gm_n45, in_19, in_18, gm_n2643, in_21);
	nand (gm_n2645, in_8, in_7, gm_n82, gm_n757, in_9);
	nor (gm_n2646, in_12, gm_n53, gm_n52, gm_n2645, gm_n49);
	nand (gm_n2647, gm_n46, gm_n63, gm_n50, gm_n2646, in_17);
	nor (gm_n2648, gm_n45, gm_n62, in_18, gm_n2647, gm_n71);
	nand (gm_n2649, gm_n53, in_10, gm_n51, gm_n1856, in_12);
	nor (gm_n2650, gm_n63, gm_n50, in_13, gm_n2649, gm_n46);
	nand (gm_n2651, in_19, gm_n47, in_17, gm_n2650, in_20);
	nor (gm_n2652, gm_n2651, gm_n71);
	nor (gm_n2653, in_7, gm_n82, in_5, gm_n124, gm_n64);
	and (gm_n2654, in_11, in_10, in_9, gm_n2653);
	nand (gm_n2655, gm_n50, gm_n49, gm_n48, gm_n2654, in_15);
	nor (gm_n2656, gm_n2655, in_17, in_16);
	nand (gm_n2657, in_20, in_19, in_18, gm_n2656, gm_n71);
	nor (gm_n2658, in_12, gm_n53, in_10, gm_n1723, in_13);
	and (gm_n2659, gm_n46, gm_n63, in_14, gm_n2658, gm_n81);
	nand (gm_n2660, in_20, gm_n62, in_18, gm_n2659, gm_n71);
	and (gm_n2661, gm_n64, in_7, gm_n82, gm_n374, gm_n51);
	nand (gm_n2662, in_12, gm_n53, gm_n52, gm_n2661, gm_n49);
	nor (gm_n2663, gm_n46, in_15, in_14, gm_n2662, in_17);
	nand (gm_n2664, gm_n45, gm_n62, in_18, gm_n2663, gm_n71);
	and (gm_n2665, gm_n53, gm_n52, in_9, gm_n494, in_12);
	nand (gm_n2666, gm_n63, gm_n50, gm_n49, gm_n2665, in_16);
	nor (gm_n2667, in_19, in_18, gm_n81, gm_n2666, in_20);
	nand (gm_n2668, gm_n2667, gm_n71);
	and (gm_n2669, gm_n49, in_12, in_11, gm_n526, in_14);
	nand (gm_n2670, gm_n81, in_16, in_15, gm_n2669, gm_n47);
	nor (gm_n2671, in_21, in_20, in_19, gm_n2670);
	and (gm_n2672, in_8, in_7, in_6, gm_n638, in_9);
	and (gm_n2673, gm_n48, gm_n53, gm_n52, gm_n2672, gm_n49);
	nand (gm_n2674, in_16, in_15, gm_n50, gm_n2673, in_17);
	nor (gm_n2675, gm_n45, gm_n62, in_18, gm_n2674, in_21);
	nor (gm_n2676, in_7, in_6, gm_n72, gm_n188, gm_n64);
	nand (gm_n2677, gm_n2676, gm_n52, gm_n51);
	nor (gm_n2678, gm_n49, in_12, in_11, gm_n2677, gm_n50);
	nand (gm_n2679, in_17, gm_n46, gm_n63, gm_n2678, in_18);
	nor (gm_n2680, gm_n71, in_20, gm_n62, gm_n2679);
	and (gm_n2681, in_8, in_7, gm_n82, gm_n638, gm_n51);
	and (gm_n2682, in_12, in_11, in_10, gm_n2681, in_13);
	nand (gm_n2683, gm_n46, in_15, in_14, gm_n2682, in_17);
	nor (gm_n2684, gm_n45, in_19, gm_n47, gm_n2683, in_21);
	nor (gm_n2685, gm_n64, gm_n55, gm_n82, gm_n103, gm_n51);
	nand (gm_n2686, in_12, in_11, gm_n52, gm_n2685, in_13);
	nor (gm_n2687, in_16, gm_n63, gm_n50, gm_n2686, in_17);
	nand (gm_n2688, gm_n45, in_19, in_18, gm_n2687, in_21);
	or (gm_n2689, gm_n53, gm_n52, gm_n51, gm_n1879, in_12);
	or (gm_n2690, in_15, gm_n50, in_13, gm_n2689, in_16);
	nor (gm_n2691, gm_n62, in_18, gm_n81, gm_n2690, in_20);
	nand (gm_n2692, gm_n2691, in_21);
	nor (gm_n2693, gm_n64, gm_n55, in_6, gm_n199, in_9);
	nand (gm_n2694, gm_n48, in_11, in_10, gm_n2693, gm_n49);
	nor (gm_n2695, in_16, gm_n63, gm_n50, gm_n2694, gm_n81);
	nand (gm_n2696, in_20, gm_n62, gm_n47, gm_n2695, in_21);
	and (gm_n2697, gm_n81, gm_n46, in_15, gm_n318, gm_n47);
	nand (gm_n2698, in_21, in_20, gm_n62, gm_n2697);
	nor (gm_n2699, gm_n55, in_6, gm_n72, gm_n867, in_8);
	nand (gm_n2700, gm_n2699, gm_n52, gm_n51);
	nor (gm_n2701, in_13, in_12, gm_n53, gm_n2700, in_14);
	nand (gm_n2702, in_17, in_16, in_15, gm_n2701, gm_n47);
	nor (gm_n2703, in_21, in_20, in_19, gm_n2702);
	nand (gm_n2704, in_11, in_10, in_9, gm_n1634, in_12);
	nor (gm_n2705, in_15, gm_n50, gm_n49, gm_n2704, in_16);
	nand (gm_n2706, in_19, gm_n47, in_17, gm_n2705, gm_n45);
	nor (gm_n2707, gm_n2706, in_21);
	nor (gm_n2708, in_6, in_5, in_4, gm_n315, gm_n55);
	nand (gm_n2709, in_10, in_9, gm_n64, gm_n2708, in_11);
	nor (gm_n2710, in_14, in_13, in_12, gm_n2709, in_15);
	nand (gm_n2711, gm_n47, in_17, gm_n46, gm_n2710, in_19);
	nor (gm_n2712, gm_n2711, gm_n71, in_20);
	nand (gm_n2713, gm_n53, gm_n52, gm_n51, gm_n1192, in_12);
	nor (gm_n2714, gm_n63, in_14, in_13, gm_n2713, gm_n46);
	nand (gm_n2715, gm_n62, gm_n47, gm_n81, gm_n2714, gm_n45);
	nor (gm_n2716, gm_n2715, gm_n71);
	nand (gm_n2717, gm_n63, gm_n50, in_13, gm_n356, gm_n46);
	nor (gm_n2718, in_19, in_18, gm_n81, gm_n2717, in_20);
	nand (gm_n2719, gm_n2718, in_21);
	or (gm_n2720, in_8, in_7, in_6, gm_n204, gm_n51);
	nor (gm_n2721, gm_n2720, in_10);
	nand (gm_n2722, gm_n49, in_12, in_11, gm_n2721, gm_n50);
	nor (gm_n2723, gm_n81, in_16, in_15, gm_n2722, gm_n47);
	nand (gm_n2724, gm_n71, gm_n45, in_19, gm_n2723);
	nor (gm_n2725, gm_n2397, gm_n52, gm_n51);
	nand (gm_n2726, in_13, gm_n48, in_11, gm_n2725, gm_n50);
	nor (gm_n2727, gm_n81, in_16, gm_n63, gm_n2726, in_18);
	nand (gm_n2728, gm_n71, gm_n45, in_19, gm_n2727);
	and (gm_n2729, gm_n64, gm_n55, in_6, gm_n379, in_9);
	nand (gm_n2730, gm_n48, in_11, gm_n52, gm_n2729, gm_n49);
	nor (gm_n2731, gm_n46, gm_n63, in_14, gm_n2730, in_17);
	nand (gm_n2732, in_20, gm_n62, gm_n47, gm_n2731, gm_n71);
	nor (gm_n2733, gm_n49, gm_n48, gm_n53, gm_n2359, gm_n50);
	nand (gm_n2734, gm_n81, gm_n46, in_15, gm_n2733, in_18);
	nor (gm_n2735, in_21, gm_n45, in_19, gm_n2734);
	nor (gm_n2736, in_12, gm_n53, gm_n52, gm_n1372, in_13);
	nand (gm_n2737, gm_n46, gm_n63, in_14, gm_n2736, gm_n81);
	nor (gm_n2738, gm_n45, gm_n62, in_18, gm_n2737, in_21);
	nand (gm_n2739, in_11, in_10, gm_n51, gm_n1057);
	nor (gm_n2740, in_14, in_13, in_12, gm_n2739, gm_n63);
	nand (gm_n2741, in_18, in_17, in_16, gm_n2740, in_19);
	nor (gm_n2742, gm_n2741, gm_n71, in_20);
	nand (gm_n2743, gm_n64, in_7, in_6, gm_n2640, in_9);
	nor (gm_n2744, in_12, gm_n53, gm_n52, gm_n2743, in_13);
	nand (gm_n2745, in_16, gm_n63, in_14, gm_n2744, in_17);
	nor (gm_n2746, in_20, in_19, gm_n47, gm_n2745, gm_n71);
	nor (gm_n2747, gm_n46, gm_n63, in_14, gm_n913, in_17);
	nand (gm_n2748, in_20, gm_n62, in_18, gm_n2747, gm_n71);
	nor (gm_n2749, gm_n64, in_7, gm_n82, gm_n119, in_9);
	nand (gm_n2750, gm_n48, in_11, gm_n52, gm_n2749, gm_n49);
	nor (gm_n2751, gm_n46, in_15, gm_n50, gm_n2750, gm_n81);
	nand (gm_n2752, in_20, in_19, in_18, gm_n2751, in_21);
	nor (gm_n2753, gm_n64, gm_n55, gm_n82, gm_n141, gm_n51);
	nand (gm_n2754, in_12, gm_n53, gm_n52, gm_n2753, in_13);
	nor (gm_n2755, gm_n46, gm_n63, gm_n50, gm_n2754, gm_n81);
	nand (gm_n2756, gm_n45, in_19, gm_n47, gm_n2755, in_21);
	nand (gm_n2757, in_12, gm_n53, gm_n52, gm_n678, in_13);
	nor (gm_n2758, in_16, gm_n63, gm_n50, gm_n2757, in_17);
	nand (gm_n2759, in_20, in_19, in_18, gm_n2758, gm_n71);
	nor (gm_n2760, in_8, gm_n55, in_6, gm_n530, gm_n51);
	nand (gm_n2761, gm_n48, gm_n53, in_10, gm_n2760, in_13);
	nor (gm_n2762, in_16, gm_n63, in_14, gm_n2761, in_17);
	nand (gm_n2763, gm_n45, gm_n62, gm_n47, gm_n2762, in_21);
	nand (gm_n2764, gm_n2756, gm_n2752, gm_n2748, gm_n2763, gm_n2759);
	nor (gm_n2765, gm_n2742, gm_n2738, gm_n2735, gm_n2764, gm_n2746);
	nand (gm_n2766, gm_n2728, gm_n2724, gm_n2719, gm_n2765, gm_n2732);
	nor (gm_n2767, gm_n2712, gm_n2707, gm_n2703, gm_n2766, gm_n2716);
	nand (gm_n2768, gm_n2696, gm_n2692, gm_n2688, gm_n2767, gm_n2698);
	nor (gm_n2769, gm_n2680, gm_n2675, gm_n2671, gm_n2768, gm_n2684);
	nand (gm_n2770, gm_n2664, gm_n2660, gm_n2657, gm_n2769, gm_n2668);
	nor (gm_n2771, gm_n2648, gm_n2644, gm_n2639, gm_n2770, gm_n2652);
	nand (gm_n2772, gm_n2630, gm_n2626, gm_n2622, gm_n2771, gm_n2635);
	nor (gm_n2773, gm_n2614, gm_n2609, gm_n2605, gm_n2772, gm_n2618);
	nand (gm_n2774, gm_n2596, gm_n2592, gm_n2588, gm_n2773, gm_n2600);
	nor (gm_n2775, gm_n2581, gm_n2578, gm_n2574, gm_n2774, gm_n2585);
	nand (gm_n2776, gm_n2568, gm_n2563, gm_n2558, gm_n2775, gm_n2571);
	nor (gm_n2777, gm_n2550, gm_n2545, gm_n2541, gm_n2776, gm_n2554);
	nand (gm_n2778, gm_n2533, gm_n2530, gm_n2525, gm_n2777, gm_n2537);
	nor (gm_n2779, gm_n2517, gm_n2512, gm_n2507, gm_n2778, gm_n2521);
	nand (gm_n2780, gm_n2498, gm_n2494, gm_n2491, gm_n2779, gm_n2502);
	nor (gm_n2781, gm_n2485, gm_n2480, gm_n2476, gm_n2780, gm_n2488);
	nand (gm_n2782, gm_n2467, gm_n2463, gm_n2459, gm_n2781, gm_n2471);
	nor (gm_n2783, gm_n2453, gm_n2449, gm_n2444, gm_n2782, gm_n2456);
	nand (gm_n2784, gm_n2436, gm_n2431, gm_n2427, gm_n2783, gm_n2440);
	nor (gm_n2785, gm_n2418, gm_n2414, gm_n2411, gm_n2784, gm_n2423);
	nand (gm_n2786, gm_n2404, gm_n2401, gm_n2396, gm_n2785, gm_n2408);
	nor (gm_n2787, gm_n2388, gm_n2385, gm_n2381, gm_n2786, gm_n2392);
	nand (gm_n2788, gm_n2374, gm_n2369, gm_n2365, gm_n2787, gm_n2378);
	nor (gm_n2789, gm_n2358, gm_n2354, gm_n2351, gm_n2788, gm_n2362);
	nand (gm_n2790, gm_n2344, gm_n2340, gm_n2337, gm_n2789, gm_n2349);
	nor (gm_n2791, gm_n2330, gm_n2326, gm_n2323, gm_n2790, gm_n2333);
	nand (gm_n2792, gm_n2315, gm_n2311, gm_n2308, gm_n2791, gm_n2319);
	nor (gm_n2793, gm_n2299, gm_n2295, gm_n2291, gm_n2792, gm_n2304);
	nand (gm_n2794, gm_n2283, gm_n2279, gm_n2274, gm_n2793, gm_n2287);
	nor (gm_n2795, gm_n2265, gm_n2261, gm_n2258, gm_n2794, gm_n2270);
	nand (gm_n2796, gm_n2250, gm_n2247, gm_n2243, gm_n2795, gm_n2253);
	nor (gm_n2797, gm_n2233, gm_n2228, gm_n2224, gm_n2796, gm_n2238);
	nand (gm_n2798, gm_n2217, gm_n2213, gm_n2209, gm_n2797, gm_n2221);
	nor (gm_n2799, gm_n2202, gm_n2198, gm_n2193, gm_n2798, gm_n2206);
	nand (gm_n2800, gm_n2185, gm_n2180, gm_n2177, gm_n2799, gm_n2189);
	nor (out_3, gm_n2800, gm_n2174);
	nor (gm_n2802, gm_n1316, gm_n50, in_13);
	nand (gm_n2803, in_17, in_16, in_15, gm_n2802, gm_n47);
	nor (gm_n2804, gm_n71, gm_n45, gm_n62, gm_n2803);
	nor (gm_n2805, gm_n49, in_12, gm_n53, gm_n2518, in_14);
	nand (gm_n2806, gm_n81, in_16, in_15, gm_n2805, gm_n47);
	nor (gm_n2807, in_21, gm_n45, gm_n62, gm_n2806);
	and (gm_n2808, gm_n50, in_13, gm_n48, gm_n567, in_15);
	nand (gm_n2809, in_18, gm_n81, gm_n46, gm_n2808, gm_n62);
	nor (gm_n2810, gm_n2809, gm_n71, gm_n45);
	nand (gm_n2811, in_9, in_8, gm_n55, gm_n1007, gm_n52);
	nor (gm_n2812, in_13, in_12, gm_n53, gm_n2811, gm_n50);
	nand (gm_n2813, gm_n81, gm_n46, gm_n63, gm_n2812, gm_n47);
	nor (gm_n2814, in_21, gm_n45, in_19, gm_n2813);
	nor (gm_n2815, gm_n90, gm_n52, gm_n51);
	nand (gm_n2816, gm_n49, in_12, in_11, gm_n2815, in_14);
	nor (gm_n2817, gm_n81, in_16, gm_n63, gm_n2816, gm_n47);
	nand (gm_n2818, gm_n71, in_20, gm_n62, gm_n2817);
	and (gm_n2819, in_8, in_7, in_6, gm_n1075, gm_n51);
	nand (gm_n2820, in_12, gm_n53, gm_n52, gm_n2819, gm_n49);
	nor (gm_n2821, in_16, in_15, gm_n50, gm_n2820, in_17);
	nand (gm_n2822, in_20, in_19, gm_n47, gm_n2821, gm_n71);
	nand (gm_n2823, in_7, in_6, gm_n72, gm_n252, gm_n64);
	nor (gm_n2824, gm_n53, gm_n52, gm_n51, gm_n2823);
	nand (gm_n2825, gm_n50, in_13, gm_n48, gm_n2824, in_15);
	nor (gm_n2826, gm_n47, gm_n81, in_16, gm_n2825, gm_n62);
	nand (gm_n2827, gm_n2826, gm_n71, gm_n45);
	and (gm_n2828, gm_n1704, gm_n52, in_9);
	nand (gm_n2829, gm_n49, in_12, in_11, gm_n2828, in_14);
	nor (gm_n2830, in_17, in_16, in_15, gm_n2829, in_18);
	nand (gm_n2831, in_21, in_20, in_19, gm_n2830);
	nand (gm_n2832, gm_n52, in_9, in_8, gm_n316, in_11);
	nor (gm_n2833, in_14, gm_n49, gm_n48, gm_n2832, gm_n63);
	nand (gm_n2834, gm_n47, in_17, gm_n46, gm_n2833, in_19);
	nor (gm_n2835, gm_n2834, in_21, in_20);
	nand (gm_n2836, gm_n55, in_6, in_5, gm_n519, gm_n64);
	or (gm_n2837, gm_n2836, in_9);
	nor (gm_n2838, in_12, gm_n53, gm_n52, gm_n2837, in_13);
	nand (gm_n2839, in_16, gm_n63, in_14, gm_n2838, gm_n81);
	nor (gm_n2840, in_20, in_19, gm_n47, gm_n2839, in_21);
	nand (gm_n2841, gm_n64, in_7, in_6, gm_n379, gm_n51);
	nor (gm_n2842, in_12, gm_n53, gm_n52, gm_n2841, in_13);
	nand (gm_n2843, in_16, in_15, in_14, gm_n2842, gm_n81);
	nor (gm_n2844, in_20, gm_n62, in_18, gm_n2843, in_21);
	or (gm_n2845, gm_n64, gm_n55, in_6, gm_n1429, in_9);
	nor (gm_n2846, gm_n48, in_11, gm_n52, gm_n2845, in_13);
	nand (gm_n2847, gm_n46, in_15, gm_n50, gm_n2846, gm_n81);
	nor (gm_n2848, in_20, in_19, in_18, gm_n2847, gm_n71);
	nand (gm_n2849, gm_n55, in_6, in_5, gm_n241, gm_n64);
	nor (gm_n2850, in_11, gm_n52, gm_n51, gm_n2849);
	nand (gm_n2851, gm_n50, in_13, in_12, gm_n2850, gm_n63);
	nor (gm_n2852, in_18, in_17, gm_n46, gm_n2851, in_19);
	nand (gm_n2853, gm_n2852, gm_n71, gm_n45);
	nand (gm_n2854, gm_n48, in_11, in_10, gm_n1332, gm_n49);
	nor (gm_n2855, gm_n46, gm_n63, in_14, gm_n2854, gm_n81);
	nand (gm_n2856, gm_n45, gm_n62, gm_n47, gm_n2855, in_21);
	nor (gm_n2857, in_11, gm_n52, in_9, gm_n285, gm_n48);
	nand (gm_n2858, in_15, gm_n50, in_13, gm_n2857, gm_n46);
	nor (gm_n2859, in_19, gm_n47, in_17, gm_n2858, in_20);
	nand (gm_n2860, gm_n2859, gm_n71);
	nand (gm_n2861, in_13, in_12, in_11, gm_n1538, gm_n50);
	nor (gm_n2862, gm_n81, in_16, in_15, gm_n2861, gm_n47);
	nand (gm_n2863, gm_n71, gm_n45, gm_n62, gm_n2862);
	or (gm_n2864, in_8, gm_n55, in_6, gm_n199, gm_n51);
	nor (gm_n2865, gm_n48, gm_n53, gm_n52, gm_n2864, gm_n49);
	nand (gm_n2866, gm_n46, gm_n63, in_14, gm_n2865, gm_n81);
	nor (gm_n2867, in_20, in_19, in_18, gm_n2866, gm_n71);
	nand (gm_n2868, in_10, in_9, in_8, gm_n838, gm_n53);
	nor (gm_n2869, in_14, in_13, gm_n48, gm_n2868);
	nand (gm_n2870, gm_n81, gm_n46, in_15, gm_n2869, in_18);
	nor (gm_n2871, in_21, in_20, in_19, gm_n2870);
	nand (gm_n2872, gm_n55, gm_n82, gm_n72, gm_n241, in_8);
	nor (gm_n2873, gm_n2872, in_9);
	and (gm_n2874, in_12, in_11, gm_n52, gm_n2873, gm_n49);
	nand (gm_n2875, gm_n46, in_15, gm_n50, gm_n2874, gm_n81);
	nor (gm_n2876, gm_n45, in_19, in_18, gm_n2875, in_21);
	and (gm_n2877, in_8, in_7, gm_n82, gm_n2640, gm_n51);
	and (gm_n2878, gm_n48, in_11, in_10, gm_n2877, gm_n49);
	nand (gm_n2879, in_16, in_15, gm_n50, gm_n2878, in_17);
	nor (gm_n2880, gm_n45, in_19, in_18, gm_n2879, in_21);
	nor (gm_n2881, in_11, gm_n52, in_9, gm_n2266);
	nand (gm_n2882, gm_n50, in_13, gm_n48, gm_n2881, gm_n63);
	nor (gm_n2883, gm_n47, gm_n81, in_16, gm_n2882, gm_n62);
	nand (gm_n2884, gm_n2883, gm_n71, in_20);
	nand (gm_n2885, gm_n55, in_6, gm_n72, gm_n1126, gm_n64);
	nor (gm_n2886, in_11, in_10, gm_n51, gm_n2885, gm_n48);
	nand (gm_n2887, gm_n63, gm_n50, in_13, gm_n2886, gm_n46);
	nor (gm_n2888, gm_n62, gm_n47, gm_n81, gm_n2887, in_20);
	nand (gm_n2889, gm_n2888, in_21);
	nor (gm_n2890, gm_n64, in_7, in_6, gm_n103, gm_n51);
	nand (gm_n2891, in_12, in_11, gm_n52, gm_n2890, gm_n49);
	nor (gm_n2892, in_16, in_15, in_14, gm_n2891, gm_n81);
	nand (gm_n2893, gm_n45, in_19, in_18, gm_n2892, gm_n71);
	nor (gm_n2894, in_11, gm_n52, gm_n51, gm_n1763, in_12);
	nand (gm_n2895, in_15, in_14, gm_n49, gm_n2894, gm_n46);
	nor (gm_n2896, gm_n62, in_18, in_17, gm_n2895, gm_n45);
	nand (gm_n2897, gm_n2896, gm_n71);
	or (gm_n2898, gm_n53, gm_n52, in_9, gm_n2564);
	nor (gm_n2899, in_14, gm_n49, gm_n48, gm_n2898, gm_n63);
	nand (gm_n2900, in_18, gm_n81, in_16, gm_n2899, in_19);
	nor (gm_n2901, gm_n2900, in_21, in_20);
	or (gm_n2902, in_7, gm_n82, gm_n72, gm_n75, in_8);
	nor (gm_n2903, gm_n53, gm_n52, gm_n51, gm_n2902, in_12);
	and (gm_n2904, in_15, gm_n50, gm_n49, gm_n2903, in_16);
	nand (gm_n2905, gm_n62, in_18, in_17, gm_n2904, in_20);
	nor (gm_n2906, gm_n2905, in_21);
	nor (gm_n2907, gm_n55, gm_n82, in_5, gm_n643, gm_n64);
	nand (gm_n2908, gm_n53, gm_n52, in_9, gm_n2907, gm_n48);
	nor (gm_n2909, gm_n63, in_14, gm_n49, gm_n2908, in_16);
	nand (gm_n2910, in_19, in_18, gm_n81, gm_n2909, gm_n45);
	nor (gm_n2911, gm_n2910, gm_n71);
	nand (gm_n2912, gm_n46, in_15, in_14, gm_n1336, in_17);
	nor (gm_n2913, in_20, gm_n62, in_18, gm_n2912, gm_n71);
	nand (gm_n2914, in_7, gm_n82, gm_n72, gm_n327, in_8);
	nor (gm_n2915, gm_n2914, gm_n51);
	nand (gm_n2916, gm_n48, in_11, in_10, gm_n2915, gm_n49);
	nor (gm_n2917, in_16, gm_n63, in_14, gm_n2916, in_17);
	nand (gm_n2918, gm_n45, gm_n62, in_18, gm_n2917, gm_n71);
	nand (gm_n2919, in_12, gm_n53, gm_n52, gm_n2915, gm_n49);
	nor (gm_n2920, in_16, gm_n63, in_14, gm_n2919, gm_n81);
	nand (gm_n2921, gm_n45, gm_n62, gm_n47, gm_n2920, in_21);
	nor (gm_n2922, in_9, gm_n64, gm_n55, gm_n1256);
	nand (gm_n2923, in_12, in_11, in_10, gm_n2922, gm_n49);
	nor (gm_n2924, in_16, gm_n63, in_14, gm_n2923, gm_n81);
	nand (gm_n2925, in_20, gm_n62, gm_n47, gm_n2924, gm_n71);
	nand (gm_n2926, gm_n55, in_6, gm_n72, gm_n89, in_8);
	nor (gm_n2927, in_11, gm_n52, gm_n51, gm_n2926, gm_n48);
	nand (gm_n2928, gm_n2927, gm_n49);
	nor (gm_n2929, in_16, gm_n63, gm_n50, gm_n2928, gm_n81);
	nand (gm_n2930, in_20, in_19, gm_n47, gm_n2929, gm_n71);
	nand (gm_n2931, in_8, in_7, in_6, gm_n374, in_9);
	nor (gm_n2932, gm_n48, gm_n53, gm_n52, gm_n2931, gm_n49);
	nand (gm_n2933, gm_n46, gm_n63, gm_n50, gm_n2932, in_17);
	nor (gm_n2934, in_20, gm_n62, in_18, gm_n2933, in_21);
	nand (gm_n2935, in_11, gm_n52, gm_n51, gm_n543);
	nor (gm_n2936, gm_n2935, gm_n49, gm_n48);
	nand (gm_n2937, gm_n46, gm_n63, in_14, gm_n2936, in_17);
	nor (gm_n2938, in_20, in_19, gm_n47, gm_n2937, gm_n71);
	nand (gm_n2939, in_11, gm_n52, gm_n51, gm_n1555, in_12);
	nor (gm_n2940, in_15, gm_n50, gm_n49, gm_n2939, gm_n46);
	nand (gm_n2941, in_19, gm_n47, gm_n81, gm_n2940, gm_n45);
	nor (gm_n2942, gm_n2941, in_21);
	or (gm_n2943, gm_n53, gm_n52, gm_n51, gm_n950, gm_n48);
	nor (gm_n2944, gm_n63, in_14, gm_n49, gm_n2943, in_16);
	nand (gm_n2945, in_19, gm_n47, gm_n81, gm_n2944, in_20);
	nor (gm_n2946, gm_n2945, gm_n71);
	and (gm_n2947, in_9, in_8, in_7, gm_n136, gm_n52);
	nand (gm_n2948, gm_n49, in_12, in_11, gm_n2947, gm_n50);
	nor (gm_n2949, gm_n81, in_16, in_15, gm_n2948, gm_n47);
	nand (gm_n2950, in_21, in_20, in_19, gm_n2949);
	nand (gm_n2951, in_7, gm_n82, gm_n72, gm_n519, in_8);
	nor (gm_n2952, in_11, in_10, gm_n51, gm_n2951, in_12);
	nand (gm_n2953, in_15, in_14, in_13, gm_n2952, in_16);
	nor (gm_n2954, gm_n62, gm_n47, in_17, gm_n2953, in_20);
	nand (gm_n2955, gm_n2954, gm_n71);
	nor (gm_n2956, gm_n64, gm_n55, gm_n82, gm_n530, gm_n51);
	nand (gm_n2957, gm_n48, gm_n53, in_10, gm_n2956, in_13);
	nor (gm_n2958, gm_n46, gm_n63, gm_n50, gm_n2957, gm_n81);
	nand (gm_n2959, in_20, gm_n62, gm_n47, gm_n2958, gm_n71);
	nor (gm_n2960, in_11, in_10, in_9, gm_n2564, gm_n48);
	nand (gm_n2961, in_15, in_14, gm_n49, gm_n2960, gm_n46);
	nor (gm_n2962, in_19, gm_n47, in_17, gm_n2961, in_20);
	nand (gm_n2963, gm_n2962, gm_n71);
	and (gm_n2964, gm_n49, in_12, in_11, gm_n1062, in_14);
	nand (gm_n2965, in_17, in_16, gm_n63, gm_n2964, in_18);
	nor (gm_n2966, gm_n71, gm_n45, gm_n62, gm_n2965);
	nor (gm_n2967, gm_n63, in_14, in_13, gm_n115, in_16);
	nand (gm_n2968, in_19, gm_n47, gm_n81, gm_n2967, in_20);
	nor (gm_n2969, gm_n2968, gm_n71);
	and (gm_n2970, in_10, in_9, in_8, gm_n2708, gm_n53);
	and (gm_n2971, in_14, in_13, in_12, gm_n2970);
	nand (gm_n2972, gm_n81, in_16, in_15, gm_n2971, in_18);
	nor (gm_n2973, in_21, in_20, in_19, gm_n2972);
	and (gm_n2974, gm_n48, gm_n53, gm_n52, gm_n1755, gm_n49);
	nand (gm_n2975, gm_n46, in_15, gm_n50, gm_n2974, in_17);
	nor (gm_n2976, in_20, gm_n62, in_18, gm_n2975, in_21);
	nor (gm_n2977, in_11, in_10, gm_n51, gm_n2445, gm_n48);
	nand (gm_n2978, in_15, in_14, gm_n49, gm_n2977, gm_n46);
	nor (gm_n2979, gm_n62, in_18, in_17, gm_n2978, in_20);
	nand (gm_n2980, gm_n2979, in_21);
	nand (gm_n2981, gm_n48, gm_n53, in_10, gm_n1385, gm_n49);
	nor (gm_n2982, gm_n46, gm_n63, gm_n50, gm_n2981, gm_n81);
	nand (gm_n2983, in_20, gm_n62, in_18, gm_n2982, gm_n71);
	and (gm_n2984, gm_n64, in_7, in_6, gm_n374, gm_n51);
	nand (gm_n2985, in_12, in_11, gm_n52, gm_n2984, in_13);
	nor (gm_n2986, in_16, in_15, in_14, gm_n2985, in_17);
	nand (gm_n2987, in_20, in_19, in_18, gm_n2986, in_21);
	nand (gm_n2988, in_12, gm_n53, in_10, gm_n1975, in_13);
	nor (gm_n2989, gm_n46, in_15, in_14, gm_n2988, in_17);
	nand (gm_n2990, gm_n45, gm_n62, in_18, gm_n2989, gm_n71);
	and (gm_n2991, in_12, in_11, in_10, gm_n1840, in_13);
	nand (gm_n2992, gm_n46, gm_n63, gm_n50, gm_n2991, in_17);
	nor (gm_n2993, in_20, in_19, in_18, gm_n2992, in_21);
	nand (gm_n2994, in_11, gm_n52, gm_n51, gm_n1459, in_12);
	nor (gm_n2995, gm_n63, gm_n50, gm_n49, gm_n2994, in_16);
	nand (gm_n2996, in_19, in_18, gm_n81, gm_n2995, gm_n45);
	nor (gm_n2997, gm_n2996, in_21);
	nand (gm_n2998, gm_n52, in_9, gm_n64, gm_n2708, in_11);
	nor (gm_n2999, in_14, in_13, in_12, gm_n2998, gm_n63);
	nand (gm_n3000, in_18, gm_n81, in_16, gm_n2999, gm_n62);
	nor (gm_n3001, gm_n3000, in_21, gm_n45);
	nand (gm_n3002, gm_n52, gm_n51, gm_n64, gm_n57, in_11);
	nor (gm_n3003, gm_n50, gm_n49, in_12, gm_n3002, gm_n63);
	nand (gm_n3004, gm_n47, in_17, in_16, gm_n3003, gm_n62);
	nor (gm_n3005, gm_n3004, in_21, gm_n45);
	nand (gm_n3006, in_13, in_12, gm_n53, gm_n1099, in_14);
	nor (gm_n3007, in_17, in_16, in_15, gm_n3006, in_18);
	nand (gm_n3008, in_21, gm_n45, in_19, gm_n3007);
	nand (gm_n3009, gm_n48, in_11, gm_n52, gm_n747, in_13);
	nor (gm_n3010, gm_n46, in_15, gm_n50, gm_n3009, gm_n81);
	nand (gm_n3011, gm_n45, gm_n62, gm_n47, gm_n3010, in_21);
	nand (gm_n3012, gm_n1572, gm_n51);
	or (gm_n3013, in_12, gm_n53, in_10, gm_n3012, gm_n49);
	nor (gm_n3014, gm_n46, in_15, gm_n50, gm_n3013, in_17);
	nand (gm_n3015, gm_n45, in_19, gm_n47, gm_n3014, gm_n71);
	nand (gm_n3016, gm_n48, in_11, gm_n52, gm_n2922, in_13);
	nor (gm_n3017, in_16, gm_n63, gm_n50, gm_n3016, gm_n81);
	nand (gm_n3018, in_20, gm_n62, gm_n47, gm_n3017, gm_n71);
	nor (gm_n3019, in_14, gm_n49, gm_n48, gm_n1875, gm_n63);
	nand (gm_n3020, gm_n47, in_17, in_16, gm_n3019, in_19);
	nor (gm_n3021, gm_n3020, gm_n71, gm_n45);
	or (gm_n3022, in_9, in_8, gm_n55, gm_n525, gm_n52);
	nor (gm_n3023, in_13, in_12, gm_n53, gm_n3022, in_14);
	nand (gm_n3024, in_17, in_16, gm_n63, gm_n3023, in_18);
	nor (gm_n3025, gm_n71, in_20, in_19, gm_n3024);
	nand (gm_n3026, in_16, gm_n63, gm_n50, gm_n789, in_17);
	nor (gm_n3027, in_20, gm_n62, gm_n47, gm_n3026, in_21);
	nor (gm_n3028, gm_n48, in_11, gm_n52, gm_n2280, in_13);
	nand (gm_n3029, gm_n46, gm_n63, gm_n50, gm_n3028, gm_n81);
	nor (gm_n3030, in_20, in_19, gm_n47, gm_n3029, gm_n71);
	nand (gm_n3031, gm_n53, in_10, gm_n51, gm_n868, gm_n48);
	nor (gm_n3032, gm_n3031, in_13);
	and (gm_n3033, gm_n46, in_15, in_14, gm_n3032, gm_n81);
	nand (gm_n3034, in_20, in_19, gm_n47, gm_n3033, in_21);
	and (gm_n3035, gm_n168, in_10, gm_n51);
	nand (gm_n3036, gm_n49, in_12, in_11, gm_n3035, gm_n50);
	nor (gm_n3037, gm_n81, gm_n46, in_15, gm_n3036, in_18);
	nand (gm_n3038, in_21, in_20, gm_n62, gm_n3037);
	and (gm_n3039, in_8, gm_n55, gm_n82, gm_n2640, in_9);
	and (gm_n3040, in_12, gm_n53, in_10, gm_n3039, gm_n49);
	and (gm_n3041, in_16, gm_n63, gm_n50, gm_n3040, gm_n81);
	nand (gm_n3042, in_20, gm_n62, gm_n47, gm_n3041, in_21);
	nor (gm_n3043, gm_n55, in_6, gm_n72, gm_n321, gm_n64);
	and (gm_n3044, in_11, gm_n52, gm_n51, gm_n3043);
	nand (gm_n3045, gm_n3044, in_13, in_12);
	nor (gm_n3046, in_16, gm_n63, gm_n50, gm_n3045, gm_n81);
	nand (gm_n3047, in_20, in_19, in_18, gm_n3046, in_21);
	nor (gm_n3048, gm_n53, in_10, in_9, gm_n1879);
	and (gm_n3049, in_14, in_13, in_12, gm_n3048, in_15);
	nand (gm_n3050, in_18, gm_n81, in_16, gm_n3049, gm_n62);
	nor (gm_n3051, gm_n3050, in_21, in_20);
	nand (gm_n3052, gm_n53, gm_n52, gm_n51, gm_n291, in_12);
	nor (gm_n3053, in_15, in_14, in_13, gm_n3052, gm_n46);
	nand (gm_n3054, gm_n62, gm_n47, in_17, gm_n3053, in_20);
	nor (gm_n3055, gm_n3054, gm_n71);
	nand (gm_n3056, in_9, gm_n64, gm_n55, gm_n1007, in_10);
	nor (gm_n3057, in_13, gm_n48, in_11, gm_n3056, gm_n50);
	nand (gm_n3058, gm_n81, in_16, gm_n63, gm_n3057, gm_n47);
	nor (gm_n3059, gm_n71, in_20, gm_n62, gm_n3058);
	and (gm_n3060, gm_n1088, in_9, in_8);
	and (gm_n3061, in_12, gm_n53, in_10, gm_n3060, gm_n49);
	nand (gm_n3062, in_16, in_15, gm_n50, gm_n3061, gm_n81);
	nor (gm_n3063, gm_n45, in_19, in_18, gm_n3062, in_21);
	nor (gm_n3064, gm_n55, in_6, in_5, gm_n290, gm_n64);
	and (gm_n3065, gm_n53, in_10, gm_n51, gm_n3064);
	nand (gm_n3066, gm_n50, gm_n49, in_12, gm_n3065, in_15);
	nor (gm_n3067, in_18, gm_n81, gm_n46, gm_n3066, in_19);
	nand (gm_n3068, gm_n3067, gm_n71, in_20);
	nor (gm_n3069, gm_n64, gm_n55, gm_n82, gm_n161, gm_n51);
	nand (gm_n3070, in_12, in_11, gm_n52, gm_n3069, gm_n49);
	nor (gm_n3071, in_16, gm_n63, gm_n50, gm_n3070, in_17);
	nand (gm_n3072, gm_n45, in_19, in_18, gm_n3071, in_21);
	and (gm_n3073, in_11, gm_n52, in_9, gm_n2229, gm_n48);
	nand (gm_n3074, gm_n3073, gm_n50, gm_n49);
	nor (gm_n3075, in_17, in_16, gm_n63, gm_n3074, in_18);
	nand (gm_n3076, gm_n71, in_20, gm_n62, gm_n3075);
	nand (gm_n3077, in_6, gm_n72, gm_n54, gm_n389, gm_n55);
	nor (gm_n3078, gm_n52, in_9, gm_n64, gm_n3077, in_11);
	nand (gm_n3079, gm_n50, gm_n49, gm_n48, gm_n3078, gm_n63);
	nor (gm_n3080, in_18, gm_n81, gm_n46, gm_n3079, in_19);
	nand (gm_n3081, gm_n3080, in_21, gm_n45);
	nor (gm_n3082, gm_n440, gm_n52, gm_n51);
	and (gm_n3083, in_13, gm_n48, gm_n53, gm_n3082, in_14);
	nand (gm_n3084, in_17, gm_n46, in_15, gm_n3083, in_18);
	nor (gm_n3085, in_21, gm_n45, gm_n62, gm_n3084);
	nor (gm_n3086, in_7, in_6, gm_n72, gm_n643, in_8);
	nand (gm_n3087, gm_n53, in_10, in_9, gm_n3086);
	nor (gm_n3088, in_14, gm_n49, gm_n48, gm_n3087, gm_n63);
	nand (gm_n3089, in_18, gm_n81, in_16, gm_n3088, in_19);
	nor (gm_n3090, gm_n3089, gm_n71, gm_n45);
	and (gm_n3091, gm_n55, gm_n82, gm_n72, gm_n420, in_8);
	nand (gm_n3092, in_11, gm_n52, gm_n51, gm_n3091);
	nor (gm_n3093, gm_n50, in_13, in_12, gm_n3092, in_15);
	nand (gm_n3094, gm_n47, in_17, in_16, gm_n3093, in_19);
	nor (gm_n3095, gm_n3094, gm_n71, in_20);
	nand (gm_n3096, gm_n53, in_10, gm_n51, gm_n700, gm_n48);
	nor (gm_n3097, gm_n3096, in_13);
	nand (gm_n3098, gm_n46, gm_n63, gm_n50, gm_n3097, in_17);
	nor (gm_n3099, in_20, in_19, in_18, gm_n3098, gm_n71);
	nand (gm_n3100, gm_n48, gm_n53, in_10, gm_n3039, in_13);
	nor (gm_n3101, in_16, in_15, gm_n50, gm_n3100, gm_n81);
	nand (gm_n3102, gm_n45, gm_n62, in_18, gm_n3101, gm_n71);
	nor (gm_n3103, in_11, gm_n52, gm_n51, gm_n2445, gm_n48);
	nand (gm_n3104, gm_n63, gm_n50, gm_n49, gm_n3103, in_16);
	nor (gm_n3105, in_19, in_18, in_17, gm_n3104, in_20);
	nand (gm_n3106, gm_n3105, in_21);
	nand (gm_n3107, in_12, gm_n53, in_10, gm_n2749, in_13);
	nor (gm_n3108, in_16, in_15, in_14, gm_n3107, gm_n81);
	nand (gm_n3109, in_20, in_19, in_18, gm_n3108, gm_n71);
	nand (gm_n3110, gm_n53, gm_n52, gm_n51, gm_n543, in_12);
	nor (gm_n3111, gm_n3110, in_13);
	and (gm_n3112, gm_n46, gm_n63, in_14, gm_n3111, gm_n81);
	nand (gm_n3113, in_20, gm_n62, gm_n47, gm_n3112, in_21);
	nand (gm_n3114, in_11, gm_n52, gm_n51, gm_n3086, gm_n48);
	or (gm_n3115, gm_n63, in_14, in_13, gm_n3114, gm_n46);
	or (gm_n3116, in_19, in_18, gm_n81, gm_n3115, in_20);
	nor (gm_n3117, gm_n3116, gm_n71);
	nand (gm_n3118, gm_n53, in_10, gm_n51, gm_n3043, in_12);
	nor (gm_n3119, in_15, gm_n50, gm_n49, gm_n3118, gm_n46);
	nand (gm_n3120, in_19, gm_n47, gm_n81, gm_n3119, in_20);
	nor (gm_n3121, gm_n3120, gm_n71);
	nor (gm_n3122, in_15, gm_n50, gm_n49, gm_n2010, gm_n46);
	nand (gm_n3123, in_19, in_18, in_17, gm_n3122, in_20);
	nor (gm_n3124, gm_n3123, in_21);
	and (gm_n3125, in_12, gm_n53, in_10, gm_n2001, in_13);
	nand (gm_n3126, gm_n46, in_15, gm_n50, gm_n3125, gm_n81);
	nor (gm_n3127, in_20, gm_n62, in_18, gm_n3126, gm_n71);
	nor (gm_n3128, gm_n52, gm_n51, gm_n64, gm_n390, in_11);
	nand (gm_n3129, gm_n50, gm_n49, gm_n48, gm_n3128, gm_n63);
	nor (gm_n3130, gm_n47, in_17, gm_n46, gm_n3129, gm_n62);
	nand (gm_n3131, gm_n3130, in_21, gm_n45);
	nand (gm_n3132, gm_n48, in_11, in_10, gm_n2922, in_13);
	nor (gm_n3133, gm_n46, gm_n63, gm_n50, gm_n3132, gm_n81);
	nand (gm_n3134, gm_n45, gm_n62, gm_n47, gm_n3133, in_21);
	nor (gm_n3135, in_11, gm_n52, in_9, gm_n873, in_12);
	nand (gm_n3136, gm_n63, in_14, in_13, gm_n3135);
	nor (gm_n3137, in_18, gm_n81, in_16, gm_n3136, gm_n62);
	nand (gm_n3138, gm_n3137, in_21, in_20);
	nor (gm_n3139, gm_n53, in_10, gm_n51, gm_n1247, in_12);
	nand (gm_n3140, in_15, gm_n50, gm_n49, gm_n3139, gm_n46);
	nor (gm_n3141, in_19, in_18, gm_n81, gm_n3140, gm_n45);
	nand (gm_n3142, gm_n3141, gm_n71);
	nor (gm_n3143, gm_n50, gm_n49, gm_n48, gm_n2292, in_15);
	nand (gm_n3144, gm_n47, gm_n81, in_16, gm_n3143, gm_n62);
	nor (gm_n3145, gm_n3144, gm_n71, in_20);
	or (gm_n3146, gm_n55, gm_n82, gm_n72, gm_n167, in_8);
	nor (gm_n3147, in_11, in_10, gm_n51, gm_n3146, in_12);
	and (gm_n3148, in_15, in_14, in_13, gm_n3147);
	nand (gm_n3149, in_18, gm_n81, in_16, gm_n3148, in_19);
	nor (gm_n3150, gm_n3149, gm_n71, gm_n45);
	nand (gm_n3151, gm_n53, in_10, in_9, gm_n2088, in_12);
	nor (gm_n3152, gm_n3151, in_13);
	nand (gm_n3153, gm_n46, gm_n63, gm_n50, gm_n3152, gm_n81);
	nor (gm_n3154, gm_n45, in_19, in_18, gm_n3153, in_21);
	nand (gm_n3155, gm_n53, in_10, in_9, gm_n566, gm_n48);
	nor (gm_n3156, gm_n63, gm_n50, in_13, gm_n3155, gm_n46);
	nand (gm_n3157, gm_n62, in_18, in_17, gm_n3156, in_20);
	nor (gm_n3158, gm_n3157, in_21);
	or (gm_n3159, in_8, gm_n55, in_6, gm_n119, gm_n51);
	or (gm_n3160, gm_n48, in_11, gm_n52, gm_n3159, in_13);
	nor (gm_n3161, gm_n46, in_15, in_14, gm_n3160, in_17);
	nand (gm_n3162, in_20, in_19, gm_n47, gm_n3161, in_21);
	nor (gm_n3163, in_8, gm_n55, gm_n82, gm_n96, gm_n51);
	nand (gm_n3164, gm_n48, gm_n53, in_10, gm_n3163, gm_n49);
	nor (gm_n3165, gm_n46, gm_n63, in_14, gm_n3164, gm_n81);
	nand (gm_n3166, in_20, in_19, gm_n47, gm_n3165, gm_n71);
	nand (gm_n3167, gm_n48, in_11, gm_n52, gm_n972, gm_n49);
	nor (gm_n3168, in_16, gm_n63, gm_n50, gm_n3167, gm_n81);
	nand (gm_n3169, gm_n45, in_19, in_18, gm_n3168, in_21);
	and (gm_n3170, in_10, gm_n51, gm_n64, gm_n57);
	nand (gm_n3171, in_13, in_12, in_11, gm_n3170, gm_n50);
	nor (gm_n3172, gm_n81, in_16, gm_n63, gm_n3171, gm_n47);
	nand (gm_n3173, in_21, gm_n45, in_19, gm_n3172);
	or (gm_n3174, in_6, gm_n72, gm_n54, gm_n56, gm_n55);
	or (gm_n3175, gm_n52, gm_n51, gm_n64, gm_n3174, in_11);
	nor (gm_n3176, in_14, in_13, in_12, gm_n3175, gm_n63);
	nand (gm_n3177, in_18, gm_n81, gm_n46, gm_n3176, in_19);
	nor (gm_n3178, gm_n3177, in_21, gm_n45);
	and (gm_n3179, gm_n53, in_10, in_9, gm_n1360, gm_n48);
	and (gm_n3180, in_15, in_14, in_13, gm_n3179, in_16);
	nand (gm_n3181, gm_n62, in_18, in_17, gm_n3180, gm_n45);
	nor (gm_n3182, gm_n3181, in_21);
	nor (gm_n3183, in_7, in_6, gm_n72, gm_n188, in_8);
	nand (gm_n3184, gm_n3183, in_10, gm_n51);
	nor (gm_n3185, gm_n49, in_12, gm_n53, gm_n3184);
	nand (gm_n3186, gm_n46, in_15, gm_n50, gm_n3185, gm_n81);
	nor (gm_n3187, in_20, in_19, gm_n47, gm_n3186, gm_n71);
	or (gm_n3188, gm_n64, in_7, gm_n82, gm_n199, in_9);
	nor (gm_n3189, gm_n3188, gm_n52);
	and (gm_n3190, gm_n49, gm_n48, gm_n53, gm_n3189, gm_n50);
	nand (gm_n3191, gm_n81, gm_n46, in_15, gm_n3190, gm_n47);
	nor (gm_n3192, gm_n71, gm_n45, in_19, gm_n3191);
	nor (gm_n3193, gm_n55, in_6, gm_n72, gm_n75, in_8);
	and (gm_n3194, gm_n53, gm_n52, in_9, gm_n3193);
	nand (gm_n3195, gm_n50, gm_n49, gm_n48, gm_n3194, gm_n63);
	nor (gm_n3196, in_18, gm_n81, in_16, gm_n3195, gm_n62);
	nand (gm_n3197, gm_n3196, gm_n71, in_20);
	or (gm_n3198, gm_n55, in_6, gm_n72, gm_n167, gm_n64);
	nor (gm_n3199, in_11, in_10, gm_n51, gm_n3198, gm_n48);
	nand (gm_n3200, in_15, gm_n50, gm_n49, gm_n3199, in_16);
	nor (gm_n3201, in_19, gm_n47, gm_n81, gm_n3200, in_20);
	nand (gm_n3202, gm_n3201, in_21);
	nand (gm_n3203, in_12, gm_n53, in_10, gm_n2097, in_13);
	nor (gm_n3204, gm_n46, in_15, in_14, gm_n3203, gm_n81);
	nand (gm_n3205, in_20, in_19, gm_n47, gm_n3204, in_21);
	and (gm_n3206, gm_n53, gm_n52, in_9, gm_n1469, gm_n48);
	nand (gm_n3207, in_15, gm_n50, gm_n49, gm_n3206, gm_n46);
	nor (gm_n3208, in_19, gm_n47, gm_n81, gm_n3207, in_20);
	nand (gm_n3209, gm_n3208, in_21);
	and (gm_n3210, in_10, in_9, in_8, gm_n431, in_11);
	and (gm_n3211, in_14, in_13, gm_n48, gm_n3210, in_15);
	nand (gm_n3212, in_18, in_17, in_16, gm_n3211, gm_n62);
	nor (gm_n3213, gm_n3212, in_21, gm_n45);
	and (gm_n3214, in_7, gm_n82, in_5, gm_n209, gm_n64);
	nand (gm_n3215, gm_n53, in_10, in_9, gm_n3214, in_12);
	nor (gm_n3216, gm_n63, in_14, gm_n49, gm_n3215, in_16);
	nand (gm_n3217, gm_n62, gm_n47, gm_n81, gm_n3216, gm_n45);
	nor (gm_n3218, gm_n3217, in_21);
	or (gm_n3219, in_11, in_10, in_9, gm_n2397, gm_n48);
	nor (gm_n3220, gm_n63, gm_n50, in_13, gm_n3219, gm_n46);
	nand (gm_n3221, gm_n62, in_18, in_17, gm_n3220, gm_n45);
	nor (gm_n3222, gm_n3221, in_21);
	nor (gm_n3223, gm_n48, in_11, in_10, gm_n2845, in_13);
	nand (gm_n3224, gm_n46, in_15, in_14, gm_n3223, gm_n81);
	nor (gm_n3225, in_20, in_19, gm_n47, gm_n3224, gm_n71);
	nor (gm_n3226, gm_n51, in_8, in_7, gm_n553, gm_n52);
	nand (gm_n3227, gm_n49, in_12, gm_n53, gm_n3226, gm_n50);
	nor (gm_n3228, in_17, gm_n46, gm_n63, gm_n3227, gm_n47);
	nand (gm_n3229, gm_n71, in_20, in_19, gm_n3228);
	nand (gm_n3230, in_12, gm_n53, in_10, gm_n375, gm_n49);
	nor (gm_n3231, in_16, in_15, gm_n50, gm_n3230, gm_n81);
	nand (gm_n3232, gm_n45, in_19, in_18, gm_n3231, in_21);
	or (gm_n3233, gm_n50, in_13, in_12, gm_n770, in_15);
	nor (gm_n3234, gm_n47, in_17, gm_n46, gm_n3233, gm_n62);
	nand (gm_n3235, gm_n3234, gm_n71, gm_n45);
	nand (gm_n3236, gm_n48, in_11, gm_n52, gm_n2641, in_13);
	nor (gm_n3237, in_16, gm_n63, gm_n50, gm_n3236, gm_n81);
	nand (gm_n3238, in_20, gm_n62, gm_n47, gm_n3237, in_21);
	and (gm_n3239, gm_n51, gm_n64, gm_n55, gm_n151);
	and (gm_n3240, gm_n48, gm_n53, in_10, gm_n3239, gm_n49);
	nand (gm_n3241, gm_n46, gm_n63, gm_n50, gm_n3240, in_17);
	nor (gm_n3242, gm_n45, gm_n62, in_18, gm_n3241, in_21);
	nand (gm_n3243, in_17, in_16, gm_n63, gm_n2548, gm_n47);
	nor (gm_n3244, in_21, in_20, in_19, gm_n3243);
	nand (gm_n3245, in_8, in_7, gm_n82, gm_n638, in_9);
	nor (gm_n3246, in_12, in_11, gm_n52, gm_n3245, gm_n49);
	nand (gm_n3247, in_16, gm_n63, in_14, gm_n3246, in_17);
	nor (gm_n3248, gm_n45, in_19, in_18, gm_n3247, in_21);
	nand (gm_n3249, in_8, gm_n55, gm_n82, gm_n1075, in_9);
	nor (gm_n3250, gm_n48, in_11, gm_n52, gm_n3249, in_13);
	nand (gm_n3251, gm_n46, in_15, in_14, gm_n3250, in_17);
	nor (gm_n3252, gm_n45, gm_n62, in_18, gm_n3251, gm_n71);
	nor (gm_n3253, gm_n51, in_8, in_7, gm_n525, in_10);
	nand (gm_n3254, in_13, gm_n48, in_11, gm_n3253, gm_n50);
	nor (gm_n3255, gm_n81, gm_n46, in_15, gm_n3254, gm_n47);
	nand (gm_n3256, gm_n71, gm_n45, gm_n62, gm_n3255);
	nand (gm_n3257, in_7, in_6, gm_n72, gm_n519, gm_n64);
	nor (gm_n3258, gm_n53, gm_n52, in_9, gm_n3257, gm_n48);
	nand (gm_n3259, in_15, gm_n50, in_13, gm_n3258, in_16);
	nor (gm_n3260, in_19, in_18, in_17, gm_n3259, gm_n45);
	nand (gm_n3261, gm_n3260, in_21);
	and (gm_n3262, gm_n51, gm_n64, gm_n55, gm_n404, gm_n52);
	and (gm_n3263, in_13, gm_n48, gm_n53, gm_n3262, gm_n50);
	and (gm_n3264, in_17, gm_n46, in_15, gm_n3263, gm_n47);
	nand (gm_n3265, in_21, in_20, gm_n62, gm_n3264);
	and (gm_n3266, in_16, gm_n63, gm_n50, gm_n935, gm_n81);
	nand (gm_n3267, in_20, gm_n62, gm_n47, gm_n3266, gm_n71);
	and (gm_n3268, gm_n64, gm_n55, in_6, gm_n2640, in_9);
	and (gm_n3269, gm_n48, in_11, in_10, gm_n3268, in_13);
	nand (gm_n3270, in_16, gm_n63, gm_n50, gm_n3269, gm_n81);
	nor (gm_n3271, in_20, in_19, gm_n47, gm_n3270, in_21);
	and (gm_n3272, in_11, gm_n52, in_9, gm_n3064, gm_n48);
	and (gm_n3273, gm_n63, in_14, gm_n49, gm_n3272, in_16);
	nand (gm_n3274, gm_n62, in_18, in_17, gm_n3273, gm_n45);
	nor (gm_n3275, gm_n3274, in_21);
	and (gm_n3276, gm_n53, gm_n52, gm_n51, gm_n1212);
	and (gm_n3277, in_14, gm_n49, gm_n48, gm_n3276, gm_n63);
	nand (gm_n3278, gm_n47, gm_n81, in_16, gm_n3277, in_19);
	nor (gm_n3279, gm_n3278, in_21, gm_n45);
	and (gm_n3280, in_12, in_11, in_10, gm_n1365, gm_n49);
	nand (gm_n3281, gm_n46, gm_n63, in_14, gm_n3280, in_17);
	nor (gm_n3282, gm_n45, gm_n62, in_18, gm_n3281, gm_n71);
	nor (gm_n3283, gm_n52, in_9, in_8, gm_n907, in_11);
	nand (gm_n3284, gm_n50, in_13, gm_n48, gm_n3283, gm_n63);
	nor (gm_n3285, gm_n47, in_17, gm_n46, gm_n3284, in_19);
	nand (gm_n3286, gm_n3285, gm_n71, gm_n45);
	nor (gm_n3287, in_8, gm_n55, in_6, gm_n141, gm_n51);
	nand (gm_n3288, gm_n48, in_11, gm_n52, gm_n3287, in_13);
	nor (gm_n3289, gm_n46, gm_n63, gm_n50, gm_n3288, in_17);
	nand (gm_n3290, gm_n45, gm_n62, in_18, gm_n3289, gm_n71);
	nor (gm_n3291, in_9, in_8, gm_n55, gm_n223, in_10);
	nand (gm_n3292, in_13, gm_n48, in_11, gm_n3291, gm_n50);
	nor (gm_n3293, gm_n81, in_16, gm_n63, gm_n3292, in_18);
	nand (gm_n3294, gm_n71, gm_n45, in_19, gm_n3293);
	nor (gm_n3295, in_11, gm_n52, in_9, gm_n2397);
	nand (gm_n3296, gm_n50, in_13, gm_n48, gm_n3295, in_15);
	nor (gm_n3297, gm_n47, gm_n81, in_16, gm_n3296, gm_n62);
	nand (gm_n3298, gm_n3297, gm_n71, gm_n45);
	nor (gm_n3299, in_7, gm_n82, in_5, gm_n188, in_8);
	nand (gm_n3300, gm_n3299, in_10, gm_n51);
	nor (gm_n3301, in_13, gm_n48, gm_n53, gm_n3300, in_14);
	nand (gm_n3302, gm_n81, gm_n46, gm_n63, gm_n3301, gm_n47);
	nor (gm_n3303, in_21, gm_n45, gm_n62, gm_n3302);
	or (gm_n3304, in_17, in_16, in_15, gm_n1471, in_18);
	nor (gm_n3305, in_21, gm_n45, in_19, gm_n3304);
	nor (gm_n3306, in_13, in_12, gm_n53, gm_n2514, in_14);
	nand (gm_n3307, gm_n81, in_16, in_15, gm_n3306, gm_n47);
	nor (gm_n3308, gm_n71, in_20, gm_n62, gm_n3307);
	and (gm_n3309, gm_n64, in_7, gm_n82, gm_n638, gm_n51);
	and (gm_n3310, in_12, gm_n53, in_10, gm_n3309, in_13);
	nand (gm_n3311, gm_n46, in_15, gm_n50, gm_n3310, in_17);
	nor (gm_n3312, gm_n45, gm_n62, gm_n47, gm_n3311, in_21);
	nand (gm_n3313, in_12, gm_n53, gm_n52, gm_n2890, gm_n49);
	nor (gm_n3314, in_16, gm_n63, gm_n50, gm_n3313, in_17);
	nand (gm_n3315, gm_n45, in_19, in_18, gm_n3314, gm_n71);
	and (gm_n3316, gm_n53, gm_n52, in_9, gm_n1315);
	nand (gm_n3317, gm_n50, in_13, in_12, gm_n3316, gm_n63);
	nor (gm_n3318, in_18, in_17, in_16, gm_n3317, gm_n62);
	nand (gm_n3319, gm_n3318, in_21, in_20);
	nor (gm_n3320, gm_n2823, gm_n52, in_9);
	nand (gm_n3321, in_13, in_12, in_11, gm_n3320, gm_n50);
	nor (gm_n3322, gm_n81, gm_n46, in_15, gm_n3321, in_18);
	nand (gm_n3323, gm_n71, in_20, in_19, gm_n3322);
	and (gm_n3324, gm_n1284, gm_n51);
	nand (gm_n3325, in_12, gm_n53, in_10, gm_n3324, gm_n49);
	nor (gm_n3326, in_16, in_15, gm_n50, gm_n3325, in_17);
	nand (gm_n3327, in_20, in_19, in_18, gm_n3326, in_21);
	nand (gm_n3328, gm_n53, in_10, gm_n51, gm_n1302);
	nor (gm_n3329, in_14, in_13, in_12, gm_n3328, in_15);
	nand (gm_n3330, in_18, in_17, gm_n46, gm_n3329, in_19);
	nor (gm_n3331, gm_n3330, in_21, gm_n45);
	or (gm_n3332, gm_n1239, gm_n52, in_9);
	nor (gm_n3333, gm_n49, gm_n48, gm_n53, gm_n3332, gm_n50);
	nand (gm_n3334, in_17, gm_n46, gm_n63, gm_n3333, in_18);
	nor (gm_n3335, in_21, in_20, in_19, gm_n3334);
	nand (gm_n3336, in_11, gm_n52, gm_n51, gm_n1469, in_12);
	nor (gm_n3337, in_15, gm_n50, gm_n49, gm_n3336, in_16);
	nand (gm_n3338, in_19, gm_n47, gm_n81, gm_n3337, in_20);
	nor (gm_n3339, gm_n3338, gm_n71);
	nand (gm_n3340, gm_n55, in_6, gm_n72, gm_n252, in_8);
	or (gm_n3341, gm_n53, in_10, in_9, gm_n3340);
	nor (gm_n3342, gm_n50, gm_n49, in_12, gm_n3341, gm_n63);
	nand (gm_n3343, in_18, in_17, in_16, gm_n3342, gm_n62);
	nor (gm_n3344, gm_n3343, gm_n71, gm_n45);
	nand (gm_n3345, gm_n48, gm_n53, gm_n52, gm_n1671, gm_n49);
	nor (gm_n3346, in_16, in_15, gm_n50, gm_n3345, in_17);
	nand (gm_n3347, in_20, in_19, gm_n47, gm_n3346, in_21);
	nor (gm_n3348, in_17, gm_n46, gm_n63, gm_n994, in_18);
	nand (gm_n3349, in_21, in_20, in_19, gm_n3348);
	nor (gm_n3350, gm_n51, in_8, in_7, gm_n279, in_10);
	nand (gm_n3351, in_13, gm_n48, gm_n53, gm_n3350, gm_n50);
	nor (gm_n3352, in_17, gm_n46, in_15, gm_n3351, in_18);
	nand (gm_n3353, gm_n71, in_20, in_19, gm_n3352);
	nor (gm_n3354, in_8, gm_n55, in_6, gm_n96, gm_n51);
	nand (gm_n3355, in_12, in_11, in_10, gm_n3354, in_13);
	nor (gm_n3356, in_16, in_15, gm_n50, gm_n3355, in_17);
	nand (gm_n3357, gm_n45, in_19, in_18, gm_n3356, in_21);
	or (gm_n3358, gm_n46, gm_n63, in_14, gm_n2919, gm_n81);
	nor (gm_n3359, in_20, gm_n62, in_18, gm_n3358, in_21);
	or (gm_n3360, in_9, gm_n64, in_7, gm_n843, in_10);
	nor (gm_n3361, gm_n49, in_12, gm_n53, gm_n3360, gm_n50);
	nand (gm_n3362, in_17, in_16, in_15, gm_n3361, in_18);
	nor (gm_n3363, gm_n71, in_20, in_19, gm_n3362);
	or (gm_n3364, gm_n46, gm_n63, gm_n50, gm_n2406, gm_n81);
	nor (gm_n3365, gm_n45, in_19, in_18, gm_n3364, in_21);
	nor (gm_n3366, gm_n50, in_13, in_12, gm_n3087, in_15);
	nand (gm_n3367, in_18, gm_n81, in_16, gm_n3366, in_19);
	nor (gm_n3368, gm_n3367, in_21, gm_n45);
	nand (gm_n3369, in_12, in_11, gm_n52, gm_n2284, gm_n49);
	nor (gm_n3370, gm_n46, gm_n63, gm_n50, gm_n3369, in_17);
	nand (gm_n3371, gm_n45, gm_n62, in_18, gm_n3370, in_21);
	nand (gm_n3372, gm_n48, gm_n53, gm_n52, gm_n980, gm_n49);
	nor (gm_n3373, gm_n46, in_15, in_14, gm_n3372, in_17);
	nand (gm_n3374, gm_n45, in_19, in_18, gm_n3373, gm_n71);
	nand (gm_n3375, gm_n3374, gm_n3371);
	nor (gm_n3376, gm_n3365, gm_n3363, gm_n3359, gm_n3375, gm_n3368);
	nand (gm_n3377, gm_n3353, gm_n3349, gm_n3347, gm_n3376, gm_n3357);
	nor (gm_n3378, gm_n3339, gm_n3335, gm_n3331, gm_n3377, gm_n3344);
	nand (gm_n3379, gm_n3323, gm_n3319, gm_n3315, gm_n3378, gm_n3327);
	nor (gm_n3380, gm_n3308, gm_n3305, gm_n3303, gm_n3379, gm_n3312);
	nand (gm_n3381, gm_n3294, gm_n3290, gm_n3286, gm_n3380, gm_n3298);
	nor (gm_n3382, gm_n3279, gm_n3275, gm_n3271, gm_n3381, gm_n3282);
	nand (gm_n3383, gm_n3265, gm_n3261, gm_n3256, gm_n3382, gm_n3267);
	nor (gm_n3384, gm_n3248, gm_n3244, gm_n3242, gm_n3383, gm_n3252);
	nand (gm_n3385, gm_n3235, gm_n3232, gm_n3229, gm_n3384, gm_n3238);
	nor (gm_n3386, gm_n3222, gm_n3218, gm_n3213, gm_n3385, gm_n3225);
	nand (gm_n3387, gm_n3205, gm_n3202, gm_n3197, gm_n3386, gm_n3209);
	nor (gm_n3388, gm_n3187, gm_n3182, gm_n3178, gm_n3387, gm_n3192);
	nand (gm_n3389, gm_n3169, gm_n3166, gm_n3162, gm_n3388, gm_n3173);
	nor (gm_n3390, gm_n3154, gm_n3150, gm_n3145, gm_n3389, gm_n3158);
	nand (gm_n3391, gm_n3138, gm_n3134, gm_n3131, gm_n3390, gm_n3142);
	nor (gm_n3392, gm_n3124, gm_n3121, gm_n3117, gm_n3391, gm_n3127);
	nand (gm_n3393, gm_n3109, gm_n3106, gm_n3102, gm_n3392, gm_n3113);
	nor (gm_n3394, gm_n3095, gm_n3090, gm_n3085, gm_n3393, gm_n3099);
	nand (gm_n3395, gm_n3076, gm_n3072, gm_n3068, gm_n3394, gm_n3081);
	nor (gm_n3396, gm_n3059, gm_n3055, gm_n3051, gm_n3395, gm_n3063);
	nand (gm_n3397, gm_n3042, gm_n3038, gm_n3034, gm_n3396, gm_n3047);
	nor (gm_n3398, gm_n3027, gm_n3025, gm_n3021, gm_n3397, gm_n3030);
	nand (gm_n3399, gm_n3015, gm_n3011, gm_n3008, gm_n3398, gm_n3018);
	nor (gm_n3400, gm_n3001, gm_n2997, gm_n2993, gm_n3399, gm_n3005);
	nand (gm_n3401, gm_n2987, gm_n2983, gm_n2980, gm_n3400, gm_n2990);
	nor (gm_n3402, gm_n2973, gm_n2969, gm_n2966, gm_n3401, gm_n2976);
	nand (gm_n3403, gm_n2959, gm_n2955, gm_n2950, gm_n3402, gm_n2963);
	nor (gm_n3404, gm_n2942, gm_n2938, gm_n2934, gm_n3403, gm_n2946);
	nand (gm_n3405, gm_n2925, gm_n2921, gm_n2918, gm_n3404, gm_n2930);
	nor (gm_n3406, gm_n2911, gm_n2906, gm_n2901, gm_n3405, gm_n2913);
	nand (gm_n3407, gm_n2893, gm_n2889, gm_n2884, gm_n3406, gm_n2897);
	nor (gm_n3408, gm_n2876, gm_n2871, gm_n2867, gm_n3407, gm_n2880);
	nand (gm_n3409, gm_n2860, gm_n2856, gm_n2853, gm_n3408, gm_n2863);
	nor (gm_n3410, gm_n2844, gm_n2840, gm_n2835, gm_n3409, gm_n2848);
	nand (gm_n3411, gm_n2827, gm_n2822, gm_n2818, gm_n3410, gm_n2831);
	nor (out_4, gm_n2810, gm_n2807, gm_n2804, gm_n3411, gm_n2814);
	and (gm_n3413, gm_n48, in_11, gm_n52, gm_n280, in_13);
	nand (gm_n3414, gm_n46, in_15, in_14, gm_n3413, in_17);
	nor (gm_n3415, gm_n45, gm_n62, gm_n47, gm_n3414, in_21);
	nor (gm_n3416, in_8, in_7, gm_n82, gm_n103, in_9);
	nand (gm_n3417, gm_n48, in_11, gm_n52, gm_n3416, gm_n49);
	nor (gm_n3418, in_16, in_15, in_14, gm_n3417, gm_n81);
	nand (gm_n3419, gm_n45, in_19, in_18, gm_n3418, in_21);
	nor (gm_n3420, in_10, gm_n51, gm_n64, gm_n853);
	nand (gm_n3421, in_13, gm_n48, gm_n53, gm_n3420, gm_n50);
	nor (gm_n3422, gm_n81, in_16, gm_n63, gm_n3421, gm_n47);
	nand (gm_n3423, in_21, gm_n45, gm_n62, gm_n3422);
	nor (gm_n3424, in_11, gm_n52, gm_n51, gm_n514, in_12);
	nand (gm_n3425, gm_n63, in_14, in_13, gm_n3424, gm_n46);
	nor (gm_n3426, in_19, in_18, gm_n81, gm_n3425, gm_n45);
	nand (gm_n3427, gm_n3426, gm_n71);
	or (gm_n3428, gm_n55, gm_n82, in_5, gm_n124, in_8);
	nor (gm_n3429, gm_n3428, gm_n52, gm_n51);
	nand (gm_n3430, gm_n49, gm_n48, gm_n53, gm_n3429, gm_n50);
	nor (gm_n3431, in_17, in_16, gm_n63, gm_n3430, gm_n47);
	nand (gm_n3432, in_21, gm_n45, gm_n62, gm_n3431);
	nand (gm_n3433, gm_n51, in_8, gm_n55, gm_n136, gm_n52);
	nor (gm_n3434, gm_n49, in_12, in_11, gm_n3433, in_14);
	nand (gm_n3435, in_17, gm_n46, gm_n63, gm_n3434, in_18);
	nor (gm_n3436, in_21, in_20, in_19, gm_n3435);
	nor (gm_n3437, in_14, gm_n49, gm_n48, gm_n369, gm_n63);
	nand (gm_n3438, in_18, gm_n81, in_16, gm_n3437, in_19);
	nor (gm_n3439, gm_n3438, gm_n71, in_20);
	nor (gm_n3440, gm_n49, gm_n48, gm_n53, gm_n2575, gm_n50);
	nand (gm_n3441, gm_n81, gm_n46, in_15, gm_n3440, gm_n47);
	nor (gm_n3442, in_21, in_20, in_19, gm_n3441);
	and (gm_n3443, gm_n673, in_9);
	and (gm_n3444, gm_n48, in_11, gm_n52, gm_n3443, in_13);
	nand (gm_n3445, in_16, gm_n63, gm_n50, gm_n3444, gm_n81);
	nor (gm_n3446, in_20, in_19, in_18, gm_n3445, in_21);
	and (gm_n3447, gm_n53, gm_n52, in_9, gm_n593, gm_n48);
	nand (gm_n3448, in_15, in_14, gm_n49, gm_n3447, gm_n46);
	nor (gm_n3449, gm_n62, gm_n47, gm_n81, gm_n3448, in_20);
	nand (gm_n3450, gm_n3449, in_21);
	and (gm_n3451, gm_n55, in_6, gm_n72, gm_n241, gm_n64);
	and (gm_n3452, gm_n53, in_10, in_9, gm_n3451, gm_n48);
	nand (gm_n3453, gm_n63, gm_n50, in_13, gm_n3452, in_16);
	nor (gm_n3454, in_19, in_18, in_17, gm_n3453, in_20);
	nand (gm_n3455, gm_n3454, gm_n71);
	and (gm_n3456, in_11, in_10, gm_n51, gm_n2234);
	nand (gm_n3457, gm_n50, gm_n49, in_12, gm_n3456, in_15);
	nor (gm_n3458, in_18, gm_n81, gm_n46, gm_n3457, gm_n62);
	nand (gm_n3459, gm_n3458, in_21, in_20);
	nor (gm_n3460, gm_n51, gm_n64, gm_n55, gm_n463, in_10);
	nand (gm_n3461, in_13, in_12, in_11, gm_n3460, in_14);
	nor (gm_n3462, in_17, gm_n46, in_15, gm_n3461, in_18);
	nand (gm_n3463, in_21, gm_n45, in_19, gm_n3462);
	nand (gm_n3464, in_11, in_10, in_9, gm_n1643, gm_n48);
	nor (gm_n3465, gm_n63, in_14, gm_n49, gm_n3464, in_16);
	nand (gm_n3466, gm_n62, in_18, in_17, gm_n3465, gm_n45);
	nor (gm_n3467, gm_n3466, in_21);
	nor (gm_n3468, gm_n49, gm_n48, in_11, gm_n2473, in_14);
	nand (gm_n3469, gm_n81, in_16, in_15, gm_n3468, gm_n47);
	nor (gm_n3470, in_21, gm_n45, gm_n62, gm_n3469);
	nor (gm_n3471, in_11, gm_n52, in_9, gm_n2445);
	and (gm_n3472, in_14, gm_n49, in_12, gm_n3471, in_15);
	nand (gm_n3473, gm_n47, gm_n81, in_16, gm_n3472, in_19);
	nor (gm_n3474, gm_n3473, in_21, gm_n45);
	nand (gm_n3475, in_7, in_6, gm_n72, gm_n241, gm_n64);
	or (gm_n3476, gm_n53, gm_n52, in_9, gm_n3475);
	nor (gm_n3477, in_14, in_13, in_12, gm_n3476, gm_n63);
	nand (gm_n3478, gm_n47, in_17, gm_n46, gm_n3477, in_19);
	nor (gm_n3479, gm_n3478, in_21, gm_n45);
	nor (gm_n3480, gm_n51, gm_n64, in_7, gm_n463, in_10);
	nand (gm_n3481, gm_n49, gm_n48, in_11, gm_n3480, gm_n50);
	nor (gm_n3482, in_17, gm_n46, gm_n63, gm_n3481, gm_n47);
	nand (gm_n3483, gm_n71, gm_n45, in_19, gm_n3482);
	nand (gm_n3484, gm_n55, gm_n82, gm_n72, gm_n519, in_8);
	nor (gm_n3485, gm_n53, gm_n52, gm_n51, gm_n3484, gm_n48);
	nand (gm_n3486, gm_n63, in_14, in_13, gm_n3485);
	nor (gm_n3487, in_18, gm_n81, gm_n46, gm_n3486, in_19);
	nand (gm_n3488, gm_n3487, gm_n71, in_20);
	and (gm_n3489, in_7, in_6, in_5, gm_n284, in_8);
	and (gm_n3490, in_11, gm_n52, in_9, gm_n3489, gm_n48);
	nand (gm_n3491, gm_n63, in_14, in_13, gm_n3490, in_16);
	nor (gm_n3492, gm_n62, in_18, in_17, gm_n3491, in_20);
	nand (gm_n3493, gm_n3492, gm_n71);
	or (gm_n3494, gm_n51, gm_n64, in_7, gm_n279, gm_n52);
	nor (gm_n3495, gm_n49, in_12, in_11, gm_n3494);
	and (gm_n3496, gm_n46, in_15, in_14, gm_n3495, gm_n81);
	nand (gm_n3497, gm_n45, gm_n62, in_18, gm_n3496, in_21);
	nor (gm_n3498, in_12, in_11, in_10, gm_n1784, gm_n49);
	nand (gm_n3499, in_16, in_15, in_14, gm_n3498, in_17);
	nor (gm_n3500, gm_n45, gm_n62, in_18, gm_n3499, gm_n71);
	or (gm_n3501, gm_n53, gm_n52, in_9, gm_n1261, gm_n48);
	nor (gm_n3502, in_15, gm_n50, gm_n49, gm_n3501, gm_n46);
	nand (gm_n3503, gm_n62, gm_n47, in_17, gm_n3502, gm_n45);
	nor (gm_n3504, gm_n3503, in_21);
	nor (gm_n3505, gm_n48, gm_n53, gm_n52, gm_n3159, in_13);
	nand (gm_n3506, in_16, in_15, in_14, gm_n3505, gm_n81);
	nor (gm_n3507, in_20, in_19, in_18, gm_n3506, in_21);
	or (gm_n3508, gm_n51, in_8, gm_n55, gm_n463);
	nor (gm_n3509, in_12, in_11, gm_n52, gm_n3508, in_13);
	nand (gm_n3510, gm_n46, gm_n63, in_14, gm_n3509, gm_n81);
	nor (gm_n3511, gm_n45, gm_n62, gm_n47, gm_n3510, in_21);
	nand (gm_n3512, in_14, gm_n49, in_12, gm_n1444, gm_n63);
	nor (gm_n3513, gm_n47, gm_n81, in_16, gm_n3512, gm_n62);
	nand (gm_n3514, gm_n3513, gm_n71, in_20);
	nand (gm_n3515, in_8, in_7, gm_n82, gm_n2640, in_9);
	or (gm_n3516, gm_n48, in_11, in_10, gm_n3515, in_13);
	nor (gm_n3517, gm_n46, in_15, gm_n50, gm_n3516, gm_n81);
	nand (gm_n3518, gm_n45, in_19, gm_n47, gm_n3517, gm_n71);
	nor (gm_n3519, in_7, gm_n82, gm_n72, gm_n643, gm_n64);
	and (gm_n3520, gm_n53, gm_n52, in_9, gm_n3519, gm_n48);
	nand (gm_n3521, gm_n63, gm_n50, in_13, gm_n3520, gm_n46);
	nor (gm_n3522, in_19, gm_n47, in_17, gm_n3521, gm_n45);
	nand (gm_n3523, gm_n3522, gm_n71);
	nor (gm_n3524, in_11, gm_n52, gm_n51, gm_n2345);
	nand (gm_n3525, gm_n50, in_13, in_12, gm_n3524, in_15);
	nor (gm_n3526, gm_n47, in_17, in_16, gm_n3525, in_19);
	nand (gm_n3527, gm_n3526, in_21, in_20);
	nor (gm_n3528, gm_n51, gm_n64, gm_n55, gm_n553, in_10);
	and (gm_n3529, in_13, gm_n48, in_11, gm_n3528, in_14);
	nand (gm_n3530, in_17, in_16, in_15, gm_n3529, gm_n47);
	nor (gm_n3531, gm_n71, gm_n45, gm_n62, gm_n3530);
	nand (gm_n3532, gm_n46, in_15, gm_n50, gm_n2598, gm_n81);
	nor (gm_n3533, gm_n45, gm_n62, gm_n47, gm_n3532, in_21);
	nand (gm_n3534, gm_n2907, gm_n52, gm_n51);
	nor (gm_n3535, in_13, in_12, in_11, gm_n3534, in_14);
	nand (gm_n3536, gm_n81, gm_n46, in_15, gm_n3535, gm_n47);
	nor (gm_n3537, in_21, in_20, gm_n62, gm_n3536);
	nand (gm_n3538, gm_n53, in_10, gm_n51, gm_n194, gm_n48);
	nor (gm_n3539, in_15, in_14, in_13, gm_n3538, in_16);
	nand (gm_n3540, in_19, gm_n47, gm_n81, gm_n3539, in_20);
	nor (gm_n3541, gm_n3540, in_21);
	nand (gm_n3542, in_7, in_6, gm_n72, gm_n209, gm_n64);
	nor (gm_n3543, gm_n3542, in_10, in_9);
	nand (gm_n3544, gm_n49, in_12, gm_n53, gm_n3543, in_14);
	nor (gm_n3545, in_17, gm_n46, gm_n63, gm_n3544, gm_n47);
	nand (gm_n3546, gm_n71, gm_n45, gm_n62, gm_n3545);
	and (gm_n3547, in_11, gm_n52, gm_n51, gm_n1563);
	nand (gm_n3548, gm_n50, in_13, in_12, gm_n3547, gm_n63);
	nor (gm_n3549, in_18, gm_n81, gm_n46, gm_n3548, gm_n62);
	nand (gm_n3550, gm_n3549, in_21, in_20);
	nor (gm_n3551, in_16, in_15, gm_n50, gm_n2919, gm_n81);
	nand (gm_n3552, gm_n45, gm_n62, in_18, gm_n3551, in_21);
	nor (gm_n3553, gm_n64, gm_n55, in_6, gm_n119, gm_n51);
	nand (gm_n3554, gm_n48, in_11, gm_n52, gm_n3553, gm_n49);
	nor (gm_n3555, gm_n46, in_15, in_14, gm_n3554, gm_n81);
	nand (gm_n3556, gm_n45, gm_n62, gm_n47, gm_n3555, gm_n71);
	nand (gm_n3557, gm_n55, gm_n82, in_5, gm_n89, gm_n64);
	nor (gm_n3558, in_11, gm_n52, gm_n51, gm_n3557, gm_n48);
	and (gm_n3559, in_15, gm_n50, in_13, gm_n3558, gm_n46);
	nand (gm_n3560, in_19, gm_n47, gm_n81, gm_n3559, gm_n45);
	nor (gm_n3561, gm_n3560, gm_n71);
	and (gm_n3562, gm_n64, in_7, gm_n82, gm_n1075, gm_n51);
	and (gm_n3563, in_12, in_11, in_10, gm_n3562, gm_n49);
	nand (gm_n3564, in_16, in_15, gm_n50, gm_n3563, in_17);
	nor (gm_n3565, gm_n45, in_19, in_18, gm_n3564, gm_n71);
	and (gm_n3566, gm_n64, gm_n55, in_6, gm_n2640, gm_n51);
	and (gm_n3567, gm_n48, in_11, in_10, gm_n3566, gm_n49);
	nand (gm_n3568, in_16, in_15, gm_n50, gm_n3567, in_17);
	nor (gm_n3569, in_20, in_19, in_18, gm_n3568, in_21);
	nor (gm_n3570, gm_n49, gm_n48, in_11, gm_n1812, in_14);
	nand (gm_n3571, in_17, gm_n46, gm_n63, gm_n3570, in_18);
	nor (gm_n3572, in_21, in_20, in_19, gm_n3571);
	nor (gm_n3573, in_9, in_8, in_7, gm_n223, in_10);
	nand (gm_n3574, gm_n49, gm_n48, in_11, gm_n3573, in_14);
	nor (gm_n3575, in_17, in_16, in_15, gm_n3574, gm_n47);
	nand (gm_n3576, gm_n71, in_20, in_19, gm_n3575);
	and (gm_n3577, in_11, in_10, in_9, gm_n2907);
	and (gm_n3578, gm_n3577, gm_n49, gm_n48);
	and (gm_n3579, gm_n46, gm_n63, gm_n50, gm_n3578, in_17);
	nand (gm_n3580, in_20, in_19, gm_n47, gm_n3579, in_21);
	nand (gm_n3581, gm_n48, gm_n53, in_10, gm_n1962, in_13);
	nor (gm_n3582, gm_n46, gm_n63, in_14, gm_n3581, gm_n81);
	nand (gm_n3583, gm_n45, in_19, gm_n47, gm_n3582, in_21);
	nand (gm_n3584, in_11, gm_n52, gm_n51, gm_n668);
	or (gm_n3585, gm_n50, in_13, gm_n48, gm_n3584, in_15);
	nor (gm_n3586, gm_n47, in_17, in_16, gm_n3585, gm_n62);
	nand (gm_n3587, gm_n3586, gm_n71, gm_n45);
	nand (gm_n3588, gm_n53, in_10, in_9, gm_n868, gm_n48);
	nor (gm_n3589, in_15, in_14, in_13, gm_n3588, in_16);
	nand (gm_n3590, in_19, gm_n47, in_17, gm_n3589, in_20);
	nor (gm_n3591, gm_n3590, in_21);
	nor (gm_n3592, gm_n50, gm_n49, in_12, gm_n1546, in_15);
	nand (gm_n3593, in_18, in_17, in_16, gm_n3592, in_19);
	nor (gm_n3594, gm_n3593, in_21, in_20);
	nand (gm_n3595, gm_n46, in_15, gm_n50, gm_n3032, gm_n81);
	nor (gm_n3596, in_20, gm_n62, in_18, gm_n3595, in_21);
	nand (gm_n3597, gm_n53, in_10, gm_n51, gm_n1704, gm_n48);
	nor (gm_n3598, gm_n63, in_14, gm_n49, gm_n3597, gm_n46);
	nand (gm_n3599, gm_n62, gm_n47, gm_n81, gm_n3598, in_20);
	nor (gm_n3600, gm_n3599, in_21);
	or (gm_n3601, in_9, gm_n64, in_7, gm_n525, gm_n52);
	nor (gm_n3602, gm_n3601, in_11);
	nand (gm_n3603, gm_n50, in_13, in_12, gm_n3602, gm_n63);
	nor (gm_n3604, gm_n47, gm_n81, gm_n46, gm_n3603, gm_n62);
	nand (gm_n3605, gm_n3604, gm_n71, gm_n45);
	nor (gm_n3606, in_7, in_6, gm_n72, gm_n290, in_8);
	nand (gm_n3607, in_11, in_10, in_9, gm_n3606, in_12);
	or (gm_n3608, gm_n63, in_14, in_13, gm_n3607, gm_n46);
	nor (gm_n3609, gm_n62, in_18, in_17, gm_n3608, in_20);
	nand (gm_n3610, gm_n3609, gm_n71);
	nor (gm_n3611, gm_n64, gm_n55, gm_n82, gm_n103, in_9);
	nand (gm_n3612, gm_n48, in_11, gm_n52, gm_n3611, gm_n49);
	nor (gm_n3613, gm_n46, in_15, in_14, gm_n3612, in_17);
	nand (gm_n3614, gm_n45, gm_n62, gm_n47, gm_n3613, in_21);
	nor (gm_n3615, gm_n2300, in_10, in_9);
	nand (gm_n3616, in_13, in_12, gm_n53, gm_n3615, gm_n50);
	nor (gm_n3617, gm_n81, in_16, in_15, gm_n3616, gm_n47);
	nand (gm_n3618, in_21, in_20, in_19, gm_n3617);
	nor (gm_n3619, gm_n50, in_13, in_12, gm_n726, gm_n63);
	nand (gm_n3620, gm_n47, gm_n81, in_16, gm_n3619, gm_n62);
	nor (gm_n3621, gm_n3620, in_21, gm_n45);
	and (gm_n3622, gm_n63, gm_n50, in_13, gm_n1928, in_16);
	nand (gm_n3623, gm_n62, in_18, in_17, gm_n3622, in_20);
	nor (gm_n3624, gm_n3623, gm_n71);
	nor (gm_n3625, in_13, in_12, in_11, gm_n385, in_14);
	nand (gm_n3626, in_17, gm_n46, gm_n63, gm_n3625, in_18);
	nor (gm_n3627, gm_n71, in_20, in_19, gm_n3626);
	and (gm_n3628, gm_n53, gm_n52, gm_n51, gm_n355, gm_n48);
	and (gm_n3629, gm_n63, gm_n50, gm_n49, gm_n3628, in_16);
	nand (gm_n3630, gm_n62, in_18, in_17, gm_n3629, gm_n45);
	nor (gm_n3631, gm_n3630, gm_n71);
	nand (gm_n3632, in_8, gm_n55, gm_n82, gm_n1075, gm_n51);
	nor (gm_n3633, gm_n3632, in_11, gm_n52);
	nand (gm_n3634, in_14, gm_n49, gm_n48, gm_n3633, gm_n63);
	nor (gm_n3635, in_18, gm_n81, gm_n46, gm_n3634, in_19);
	nand (gm_n3636, gm_n3635, in_21, gm_n45);
	nand (gm_n3637, gm_n48, gm_n53, in_10, gm_n2693, gm_n49);
	nor (gm_n3638, in_16, gm_n63, gm_n50, gm_n3637, gm_n81);
	nand (gm_n3639, in_20, gm_n62, in_18, gm_n3638, gm_n71);
	and (gm_n3640, gm_n53, gm_n52, gm_n51, gm_n621);
	and (gm_n3641, gm_n3640, in_13, in_12);
	and (gm_n3642, gm_n46, in_15, gm_n50, gm_n3641, gm_n81);
	nand (gm_n3643, in_20, in_19, gm_n47, gm_n3642, in_21);
	nand (gm_n3644, gm_n53, in_10, gm_n51, gm_n291);
	or (gm_n3645, gm_n50, gm_n49, in_12, gm_n3644, in_15);
	nor (gm_n3646, gm_n47, in_17, in_16, gm_n3645, gm_n62);
	nand (gm_n3647, gm_n3646, gm_n71, gm_n45);
	nor (gm_n3648, in_12, gm_n53, gm_n52, gm_n1900, gm_n49);
	nand (gm_n3649, gm_n46, in_15, in_14, gm_n3648, in_17);
	nor (gm_n3650, in_20, gm_n62, in_18, gm_n3649, gm_n71);
	nor (gm_n3651, in_9, gm_n64, gm_n55, gm_n223, gm_n52);
	and (gm_n3652, in_13, in_12, in_11, gm_n3651, gm_n50);
	nand (gm_n3653, in_17, gm_n46, in_15, gm_n3652, in_18);
	nor (gm_n3654, in_21, gm_n45, in_19, gm_n3653);
	nand (gm_n3655, gm_n51, gm_n64, gm_n55, gm_n504, gm_n52);
	nor (gm_n3656, gm_n49, in_12, gm_n53, gm_n3655, gm_n50);
	nand (gm_n3657, gm_n81, gm_n46, in_15, gm_n3656, gm_n47);
	nor (gm_n3658, gm_n71, gm_n45, in_19, gm_n3657);
	and (gm_n3659, gm_n64, in_7, in_6, gm_n374, in_9);
	and (gm_n3660, gm_n48, in_11, in_10, gm_n3659, in_13);
	nand (gm_n3661, gm_n46, in_15, in_14, gm_n3660, in_17);
	nor (gm_n3662, gm_n45, in_19, gm_n47, gm_n3661, gm_n71);
	nand (gm_n3663, gm_n49, gm_n48, in_11, gm_n351, gm_n50);
	nor (gm_n3664, gm_n81, gm_n46, gm_n63, gm_n3663, gm_n47);
	nand (gm_n3665, gm_n71, gm_n45, gm_n62, gm_n3664);
	nand (gm_n3666, in_11, in_10, in_9, gm_n868);
	or (gm_n3667, gm_n50, in_13, in_12, gm_n3666, gm_n63);
	nor (gm_n3668, gm_n47, gm_n81, in_16, gm_n3667, gm_n62);
	nand (gm_n3669, gm_n3668, gm_n71, gm_n45);
	nor (gm_n3670, in_11, in_10, gm_n51, gm_n218, in_12);
	nand (gm_n3671, gm_n63, gm_n50, gm_n49, gm_n3670, gm_n46);
	nor (gm_n3672, in_19, gm_n47, gm_n81, gm_n3671, in_20);
	nand (gm_n3673, gm_n3672, in_21);
	and (gm_n3674, gm_n49, in_12, gm_n53, gm_n1094, gm_n50);
	and (gm_n3675, gm_n81, gm_n46, gm_n63, gm_n3674, gm_n47);
	nand (gm_n3676, in_21, gm_n45, in_19, gm_n3675);
	and (gm_n3677, gm_n838, gm_n51, gm_n64);
	and (gm_n3678, gm_n48, in_11, gm_n52, gm_n3677, gm_n49);
	nand (gm_n3679, in_16, gm_n63, in_14, gm_n3678, gm_n81);
	nor (gm_n3680, gm_n45, in_19, in_18, gm_n3679, gm_n71);
	nand (gm_n3681, gm_n46, gm_n63, in_14, gm_n1390, in_17);
	nor (gm_n3682, gm_n45, gm_n62, in_18, gm_n3681, gm_n71);
	nand (gm_n3683, gm_n64, in_7, gm_n82, gm_n374, in_9);
	nor (gm_n3684, in_12, gm_n53, gm_n52, gm_n3683, in_13);
	nand (gm_n3685, gm_n46, gm_n63, in_14, gm_n3684, in_17);
	nor (gm_n3686, gm_n45, in_19, in_18, gm_n3685, in_21);
	nor (gm_n3687, in_9, in_8, in_7, gm_n588, in_10);
	and (gm_n3688, in_13, in_12, in_11, gm_n3687, gm_n50);
	nand (gm_n3689, in_17, in_16, gm_n63, gm_n3688, in_18);
	nor (gm_n3690, gm_n71, in_20, in_19, gm_n3689);
	nand (gm_n3691, in_12, gm_n53, gm_n52, gm_n2760, gm_n49);
	nor (gm_n3692, gm_n46, gm_n63, in_14, gm_n3691, gm_n81);
	nand (gm_n3693, gm_n45, in_19, gm_n47, gm_n3692, in_21);
	nand (gm_n3694, gm_n63, in_14, in_13, gm_n984, in_16);
	nor (gm_n3695, in_19, gm_n47, gm_n81, gm_n3694, gm_n45);
	nand (gm_n3696, gm_n3695, in_21);
	nand (gm_n3697, gm_n55, gm_n82, in_5, gm_n284, gm_n64);
	nor (gm_n3698, gm_n53, gm_n52, gm_n51, gm_n3697, in_12);
	nand (gm_n3699, in_15, gm_n50, gm_n49, gm_n3698, in_16);
	nor (gm_n3700, in_19, gm_n47, gm_n81, gm_n3699, in_20);
	nand (gm_n3701, gm_n3700, gm_n71);
	nand (gm_n3702, gm_n48, in_11, in_10, gm_n2555, in_13);
	nor (gm_n3703, in_16, in_15, gm_n50, gm_n3702, gm_n81);
	nand (gm_n3704, in_20, in_19, in_18, gm_n3703, in_21);
	and (gm_n3705, gm_n49, in_12, in_11, gm_n1344, gm_n50);
	nand (gm_n3706, in_17, gm_n46, gm_n63, gm_n3705, gm_n47);
	nor (gm_n3707, in_21, in_20, in_19, gm_n3706);
	nor (gm_n3708, in_9, gm_n64, in_7, gm_n84, gm_n52);
	and (gm_n3709, gm_n49, in_12, in_11, gm_n3708, gm_n50);
	nand (gm_n3710, in_17, in_16, gm_n63, gm_n3709, in_18);
	nor (gm_n3711, gm_n71, gm_n45, in_19, gm_n3710);
	nor (gm_n3712, gm_n2564, gm_n52, gm_n51);
	and (gm_n3713, gm_n49, in_12, in_11, gm_n3712, gm_n50);
	nand (gm_n3714, gm_n81, gm_n46, in_15, gm_n3713, in_18);
	nor (gm_n3715, gm_n71, gm_n45, gm_n62, gm_n3714);
	nand (gm_n3716, in_16, in_15, in_14, gm_n3185, gm_n81);
	nor (gm_n3717, gm_n45, gm_n62, in_18, gm_n3716, gm_n71);
	nand (gm_n3718, gm_n55, in_6, gm_n72, gm_n493);
	nor (gm_n3719, gm_n52, gm_n51, gm_n64, gm_n3718, gm_n53);
	nand (gm_n3720, in_14, in_13, in_12, gm_n3719, in_15);
	nor (gm_n3721, in_18, gm_n81, gm_n46, gm_n3720, gm_n62);
	nand (gm_n3722, gm_n3721, gm_n71, in_20);
	and (gm_n3723, gm_n51, gm_n64, in_7, gm_n136);
	nand (gm_n3724, in_12, gm_n53, in_10, gm_n3723, gm_n49);
	nor (gm_n3725, gm_n46, gm_n63, gm_n50, gm_n3724, in_17);
	nand (gm_n3726, gm_n45, in_19, gm_n47, gm_n3725, gm_n71);
	and (gm_n3727, gm_n51, in_8, gm_n55, gm_n151);
	nand (gm_n3728, gm_n48, in_11, in_10, gm_n3727, gm_n49);
	nor (gm_n3729, in_16, in_15, gm_n50, gm_n3728, in_17);
	nand (gm_n3730, gm_n45, in_19, in_18, gm_n3729, in_21);
	and (gm_n3731, in_8, gm_n55, in_6, gm_n1075, gm_n51);
	nand (gm_n3732, gm_n48, in_11, in_10, gm_n3731, gm_n49);
	nor (gm_n3733, in_16, in_15, in_14, gm_n3732, gm_n81);
	nand (gm_n3734, gm_n45, in_19, in_18, gm_n3733, gm_n71);
	and (gm_n3735, gm_n53, in_10, gm_n51, gm_n3193, in_12);
	and (gm_n3736, gm_n63, in_14, gm_n49, gm_n3735, gm_n46);
	nand (gm_n3737, in_19, gm_n47, gm_n81, gm_n3736, in_20);
	nor (gm_n3738, gm_n3737, in_21);
	nand (gm_n3739, gm_n53, in_10, gm_n51, gm_n1070, gm_n48);
	nor (gm_n3740, in_15, gm_n50, gm_n49, gm_n3739, gm_n46);
	nand (gm_n3741, gm_n62, in_18, gm_n81, gm_n3740, gm_n45);
	nor (gm_n3742, gm_n3741, gm_n71);
	nand (gm_n3743, in_7, gm_n82, in_5, gm_n241, in_8);
	nor (gm_n3744, gm_n3743, in_9);
	and (gm_n3745, gm_n48, gm_n53, in_10, gm_n3744, gm_n49);
	nand (gm_n3746, gm_n46, gm_n63, gm_n50, gm_n3745, gm_n81);
	nor (gm_n3747, in_20, gm_n62, in_18, gm_n3746, gm_n71);
	nor (gm_n3748, gm_n64, in_7, gm_n82, gm_n1429, in_9);
	and (gm_n3749, in_12, gm_n53, gm_n52, gm_n3748, in_13);
	nand (gm_n3750, gm_n46, gm_n63, gm_n50, gm_n3749, in_17);
	nor (gm_n3751, in_20, in_19, in_18, gm_n3750, gm_n71);
	nor (gm_n3752, gm_n53, gm_n52, in_9, gm_n583, gm_n48);
	nand (gm_n3753, in_15, gm_n50, in_13, gm_n3752, in_16);
	nor (gm_n3754, in_19, gm_n47, in_17, gm_n3753, gm_n45);
	nand (gm_n3755, gm_n3754, in_21);
	nor (gm_n3756, in_9, in_8, in_7, gm_n1256, gm_n52);
	nand (gm_n3757, in_13, gm_n48, in_11, gm_n3756, in_14);
	nor (gm_n3758, in_17, gm_n46, in_15, gm_n3757, in_18);
	nand (gm_n3759, in_21, gm_n45, in_19, gm_n3758);
	nor (gm_n3760, gm_n53, in_10, in_9, gm_n333);
	nand (gm_n3761, gm_n50, in_13, in_12, gm_n3760, in_15);
	nor (gm_n3762, in_18, in_17, in_16, gm_n3761, gm_n62);
	nand (gm_n3763, gm_n3762, in_21, in_20);
	or (gm_n3764, in_8, in_7, gm_n82, gm_n1429, in_9);
	nor (gm_n3765, gm_n48, in_11, in_10, gm_n3764, in_13);
	nand (gm_n3766, gm_n46, in_15, gm_n50, gm_n3765, gm_n81);
	or (gm_n3767, in_20, in_19, in_18, gm_n3766, in_21);
	nor (gm_n3768, gm_n55, gm_n82, gm_n72, gm_n483, in_8);
	nand (gm_n3769, in_11, in_10, in_9, gm_n3768, in_12);
	nor (gm_n3770, in_15, in_14, gm_n49, gm_n3769, in_16);
	nand (gm_n3771, gm_n62, gm_n47, in_17, gm_n3770, gm_n45);
	nor (gm_n3772, gm_n3771, in_21);
	or (gm_n3773, in_9, in_8, gm_n55, gm_n259);
	nor (gm_n3774, in_12, in_11, in_10, gm_n3773, gm_n49);
	nand (gm_n3775, in_16, gm_n63, gm_n50, gm_n3774, gm_n81);
	nor (gm_n3776, gm_n45, in_19, gm_n47, gm_n3775, in_21);
	nand (gm_n3777, in_11, in_10, in_9, gm_n494, gm_n48);
	nor (gm_n3778, gm_n63, in_14, in_13, gm_n3777, gm_n46);
	nand (gm_n3779, in_19, gm_n47, in_17, gm_n3778, in_20);
	nor (gm_n3780, gm_n3779, in_21);
	nand (gm_n3781, in_8, in_7, in_6, gm_n374, gm_n51);
	nor (gm_n3782, in_12, gm_n53, gm_n52, gm_n3781, gm_n49);
	nand (gm_n3783, gm_n46, gm_n63, gm_n50, gm_n3782, gm_n81);
	nor (gm_n3784, in_20, gm_n62, in_18, gm_n3783, in_21);
	nor (gm_n3785, in_8, in_7, in_6, gm_n156, in_9);
	and (gm_n3786, in_12, in_11, gm_n52, gm_n3785, gm_n49);
	and (gm_n3787, in_16, in_15, in_14, gm_n3786, in_17);
	nand (gm_n3788, in_20, in_19, gm_n47, gm_n3787, in_21);
	nor (gm_n3789, gm_n51, in_8, gm_n55, gm_n525, gm_n52);
	nand (gm_n3790, in_13, gm_n48, in_11, gm_n3789, in_14);
	nor (gm_n3791, in_17, gm_n46, gm_n63, gm_n3790, gm_n47);
	nand (gm_n3792, gm_n71, in_20, gm_n62, gm_n3791);
	nand (gm_n3793, in_14, gm_n49, in_12, gm_n1089, in_15);
	nor (gm_n3794, gm_n47, gm_n81, gm_n46, gm_n3793, in_19);
	nand (gm_n3795, gm_n3794, in_21, in_20);
	nand (gm_n3796, gm_n48, in_11, in_10, gm_n200, gm_n49);
	nor (gm_n3797, gm_n46, gm_n63, gm_n50, gm_n3796, in_17);
	nand (gm_n3798, in_20, gm_n62, gm_n47, gm_n3797, gm_n71);
	or (gm_n3799, gm_n46, in_15, gm_n50, gm_n3070, in_17);
	nor (gm_n3800, gm_n45, in_19, in_18, gm_n3799, gm_n71);
	nor (gm_n3801, in_13, in_12, gm_n53, gm_n3534, in_14);
	nand (gm_n3802, gm_n81, in_16, gm_n63, gm_n3801, in_18);
	nor (gm_n3803, in_21, gm_n45, gm_n62, gm_n3802);
	and (gm_n3804, in_7, gm_n82, gm_n72, gm_n241, gm_n64);
	and (gm_n3805, in_11, in_10, in_9, gm_n3804);
	and (gm_n3806, gm_n50, gm_n49, in_12, gm_n3805, gm_n63);
	nand (gm_n3807, in_18, gm_n81, gm_n46, gm_n3806, gm_n62);
	nor (gm_n3808, gm_n3807, in_21, in_20);
	nand (gm_n3809, in_8, in_7, gm_n82, gm_n757, gm_n51);
	nor (gm_n3810, gm_n48, in_11, in_10, gm_n3809, gm_n49);
	nand (gm_n3811, in_16, in_15, gm_n50, gm_n3810, gm_n81);
	nor (gm_n3812, in_20, in_19, in_18, gm_n3811, gm_n71);
	and (gm_n3813, gm_n53, gm_n52, gm_n51, gm_n1874, in_12);
	nand (gm_n3814, in_15, gm_n50, gm_n49, gm_n3813, in_16);
	nor (gm_n3815, in_19, in_18, gm_n81, gm_n3814, in_20);
	nand (gm_n3816, gm_n3815, in_21);
	nor (gm_n3817, gm_n53, in_10, gm_n51, gm_n873, in_12);
	nand (gm_n3818, in_15, gm_n50, in_13, gm_n3817, gm_n46);
	nor (gm_n3819, gm_n62, in_18, gm_n81, gm_n3818, in_20);
	nand (gm_n3820, gm_n3819, in_21);
	nand (gm_n3821, gm_n55, gm_n82, in_5, gm_n209);
	nor (gm_n3822, gm_n52, gm_n51, in_8, gm_n3821, gm_n53);
	nand (gm_n3823, in_14, in_13, in_12, gm_n3822, in_15);
	nor (gm_n3824, gm_n47, in_17, gm_n46, gm_n3823, gm_n62);
	nand (gm_n3825, gm_n3824, gm_n71, in_20);
	nand (gm_n3826, in_11, in_10, gm_n51, gm_n484);
	or (gm_n3827, gm_n50, gm_n49, in_12, gm_n3826, in_15);
	nor (gm_n3828, in_18, in_17, gm_n46, gm_n3827, in_19);
	nand (gm_n3829, gm_n3828, in_21, in_20);
	nor (gm_n3830, in_12, in_11, in_10, gm_n1684, in_13);
	nand (gm_n3831, in_16, gm_n63, gm_n50, gm_n3830, gm_n81);
	nor (gm_n3832, gm_n45, in_19, in_18, gm_n3831, gm_n71);
	nand (gm_n3833, gm_n868, gm_n52, gm_n51);
	nor (gm_n3834, in_13, gm_n48, in_11, gm_n3833, gm_n50);
	nand (gm_n3835, in_17, in_16, in_15, gm_n3834, in_18);
	nor (gm_n3836, gm_n71, in_20, in_19, gm_n3835);
	and (gm_n3837, in_13, in_12, gm_n53, gm_n1058, in_14);
	nand (gm_n3838, in_17, gm_n46, gm_n63, gm_n3837, gm_n47);
	nor (gm_n3839, in_21, in_20, gm_n62, gm_n3838);
	nand (gm_n3840, gm_n53, in_10, in_9, gm_n484, gm_n48);
	nor (gm_n3841, gm_n63, gm_n50, in_13, gm_n3840, in_16);
	nand (gm_n3842, gm_n62, in_18, gm_n81, gm_n3841, in_20);
	nor (gm_n3843, gm_n3842, in_21);
	or (gm_n3844, in_7, gm_n82, gm_n72, gm_n321, in_8);
	nor (gm_n3845, gm_n53, in_10, gm_n51, gm_n3844, gm_n48);
	nand (gm_n3846, in_15, gm_n50, in_13, gm_n3845, in_16);
	nor (gm_n3847, gm_n62, gm_n47, in_17, gm_n3846, in_20);
	nand (gm_n3848, gm_n3847, in_21);
	and (gm_n3849, gm_n53, in_10, gm_n51, gm_n3768, gm_n48);
	nand (gm_n3850, gm_n63, gm_n50, in_13, gm_n3849, in_16);
	nor (gm_n3851, in_19, gm_n47, in_17, gm_n3850, in_20);
	nand (gm_n3852, gm_n3851, gm_n71);
	nand (gm_n3853, in_15, in_14, in_13, gm_n459, in_16);
	nor (gm_n3854, in_19, in_18, gm_n81, gm_n3853, in_20);
	nand (gm_n3855, gm_n3854, gm_n71);
	nor (gm_n3856, in_7, in_6, gm_n72, gm_n321, in_8);
	and (gm_n3857, gm_n3856, in_10, gm_n51);
	nand (gm_n3858, gm_n49, in_12, gm_n53, gm_n3857, gm_n50);
	nor (gm_n3859, gm_n81, gm_n46, in_15, gm_n3858, gm_n47);
	nand (gm_n3860, gm_n71, in_20, in_19, gm_n3859);
	nand (gm_n3861, in_11, gm_n52, gm_n51, gm_n1683, gm_n48);
	nor (gm_n3862, in_15, in_14, in_13, gm_n3861, gm_n46);
	nand (gm_n3863, gm_n62, gm_n47, gm_n81, gm_n3862, in_20);
	nor (gm_n3864, gm_n3863, gm_n71);
	nor (gm_n3865, gm_n63, gm_n50, in_13, gm_n2939, in_16);
	nand (gm_n3866, gm_n62, gm_n47, gm_n81, gm_n3865, in_20);
	nor (gm_n3867, gm_n3866, in_21);
	nand (gm_n3868, gm_n53, in_10, gm_n51, gm_n538, in_12);
	nor (gm_n3869, gm_n63, gm_n50, gm_n49, gm_n3868, gm_n46);
	nand (gm_n3870, in_19, gm_n47, in_17, gm_n3869, gm_n45);
	nor (gm_n3871, gm_n3870, in_21);
	nand (gm_n3872, gm_n53, gm_n52, gm_n51, gm_n1178, in_12);
	nor (gm_n3873, in_15, in_14, gm_n49, gm_n3872, in_16);
	nand (gm_n3874, in_19, gm_n47, gm_n81, gm_n3873, gm_n45);
	nor (gm_n3875, gm_n3874, gm_n71);
	and (gm_n3876, gm_n53, in_10, gm_n51, gm_n1895, gm_n48);
	nand (gm_n3877, gm_n63, gm_n50, gm_n49, gm_n3876, gm_n46);
	nor (gm_n3878, in_19, in_18, gm_n81, gm_n3877, gm_n45);
	nand (gm_n3879, gm_n3878, gm_n71);
	nor (gm_n3880, gm_n53, in_10, in_9, gm_n520, in_12);
	nand (gm_n3881, in_15, gm_n50, in_13, gm_n3880, in_16);
	nor (gm_n3882, in_19, in_18, in_17, gm_n3881, in_20);
	nand (gm_n3883, gm_n3882, in_21);
	nand (gm_n3884, gm_n55, gm_n82, in_5, gm_n241, in_8);
	nor (gm_n3885, gm_n3884, in_10, gm_n51);
	nand (gm_n3886, in_13, in_12, in_11, gm_n3885, gm_n50);
	nor (gm_n3887, in_17, in_16, in_15, gm_n3886, in_18);
	nand (gm_n3888, in_21, in_20, in_19, gm_n3887);
	nor (gm_n3889, gm_n183, gm_n52, in_9);
	nand (gm_n3890, gm_n49, in_12, gm_n53, gm_n3889, gm_n50);
	nor (gm_n3891, in_17, in_16, in_15, gm_n3890, gm_n47);
	nand (gm_n3892, gm_n71, gm_n45, gm_n62, gm_n3891);
	nand (gm_n3893, gm_n3193, in_10, in_9);
	nor (gm_n3894, in_13, gm_n48, in_11, gm_n3893, gm_n50);
	nand (gm_n3895, gm_n81, gm_n46, in_15, gm_n3894, in_18);
	nor (gm_n3896, gm_n71, in_20, gm_n62, gm_n3895);
	nand (gm_n3897, in_11, in_10, in_9, gm_n858, gm_n48);
	nor (gm_n3898, gm_n63, in_14, in_13, gm_n3897, gm_n46);
	nand (gm_n3899, gm_n62, in_18, in_17, gm_n3898, gm_n45);
	nor (gm_n3900, gm_n3899, in_21);
	and (gm_n3901, gm_n48, gm_n53, in_10, gm_n980, gm_n49);
	nand (gm_n3902, gm_n46, gm_n63, in_14, gm_n3901, in_17);
	nor (gm_n3903, in_20, in_19, gm_n47, gm_n3902, gm_n71);
	and (gm_n3904, in_7, gm_n82, in_5, gm_n89, gm_n64);
	and (gm_n3905, gm_n3904, in_10, gm_n51);
	and (gm_n3906, gm_n49, in_12, in_11, gm_n3905, in_14);
	nand (gm_n3907, in_17, in_16, gm_n63, gm_n3906, in_18);
	nor (gm_n3908, gm_n71, gm_n45, in_19, gm_n3907);
	nor (gm_n3909, in_8, gm_n55, gm_n82, gm_n204, gm_n51);
	nand (gm_n3910, gm_n48, gm_n53, gm_n52, gm_n3909, in_13);
	nor (gm_n3911, in_16, in_15, in_14, gm_n3910, in_17);
	nand (gm_n3912, gm_n45, in_19, gm_n47, gm_n3911, in_21);
	nand (gm_n3913, in_12, gm_n53, in_10, gm_n2551, gm_n49);
	nor (gm_n3914, gm_n46, gm_n63, in_14, gm_n3913, gm_n81);
	nand (gm_n3915, in_20, gm_n62, in_18, gm_n3914, in_21);
	nor (gm_n3916, in_9, gm_n64, in_7, gm_n259, in_10);
	nand (gm_n3917, gm_n49, gm_n48, in_11, gm_n3916, in_14);
	nor (gm_n3918, in_17, gm_n46, in_15, gm_n3917, in_18);
	nand (gm_n3919, in_21, gm_n45, gm_n62, gm_n3918);
	nor (gm_n3920, gm_n1970, in_10, gm_n51);
	nand (gm_n3921, in_13, in_12, gm_n53, gm_n3920, in_14);
	nor (gm_n3922, in_17, gm_n46, gm_n63, gm_n3921, in_18);
	nand (gm_n3923, in_21, in_20, in_19, gm_n3922);
	nand (gm_n3924, gm_n64, gm_n55, gm_n82, gm_n757, in_9);
	nor (gm_n3925, in_12, in_11, in_10, gm_n3924, gm_n49);
	nand (gm_n3926, in_16, in_15, in_14, gm_n3925, gm_n81);
	nor (gm_n3927, in_20, gm_n62, gm_n47, gm_n3926, gm_n71);
	nor (gm_n3928, in_12, in_11, in_10, gm_n766, in_13);
	nand (gm_n3929, gm_n46, in_15, gm_n50, gm_n3928, in_17);
	nor (gm_n3930, gm_n45, in_19, gm_n47, gm_n3929, gm_n71);
	or (gm_n3931, in_9, in_8, gm_n55, gm_n84);
	nor (gm_n3932, in_12, gm_n53, gm_n52, gm_n3931, in_13);
	nand (gm_n3933, gm_n46, gm_n63, in_14, gm_n3932, gm_n81);
	nor (gm_n3934, gm_n45, in_19, in_18, gm_n3933, in_21);
	nand (gm_n3935, in_17, gm_n46, gm_n63, gm_n293, gm_n47);
	nor (gm_n3936, in_21, gm_n45, in_19, gm_n3935);
	and (gm_n3937, gm_n52, gm_n51, in_8, gm_n316);
	nand (gm_n3938, in_13, in_12, gm_n53, gm_n3937, gm_n50);
	nor (gm_n3939, in_17, gm_n46, in_15, gm_n3938, gm_n47);
	nand (gm_n3940, gm_n71, gm_n45, gm_n62, gm_n3939);
	nor (gm_n3941, in_8, gm_n55, in_6, gm_n204, gm_n51);
	nand (gm_n3942, in_12, gm_n53, gm_n52, gm_n3941, in_13);
	nor (gm_n3943, gm_n46, in_15, gm_n50, gm_n3942, gm_n81);
	nand (gm_n3944, gm_n45, gm_n62, gm_n47, gm_n3943, in_21);
	nor (gm_n3945, gm_n53, gm_n52, in_9, gm_n1023, gm_n48);
	nand (gm_n3946, gm_n63, in_14, gm_n49, gm_n3945);
	nor (gm_n3947, gm_n47, in_17, in_16, gm_n3946, in_19);
	nand (gm_n3948, gm_n3947, gm_n71, gm_n45);
	nand (gm_n3949, in_7, gm_n82, in_5, gm_n420, gm_n64);
	nor (gm_n3950, gm_n3949, in_9);
	nand (gm_n3951, in_12, gm_n53, in_10, gm_n3950, in_13);
	nor (gm_n3952, in_16, gm_n63, in_14, gm_n3951, gm_n81);
	nand (gm_n3953, in_20, gm_n62, gm_n47, gm_n3952, gm_n71);
	or (gm_n3954, gm_n51, gm_n64, in_7, gm_n279, in_10);
	nor (gm_n3955, gm_n49, gm_n48, in_11, gm_n3954, in_14);
	nand (gm_n3956, gm_n81, in_16, in_15, gm_n3955, gm_n47);
	nor (gm_n3957, gm_n71, gm_n45, gm_n62, gm_n3956);
	or (gm_n3958, gm_n53, gm_n52, gm_n51, gm_n2849, gm_n48);
	nor (gm_n3959, gm_n63, gm_n50, gm_n49, gm_n3958, in_16);
	nand (gm_n3960, in_19, in_18, in_17, gm_n3959, in_20);
	nor (gm_n3961, gm_n3960, gm_n71);
	or (gm_n3962, in_11, in_10, gm_n51, gm_n1098);
	nor (gm_n3963, gm_n50, in_13, in_12, gm_n3962, in_15);
	nand (gm_n3964, gm_n47, gm_n81, gm_n46, gm_n3963, in_19);
	nor (gm_n3965, gm_n3964, in_21, gm_n45);
	nand (gm_n3966, gm_n52, gm_n51, in_8, gm_n57, in_11);
	nor (gm_n3967, in_14, gm_n49, gm_n48, gm_n3966, in_15);
	nand (gm_n3968, in_18, gm_n81, in_16, gm_n3967, in_19);
	nor (gm_n3969, gm_n3968, gm_n71, in_20);
	and (gm_n3970, in_9, gm_n64, in_7, gm_n66, gm_n52);
	nand (gm_n3971, gm_n49, in_12, in_11, gm_n3970, in_14);
	nor (gm_n3972, gm_n81, in_16, in_15, gm_n3971, in_18);
	nand (gm_n3973, in_21, in_20, in_19, gm_n3972);
	nor (gm_n3974, gm_n64, gm_n55, in_6, gm_n1429, gm_n51);
	nand (gm_n3975, in_12, in_11, gm_n52, gm_n3974, in_13);
	nor (gm_n3976, in_16, in_15, in_14, gm_n3975, gm_n81);
	nand (gm_n3977, in_20, in_19, in_18, gm_n3976, gm_n71);
	nor (gm_n3978, in_11, in_10, in_9, gm_n3557, in_12);
	nand (gm_n3979, gm_n63, in_14, in_13, gm_n3978, in_16);
	nor (gm_n3980, in_19, gm_n47, gm_n81, gm_n3979, in_20);
	nand (gm_n3981, gm_n3980, gm_n71);
	nand (gm_n3982, gm_n489, gm_n50, in_13);
	nor (gm_n3983, in_17, in_16, in_15, gm_n3982, in_18);
	nand (gm_n3984, gm_n71, in_20, gm_n62, gm_n3983);
	nand (gm_n3985, in_14, in_13, in_12, gm_n1213, in_15);
	nor (gm_n3986, gm_n47, gm_n81, in_16, gm_n3985, in_19);
	nand (gm_n3987, gm_n3986, gm_n71, gm_n45);
	nand (gm_n3988, gm_n3981, gm_n3977, gm_n3973, gm_n3987, gm_n3984);
	nor (gm_n3989, gm_n3965, gm_n3961, gm_n3957, gm_n3988, gm_n3969);
	nand (gm_n3990, gm_n3948, gm_n3944, gm_n3940, gm_n3989, gm_n3953);
	nor (gm_n3991, gm_n3934, gm_n3930, gm_n3927, gm_n3990, gm_n3936);
	nand (gm_n3992, gm_n3919, gm_n3915, gm_n3912, gm_n3991, gm_n3923);
	nor (gm_n3993, gm_n3903, gm_n3900, gm_n3896, gm_n3992, gm_n3908);
	nand (gm_n3994, gm_n3888, gm_n3883, gm_n3879, gm_n3993, gm_n3892);
	nor (gm_n3995, gm_n3871, gm_n3867, gm_n3864, gm_n3994, gm_n3875);
	nand (gm_n3996, gm_n3855, gm_n3852, gm_n3848, gm_n3995, gm_n3860);
	nor (gm_n3997, gm_n3839, gm_n3836, gm_n3832, gm_n3996, gm_n3843);
	nand (gm_n3998, gm_n3825, gm_n3820, gm_n3816, gm_n3997, gm_n3829);
	nor (gm_n3999, gm_n3808, gm_n3803, gm_n3800, gm_n3998, gm_n3812);
	nand (gm_n4000, gm_n3795, gm_n3792, gm_n3788, gm_n3999, gm_n3798);
	nor (gm_n4001, gm_n3780, gm_n3776, gm_n3772, gm_n4000, gm_n3784);
	nand (gm_n4002, gm_n3763, gm_n3759, gm_n3755, gm_n4001, gm_n3767);
	nor (gm_n4003, gm_n3747, gm_n3742, gm_n3738, gm_n4002, gm_n3751);
	nand (gm_n4004, gm_n3730, gm_n3726, gm_n3722, gm_n4003, gm_n3734);
	nor (gm_n4005, gm_n3715, gm_n3711, gm_n3707, gm_n4004, gm_n3717);
	nand (gm_n4006, gm_n3701, gm_n3696, gm_n3693, gm_n4005, gm_n3704);
	nor (gm_n4007, gm_n3686, gm_n3682, gm_n3680, gm_n4006, gm_n3690);
	nand (gm_n4008, gm_n3673, gm_n3669, gm_n3665, gm_n4007, gm_n3676);
	nor (gm_n4009, gm_n3658, gm_n3654, gm_n3650, gm_n4008, gm_n3662);
	nand (gm_n4010, gm_n3643, gm_n3639, gm_n3636, gm_n4009, gm_n3647);
	nor (gm_n4011, gm_n3627, gm_n3624, gm_n3621, gm_n4010, gm_n3631);
	nand (gm_n4012, gm_n3614, gm_n3610, gm_n3605, gm_n4011, gm_n3618);
	nor (gm_n4013, gm_n3596, gm_n3594, gm_n3591, gm_n4012, gm_n3600);
	nand (gm_n4014, gm_n3583, gm_n3580, gm_n3576, gm_n4013, gm_n3587);
	nor (gm_n4015, gm_n3569, gm_n3565, gm_n3561, gm_n4014, gm_n3572);
	nand (gm_n4016, gm_n3552, gm_n3550, gm_n3546, gm_n4015, gm_n3556);
	nor (gm_n4017, gm_n3537, gm_n3533, gm_n3531, gm_n4016, gm_n3541);
	nand (gm_n4018, gm_n3523, gm_n3518, gm_n3514, gm_n4017, gm_n3527);
	nor (gm_n4019, gm_n3507, gm_n3504, gm_n3500, gm_n4018, gm_n3511);
	nand (gm_n4020, gm_n3493, gm_n3488, gm_n3483, gm_n4019, gm_n3497);
	nor (gm_n4021, gm_n3474, gm_n3470, gm_n3467, gm_n4020, gm_n3479);
	nand (gm_n4022, gm_n3459, gm_n3455, gm_n3450, gm_n4021, gm_n3463);
	nor (gm_n4023, gm_n3442, gm_n3439, gm_n3436, gm_n4022, gm_n3446);
	nand (gm_n4024, gm_n3427, gm_n3423, gm_n3419, gm_n4023, gm_n3432);
	nor (out_5, gm_n4024, gm_n3415);
	nand (gm_n4026, in_8, gm_n55, in_6, gm_n379, in_9);
	nor (gm_n4027, gm_n4026, in_10);
	and (gm_n4028, in_13, gm_n48, in_11, gm_n4027, in_14);
	nand (gm_n4029, gm_n81, gm_n46, in_15, gm_n4028, gm_n47);
	nor (gm_n4030, in_21, in_20, gm_n62, gm_n4029);
	nor (gm_n4031, gm_n53, gm_n52, gm_n51, gm_n2275, in_12);
	nand (gm_n4032, gm_n63, gm_n50, in_13, gm_n4031, in_16);
	nor (gm_n4033, in_19, gm_n47, in_17, gm_n4032, in_20);
	nand (gm_n4034, gm_n4033, gm_n71);
	nand (gm_n4035, in_13, gm_n48, in_11, gm_n3857, gm_n50);
	nor (gm_n4036, gm_n81, gm_n46, in_15, gm_n4035, gm_n47);
	nand (gm_n4037, in_21, gm_n45, gm_n62, gm_n4036);
	and (gm_n4038, in_11, gm_n52, in_9, gm_n3768, in_12);
	nand (gm_n4039, in_15, gm_n50, gm_n49, gm_n4038, gm_n46);
	nor (gm_n4040, in_19, gm_n47, in_17, gm_n4039, gm_n45);
	nand (gm_n4041, gm_n4040, in_21);
	nor (gm_n4042, gm_n55, in_6, gm_n72, gm_n643, in_8);
	and (gm_n4043, gm_n4042, gm_n52, in_9);
	nand (gm_n4044, gm_n49, in_12, in_11, gm_n4043, gm_n50);
	nor (gm_n4045, gm_n81, in_16, in_15, gm_n4044, in_18);
	nand (gm_n4046, in_21, in_20, gm_n62, gm_n4045);
	nor (gm_n4047, in_12, gm_n53, in_10, gm_n3245, gm_n49);
	nand (gm_n4048, gm_n46, in_15, gm_n50, gm_n4047, in_17);
	nor (gm_n4049, gm_n45, gm_n62, in_18, gm_n4048, in_21);
	nor (gm_n4050, in_7, gm_n82, gm_n72, gm_n483, gm_n64);
	and (gm_n4051, in_11, gm_n52, gm_n51, gm_n4050);
	and (gm_n4052, in_14, in_13, gm_n48, gm_n4051, gm_n63);
	nand (gm_n4053, gm_n47, gm_n81, in_16, gm_n4052, in_19);
	nor (gm_n4054, gm_n4053, in_21, in_20);
	and (gm_n4055, in_11, in_10, in_9, gm_n1212, in_12);
	and (gm_n4056, in_15, gm_n50, gm_n49, gm_n4055, in_16);
	nand (gm_n4057, gm_n62, gm_n47, gm_n81, gm_n4056, gm_n45);
	nor (gm_n4058, gm_n4057, in_21);
	nor (gm_n4059, gm_n50, gm_n49, in_12, gm_n1625, in_15);
	nand (gm_n4060, gm_n47, gm_n81, gm_n46, gm_n4059, gm_n62);
	nor (gm_n4061, gm_n4060, gm_n71, in_20);
	nand (gm_n4062, gm_n48, in_11, gm_n52, gm_n1962, in_13);
	nor (gm_n4063, gm_n46, in_15, in_14, gm_n4062, in_17);
	nand (gm_n4064, gm_n45, gm_n62, in_18, gm_n4063, in_21);
	nor (gm_n4065, in_11, in_10, in_9, gm_n131, in_12);
	nand (gm_n4066, gm_n63, gm_n50, in_13, gm_n4065, gm_n46);
	nor (gm_n4067, gm_n62, gm_n47, gm_n81, gm_n4066, gm_n45);
	nand (gm_n4068, gm_n4067, gm_n71);
	nand (gm_n4069, in_12, gm_n53, in_10, gm_n3748, gm_n49);
	nor (gm_n4070, in_16, gm_n63, gm_n50, gm_n4069, in_17);
	nand (gm_n4071, in_20, gm_n62, in_18, gm_n4070, gm_n71);
	nor (gm_n4072, in_8, gm_n55, in_6, gm_n204, in_9);
	nand (gm_n4073, gm_n48, in_11, gm_n52, gm_n4072, gm_n49);
	nor (gm_n4074, gm_n46, in_15, gm_n50, gm_n4073, gm_n81);
	nand (gm_n4075, in_20, gm_n62, gm_n47, gm_n4074, in_21);
	and (gm_n4076, in_12, gm_n53, gm_n52, gm_n946, gm_n49);
	nand (gm_n4077, in_16, in_15, gm_n50, gm_n4076, gm_n81);
	nor (gm_n4078, gm_n45, gm_n62, gm_n47, gm_n4077, in_21);
	nand (gm_n4079, in_7, in_6, gm_n72, gm_n598);
	nor (gm_n4080, in_10, in_9, gm_n64, gm_n4079, gm_n53);
	and (gm_n4081, gm_n50, in_13, in_12, gm_n4080, gm_n63);
	nand (gm_n4082, gm_n47, in_17, gm_n46, gm_n4081, gm_n62);
	nor (gm_n4083, gm_n4082, in_21, in_20);
	nor (gm_n4084, in_12, gm_n53, gm_n52, gm_n3924, in_13);
	nand (gm_n4085, gm_n46, gm_n63, gm_n50, gm_n4084, in_17);
	nor (gm_n4086, gm_n45, gm_n62, in_18, gm_n4085, in_21);
	and (gm_n4087, in_14, gm_n49, in_12, gm_n1604, gm_n63);
	nand (gm_n4088, gm_n47, gm_n81, in_16, gm_n4087, in_19);
	nor (gm_n4089, gm_n4088, in_21, in_20);
	and (gm_n4090, gm_n52, in_9, gm_n64, gm_n1088, gm_n53);
	nand (gm_n4091, gm_n50, gm_n49, gm_n48, gm_n4090);
	nor (gm_n4092, gm_n81, gm_n46, in_15, gm_n4091, in_18);
	nand (gm_n4093, in_21, in_20, in_19, gm_n4092);
	nand (gm_n4094, in_12, gm_n53, gm_n52, gm_n380, gm_n49);
	nor (gm_n4095, in_16, in_15, gm_n50, gm_n4094, in_17);
	nand (gm_n4096, gm_n45, gm_n62, in_18, gm_n4095, in_21);
	nand (gm_n4097, gm_n64, gm_n55, in_6, gm_n379, gm_n51);
	or (gm_n4098, gm_n48, in_11, gm_n52, gm_n4097, in_13);
	nor (gm_n4099, in_16, in_15, in_14, gm_n4098, in_17);
	nand (gm_n4100, gm_n45, in_19, in_18, gm_n4099, in_21);
	nand (gm_n4101, in_12, gm_n53, in_10, gm_n1941, gm_n49);
	nor (gm_n4102, gm_n46, gm_n63, gm_n50, gm_n4101, in_17);
	nand (gm_n4103, gm_n45, in_19, gm_n47, gm_n4102, gm_n71);
	nand (gm_n4104, gm_n2526, gm_n51);
	nor (gm_n4105, in_12, gm_n53, in_10, gm_n4104, in_13);
	nand (gm_n4106, in_16, gm_n63, gm_n50, gm_n4105, in_17);
	nor (gm_n4107, gm_n45, in_19, in_18, gm_n4106, gm_n71);
	nor (gm_n4108, gm_n53, gm_n52, in_9, gm_n1035, in_12);
	and (gm_n4109, gm_n63, gm_n50, gm_n49, gm_n4108, in_16);
	nand (gm_n4110, in_19, in_18, in_17, gm_n4109, gm_n45);
	nor (gm_n4111, gm_n4110, in_21);
	and (gm_n4112, in_14, in_13, gm_n48, gm_n3078, in_15);
	nand (gm_n4113, gm_n47, in_17, gm_n46, gm_n4112, in_19);
	nor (gm_n4114, gm_n4113, in_21, gm_n45);
	or (gm_n4115, in_11, gm_n52, gm_n51, gm_n253, gm_n48);
	nor (gm_n4116, in_15, in_14, gm_n49, gm_n4115, gm_n46);
	nand (gm_n4117, in_19, in_18, in_17, gm_n4116, gm_n45);
	nor (gm_n4118, gm_n4117, gm_n71);
	nor (gm_n4119, in_7, gm_n82, gm_n72, gm_n290, gm_n64);
	and (gm_n4120, gm_n4119, in_10, gm_n51);
	nand (gm_n4121, in_13, gm_n48, gm_n53, gm_n4120, gm_n50);
	nor (gm_n4122, gm_n81, in_16, gm_n63, gm_n4121, in_18);
	nand (gm_n4123, gm_n71, in_20, in_19, gm_n4122);
	nand (gm_n4124, in_12, in_11, gm_n52, gm_n3748, in_13);
	nor (gm_n4125, gm_n46, in_15, in_14, gm_n4124, gm_n81);
	nand (gm_n4126, gm_n45, in_19, gm_n47, gm_n4125, gm_n71);
	and (gm_n4127, gm_n64, in_7, in_6, gm_n1075, gm_n51);
	nand (gm_n4128, in_12, in_11, in_10, gm_n4127, gm_n49);
	nor (gm_n4129, gm_n46, in_15, in_14, gm_n4128, in_17);
	nand (gm_n4130, gm_n45, in_19, in_18, gm_n4129, gm_n71);
	nand (gm_n4131, in_12, gm_n53, in_10, gm_n1719, in_13);
	nor (gm_n4132, in_16, gm_n63, in_14, gm_n4131, gm_n81);
	nand (gm_n4133, gm_n45, gm_n62, in_18, gm_n4132, gm_n71);
	nand (gm_n4134, in_11, gm_n52, in_9, gm_n2653, in_12);
	nor (gm_n4135, in_15, in_14, in_13, gm_n4134, gm_n46);
	nand (gm_n4136, in_19, gm_n47, in_17, gm_n4135, in_20);
	nor (gm_n4137, gm_n4136, gm_n71);
	nand (gm_n4138, in_16, gm_n63, in_14, gm_n981, gm_n81);
	nor (gm_n4139, gm_n45, in_19, in_18, gm_n4138, gm_n71);
	and (gm_n4140, in_12, in_11, in_10, gm_n142, in_13);
	nand (gm_n4141, in_16, gm_n63, in_14, gm_n4140, in_17);
	nor (gm_n4142, in_20, in_19, in_18, gm_n4141, gm_n71);
	and (gm_n4143, gm_n53, in_10, gm_n51, gm_n125, in_12);
	and (gm_n4144, gm_n4143, gm_n49);
	nand (gm_n4145, gm_n46, gm_n63, in_14, gm_n4144, in_17);
	nor (gm_n4146, gm_n45, in_19, gm_n47, gm_n4145, gm_n71);
	nor (gm_n4147, gm_n46, gm_n63, in_14, gm_n2121, in_17);
	nand (gm_n4148, gm_n45, in_19, in_18, gm_n4147, gm_n71);
	and (gm_n4149, in_10, in_9, gm_n64, gm_n338);
	nand (gm_n4150, in_13, in_12, gm_n53, gm_n4149, in_14);
	nor (gm_n4151, gm_n81, gm_n46, gm_n63, gm_n4150, in_18);
	nand (gm_n4152, gm_n71, gm_n45, in_19, gm_n4151);
	nand (gm_n4153, in_7, gm_n82, gm_n72, gm_n493, gm_n64);
	nor (gm_n4154, gm_n53, gm_n52, in_9, gm_n4153);
	nand (gm_n4155, in_14, gm_n49, gm_n48, gm_n4154, gm_n63);
	nor (gm_n4156, gm_n47, in_17, gm_n46, gm_n4155, in_19);
	nand (gm_n4157, gm_n4156, in_21, gm_n45);
	nand (gm_n4158, in_12, in_11, in_10, gm_n544, in_13);
	nor (gm_n4159, gm_n46, gm_n63, in_14, gm_n4158, in_17);
	nand (gm_n4160, in_20, in_19, gm_n47, gm_n4159, gm_n71);
	nand (gm_n4161, in_11, in_10, in_9, gm_n3091, gm_n48);
	nor (gm_n4162, gm_n63, in_14, in_13, gm_n4161, gm_n46);
	nand (gm_n4163, gm_n62, gm_n47, gm_n81, gm_n4162, in_20);
	nor (gm_n4164, gm_n4163, in_21);
	nor (gm_n4165, in_14, in_13, gm_n48, gm_n3092, gm_n63);
	nand (gm_n4166, in_18, in_17, in_16, gm_n4165, gm_n62);
	nor (gm_n4167, gm_n4166, gm_n71, in_20);
	nor (gm_n4168, in_7, in_6, in_5, gm_n124, in_8);
	nand (gm_n4169, gm_n4168, gm_n51);
	nor (gm_n4170, in_12, in_11, in_10, gm_n4169, gm_n49);
	nand (gm_n4171, in_16, gm_n63, in_14, gm_n4170, in_17);
	nor (gm_n4172, in_20, gm_n62, in_18, gm_n4171, gm_n71);
	or (gm_n4173, in_11, in_10, in_9, gm_n1464, gm_n48);
	nor (gm_n4174, gm_n63, in_14, in_13, gm_n4173, gm_n46);
	nand (gm_n4175, gm_n62, gm_n47, in_17, gm_n4174, gm_n45);
	nor (gm_n4176, gm_n4175, in_21);
	nand (gm_n4177, gm_n55, gm_n82, gm_n72, gm_n327, gm_n64);
	nor (gm_n4178, in_11, in_10, gm_n51, gm_n4177, in_12);
	nand (gm_n4179, in_15, in_14, in_13, gm_n4178, in_16);
	nor (gm_n4180, gm_n62, in_18, in_17, gm_n4179, gm_n45);
	nand (gm_n4181, gm_n4180, gm_n71);
	nand (gm_n4182, gm_n48, gm_n53, in_10, gm_n968, gm_n49);
	nor (gm_n4183, gm_n46, in_15, gm_n50, gm_n4182, gm_n81);
	nand (gm_n4184, gm_n45, gm_n62, gm_n47, gm_n4183, gm_n71);
	nand (gm_n4185, in_12, gm_n53, gm_n52, gm_n1170, gm_n49);
	nor (gm_n4186, in_16, gm_n63, in_14, gm_n4185, gm_n81);
	nand (gm_n4187, gm_n45, gm_n62, in_18, gm_n4186, in_21);
	or (gm_n4188, in_13, in_12, in_11, gm_n1844, in_14);
	nor (gm_n4189, gm_n81, gm_n46, gm_n63, gm_n4188, in_18);
	nand (gm_n4190, in_21, in_20, in_19, gm_n4189);
	nand (gm_n4191, in_11, gm_n52, in_9, gm_n997, in_12);
	nor (gm_n4192, in_15, gm_n50, in_13, gm_n4191, in_16);
	nand (gm_n4193, gm_n62, in_18, in_17, gm_n4192, in_20);
	nor (gm_n4194, gm_n4193, gm_n71);
	nand (gm_n4195, gm_n64, gm_n55, gm_n82, gm_n2640, gm_n51);
	nor (gm_n4196, gm_n4195, in_11, gm_n52);
	and (gm_n4197, in_14, gm_n49, gm_n48, gm_n4196, in_15);
	nand (gm_n4198, gm_n47, in_17, gm_n46, gm_n4197, in_19);
	nor (gm_n4199, gm_n4198, gm_n71, in_20);
	nor (gm_n4200, in_7, in_6, gm_n72, gm_n167, gm_n64);
	nand (gm_n4201, gm_n53, in_10, in_9, gm_n4200, gm_n48);
	nor (gm_n4202, gm_n63, gm_n50, gm_n49, gm_n4201, in_16);
	nand (gm_n4203, gm_n62, in_18, in_17, gm_n4202, gm_n45);
	nor (gm_n4204, gm_n4203, in_21);
	or (gm_n4205, gm_n51, in_8, gm_n55, gm_n1256);
	nor (gm_n4206, gm_n48, in_11, gm_n52, gm_n4205, in_13);
	nand (gm_n4207, gm_n46, gm_n63, in_14, gm_n4206, gm_n81);
	nor (gm_n4208, in_20, in_19, gm_n47, gm_n4207, in_21);
	nor (gm_n4209, gm_n2951, gm_n52, gm_n51);
	nand (gm_n4210, in_13, gm_n48, in_11, gm_n4209);
	nor (gm_n4211, gm_n46, in_15, in_14, gm_n4210, in_17);
	nand (gm_n4212, gm_n45, in_19, gm_n47, gm_n4211, gm_n71);
	nor (gm_n4213, gm_n55, in_6, in_5, gm_n124);
	and (gm_n4214, gm_n52, gm_n51, gm_n64, gm_n4213, gm_n53);
	nand (gm_n4215, gm_n50, in_13, in_12, gm_n4214, in_15);
	nor (gm_n4216, gm_n47, gm_n81, in_16, gm_n4215, in_19);
	nand (gm_n4217, gm_n4216, in_21, in_20);
	nand (gm_n4218, in_14, gm_n49, gm_n48, gm_n3640, gm_n63);
	nor (gm_n4219, in_18, gm_n81, gm_n46, gm_n4218, in_19);
	nand (gm_n4220, gm_n4219, in_21, in_20);
	nand (gm_n4221, gm_n50, in_13, gm_n48, gm_n1751, gm_n63);
	nor (gm_n4222, in_18, gm_n81, in_16, gm_n4221, gm_n62);
	nand (gm_n4223, gm_n4222, gm_n71, in_20);
	nor (gm_n4224, gm_n48, in_11, in_10, gm_n4205, in_13);
	nand (gm_n4225, in_16, gm_n63, in_14, gm_n4224, in_17);
	nor (gm_n4226, in_20, gm_n62, in_18, gm_n4225, in_21);
	nor (gm_n4227, in_13, gm_n48, in_11, gm_n2296, in_14);
	nand (gm_n4228, in_17, gm_n46, gm_n63, gm_n4227, in_18);
	nor (gm_n4229, in_21, gm_n45, gm_n62, gm_n4228);
	and (gm_n4230, gm_n48, gm_n53, gm_n52, gm_n1962, gm_n49);
	nand (gm_n4231, gm_n46, in_15, in_14, gm_n4230, gm_n81);
	nor (gm_n4232, in_20, in_19, gm_n47, gm_n4231, in_21);
	nand (gm_n4233, gm_n52, gm_n51, in_8, gm_n302, gm_n53);
	nor (gm_n4234, gm_n50, in_13, in_12, gm_n4233, gm_n63);
	nand (gm_n4235, in_18, gm_n81, gm_n46, gm_n4234, in_19);
	nor (gm_n4236, gm_n4235, in_21, gm_n45);
	nor (gm_n4237, gm_n49, gm_n48, in_11, gm_n2700, in_14);
	and (gm_n4238, gm_n81, in_16, in_15, gm_n4237, gm_n47);
	nand (gm_n4239, gm_n71, in_20, gm_n62, gm_n4238);
	nand (gm_n4240, gm_n49, in_12, in_11, gm_n881, gm_n50);
	nor (gm_n4241, in_17, gm_n46, gm_n63, gm_n4240, in_18);
	nand (gm_n4242, gm_n71, gm_n45, in_19, gm_n4241);
	nor (gm_n4243, in_11, gm_n52, gm_n51, gm_n322, gm_n48);
	nand (gm_n4244, gm_n63, in_14, in_13, gm_n4243, in_16);
	nor (gm_n4245, gm_n62, in_18, gm_n81, gm_n4244, in_20);
	nand (gm_n4246, gm_n4245, in_21);
	nand (gm_n4247, gm_n48, gm_n53, in_10, gm_n2672, in_13);
	nor (gm_n4248, in_16, gm_n63, gm_n50, gm_n4247, gm_n81);
	nand (gm_n4249, gm_n45, in_19, gm_n47, gm_n4248, gm_n71);
	or (gm_n4250, gm_n53, in_10, in_9, gm_n1709, in_12);
	nor (gm_n4251, in_15, in_14, in_13, gm_n4250, gm_n46);
	nand (gm_n4252, gm_n62, in_18, gm_n81, gm_n4251, gm_n45);
	nor (gm_n4253, gm_n4252, gm_n71);
	nand (gm_n4254, gm_n53, in_10, gm_n51, gm_n484, in_12);
	nor (gm_n4255, in_15, gm_n50, in_13, gm_n4254, in_16);
	nand (gm_n4256, gm_n62, gm_n47, gm_n81, gm_n4255, gm_n45);
	nor (gm_n4257, gm_n4256, in_21);
	nand (gm_n4258, gm_n53, gm_n52, gm_n51, gm_n3193);
	nor (gm_n4259, in_14, in_13, gm_n48, gm_n4258, in_15);
	nand (gm_n4260, gm_n47, gm_n81, gm_n46, gm_n4259, gm_n62);
	nor (gm_n4261, gm_n4260, gm_n71, in_20);
	or (gm_n4262, gm_n64, gm_n55, gm_n82, gm_n530, in_9);
	nor (gm_n4263, gm_n48, in_11, in_10, gm_n4262, in_13);
	nand (gm_n4264, gm_n46, in_15, in_14, gm_n4263, in_17);
	nor (gm_n4265, in_20, in_19, gm_n47, gm_n4264, gm_n71);
	and (gm_n4266, in_8, gm_n55, gm_n82, gm_n638, gm_n51);
	nand (gm_n4267, in_12, in_11, gm_n52, gm_n4266, gm_n49);
	nor (gm_n4268, in_16, gm_n63, in_14, gm_n4267, in_17);
	nand (gm_n4269, gm_n45, in_19, in_18, gm_n4268, in_21);
	nand (gm_n4270, gm_n63, in_14, in_13, gm_n1727, in_16);
	nor (gm_n4271, in_19, gm_n47, in_17, gm_n4270, gm_n45);
	nand (gm_n4272, gm_n4271, gm_n71);
	and (gm_n4273, gm_n55, in_6, gm_n72, gm_n241, in_8);
	and (gm_n4274, in_11, in_10, in_9, gm_n4273, gm_n48);
	nand (gm_n4275, gm_n63, gm_n50, in_13, gm_n4274, in_16);
	nor (gm_n4276, in_19, gm_n47, in_17, gm_n4275, gm_n45);
	nand (gm_n4277, gm_n4276, in_21);
	nand (gm_n4278, gm_n53, gm_n52, in_9, gm_n2631, gm_n48);
	nor (gm_n4279, gm_n4278, in_13);
	and (gm_n4280, gm_n46, in_15, gm_n50, gm_n4279, gm_n81);
	nand (gm_n4281, gm_n45, in_19, in_18, gm_n4280, gm_n71);
	nor (gm_n4282, gm_n48, gm_n53, in_10, gm_n2597, in_13);
	nand (gm_n4283, in_16, gm_n63, in_14, gm_n4282, gm_n81);
	nor (gm_n4284, gm_n45, in_19, in_18, gm_n4283, in_21);
	nor (gm_n4285, gm_n55, in_6, in_5, gm_n75, gm_n64);
	nand (gm_n4286, in_11, gm_n52, gm_n51, gm_n4285, gm_n48);
	nor (gm_n4287, gm_n63, gm_n50, in_13, gm_n4286, gm_n46);
	nand (gm_n4288, in_19, gm_n47, in_17, gm_n4287, in_20);
	nor (gm_n4289, gm_n4288, in_21);
	nor (gm_n4290, in_15, in_14, in_13, gm_n2606, gm_n46);
	nand (gm_n4291, in_19, in_18, gm_n81, gm_n4290, in_20);
	nor (gm_n4292, gm_n4291, in_21);
	nor (gm_n4293, gm_n55, in_6, in_5, gm_n188, in_8);
	nand (gm_n4294, gm_n4293, in_9);
	nor (gm_n4295, in_12, gm_n53, gm_n52, gm_n4294, gm_n49);
	nand (gm_n4296, gm_n46, in_15, in_14, gm_n4295, in_17);
	nor (gm_n4297, gm_n45, in_19, gm_n47, gm_n4296, gm_n71);
	and (gm_n4298, in_11, in_10, in_9, gm_n1459);
	nand (gm_n4299, in_14, in_13, in_12, gm_n4298, gm_n63);
	nor (gm_n4300, in_18, in_17, gm_n46, gm_n4299, gm_n62);
	nand (gm_n4301, gm_n4300, gm_n71, in_20);
	nor (gm_n4302, in_11, gm_n52, in_9, gm_n2345, in_12);
	nand (gm_n4303, gm_n63, gm_n50, gm_n49, gm_n4302, in_16);
	nor (gm_n4304, in_19, gm_n47, in_17, gm_n4303, gm_n45);
	nand (gm_n4305, gm_n4304, in_21);
	nand (gm_n4306, gm_n53, in_10, in_9, gm_n1555, gm_n48);
	nor (gm_n4307, gm_n4306, in_13);
	and (gm_n4308, in_16, gm_n63, in_14, gm_n4307, gm_n81);
	nand (gm_n4309, gm_n45, gm_n62, gm_n47, gm_n4308, gm_n71);
	and (gm_n4310, gm_n1274, in_10, in_9);
	nand (gm_n4311, gm_n49, gm_n48, in_11, gm_n4310, in_14);
	nor (gm_n4312, gm_n81, in_16, in_15, gm_n4311, in_18);
	nand (gm_n4313, in_21, gm_n45, gm_n62, gm_n4312);
	nand (gm_n4314, gm_n55, in_6, in_5, gm_n598, gm_n64);
	nor (gm_n4315, in_11, in_10, gm_n51, gm_n4314);
	and (gm_n4316, gm_n4315, gm_n49, gm_n48);
	nand (gm_n4317, in_16, in_15, in_14, gm_n4316, in_17);
	nor (gm_n4318, in_20, gm_n62, in_18, gm_n4317, in_21);
	nor (gm_n4319, in_8, gm_n55, in_6, gm_n96, in_9);
	and (gm_n4320, in_12, in_11, in_10, gm_n4319, gm_n49);
	nand (gm_n4321, gm_n46, gm_n63, gm_n50, gm_n4320, gm_n81);
	nor (gm_n4322, in_20, in_19, in_18, gm_n4321, gm_n71);
	nand (gm_n4323, in_16, in_15, gm_n50, gm_n1574, gm_n81);
	nor (gm_n4324, in_20, gm_n62, gm_n47, gm_n4323, in_21);
	nand (gm_n4325, gm_n1165, gm_n52, gm_n51);
	nor (gm_n4326, gm_n49, gm_n48, in_11, gm_n4325, in_14);
	nand (gm_n4327, in_17, in_16, in_15, gm_n4326, gm_n47);
	nor (gm_n4328, gm_n71, in_20, gm_n62, gm_n4327);
	nor (gm_n4329, gm_n64, in_7, in_6, gm_n204, gm_n51);
	nand (gm_n4330, gm_n48, gm_n53, in_10, gm_n4329, in_13);
	nor (gm_n4331, gm_n46, in_15, in_14, gm_n4330, in_17);
	nand (gm_n4332, gm_n45, gm_n62, gm_n47, gm_n4331, in_21);
	and (gm_n4333, in_17, gm_n46, gm_n63, gm_n2971, in_18);
	nand (gm_n4334, in_21, in_20, in_19, gm_n4333);
	nand (gm_n4335, in_12, gm_n53, in_10, gm_n4072, in_13);
	nor (gm_n4336, gm_n46, gm_n63, in_14, gm_n4335, in_17);
	nand (gm_n4337, in_20, in_19, gm_n47, gm_n4336, gm_n71);
	nand (gm_n4338, in_14, gm_n49, gm_n48, gm_n4080, gm_n63);
	nor (gm_n4339, in_18, gm_n81, gm_n46, gm_n4338, gm_n62);
	nand (gm_n4340, gm_n4339, in_21, gm_n45);
	nor (gm_n4341, gm_n49, in_12, gm_n53, gm_n3893, gm_n50);
	nand (gm_n4342, in_17, gm_n46, gm_n63, gm_n4341, in_18);
	nor (gm_n4343, in_21, gm_n45, gm_n62, gm_n4342);
	nor (gm_n4344, gm_n48, in_11, in_10, gm_n228, gm_n49);
	nand (gm_n4345, in_16, gm_n63, in_14, gm_n4344, in_17);
	nor (gm_n4346, in_20, gm_n62, gm_n47, gm_n4345, gm_n71);
	or (gm_n4347, in_9, gm_n64, gm_n55, gm_n588, gm_n52);
	nor (gm_n4348, gm_n49, gm_n48, in_11, gm_n4347, gm_n50);
	nand (gm_n4349, in_17, gm_n46, in_15, gm_n4348, in_18);
	nor (gm_n4350, gm_n71, in_20, gm_n62, gm_n4349);
	or (gm_n4351, gm_n51, in_8, in_7, gm_n84, in_10);
	nor (gm_n4352, in_13, in_12, in_11, gm_n4351, in_14);
	nand (gm_n4353, in_17, gm_n46, in_15, gm_n4352, gm_n47);
	nor (gm_n4354, in_21, gm_n45, gm_n62, gm_n4353);
	and (gm_n4355, gm_n2424, gm_n49);
	and (gm_n4356, in_16, in_15, in_14, gm_n4355, in_17);
	nand (gm_n4357, gm_n45, gm_n62, in_18, gm_n4356, in_21);
	and (gm_n4358, gm_n51, gm_n64, in_7, gm_n404, in_10);
	nand (gm_n4359, in_13, in_12, in_11, gm_n4358, in_14);
	nor (gm_n4360, in_17, in_16, gm_n63, gm_n4359, gm_n47);
	nand (gm_n4361, gm_n71, in_20, in_19, gm_n4360);
	or (gm_n4362, in_8, gm_n55, gm_n82, gm_n1429, gm_n51);
	or (gm_n4363, in_12, gm_n53, in_10, gm_n4362, gm_n49);
	nor (gm_n4364, gm_n46, gm_n63, gm_n50, gm_n4363, gm_n81);
	nand (gm_n4365, gm_n45, in_19, in_18, gm_n4364, gm_n71);
	or (gm_n4366, in_8, in_7, gm_n82, gm_n199, in_9);
	or (gm_n4367, gm_n48, gm_n53, gm_n52, gm_n4366, in_13);
	nor (gm_n4368, in_16, in_15, gm_n50, gm_n4367, in_17);
	nand (gm_n4369, gm_n45, in_19, gm_n47, gm_n4368, gm_n71);
	nor (gm_n4370, gm_n53, in_10, gm_n51, gm_n1127);
	and (gm_n4371, gm_n50, in_13, in_12, gm_n4370, gm_n63);
	nand (gm_n4372, in_18, in_17, in_16, gm_n4371, in_19);
	nor (gm_n4373, gm_n4372, in_21, in_20);
	and (gm_n4374, in_12, gm_n53, gm_n52, gm_n3950, gm_n49);
	nand (gm_n4375, gm_n46, gm_n63, in_14, gm_n4374, gm_n81);
	nor (gm_n4376, in_20, in_19, in_18, gm_n4375, gm_n71);
	nor (gm_n4377, gm_n53, gm_n52, gm_n51, gm_n3146);
	and (gm_n4378, gm_n50, in_13, gm_n48, gm_n4377, gm_n63);
	nand (gm_n4379, gm_n47, in_17, in_16, gm_n4378, gm_n62);
	nor (gm_n4380, gm_n4379, gm_n71, gm_n45);
	nand (gm_n4381, gm_n4200, gm_n51);
	nor (gm_n4382, in_12, in_11, in_10, gm_n4381, gm_n49);
	nand (gm_n4383, gm_n46, in_15, in_14, gm_n4382, in_17);
	nor (gm_n4384, in_20, gm_n62, in_18, gm_n4383, gm_n71);
	nand (gm_n4385, gm_n49, in_12, gm_n53, gm_n500, in_14);
	nor (gm_n4386, in_17, gm_n46, gm_n63, gm_n4385, gm_n47);
	nand (gm_n4387, gm_n71, in_20, in_19, gm_n4386);
	nor (gm_n4388, in_7, gm_n82, in_5, gm_n75, in_8);
	and (gm_n4389, gm_n53, in_10, in_9, gm_n4388, in_12);
	nand (gm_n4390, gm_n63, gm_n50, in_13, gm_n4389, in_16);
	nor (gm_n4391, in_19, gm_n47, in_17, gm_n4390, in_20);
	nand (gm_n4392, gm_n4391, in_21);
	nand (gm_n4393, in_7, gm_n82, in_5, gm_n1126, gm_n64);
	nor (gm_n4394, in_11, gm_n52, gm_n51, gm_n4393, gm_n48);
	nand (gm_n4395, in_15, gm_n50, gm_n49, gm_n4394, in_16);
	nor (gm_n4396, gm_n62, in_18, in_17, gm_n4395, in_20);
	nand (gm_n4397, gm_n4396, in_21);
	or (gm_n4398, in_9, gm_n64, in_7, gm_n259, gm_n52);
	nor (gm_n4399, in_13, in_12, in_11, gm_n4398, in_14);
	and (gm_n4400, in_17, in_16, gm_n63, gm_n4399, in_18);
	nand (gm_n4401, gm_n71, in_20, gm_n62, gm_n4400);
	nand (gm_n4402, in_11, in_10, gm_n51, gm_n2432);
	nor (gm_n4403, gm_n50, in_13, in_12, gm_n4402, in_15);
	nand (gm_n4404, gm_n47, gm_n81, gm_n46, gm_n4403, in_19);
	nor (gm_n4405, gm_n4404, gm_n71, gm_n45);
	nand (gm_n4406, in_11, in_10, in_9, gm_n2508, in_12);
	nor (gm_n4407, gm_n63, gm_n50, in_13, gm_n4406, in_16);
	nand (gm_n4408, gm_n62, gm_n47, in_17, gm_n4407, in_20);
	nor (gm_n4409, gm_n4408, in_21);
	nand (gm_n4410, in_10, gm_n51, gm_n64, gm_n1088);
	nor (gm_n4411, in_13, gm_n48, gm_n53, gm_n4410, in_14);
	nand (gm_n4412, in_17, gm_n46, in_15, gm_n4411, gm_n47);
	nor (gm_n4413, gm_n71, in_20, in_19, gm_n4412);
	or (gm_n4414, gm_n415, gm_n52, gm_n51);
	nor (gm_n4415, in_13, gm_n48, in_11, gm_n4414, in_14);
	nand (gm_n4416, gm_n81, gm_n46, gm_n63, gm_n4415, gm_n47);
	nor (gm_n4417, gm_n71, gm_n45, gm_n62, gm_n4416);
	nor (gm_n4418, gm_n64, in_7, in_6, gm_n199, in_9);
	nand (gm_n4419, gm_n48, gm_n53, gm_n52, gm_n4418, gm_n49);
	nor (gm_n4420, gm_n46, in_15, gm_n50, gm_n4419, gm_n81);
	nand (gm_n4421, gm_n45, gm_n62, in_18, gm_n4420, gm_n71);
	nand (gm_n4422, in_12, in_11, gm_n52, gm_n912, gm_n49);
	nor (gm_n4423, gm_n46, in_15, gm_n50, gm_n4422, gm_n81);
	nand (gm_n4424, gm_n45, in_19, gm_n47, gm_n4423, gm_n71);
	nand (gm_n4425, in_13, gm_n48, in_11, gm_n3651, gm_n50);
	nor (gm_n4426, gm_n81, in_16, gm_n63, gm_n4425, in_18);
	nand (gm_n4427, in_21, in_20, gm_n62, gm_n4426);
	nor (gm_n4428, gm_n53, in_10, gm_n51, gm_n2300, in_12);
	nand (gm_n4429, gm_n63, gm_n50, in_13, gm_n4428, gm_n46);
	nor (gm_n4430, gm_n62, gm_n47, gm_n81, gm_n4429, in_20);
	nand (gm_n4431, gm_n4430, gm_n71);
	nand (gm_n4432, gm_n51, gm_n64, gm_n55, gm_n404, in_10);
	nor (gm_n4433, in_13, gm_n48, gm_n53, gm_n4432, in_14);
	nand (gm_n4434, in_17, gm_n46, gm_n63, gm_n4433, in_18);
	nor (gm_n4435, in_21, in_20, gm_n62, gm_n4434);
	nor (gm_n4436, gm_n53, in_10, in_9, gm_n2445, gm_n48);
	and (gm_n4437, in_15, in_14, in_13, gm_n4436, in_16);
	nand (gm_n4438, gm_n62, in_18, gm_n81, gm_n4437, in_20);
	nor (gm_n4439, gm_n4438, gm_n71);
	and (gm_n4440, in_12, in_11, gm_n52, gm_n3163, in_13);
	nand (gm_n4441, in_16, in_15, gm_n50, gm_n4440, in_17);
	nor (gm_n4442, in_20, gm_n62, in_18, gm_n4441, gm_n71);
	nand (gm_n4443, gm_n53, in_10, in_9, gm_n1147, gm_n48);
	nor (gm_n4444, in_15, in_14, gm_n49, gm_n4443, in_16);
	nand (gm_n4445, in_19, gm_n47, in_17, gm_n4444, in_20);
	nor (gm_n4446, gm_n4445, gm_n71);
	nor (gm_n4447, gm_n2345, in_10, gm_n51);
	nand (gm_n4448, in_13, in_12, gm_n53, gm_n4447, gm_n50);
	nor (gm_n4449, in_17, gm_n46, in_15, gm_n4448, in_18);
	nand (gm_n4450, in_21, in_20, gm_n62, gm_n4449);
	nor (gm_n4451, gm_n52, gm_n51, gm_n64, gm_n390, gm_n53);
	nand (gm_n4452, in_14, gm_n49, gm_n48, gm_n4451, in_15);
	nor (gm_n4453, gm_n47, gm_n81, gm_n46, gm_n4452, gm_n62);
	nand (gm_n4454, gm_n4453, gm_n71, in_20);
	nand (gm_n4455, gm_n50, in_13, gm_n48, gm_n2850, gm_n63);
	nor (gm_n4456, gm_n47, gm_n81, gm_n46, gm_n4455, in_19);
	nand (gm_n4457, gm_n4456, gm_n71, in_20);
	nand (gm_n4458, in_13, in_12, in_11, gm_n4149, in_14);
	nor (gm_n4459, gm_n81, in_16, gm_n63, gm_n4458, gm_n47);
	nand (gm_n4460, gm_n71, in_20, in_19, gm_n4459);
	and (gm_n4461, gm_n50, gm_n49, in_12, gm_n485, in_15);
	nand (gm_n4462, in_18, in_17, in_16, gm_n4461, gm_n62);
	nor (gm_n4463, gm_n4462, in_21, in_20);
	nand (gm_n4464, in_11, in_10, gm_n51, gm_n4042, in_12);
	nor (gm_n4465, in_15, gm_n50, in_13, gm_n4464, gm_n46);
	nand (gm_n4466, in_19, gm_n47, in_17, gm_n4465, in_20);
	nor (gm_n4467, gm_n4466, gm_n71);
	nor (gm_n4468, gm_n63, in_14, in_13, gm_n515, in_16);
	nand (gm_n4469, gm_n62, gm_n47, gm_n81, gm_n4468, gm_n45);
	nor (gm_n4470, gm_n4469, gm_n71);
	or (gm_n4471, gm_n52, gm_n51, gm_n64, gm_n3718, in_11);
	nor (gm_n4472, in_14, in_13, in_12, gm_n4471, in_15);
	nand (gm_n4473, gm_n47, gm_n81, in_16, gm_n4472, gm_n62);
	nor (gm_n4474, gm_n4473, gm_n71, gm_n45);
	or (gm_n4475, gm_n52, gm_n51, in_8, gm_n907, in_11);
	nor (gm_n4476, gm_n4475, in_13, in_12);
	and (gm_n4477, in_16, in_15, in_14, gm_n4476, in_17);
	nand (gm_n4478, in_20, in_19, gm_n47, gm_n4477, in_21);
	and (gm_n4479, gm_n81, gm_n46, gm_n63, gm_n1813, in_18);
	nand (gm_n4480, gm_n71, in_20, gm_n62, gm_n4479);
	nand (gm_n4481, in_13, gm_n48, gm_n53, gm_n3708, gm_n50);
	nor (gm_n4482, in_17, in_16, gm_n63, gm_n4481, in_18);
	nand (gm_n4483, in_21, in_20, in_19, gm_n4482);
	and (gm_n4484, in_7, gm_n82, gm_n72, gm_n241, in_8);
	and (gm_n4485, gm_n53, in_10, in_9, gm_n4484);
	nand (gm_n4486, in_14, in_13, in_12, gm_n4485, in_15);
	nor (gm_n4487, in_18, gm_n81, gm_n46, gm_n4486, in_19);
	nand (gm_n4488, gm_n4487, in_21, gm_n45);
	nand (gm_n4489, gm_n55, gm_n82, gm_n72, gm_n209, in_8);
	or (gm_n4490, gm_n53, gm_n52, in_9, gm_n4489, in_12);
	nor (gm_n4491, in_15, gm_n50, in_13, gm_n4490, gm_n46);
	nand (gm_n4492, gm_n62, in_18, gm_n81, gm_n4491, in_20);
	nor (gm_n4493, gm_n4492, in_21);
	or (gm_n4494, gm_n53, in_10, gm_n51, gm_n3557);
	nor (gm_n4495, gm_n50, in_13, in_12, gm_n4494, gm_n63);
	nand (gm_n4496, gm_n47, in_17, gm_n46, gm_n4495, gm_n62);
	nor (gm_n4497, gm_n4496, in_21, in_20);
	nor (gm_n4498, in_12, gm_n53, gm_n52, gm_n228, in_13);
	nand (gm_n4499, gm_n46, in_15, in_14, gm_n4498, gm_n81);
	nor (gm_n4500, gm_n45, gm_n62, in_18, gm_n4499, in_21);
	nand (gm_n4501, gm_n53, in_10, in_9, gm_n3606, in_12);
	nor (gm_n4502, gm_n4501, in_13);
	nand (gm_n4503, in_16, in_15, gm_n50, gm_n4502, gm_n81);
	nor (gm_n4504, in_20, gm_n62, in_18, gm_n4503, in_21);
	nand (gm_n4505, in_12, in_11, gm_n52, gm_n1385, gm_n49);
	nor (gm_n4506, in_16, gm_n63, in_14, gm_n4505, in_17);
	nand (gm_n4507, gm_n45, in_19, in_18, gm_n4506, gm_n71);
	and (gm_n4508, in_13, in_12, gm_n53, gm_n526, gm_n50);
	and (gm_n4509, gm_n81, gm_n46, gm_n63, gm_n4508, in_18);
	nand (gm_n4510, gm_n71, in_20, gm_n62, gm_n4509);
	nand (gm_n4511, in_12, gm_n53, in_10, gm_n1332, gm_n49);
	nor (gm_n4512, gm_n46, in_15, in_14, gm_n4511, in_17);
	nand (gm_n4513, in_20, in_19, in_18, gm_n4512, gm_n71);
	nand (gm_n4514, in_7, in_6, in_5, gm_n241);
	nor (gm_n4515, in_10, in_9, gm_n64, gm_n4514);
	nand (gm_n4516, in_13, gm_n48, gm_n53, gm_n4515, gm_n50);
	nor (gm_n4517, in_17, gm_n46, gm_n63, gm_n4516, gm_n47);
	nand (gm_n4518, in_21, gm_n45, in_19, gm_n4517);
	and (gm_n4519, gm_n48, gm_n53, in_10, gm_n1932, gm_n49);
	nand (gm_n4520, in_16, in_15, gm_n50, gm_n4519, in_17);
	nor (gm_n4521, in_20, in_19, in_18, gm_n4520, gm_n71);
	nor (gm_n4522, gm_n4471, gm_n49, gm_n48);
	nand (gm_n4523, gm_n46, gm_n63, gm_n50, gm_n4522, gm_n81);
	nor (gm_n4524, in_20, in_19, in_18, gm_n4523, gm_n71);
	nor (gm_n4525, in_7, gm_n82, in_5, gm_n321, in_8);
	nand (gm_n4526, in_11, gm_n52, in_9, gm_n4525, in_12);
	nor (gm_n4527, in_15, in_14, gm_n49, gm_n4526, in_16);
	nand (gm_n4528, in_19, in_18, gm_n81, gm_n4527, in_20);
	nor (gm_n4529, gm_n4528, in_21);
	nand (gm_n4530, gm_n4213, gm_n51, gm_n64);
	nor (gm_n4531, in_12, gm_n53, gm_n52, gm_n4530, gm_n49);
	nand (gm_n4532, in_16, gm_n63, gm_n50, gm_n4531, in_17);
	nor (gm_n4533, gm_n45, in_19, gm_n47, gm_n4532, gm_n71);
	or (gm_n4534, gm_n48, in_11, in_10, gm_n2327, gm_n49);
	nor (gm_n4535, in_16, gm_n63, in_14, gm_n4534, in_17);
	nand (gm_n4536, in_20, gm_n62, gm_n47, gm_n4535, in_21);
	or (gm_n4537, in_12, gm_n53, gm_n52, gm_n4366, in_13);
	nor (gm_n4538, gm_n46, in_15, gm_n50, gm_n4537, in_17);
	nand (gm_n4539, in_20, in_19, in_18, gm_n4538, in_21);
	nand (gm_n4540, gm_n48, in_11, in_10, gm_n4266, gm_n49);
	nor (gm_n4541, gm_n46, gm_n63, gm_n50, gm_n4540, gm_n81);
	nand (gm_n4542, gm_n45, gm_n62, in_18, gm_n4541, in_21);
	nor (gm_n4543, in_11, gm_n52, in_9, gm_n520, in_12);
	nand (gm_n4544, in_15, in_14, gm_n49, gm_n4543, in_16);
	nor (gm_n4545, in_19, in_18, gm_n81, gm_n4544, in_20);
	nand (gm_n4546, gm_n4545, in_21);
	nand (gm_n4547, gm_n189, gm_n51);
	nor (gm_n4548, in_12, in_11, gm_n52, gm_n4547, in_13);
	nand (gm_n4549, in_16, in_15, in_14, gm_n4548, gm_n81);
	nor (gm_n4550, gm_n45, in_19, in_18, gm_n4549, gm_n71);
	nor (gm_n4551, gm_n48, in_11, gm_n52, gm_n1621, in_13);
	nand (gm_n4552, in_16, gm_n63, gm_n50, gm_n4551, gm_n81);
	nor (gm_n4553, in_20, in_19, in_18, gm_n4552, gm_n71);
	or (gm_n4554, in_8, in_7, in_6, gm_n1429, in_9);
	nor (gm_n4555, gm_n48, gm_n53, in_10, gm_n4554, gm_n49);
	nand (gm_n4556, gm_n46, in_15, gm_n50, gm_n4555, in_17);
	nor (gm_n4557, in_20, gm_n62, gm_n47, gm_n4556, in_21);
	nand (gm_n4558, gm_n53, gm_n52, in_9, gm_n1360, in_12);
	nor (gm_n4559, in_15, gm_n50, in_13, gm_n4558);
	nand (gm_n4560, in_18, in_17, in_16, gm_n4559, gm_n62);
	nor (gm_n4561, gm_n4560, in_21, in_20);
	nand (gm_n4562, in_7, in_6, gm_n72, gm_n284, in_8);
	nor (gm_n4563, gm_n53, in_10, in_9, gm_n4562, gm_n48);
	nand (gm_n4564, gm_n63, in_14, in_13, gm_n4563, gm_n46);
	nor (gm_n4565, in_19, in_18, in_17, gm_n4564, gm_n45);
	nand (gm_n4566, gm_n4565, in_21);
	nand (gm_n4567, gm_n50, gm_n49, gm_n48, gm_n3719, in_15);
	nor (gm_n4568, gm_n47, gm_n81, gm_n46, gm_n4567, gm_n62);
	nand (gm_n4569, gm_n4568, gm_n71, gm_n45);
	nor (gm_n4570, gm_n51, gm_n64, gm_n55, gm_n525);
	nand (gm_n4571, gm_n48, gm_n53, gm_n52, gm_n4570, in_13);
	nor (gm_n4572, in_16, gm_n63, gm_n50, gm_n4571, gm_n81);
	nand (gm_n4573, gm_n45, in_19, gm_n47, gm_n4572, gm_n71);
	nor (gm_n4574, in_16, in_15, gm_n50, gm_n1569, in_17);
	nand (gm_n4575, in_20, gm_n62, gm_n47, gm_n4574, gm_n71);
	nand (gm_n4576, gm_n421, in_10, gm_n51);
	or (gm_n4577, gm_n49, gm_n48, in_11, gm_n4576, gm_n50);
	nor (gm_n4578, gm_n81, gm_n46, in_15, gm_n4577, gm_n47);
	nand (gm_n4579, in_21, in_20, gm_n62, gm_n4578);
	nand (gm_n4580, gm_n4573, gm_n4569, gm_n4566, gm_n4579, gm_n4575);
	nor (gm_n4581, gm_n4557, gm_n4553, gm_n4550, gm_n4580, gm_n4561);
	nand (gm_n4582, gm_n4542, gm_n4539, gm_n4536, gm_n4581, gm_n4546);
	nor (gm_n4583, gm_n4529, gm_n4524, gm_n4521, gm_n4582, gm_n4533);
	nand (gm_n4584, gm_n4513, gm_n4510, gm_n4507, gm_n4583, gm_n4518);
	nor (gm_n4585, gm_n4500, gm_n4497, gm_n4493, gm_n4584, gm_n4504);
	nand (gm_n4586, gm_n4483, gm_n4480, gm_n4478, gm_n4585, gm_n4488);
	nor (gm_n4587, gm_n4470, gm_n4467, gm_n4463, gm_n4586, gm_n4474);
	nand (gm_n4588, gm_n4457, gm_n4454, gm_n4450, gm_n4587, gm_n4460);
	nor (gm_n4589, gm_n4442, gm_n4439, gm_n4435, gm_n4588, gm_n4446);
	nand (gm_n4590, gm_n4427, gm_n4424, gm_n4421, gm_n4589, gm_n4431);
	nor (gm_n4591, gm_n4413, gm_n4409, gm_n4405, gm_n4590, gm_n4417);
	nand (gm_n4592, gm_n4397, gm_n4392, gm_n4387, gm_n4591, gm_n4401);
	nor (gm_n4593, gm_n4380, gm_n4376, gm_n4373, gm_n4592, gm_n4384);
	nand (gm_n4594, gm_n4365, gm_n4361, gm_n4357, gm_n4593, gm_n4369);
	nor (gm_n4595, gm_n4350, gm_n4346, gm_n4343, gm_n4594, gm_n4354);
	nand (gm_n4596, gm_n4337, gm_n4334, gm_n4332, gm_n4595, gm_n4340);
	nor (gm_n4597, gm_n4324, gm_n4322, gm_n4318, gm_n4596, gm_n4328);
	nand (gm_n4598, gm_n4309, gm_n4305, gm_n4301, gm_n4597, gm_n4313);
	nor (gm_n4599, gm_n4292, gm_n4289, gm_n4284, gm_n4598, gm_n4297);
	nand (gm_n4600, gm_n4277, gm_n4272, gm_n4269, gm_n4599, gm_n4281);
	nor (gm_n4601, gm_n4261, gm_n4257, gm_n4253, gm_n4600, gm_n4265);
	nand (gm_n4602, gm_n4246, gm_n4242, gm_n4239, gm_n4601, gm_n4249);
	nor (gm_n4603, gm_n4232, gm_n4229, gm_n4226, gm_n4602, gm_n4236);
	nand (gm_n4604, gm_n4220, gm_n4217, gm_n4212, gm_n4603, gm_n4223);
	nor (gm_n4605, gm_n4204, gm_n4199, gm_n4194, gm_n4604, gm_n4208);
	nand (gm_n4606, gm_n4187, gm_n4184, gm_n4181, gm_n4605, gm_n4190);
	nor (gm_n4607, gm_n4172, gm_n4167, gm_n4164, gm_n4606, gm_n4176);
	nand (gm_n4608, gm_n4157, gm_n4152, gm_n4148, gm_n4607, gm_n4160);
	nor (gm_n4609, gm_n4142, gm_n4139, gm_n4137, gm_n4608, gm_n4146);
	nand (gm_n4610, gm_n4130, gm_n4126, gm_n4123, gm_n4609, gm_n4133);
	nor (gm_n4611, gm_n4114, gm_n4111, gm_n4107, gm_n4610, gm_n4118);
	nand (gm_n4612, gm_n4100, gm_n4096, gm_n4093, gm_n4611, gm_n4103);
	nor (gm_n4613, gm_n4086, gm_n4083, gm_n4078, gm_n4612, gm_n4089);
	nand (gm_n4614, gm_n4071, gm_n4068, gm_n4064, gm_n4613, gm_n4075);
	nor (gm_n4615, gm_n4058, gm_n4054, gm_n4049, gm_n4614, gm_n4061);
	nand (gm_n4616, gm_n4041, gm_n4037, gm_n4034, gm_n4615, gm_n4046);
	nor (out_6, gm_n4616, gm_n4030);
	nor (gm_n4618, gm_n55, in_6, gm_n72, gm_n124, gm_n64);
	and (gm_n4619, gm_n53, gm_n52, in_9, gm_n4618);
	and (gm_n4620, gm_n50, in_13, gm_n48, gm_n4619, gm_n63);
	nand (gm_n4621, in_18, in_17, in_16, gm_n4620, gm_n62);
	nor (gm_n4622, gm_n4621, in_21, gm_n45);
	nand (gm_n4623, gm_n48, in_11, gm_n52, gm_n2441, in_13);
	nor (gm_n4624, gm_n46, gm_n63, gm_n50, gm_n4623, gm_n81);
	nand (gm_n4625, gm_n45, in_19, in_18, gm_n4624, gm_n71);
	nor (gm_n4626, gm_n53, in_10, gm_n51, gm_n649, in_12);
	nand (gm_n4627, in_15, gm_n50, gm_n49, gm_n4626, in_16);
	nor (gm_n4628, in_19, gm_n47, in_17, gm_n4627, gm_n45);
	nand (gm_n4629, gm_n4628, gm_n71);
	and (gm_n4630, in_8, gm_n55, gm_n82, gm_n379, in_9);
	nand (gm_n4631, gm_n48, in_11, gm_n52, gm_n4630, in_13);
	nor (gm_n4632, gm_n46, in_15, gm_n50, gm_n4631, gm_n81);
	nand (gm_n4633, gm_n45, in_19, in_18, gm_n4632, in_21);
	nand (gm_n4634, gm_n49, in_12, gm_n53, gm_n260, in_14);
	nor (gm_n4635, in_17, in_16, gm_n63, gm_n4634, in_18);
	nand (gm_n4636, in_21, in_20, in_19, gm_n4635);
	nor (gm_n4637, gm_n49, in_12, in_11, gm_n942, gm_n50);
	nand (gm_n4638, in_17, gm_n46, in_15, gm_n4637, in_18);
	nor (gm_n4639, gm_n71, in_20, gm_n62, gm_n4638);
	and (gm_n4640, gm_n1284, in_10, in_9);
	and (gm_n4641, in_13, in_12, in_11, gm_n4640, in_14);
	nand (gm_n4642, gm_n81, gm_n46, in_15, gm_n4641, gm_n47);
	nor (gm_n4643, in_21, in_20, gm_n62, gm_n4642);
	nor (gm_n4644, in_12, in_11, gm_n52, gm_n1784, in_13);
	nand (gm_n4645, in_16, gm_n63, in_14, gm_n4644, gm_n81);
	nor (gm_n4646, gm_n45, in_19, in_18, gm_n4645, in_21);
	and (gm_n4647, in_14, in_13, in_12, gm_n1303, gm_n63);
	nand (gm_n4648, in_18, in_17, in_16, gm_n4647, in_19);
	nor (gm_n4649, gm_n4648, gm_n71, gm_n45);
	nor (gm_n4650, gm_n53, in_10, in_9, gm_n3475, in_12);
	nand (gm_n4651, in_15, gm_n50, in_13, gm_n4650, in_16);
	nor (gm_n4652, gm_n62, in_18, gm_n81, gm_n4651, in_20);
	nand (gm_n4653, gm_n4652, in_21);
	nor (gm_n4654, gm_n53, in_10, gm_n51, gm_n4314, gm_n48);
	nand (gm_n4655, gm_n63, gm_n50, in_13, gm_n4654, in_16);
	nor (gm_n4656, in_19, in_18, gm_n81, gm_n4655, in_20);
	nand (gm_n4657, gm_n4656, in_21);
	nand (gm_n4658, gm_n63, in_14, in_13, gm_n2894, in_16);
	nor (gm_n4659, gm_n62, gm_n47, in_17, gm_n4658, gm_n45);
	nand (gm_n4660, gm_n4659, in_21);
	and (gm_n4661, gm_n53, gm_n52, gm_n51, gm_n1986, gm_n48);
	nand (gm_n4662, gm_n63, gm_n50, in_13, gm_n4661, in_16);
	nor (gm_n4663, gm_n62, gm_n47, gm_n81, gm_n4662, gm_n45);
	nand (gm_n4664, gm_n4663, in_21);
	nand (gm_n4665, in_19, in_18, gm_n81, gm_n2637, gm_n45);
	nor (gm_n4666, gm_n4665, in_21);
	nand (gm_n4667, gm_n53, gm_n52, gm_n51, gm_n114, gm_n48);
	nor (gm_n4668, gm_n63, gm_n50, gm_n49, gm_n4667, in_16);
	nand (gm_n4669, gm_n62, gm_n47, in_17, gm_n4668, in_20);
	nor (gm_n4670, gm_n4669, gm_n71);
	nor (gm_n4671, gm_n48, in_11, gm_n52, gm_n3159, gm_n49);
	nand (gm_n4672, gm_n46, gm_n63, gm_n50, gm_n4671, in_17);
	nor (gm_n4673, gm_n45, gm_n62, gm_n47, gm_n4672, gm_n71);
	nor (gm_n4674, gm_n49, gm_n48, gm_n53, gm_n391, in_14);
	nand (gm_n4675, in_17, gm_n46, in_15, gm_n4674, gm_n47);
	nor (gm_n4676, in_21, gm_n45, in_19, gm_n4675);
	nor (gm_n4677, in_10, in_9, gm_n64, gm_n3174);
	nand (gm_n4678, gm_n49, gm_n48, gm_n53, gm_n4677, in_14);
	nor (gm_n4679, gm_n81, gm_n46, in_15, gm_n4678, gm_n47);
	nand (gm_n4680, gm_n71, gm_n45, gm_n62, gm_n4679);
	and (gm_n4681, gm_n52, in_9, in_8, gm_n57);
	nand (gm_n4682, in_13, in_12, gm_n53, gm_n4681, gm_n50);
	nor (gm_n4683, in_17, gm_n46, in_15, gm_n4682, in_18);
	nand (gm_n4684, gm_n71, gm_n45, gm_n62, gm_n4683);
	nand (gm_n4685, in_12, gm_n53, gm_n52, gm_n3354, in_13);
	nor (gm_n4686, gm_n46, in_15, in_14, gm_n4685, gm_n81);
	nand (gm_n4687, in_20, in_19, in_18, gm_n4686, in_21);
	and (gm_n4688, gm_n51, in_8, in_7, gm_n404, gm_n52);
	nand (gm_n4689, gm_n49, in_12, gm_n53, gm_n4688, gm_n50);
	nor (gm_n4690, in_17, in_16, gm_n63, gm_n4689, in_18);
	nand (gm_n4691, in_21, gm_n45, in_19, gm_n4690);
	or (gm_n4692, in_8, in_7, in_6, gm_n199, in_9);
	nor (gm_n4693, in_12, in_11, in_10, gm_n4692, in_13);
	nand (gm_n4694, gm_n46, in_15, in_14, gm_n4693, in_17);
	nor (gm_n4695, in_20, in_19, in_18, gm_n4694, gm_n71);
	or (gm_n4696, in_8, in_7, gm_n82, gm_n204, in_9);
	nor (gm_n4697, in_12, gm_n53, in_10, gm_n4696, gm_n49);
	nand (gm_n4698, in_16, in_15, gm_n50, gm_n4697, gm_n81);
	nor (gm_n4699, in_20, gm_n62, gm_n47, gm_n4698, gm_n71);
	and (gm_n4700, gm_n48, in_11, gm_n52, gm_n3324, in_13);
	nand (gm_n4701, gm_n46, gm_n63, in_14, gm_n4700, in_17);
	nor (gm_n4702, in_20, in_19, gm_n47, gm_n4701, in_21);
	and (gm_n4703, gm_n792, gm_n52, in_9);
	and (gm_n4704, gm_n49, gm_n48, gm_n53, gm_n4703, gm_n50);
	nand (gm_n4705, in_17, in_16, in_15, gm_n4704, in_18);
	nor (gm_n4706, in_21, in_20, in_19, gm_n4705);
	nor (gm_n4707, gm_n81, gm_n46, gm_n63, gm_n4091, in_18);
	nand (gm_n4708, in_21, gm_n45, gm_n62, gm_n4707);
	nand (gm_n4709, in_15, in_14, gm_n49, gm_n4661, in_16);
	nor (gm_n4710, in_19, in_18, in_17, gm_n4709, gm_n45);
	nand (gm_n4711, gm_n4710, in_21);
	nor (gm_n4712, in_12, in_11, in_10, gm_n3508, gm_n49);
	nand (gm_n4713, gm_n46, gm_n63, gm_n50, gm_n4712, gm_n81);
	or (gm_n4714, gm_n45, gm_n62, in_18, gm_n4713, in_21);
	or (gm_n4715, gm_n468, gm_n51, in_8);
	or (gm_n4716, gm_n48, in_11, in_10, gm_n4715, gm_n49);
	nor (gm_n4717, in_16, gm_n63, in_14, gm_n4716, in_17);
	nand (gm_n4718, gm_n45, in_19, in_18, gm_n4717, in_21);
	nand (gm_n4719, in_11, gm_n52, gm_n51, gm_n494, gm_n48);
	nor (gm_n4720, gm_n63, gm_n50, in_13, gm_n4719, in_16);
	nand (gm_n4721, in_19, gm_n47, gm_n81, gm_n4720, gm_n45);
	nor (gm_n4722, gm_n4721, in_21);
	nor (gm_n4723, in_7, gm_n82, gm_n72, gm_n124, gm_n64);
	nand (gm_n4724, in_11, in_10, gm_n51, gm_n4723, gm_n48);
	nor (gm_n4725, gm_n63, in_14, gm_n49, gm_n4724, gm_n46);
	nand (gm_n4726, gm_n62, in_18, gm_n81, gm_n4725, gm_n45);
	nor (gm_n4727, gm_n4726, gm_n71);
	and (gm_n4728, in_13, in_12, gm_n53, gm_n2721, gm_n50);
	nand (gm_n4729, in_17, in_16, gm_n63, gm_n4728, in_18);
	nor (gm_n4730, gm_n71, in_20, gm_n62, gm_n4729);
	nand (gm_n4731, in_11, gm_n52, in_9, gm_n3043, in_12);
	nor (gm_n4732, in_15, in_14, in_13, gm_n4731, in_16);
	nand (gm_n4733, in_19, gm_n47, gm_n81, gm_n4732, in_20);
	nor (gm_n4734, gm_n4733, in_21);
	nand (gm_n4735, in_12, in_11, in_10, gm_n934, in_13);
	nor (gm_n4736, in_16, in_15, in_14, gm_n4735, in_17);
	nand (gm_n4737, gm_n45, in_19, gm_n47, gm_n4736, gm_n71);
	nand (gm_n4738, gm_n49, in_12, gm_n53, gm_n2611);
	nor (gm_n4739, gm_n46, gm_n63, in_14, gm_n4738, in_17);
	nand (gm_n4740, gm_n45, in_19, gm_n47, gm_n4739, gm_n71);
	and (gm_n4741, gm_n2481, gm_n52, gm_n51);
	nand (gm_n4742, gm_n49, in_12, in_11, gm_n4741, in_14);
	nor (gm_n4743, in_17, in_16, in_15, gm_n4742, in_18);
	nand (gm_n4744, gm_n71, gm_n45, in_19, gm_n4743);
	nand (gm_n4745, in_15, in_14, gm_n49, gm_n3849, gm_n46);
	nor (gm_n4746, gm_n62, gm_n47, gm_n81, gm_n4745, in_20);
	nand (gm_n4747, gm_n4746, in_21);
	nand (gm_n4748, gm_n53, gm_n52, gm_n51, gm_n1895);
	nor (gm_n4749, gm_n50, in_13, gm_n48, gm_n4748, gm_n63);
	nand (gm_n4750, in_18, in_17, gm_n46, gm_n4749, in_19);
	nor (gm_n4751, gm_n4750, in_21, in_20);
	nor (gm_n4752, in_8, in_7, in_6, gm_n204, in_9);
	and (gm_n4753, in_12, gm_n53, in_10, gm_n4752, in_13);
	nand (gm_n4754, gm_n46, gm_n63, in_14, gm_n4753, gm_n81);
	nor (gm_n4755, in_20, in_19, in_18, gm_n4754, gm_n71);
	and (gm_n4756, gm_n48, in_11, gm_n52, gm_n205, gm_n49);
	nand (gm_n4757, gm_n46, in_15, gm_n50, gm_n4756, in_17);
	nor (gm_n4758, in_20, in_19, gm_n47, gm_n4757, in_21);
	nor (gm_n4759, gm_n49, gm_n48, gm_n53, gm_n4414, gm_n50);
	nand (gm_n4760, in_17, in_16, gm_n63, gm_n4759, gm_n47);
	nor (gm_n4761, in_21, in_20, in_19, gm_n4760);
	nor (gm_n4762, gm_n53, gm_n52, in_9, gm_n1481, gm_n48);
	nand (gm_n4763, in_15, gm_n50, gm_n49, gm_n4762, in_16);
	nor (gm_n4764, in_19, gm_n47, gm_n81, gm_n4763, gm_n45);
	nand (gm_n4765, gm_n4764, gm_n71);
	nand (gm_n4766, gm_n49, in_12, gm_n53, gm_n3756, gm_n50);
	nor (gm_n4767, gm_n81, in_16, gm_n63, gm_n4766, in_18);
	nand (gm_n4768, gm_n71, in_20, gm_n62, gm_n4767);
	nor (gm_n4769, gm_n53, in_10, gm_n51, gm_n1879, gm_n48);
	nand (gm_n4770, gm_n63, gm_n50, gm_n49, gm_n4769, in_16);
	nor (gm_n4771, in_19, gm_n47, gm_n81, gm_n4770, in_20);
	nand (gm_n4772, gm_n4771, gm_n71);
	nor (gm_n4773, in_17, gm_n46, in_15, gm_n2313, in_18);
	nand (gm_n4774, in_21, in_20, gm_n62, gm_n4773);
	nor (gm_n4775, gm_n50, gm_n49, in_12, gm_n2935, gm_n63);
	nand (gm_n4776, gm_n47, gm_n81, in_16, gm_n4775, gm_n62);
	nor (gm_n4777, gm_n4776, gm_n71, in_20);
	nor (gm_n4778, gm_n49, gm_n48, in_11, gm_n445, in_14);
	nand (gm_n4779, gm_n81, gm_n46, gm_n63, gm_n4778, gm_n47);
	nor (gm_n4780, in_21, gm_n45, gm_n62, gm_n4779);
	nor (gm_n4781, in_15, gm_n50, in_13, gm_n3464, in_16);
	nand (gm_n4782, in_19, in_18, gm_n81, gm_n4781, in_20);
	nor (gm_n4783, gm_n4782, gm_n71);
	nor (gm_n4784, gm_n53, gm_n52, gm_n51, gm_n2546, in_12);
	and (gm_n4785, in_15, in_14, in_13, gm_n4784, in_16);
	nand (gm_n4786, gm_n62, in_18, in_17, gm_n4785, in_20);
	nor (gm_n4787, gm_n4786, in_21);
	and (gm_n4788, in_18, gm_n81, in_16, gm_n116, gm_n62);
	nand (gm_n4789, gm_n4788, in_21, gm_n45);
	nand (gm_n4790, in_11, gm_n52, gm_n51, gm_n3451);
	or (gm_n4791, gm_n50, in_13, gm_n48, gm_n4790, gm_n63);
	nor (gm_n4792, gm_n47, in_17, gm_n46, gm_n4791, gm_n62);
	nand (gm_n4793, gm_n4792, in_21, in_20);
	and (gm_n4794, in_10, in_9, gm_n64, gm_n1608);
	nand (gm_n4795, in_13, gm_n48, in_11, gm_n4794, in_14);
	nor (gm_n4796, gm_n81, gm_n46, in_15, gm_n4795, in_18);
	nand (gm_n4797, in_21, in_20, gm_n62, gm_n4796);
	and (gm_n4798, gm_n53, in_10, gm_n51, gm_n473, in_12);
	nand (gm_n4799, gm_n63, in_14, in_13, gm_n4798, gm_n46);
	nor (gm_n4800, gm_n62, in_18, in_17, gm_n4799, gm_n45);
	nand (gm_n4801, gm_n4800, gm_n71);
	and (gm_n4802, gm_n53, gm_n52, gm_n51, gm_n1683);
	and (gm_n4803, in_14, in_13, in_12, gm_n4802, in_15);
	nand (gm_n4804, in_18, in_17, in_16, gm_n4803, in_19);
	nor (gm_n4805, gm_n4804, gm_n71, gm_n45);
	and (gm_n4806, in_12, gm_n53, in_10, gm_n885, in_13);
	nand (gm_n4807, gm_n46, in_15, in_14, gm_n4806, in_17);
	nor (gm_n4808, in_20, in_19, in_18, gm_n4807, in_21);
	nand (gm_n4809, gm_n173, gm_n51);
	nor (gm_n4810, gm_n48, gm_n53, in_10, gm_n4809, in_13);
	nand (gm_n4811, in_16, gm_n63, gm_n50, gm_n4810, gm_n81);
	nor (gm_n4812, in_20, gm_n62, in_18, gm_n4811, in_21);
	and (gm_n4813, gm_n4050, in_10, in_9);
	and (gm_n4814, in_13, gm_n48, in_11, gm_n4813, in_14);
	nand (gm_n4815, gm_n81, in_16, in_15, gm_n4814, in_18);
	nor (gm_n4816, in_21, gm_n45, in_19, gm_n4815);
	nor (gm_n4817, gm_n53, in_10, gm_n51, gm_n774, gm_n48);
	nand (gm_n4818, gm_n63, in_14, gm_n49, gm_n4817, gm_n46);
	nor (gm_n4819, gm_n62, in_18, in_17, gm_n4818, gm_n45);
	nand (gm_n4820, gm_n4819, in_21);
	nand (gm_n4821, in_13, gm_n48, gm_n53, gm_n1344, in_14);
	nor (gm_n4822, in_17, in_16, in_15, gm_n4821, gm_n47);
	nand (gm_n4823, gm_n71, in_20, in_19, gm_n4822);
	and (gm_n4824, in_17, gm_n46, gm_n63, gm_n763, in_18);
	nand (gm_n4825, gm_n71, in_20, gm_n62, gm_n4824);
	nor (gm_n4826, in_10, gm_n51, gm_n64, gm_n468, gm_n53);
	nand (gm_n4827, in_14, in_13, in_12, gm_n4826, gm_n63);
	nor (gm_n4828, in_18, in_17, gm_n46, gm_n4827, gm_n62);
	nand (gm_n4829, gm_n4828, in_21, in_20);
	nor (gm_n4830, in_15, in_14, in_13, gm_n110, in_16);
	nand (gm_n4831, in_19, gm_n47, in_17, gm_n4830, gm_n45);
	nor (gm_n4832, gm_n4831, gm_n71);
	nor (gm_n4833, in_13, gm_n48, in_11, gm_n1208, in_14);
	nand (gm_n4834, gm_n81, gm_n46, in_15, gm_n4833, in_18);
	nor (gm_n4835, in_21, gm_n45, in_19, gm_n4834);
	nand (gm_n4836, gm_n53, in_10, in_9, gm_n2653, in_12);
	nor (gm_n4837, in_15, gm_n50, gm_n49, gm_n4836, gm_n46);
	nand (gm_n4838, gm_n62, in_18, gm_n81, gm_n4837, gm_n45);
	nor (gm_n4839, gm_n4838, gm_n71);
	and (gm_n4840, in_12, gm_n53, in_10, gm_n2760, gm_n49);
	nand (gm_n4841, in_16, gm_n63, in_14, gm_n4840, gm_n81);
	nor (gm_n4842, gm_n45, in_19, gm_n47, gm_n4841, in_21);
	nand (gm_n4843, gm_n49, gm_n48, in_11, gm_n3429, in_14);
	nor (gm_n4844, gm_n81, gm_n46, gm_n63, gm_n4843, in_18);
	nand (gm_n4845, gm_n71, gm_n45, in_19, gm_n4844);
	nor (gm_n4846, in_11, in_10, in_9, gm_n2546, gm_n48);
	nand (gm_n4847, gm_n63, in_14, gm_n49, gm_n4846, in_16);
	nor (gm_n4848, in_19, gm_n47, gm_n81, gm_n4847, in_20);
	nand (gm_n4849, gm_n4848, in_21);
	nor (gm_n4850, gm_n52, gm_n51, gm_n64, gm_n468, gm_n53);
	nand (gm_n4851, in_14, gm_n49, gm_n48, gm_n4850, gm_n63);
	nor (gm_n4852, in_18, in_17, gm_n46, gm_n4851, in_19);
	nand (gm_n4853, gm_n4852, in_21, in_20);
	nand (gm_n4854, in_14, gm_n49, gm_n48, gm_n709, in_15);
	nor (gm_n4855, in_18, in_17, in_16, gm_n4854, in_19);
	nand (gm_n4856, gm_n4855, gm_n71, in_20);
	and (gm_n4857, in_12, in_11, in_10, gm_n1804, gm_n49);
	nand (gm_n4858, gm_n46, in_15, gm_n50, gm_n4857, gm_n81);
	nor (gm_n4859, in_20, in_19, gm_n47, gm_n4858, gm_n71);
	nor (gm_n4860, in_11, gm_n52, in_9, gm_n520, gm_n48);
	and (gm_n4861, in_15, gm_n50, gm_n49, gm_n4860, in_16);
	nand (gm_n4862, gm_n62, gm_n47, in_17, gm_n4861, gm_n45);
	nor (gm_n4863, gm_n4862, gm_n71);
	nand (gm_n4864, in_11, gm_n52, in_9, gm_n473);
	nor (gm_n4865, in_14, gm_n49, in_12, gm_n4864, in_15);
	nand (gm_n4866, in_18, gm_n81, gm_n46, gm_n4865, gm_n62);
	nor (gm_n4867, gm_n4866, gm_n71, gm_n45);
	nor (gm_n4868, in_11, in_10, gm_n51, gm_n368, gm_n48);
	and (gm_n4869, in_15, gm_n50, in_13, gm_n4868, gm_n46);
	nand (gm_n4870, gm_n62, gm_n47, gm_n81, gm_n4869, in_20);
	nor (gm_n4871, gm_n4870, in_21);
	nor (gm_n4872, in_9, gm_n64, in_7, gm_n279, gm_n52);
	nand (gm_n4873, gm_n49, gm_n48, in_11, gm_n4872, gm_n50);
	nor (gm_n4874, gm_n81, gm_n46, gm_n63, gm_n4873, gm_n47);
	nand (gm_n4875, gm_n71, gm_n45, in_19, gm_n4874);
	nor (gm_n4876, in_8, in_7, in_6, gm_n530, gm_n51);
	nand (gm_n4877, in_12, gm_n53, gm_n52, gm_n4876, gm_n49);
	nor (gm_n4878, gm_n46, gm_n63, in_14, gm_n4877, gm_n81);
	nand (gm_n4879, gm_n45, gm_n62, in_18, gm_n4878, in_21);
	or (gm_n4880, in_11, gm_n52, gm_n51, gm_n178, in_12);
	nor (gm_n4881, gm_n4880, gm_n49);
	and (gm_n4882, gm_n46, gm_n63, gm_n50, gm_n4881, in_17);
	nand (gm_n4883, gm_n45, in_19, in_18, gm_n4882, gm_n71);
	nand (gm_n4884, gm_n48, in_11, in_10, gm_n311, in_13);
	nor (gm_n4885, in_16, gm_n63, in_14, gm_n4884, gm_n81);
	nand (gm_n4886, in_20, gm_n62, gm_n47, gm_n4885, in_21);
	nor (gm_n4887, gm_n53, gm_n52, in_9, gm_n218);
	and (gm_n4888, in_14, gm_n49, in_12, gm_n4887, in_15);
	nand (gm_n4889, gm_n47, gm_n81, in_16, gm_n4888, in_19);
	nor (gm_n4890, gm_n4889, in_21, gm_n45);
	nand (gm_n4891, gm_n109, in_10, gm_n51);
	nor (gm_n4892, gm_n49, in_12, in_11, gm_n4891, in_14);
	nand (gm_n4893, in_17, gm_n46, in_15, gm_n4892, in_18);
	nor (gm_n4894, gm_n71, gm_n45, gm_n62, gm_n4893);
	nand (gm_n4895, in_17, gm_n46, in_15, gm_n3674, in_18);
	nor (gm_n4896, in_21, in_20, gm_n62, gm_n4895);
	nor (gm_n4897, in_12, in_11, gm_n52, gm_n2280, in_13);
	nand (gm_n4898, in_16, gm_n63, in_14, gm_n4897, in_17);
	nor (gm_n4899, gm_n45, in_19, in_18, gm_n4898, gm_n71);
	nor (gm_n4900, in_16, in_15, in_14, gm_n446, gm_n81);
	nand (gm_n4901, gm_n45, gm_n62, in_18, gm_n4900, gm_n71);
	nor (gm_n4902, in_11, in_10, gm_n51, gm_n2114, gm_n48);
	nand (gm_n4903, gm_n63, gm_n50, in_13, gm_n4902, in_16);
	nor (gm_n4904, gm_n62, gm_n47, gm_n81, gm_n4903, gm_n45);
	nand (gm_n4905, gm_n4904, gm_n71);
	or (gm_n4906, gm_n64, in_7, gm_n82, gm_n204, gm_n51);
	nor (gm_n4907, gm_n4906, in_10);
	nand (gm_n4908, in_13, gm_n48, gm_n53, gm_n4907, in_14);
	nor (gm_n4909, gm_n81, gm_n46, in_15, gm_n4908, in_18);
	nand (gm_n4910, in_21, gm_n45, gm_n62, gm_n4909);
	nor (gm_n4911, gm_n64, gm_n55, in_6, gm_n141, in_9);
	nand (gm_n4912, gm_n48, gm_n53, gm_n52, gm_n4911, gm_n49);
	nor (gm_n4913, gm_n46, in_15, gm_n50, gm_n4912, gm_n81);
	nand (gm_n4914, in_20, in_19, in_18, gm_n4913, in_21);
	nor (gm_n4915, in_12, gm_n53, in_10, gm_n3931, gm_n49);
	nand (gm_n4916, in_16, gm_n63, in_14, gm_n4915, gm_n81);
	nor (gm_n4917, gm_n45, gm_n62, gm_n47, gm_n4916, gm_n71);
	nor (gm_n4918, gm_n1035, gm_n51);
	and (gm_n4919, gm_n48, in_11, in_10, gm_n4918, in_13);
	nand (gm_n4920, in_16, in_15, gm_n50, gm_n4919, in_17);
	nor (gm_n4921, in_20, gm_n62, gm_n47, gm_n4920, gm_n71);
	nor (gm_n4922, gm_n51, gm_n64, in_7, gm_n84, gm_n52);
	and (gm_n4923, gm_n49, in_12, gm_n53, gm_n4922, gm_n50);
	nand (gm_n4924, gm_n81, in_16, gm_n63, gm_n4923, in_18);
	nor (gm_n4925, in_21, in_20, in_19, gm_n4924);
	nor (gm_n4926, in_13, gm_n48, gm_n53, gm_n1381, in_14);
	nand (gm_n4927, gm_n81, gm_n46, gm_n63, gm_n4926, gm_n47);
	nor (gm_n4928, in_21, in_20, gm_n62, gm_n4927);
	or (gm_n4929, gm_n53, in_10, gm_n51, gm_n410, in_12);
	or (gm_n4930, gm_n63, in_14, gm_n49, gm_n4929, gm_n46);
	nor (gm_n4931, gm_n62, in_18, in_17, gm_n4930, gm_n45);
	nand (gm_n4932, gm_n4931, in_21);
	or (gm_n4933, gm_n50, in_13, gm_n48, gm_n922, in_15);
	nor (gm_n4934, in_18, gm_n81, gm_n46, gm_n4933, in_19);
	nand (gm_n4935, gm_n4934, gm_n71, gm_n45);
	and (gm_n4936, in_11, gm_n52, in_9, gm_n658);
	nand (gm_n4937, in_14, gm_n49, in_12, gm_n4936, gm_n63);
	nor (gm_n4938, in_18, in_17, gm_n46, gm_n4937, in_19);
	nand (gm_n4939, gm_n4938, in_21, in_20);
	nand (gm_n4940, gm_n48, gm_n53, gm_n52, gm_n1128, in_13);
	nor (gm_n4941, in_16, gm_n63, in_14, gm_n4940, in_17);
	nand (gm_n4942, gm_n45, in_19, gm_n47, gm_n4941, in_21);
	nand (gm_n4943, in_11, in_10, gm_n51, gm_n543);
	nor (gm_n4944, gm_n50, gm_n49, in_12, gm_n4943, gm_n63);
	nand (gm_n4945, gm_n47, in_17, in_16, gm_n4944, in_19);
	nor (gm_n4946, gm_n4945, in_21, in_20);
	nor (gm_n4947, gm_n49, gm_n48, gm_n53, gm_n3954, gm_n50);
	nand (gm_n4948, gm_n81, in_16, gm_n63, gm_n4947, gm_n47);
	nor (gm_n4949, gm_n71, gm_n45, in_19, gm_n4948);
	nor (gm_n4950, in_9, gm_n64, in_7, gm_n553);
	and (gm_n4951, gm_n48, in_11, in_10, gm_n4950, in_13);
	nand (gm_n4952, in_16, in_15, gm_n50, gm_n4951, gm_n81);
	nor (gm_n4953, in_20, in_19, gm_n47, gm_n4952, in_21);
	and (gm_n4954, gm_n48, in_11, gm_n52, gm_n2593, gm_n49);
	nand (gm_n4955, gm_n46, in_15, gm_n50, gm_n4954, gm_n81);
	nor (gm_n4956, gm_n45, gm_n62, gm_n47, gm_n4955, in_21);
	nand (gm_n4957, gm_n45, gm_n62, gm_n47, gm_n2656, gm_n71);
	nand (gm_n4958, in_13, in_12, gm_n53, gm_n4872, gm_n50);
	nor (gm_n4959, gm_n81, in_16, in_15, gm_n4958, in_18);
	nand (gm_n4960, in_21, gm_n45, in_19, gm_n4959);
	nor (gm_n4961, in_10, in_9, in_8, gm_n3077, gm_n53);
	nand (gm_n4962, gm_n50, gm_n49, gm_n48, gm_n4961, gm_n63);
	nor (gm_n4963, in_18, gm_n81, in_16, gm_n4962, gm_n62);
	nand (gm_n4964, gm_n4963, in_21, gm_n45);
	nand (gm_n4965, in_12, in_11, in_10, gm_n3163, in_13);
	nor (gm_n4966, in_16, gm_n63, gm_n50, gm_n4965, gm_n81);
	nand (gm_n4967, in_20, gm_n62, gm_n47, gm_n4966, gm_n71);
	and (gm_n4968, gm_n4484, gm_n51);
	and (gm_n4969, in_12, gm_n53, gm_n52, gm_n4968, gm_n49);
	nand (gm_n4970, in_16, in_15, in_14, gm_n4969, in_17);
	nor (gm_n4971, in_20, in_19, in_18, gm_n4970, in_21);
	or (gm_n4972, gm_n51, in_8, in_7, gm_n553, in_10);
	nor (gm_n4973, in_13, gm_n48, gm_n53, gm_n4972, gm_n50);
	nand (gm_n4974, gm_n81, gm_n46, gm_n63, gm_n4973, in_18);
	nor (gm_n4975, gm_n71, in_20, gm_n62, gm_n4974);
	nand (gm_n4976, gm_n64, in_7, gm_n82, gm_n379, gm_n51);
	nor (gm_n4977, gm_n48, in_11, gm_n52, gm_n4976, gm_n49);
	nand (gm_n4978, gm_n46, in_15, gm_n50, gm_n4977, gm_n81);
	nor (gm_n4979, gm_n45, in_19, in_18, gm_n4978, in_21);
	or (gm_n4980, gm_n51, gm_n64, gm_n55, gm_n897, gm_n52);
	nor (gm_n4981, gm_n49, in_12, gm_n53, gm_n4980, gm_n50);
	nand (gm_n4982, in_17, gm_n46, gm_n63, gm_n4981, in_18);
	nor (gm_n4983, in_21, gm_n45, gm_n62, gm_n4982);
	and (gm_n4984, in_8, in_7, gm_n82, gm_n379, in_9);
	nand (gm_n4985, in_12, gm_n53, gm_n52, gm_n4984, in_13);
	nor (gm_n4986, in_16, gm_n63, gm_n50, gm_n4985, in_17);
	nand (gm_n4987, gm_n45, in_19, gm_n47, gm_n4986, in_21);
	nand (gm_n4988, gm_n49, in_12, in_11, gm_n3291, gm_n50);
	nor (gm_n4989, gm_n81, in_16, in_15, gm_n4988, gm_n47);
	nand (gm_n4990, gm_n71, gm_n45, in_19, gm_n4989);
	or (gm_n4991, in_20, gm_n62, in_18, gm_n4713, in_21);
	nor (gm_n4992, in_11, in_10, gm_n51, gm_n3844);
	nand (gm_n4993, gm_n50, in_13, in_12, gm_n4992, in_15);
	nor (gm_n4994, in_18, gm_n81, gm_n46, gm_n4993, gm_n62);
	nand (gm_n4995, gm_n4994, in_21, in_20);
	nor (gm_n4996, gm_n48, gm_n53, in_10, gm_n3159, gm_n49);
	nand (gm_n4997, in_16, gm_n63, gm_n50, gm_n4996, gm_n81);
	nor (gm_n4998, gm_n45, in_19, gm_n47, gm_n4997, in_21);
	and (gm_n4999, gm_n53, in_10, gm_n51, gm_n1936);
	and (gm_n5000, gm_n50, in_13, gm_n48, gm_n4999, gm_n63);
	nand (gm_n5001, gm_n47, gm_n81, gm_n46, gm_n5000, in_19);
	nor (gm_n5002, gm_n5001, gm_n71, gm_n45);
	and (gm_n5003, gm_n51, in_8, in_7, gm_n66, in_10);
	and (gm_n5004, gm_n49, gm_n48, in_11, gm_n5003, gm_n50);
	nand (gm_n5005, gm_n81, in_16, gm_n63, gm_n5004, in_18);
	nor (gm_n5006, in_21, in_20, in_19, gm_n5005);
	nor (gm_n5007, in_14, gm_n49, gm_n48, gm_n1066, gm_n63);
	nand (gm_n5008, gm_n47, in_17, in_16, gm_n5007, in_19);
	nor (gm_n5009, gm_n5008, gm_n71, gm_n45);
	nor (gm_n5010, in_11, in_10, in_9, gm_n2926, gm_n48);
	nand (gm_n5011, in_15, in_14, gm_n49, gm_n5010, in_16);
	nor (gm_n5012, gm_n62, in_18, gm_n81, gm_n5011, in_20);
	nand (gm_n5013, gm_n5012, gm_n71);
	nor (gm_n5014, in_11, gm_n52, gm_n51, gm_n395, gm_n48);
	nand (gm_n5015, gm_n63, in_14, in_13, gm_n5014, in_16);
	nor (gm_n5016, in_19, in_18, gm_n81, gm_n5015, in_20);
	nand (gm_n5017, gm_n5016, in_21);
	and (gm_n5018, gm_n46, in_15, gm_n50, gm_n312, in_17);
	nand (gm_n5019, gm_n45, in_19, in_18, gm_n5018, in_21);
	nand (gm_n5020, gm_n48, in_11, gm_n52, gm_n2619, gm_n49);
	nor (gm_n5021, in_16, gm_n63, gm_n50, gm_n5020, gm_n81);
	nand (gm_n5022, in_20, in_19, in_18, gm_n5021, in_21);
	nor (gm_n5023, gm_n50, in_13, gm_n48, gm_n3002, gm_n63);
	nand (gm_n5024, in_18, gm_n81, gm_n46, gm_n5023, in_19);
	nor (gm_n5025, gm_n5024, gm_n71, in_20);
	nand (gm_n5026, in_11, in_10, gm_n51, gm_n1142, in_12);
	nor (gm_n5027, in_15, gm_n50, gm_n49, gm_n5026, gm_n46);
	nand (gm_n5028, gm_n62, gm_n47, in_17, gm_n5027, gm_n45);
	nor (gm_n5029, gm_n5028, in_21);
	or (gm_n5030, gm_n64, in_7, gm_n82, gm_n156, in_9);
	nor (gm_n5031, in_12, in_11, in_10, gm_n5030, in_13);
	nand (gm_n5032, in_16, gm_n63, gm_n50, gm_n5031, gm_n81);
	nor (gm_n5033, gm_n45, gm_n62, gm_n47, gm_n5032, gm_n71);
	nor (gm_n5034, in_11, gm_n52, gm_n51, gm_n1831);
	and (gm_n5035, gm_n50, gm_n49, in_12, gm_n5034, in_15);
	nand (gm_n5036, in_18, in_17, in_16, gm_n5035, gm_n62);
	nor (gm_n5037, gm_n5036, gm_n71, gm_n45);
	and (gm_n5038, in_12, in_11, gm_n52, gm_n4984, in_13);
	and (gm_n5039, in_16, in_15, in_14, gm_n5038, gm_n81);
	nand (gm_n5040, in_20, in_19, in_18, gm_n5039, in_21);
	or (gm_n5041, gm_n51, in_8, in_7, gm_n259, gm_n52);
	nor (gm_n5042, in_13, in_12, in_11, gm_n5041, in_14);
	and (gm_n5043, in_17, in_16, in_15, gm_n5042, gm_n47);
	nand (gm_n5044, in_21, in_20, in_19, gm_n5043);
	nand (gm_n5045, gm_n48, gm_n53, in_10, gm_n2873, in_13);
	nor (gm_n5046, gm_n46, in_15, in_14, gm_n5045, gm_n81);
	nand (gm_n5047, gm_n45, in_19, gm_n47, gm_n5046, in_21);
	nor (gm_n5048, in_9, in_8, gm_n55, gm_n553, gm_n52);
	nand (gm_n5049, in_13, gm_n48, gm_n53, gm_n5048, gm_n50);
	nor (gm_n5050, in_17, in_16, gm_n63, gm_n5049, gm_n47);
	nand (gm_n5051, in_21, gm_n45, in_19, gm_n5050);
	nand (gm_n5052, gm_n51, gm_n64, in_7, gm_n136, gm_n52);
	nor (gm_n5053, gm_n49, gm_n48, gm_n53, gm_n5052, in_14);
	nand (gm_n5054, in_17, in_16, gm_n63, gm_n5053, gm_n47);
	nor (gm_n5055, gm_n71, gm_n45, in_19, gm_n5054);
	or (gm_n5056, gm_n52, in_9, gm_n64, gm_n390);
	nor (gm_n5057, in_13, gm_n48, in_11, gm_n5056, gm_n50);
	nand (gm_n5058, in_17, in_16, in_15, gm_n5057, in_18);
	nor (gm_n5059, in_21, in_20, in_19, gm_n5058);
	or (gm_n5060, gm_n53, in_10, gm_n51, gm_n1803);
	nor (gm_n5061, gm_n5060, in_13, in_12);
	nand (gm_n5062, in_16, gm_n63, gm_n50, gm_n5061, gm_n81);
	nor (gm_n5063, gm_n45, in_19, in_18, gm_n5062, gm_n71);
	and (gm_n5064, in_11, gm_n52, gm_n51, gm_n2432);
	and (gm_n5065, in_14, in_13, gm_n48, gm_n5064, in_15);
	nand (gm_n5066, gm_n47, gm_n81, in_16, gm_n5065, gm_n62);
	nor (gm_n5067, gm_n5066, in_21, gm_n45);
	nand (gm_n5068, in_15, gm_n50, gm_n49, gm_n4274, in_16);
	nor (gm_n5069, in_19, gm_n47, gm_n81, gm_n5068, in_20);
	nand (gm_n5070, gm_n5069, gm_n71);
	nor (gm_n5071, in_11, in_10, gm_n51, gm_n2823, gm_n48);
	nand (gm_n5072, gm_n63, in_14, gm_n49, gm_n5071, gm_n46);
	nor (gm_n5073, gm_n62, in_18, gm_n81, gm_n5072, gm_n45);
	nand (gm_n5074, gm_n5073, gm_n71);
	nand (gm_n5075, in_12, gm_n53, gm_n52, gm_n4918, gm_n49);
	nor (gm_n5076, gm_n46, gm_n63, gm_n50, gm_n5075, gm_n81);
	nand (gm_n5077, gm_n45, gm_n62, gm_n47, gm_n5076, in_21);
	and (gm_n5078, in_12, in_11, gm_n52, gm_n2619, gm_n49);
	and (gm_n5079, gm_n46, in_15, gm_n50, gm_n5078, in_17);
	nand (gm_n5080, gm_n45, in_19, gm_n47, gm_n5079, in_21);
	nor (gm_n5081, in_13, gm_n48, gm_n53, gm_n4576, in_14);
	nand (gm_n5082, gm_n81, gm_n46, in_15, gm_n5081, in_18);
	nor (gm_n5083, in_21, in_20, gm_n62, gm_n5082);
	nand (gm_n5084, gm_n53, in_10, in_9, gm_n2631);
	nor (gm_n5085, in_14, gm_n49, in_12, gm_n5084, gm_n63);
	nand (gm_n5086, in_18, gm_n81, in_16, gm_n5085, in_19);
	nor (gm_n5087, gm_n5086, gm_n71, gm_n45);
	nor (gm_n5088, gm_n50, in_13, gm_n48, gm_n3666, gm_n63);
	nand (gm_n5089, gm_n47, gm_n81, gm_n46, gm_n5088, in_19);
	nor (gm_n5090, gm_n5089, gm_n71, gm_n45);
	nand (gm_n5091, in_11, in_10, in_9, gm_n210, gm_n48);
	nor (gm_n5092, in_15, in_14, in_13, gm_n5091, in_16);
	nand (gm_n5093, in_19, in_18, in_17, gm_n5092, gm_n45);
	nor (gm_n5094, gm_n5093, in_21);
	nor (gm_n5095, in_11, gm_n52, gm_n51, gm_n2419, gm_n48);
	nand (gm_n5096, gm_n63, gm_n50, gm_n49, gm_n5095, gm_n46);
	nor (gm_n5097, gm_n62, in_18, in_17, gm_n5096, in_20);
	nand (gm_n5098, gm_n5097, in_21);
	and (gm_n5099, gm_n53, in_10, gm_n51, gm_n644);
	nand (gm_n5100, gm_n50, gm_n49, in_12, gm_n5099, gm_n63);
	nor (gm_n5101, in_18, in_17, gm_n46, gm_n5100, gm_n62);
	nand (gm_n5102, gm_n5101, in_21, gm_n45);
	nand (gm_n5103, gm_n63, gm_n50, in_13, gm_n179, in_16);
	nor (gm_n5104, gm_n62, in_18, in_17, gm_n5103, gm_n45);
	nand (gm_n5105, gm_n5104, in_21);
	nand (gm_n5106, in_13, in_12, gm_n53, gm_n2815, gm_n50);
	nor (gm_n5107, gm_n81, gm_n46, in_15, gm_n5106, gm_n47);
	nand (gm_n5108, in_21, gm_n45, in_19, gm_n5107);
	nand (gm_n5109, in_11, in_10, in_9, gm_n4119, gm_n48);
	nor (gm_n5110, gm_n63, in_14, in_13, gm_n5109, in_16);
	nand (gm_n5111, in_19, in_18, in_17, gm_n5110, gm_n45);
	nor (gm_n5112, gm_n5111, in_21);
	nor (gm_n5113, gm_n48, in_11, in_10, gm_n3773, in_13);
	nand (gm_n5114, in_16, gm_n63, in_14, gm_n5113, in_17);
	nor (gm_n5115, in_20, in_19, in_18, gm_n5114, in_21);
	nor (gm_n5116, gm_n3884, gm_n52, in_9);
	and (gm_n5117, gm_n49, gm_n48, in_11, gm_n5116);
	nand (gm_n5118, in_16, in_15, gm_n50, gm_n5117, in_17);
	nor (gm_n5119, gm_n45, in_19, in_18, gm_n5118, in_21);
	nand (gm_n5120, gm_n53, in_10, in_9, gm_n3856, in_12);
	nor (gm_n5121, in_15, in_14, in_13, gm_n5120, gm_n46);
	nand (gm_n5122, in_19, in_18, in_17, gm_n5121, gm_n45);
	nor (gm_n5123, gm_n5122, in_21);
	nand (gm_n5124, in_15, in_14, in_13, gm_n1482, gm_n46);
	nor (gm_n5125, gm_n62, gm_n47, gm_n81, gm_n5124, in_20);
	nand (gm_n5126, gm_n5125, in_21);
	nand (gm_n5127, in_13, gm_n48, gm_n53, gm_n3651, in_14);
	nor (gm_n5128, in_17, in_16, gm_n63, gm_n5127, in_18);
	nand (gm_n5129, in_21, gm_n45, gm_n62, gm_n5128);
	nand (gm_n5130, gm_n63, in_14, gm_n49, gm_n4389, gm_n46);
	nor (gm_n5131, in_19, gm_n47, gm_n81, gm_n5130, gm_n45);
	nand (gm_n5132, gm_n5131, in_21);
	and (gm_n5133, in_9, gm_n64, in_7, gm_n136, in_10);
	nand (gm_n5134, gm_n49, gm_n48, in_11, gm_n5133, in_14);
	nor (gm_n5135, gm_n81, in_16, in_15, gm_n5134, in_18);
	nand (gm_n5136, gm_n71, in_20, gm_n62, gm_n5135);
	nand (gm_n5137, gm_n55, gm_n82, in_5, gm_n1126, in_8);
	nor (gm_n5138, gm_n5137, gm_n51);
	nand (gm_n5139, gm_n48, in_11, in_10, gm_n5138, in_13);
	nor (gm_n5140, in_16, in_15, gm_n50, gm_n5139, gm_n81);
	nand (gm_n5141, gm_n45, gm_n62, gm_n47, gm_n5140, in_21);
	nand (gm_n5142, gm_n5132, gm_n5129, gm_n5126, gm_n5141, gm_n5136);
	nor (gm_n5143, gm_n5119, gm_n5115, gm_n5112, gm_n5142, gm_n5123);
	nand (gm_n5144, gm_n5105, gm_n5102, gm_n5098, gm_n5143, gm_n5108);
	nor (gm_n5145, gm_n5090, gm_n5087, gm_n5083, gm_n5144, gm_n5094);
	nand (gm_n5146, gm_n5077, gm_n5074, gm_n5070, gm_n5145, gm_n5080);
	nor (gm_n5147, gm_n5063, gm_n5059, gm_n5055, gm_n5146, gm_n5067);
	nand (gm_n5148, gm_n5047, gm_n5044, gm_n5040, gm_n5147, gm_n5051);
	nor (gm_n5149, gm_n5033, gm_n5029, gm_n5025, gm_n5148, gm_n5037);
	nand (gm_n5150, gm_n5019, gm_n5017, gm_n5013, gm_n5149, gm_n5022);
	nor (gm_n5151, gm_n5006, gm_n5002, gm_n4998, gm_n5150, gm_n5009);
	nand (gm_n5152, gm_n4991, gm_n4990, gm_n4987, gm_n5151, gm_n4995);
	nor (gm_n5153, gm_n4979, gm_n4975, gm_n4971, gm_n5152, gm_n4983);
	nand (gm_n5154, gm_n4964, gm_n4960, gm_n4957, gm_n5153, gm_n4967);
	nor (gm_n5155, gm_n4953, gm_n4949, gm_n4946, gm_n5154, gm_n4956);
	nand (gm_n5156, gm_n4939, gm_n4935, gm_n4932, gm_n5155, gm_n4942);
	nor (gm_n5157, gm_n4925, gm_n4921, gm_n4917, gm_n5156, gm_n4928);
	nand (gm_n5158, gm_n4910, gm_n4905, gm_n4901, gm_n5157, gm_n4914);
	nor (gm_n5159, gm_n4896, gm_n4894, gm_n4890, gm_n5158, gm_n4899);
	nand (gm_n5160, gm_n4883, gm_n4879, gm_n4875, gm_n5159, gm_n4886);
	nor (gm_n5161, gm_n4867, gm_n4863, gm_n4859, gm_n5160, gm_n4871);
	nand (gm_n5162, gm_n4853, gm_n4849, gm_n4845, gm_n5161, gm_n4856);
	nor (gm_n5163, gm_n4839, gm_n4835, gm_n4832, gm_n5162, gm_n4842);
	nand (gm_n5164, gm_n4825, gm_n4823, gm_n4820, gm_n5163, gm_n4829);
	nor (gm_n5165, gm_n4812, gm_n4808, gm_n4805, gm_n5164, gm_n4816);
	nand (gm_n5166, gm_n4797, gm_n4793, gm_n4789, gm_n5165, gm_n4801);
	nor (gm_n5167, gm_n4783, gm_n4780, gm_n4777, gm_n5166, gm_n4787);
	nand (gm_n5168, gm_n4772, gm_n4768, gm_n4765, gm_n5167, gm_n4774);
	nor (gm_n5169, gm_n4758, gm_n4755, gm_n4751, gm_n5168, gm_n4761);
	nand (gm_n5170, gm_n4744, gm_n4740, gm_n4737, gm_n5169, gm_n4747);
	nor (gm_n5171, gm_n4730, gm_n4727, gm_n4722, gm_n5170, gm_n4734);
	nand (gm_n5172, gm_n4714, gm_n4711, gm_n4708, gm_n5171, gm_n4718);
	nor (gm_n5173, gm_n4702, gm_n4699, gm_n4695, gm_n5172, gm_n4706);
	nand (gm_n5174, gm_n4687, gm_n4684, gm_n4680, gm_n5173, gm_n4691);
	nor (gm_n5175, gm_n4673, gm_n4670, gm_n4666, gm_n5174, gm_n4676);
	nand (gm_n5176, gm_n4660, gm_n4657, gm_n4653, gm_n5175, gm_n4664);
	nor (gm_n5177, gm_n4646, gm_n4643, gm_n4639, gm_n5176, gm_n4649);
	nand (gm_n5178, gm_n4633, gm_n4629, gm_n4625, gm_n5177, gm_n4636);
	nor (out_7, gm_n5178, gm_n4622);
	nand (gm_n5180, gm_n55, in_6, gm_n72, gm_n89);
	nor (gm_n5181, gm_n52, in_9, in_8, gm_n5180);
	and (gm_n5182, gm_n49, in_12, in_11, gm_n5181, in_14);
	nand (gm_n5183, gm_n81, gm_n46, in_15, gm_n5182, gm_n47);
	nor (gm_n5184, in_21, gm_n45, in_19, gm_n5183);
	nor (gm_n5185, gm_n55, in_6, in_5, gm_n167, in_8);
	nand (gm_n5186, gm_n53, in_10, gm_n51, gm_n5185, gm_n48);
	nor (gm_n5187, gm_n63, in_14, gm_n49, gm_n5186, gm_n46);
	nand (gm_n5188, in_19, gm_n47, in_17, gm_n5187, in_20);
	nor (gm_n5189, gm_n5188, gm_n71);
	nand (gm_n5190, in_8, in_7, in_6, gm_n379, in_9);
	nor (gm_n5191, gm_n48, gm_n53, in_10, gm_n5190, in_13);
	nand (gm_n5192, in_16, in_15, in_14, gm_n5191, gm_n81);
	nor (gm_n5193, gm_n45, gm_n62, gm_n47, gm_n5192, in_21);
	nand (gm_n5194, in_11, in_10, gm_n51, gm_n3606, gm_n48);
	nor (gm_n5195, gm_n63, gm_n50, in_13, gm_n5194, gm_n46);
	nand (gm_n5196, gm_n62, in_18, in_17, gm_n5195, in_20);
	nor (gm_n5197, gm_n5196, in_21);
	nor (gm_n5198, in_11, gm_n52, in_9, gm_n1035, in_12);
	nand (gm_n5199, in_15, gm_n50, gm_n49, gm_n5198, in_16);
	nor (gm_n5200, gm_n62, gm_n47, gm_n81, gm_n5199, in_20);
	nand (gm_n5201, gm_n5200, in_21);
	nor (gm_n5202, in_9, in_8, in_7, gm_n897, gm_n52);
	nand (gm_n5203, in_13, gm_n48, gm_n53, gm_n5202, gm_n50);
	nor (gm_n5204, gm_n81, gm_n46, gm_n63, gm_n5203, in_18);
	nand (gm_n5205, in_21, in_20, gm_n62, gm_n5204);
	and (gm_n5206, gm_n64, in_7, gm_n82, gm_n2640, in_9);
	nand (gm_n5207, in_12, gm_n53, gm_n52, gm_n5206, gm_n49);
	nor (gm_n5208, in_16, gm_n63, gm_n50, gm_n5207, in_17);
	nand (gm_n5209, gm_n45, gm_n62, gm_n47, gm_n5208, in_21);
	and (gm_n5210, gm_n53, in_10, gm_n51, gm_n1459);
	nand (gm_n5211, gm_n50, in_13, in_12, gm_n5210, in_15);
	nor (gm_n5212, in_18, in_17, gm_n46, gm_n5211, in_19);
	nand (gm_n5213, gm_n5212, in_21, gm_n45);
	nor (gm_n5214, in_12, gm_n53, in_10, gm_n1430, gm_n49);
	nand (gm_n5215, in_16, gm_n63, gm_n50, gm_n5214, gm_n81);
	nor (gm_n5216, gm_n45, in_19, gm_n47, gm_n5215, gm_n71);
	nand (gm_n5217, gm_n46, in_15, in_14, gm_n3786, gm_n81);
	nor (gm_n5218, gm_n45, in_19, gm_n47, gm_n5217, gm_n71);
	and (gm_n5219, gm_n49, gm_n48, in_11, gm_n2947, gm_n50);
	nand (gm_n5220, gm_n81, gm_n46, gm_n63, gm_n5219, gm_n47);
	nor (gm_n5221, gm_n71, in_20, gm_n62, gm_n5220);
	and (gm_n5222, gm_n50, in_13, gm_n48, gm_n3602, in_15);
	nand (gm_n5223, in_18, in_17, gm_n46, gm_n5222, in_19);
	nor (gm_n5224, gm_n5223, gm_n71, in_20);
	and (gm_n5225, gm_n53, in_10, in_9, gm_n3519);
	nand (gm_n5226, gm_n50, gm_n49, gm_n48, gm_n5225, gm_n63);
	nor (gm_n5227, gm_n47, gm_n81, gm_n46, gm_n5226, gm_n62);
	nand (gm_n5228, gm_n5227, in_21, gm_n45);
	and (gm_n5229, gm_n53, in_10, gm_n51, gm_n1555, gm_n48);
	nand (gm_n5230, gm_n63, in_14, in_13, gm_n5229, gm_n46);
	nor (gm_n5231, gm_n62, gm_n47, gm_n81, gm_n5230, in_20);
	nand (gm_n5232, gm_n5231, in_21);
	nand (gm_n5233, gm_n63, in_14, gm_n49, gm_n3179, gm_n46);
	nor (gm_n5234, gm_n62, in_18, gm_n81, gm_n5233, gm_n45);
	nand (gm_n5235, gm_n5234, gm_n71);
	nand (gm_n5236, gm_n48, in_11, in_10, gm_n380, gm_n49);
	nor (gm_n5237, gm_n46, gm_n63, in_14, gm_n5236, gm_n81);
	nand (gm_n5238, gm_n45, in_19, gm_n47, gm_n5237, in_21);
	nor (gm_n5239, gm_n63, in_14, in_13, gm_n126);
	nand (gm_n5240, gm_n47, gm_n81, gm_n46, gm_n5239, in_19);
	nor (gm_n5241, gm_n5240, in_21, gm_n45);
	nor (gm_n5242, gm_n49, in_12, in_11, gm_n1848, in_14);
	nand (gm_n5243, in_17, in_16, in_15, gm_n5242, gm_n47);
	nor (gm_n5244, in_21, gm_n45, in_19, gm_n5243);
	nor (gm_n5245, in_12, gm_n53, gm_n52, gm_n4362, in_13);
	nand (gm_n5246, gm_n46, gm_n63, gm_n50, gm_n5245, gm_n81);
	nor (gm_n5247, gm_n45, in_19, in_18, gm_n5246, gm_n71);
	and (gm_n5248, in_11, in_10, gm_n51, gm_n494, gm_n48);
	and (gm_n5249, in_15, gm_n50, in_13, gm_n5248, in_16);
	nand (gm_n5250, gm_n62, in_18, in_17, gm_n5249, gm_n45);
	nor (gm_n5251, gm_n5250, in_21);
	nand (gm_n5252, gm_n55, in_6, in_5, gm_n284, gm_n64);
	nor (gm_n5253, in_11, gm_n52, gm_n51, gm_n5252, gm_n48);
	nand (gm_n5254, in_15, in_14, in_13, gm_n5253, in_16);
	nor (gm_n5255, in_19, gm_n47, in_17, gm_n5254, in_20);
	nand (gm_n5256, gm_n5255, in_21);
	nand (gm_n5257, gm_n48, in_11, in_10, gm_n427, in_13);
	nor (gm_n5258, gm_n46, in_15, in_14, gm_n5257, gm_n81);
	nand (gm_n5259, gm_n45, in_19, in_18, gm_n5258, in_21);
	nand (gm_n5260, in_12, in_11, gm_n52, gm_n2877, in_13);
	nor (gm_n5261, in_16, gm_n63, gm_n50, gm_n5260, in_17);
	nand (gm_n5262, in_20, gm_n62, gm_n47, gm_n5261, gm_n71);
	nand (gm_n5263, in_7, gm_n82, in_5, gm_n493, in_8);
	nor (gm_n5264, gm_n53, in_10, gm_n51, gm_n5263);
	nand (gm_n5265, gm_n50, gm_n49, gm_n48, gm_n5264, gm_n63);
	nor (gm_n5266, in_18, in_17, gm_n46, gm_n5265, in_19);
	nand (gm_n5267, gm_n5266, in_21, in_20);
	or (gm_n5268, gm_n64, gm_n55, gm_n82, gm_n156, gm_n51);
	nor (gm_n5269, in_12, in_11, gm_n52, gm_n5268, in_13);
	nand (gm_n5270, gm_n46, gm_n63, gm_n50, gm_n5269, in_17);
	nor (gm_n5271, gm_n45, in_19, gm_n47, gm_n5270, gm_n71);
	nand (gm_n5272, gm_n52, in_9, in_8, gm_n1608);
	nor (gm_n5273, in_13, gm_n48, in_11, gm_n5272, in_14);
	nand (gm_n5274, in_17, gm_n46, in_15, gm_n5273, gm_n47);
	nor (gm_n5275, in_21, gm_n45, gm_n62, gm_n5274);
	and (gm_n5276, in_14, gm_n49, gm_n48, gm_n4214, in_15);
	nand (gm_n5277, gm_n47, in_17, gm_n46, gm_n5276, in_19);
	nor (gm_n5278, gm_n5277, gm_n71, gm_n45);
	nor (gm_n5279, in_11, in_10, gm_n51, gm_n2546);
	and (gm_n5280, gm_n50, gm_n49, in_12, gm_n5279, in_15);
	nand (gm_n5281, gm_n47, gm_n81, gm_n46, gm_n5280, gm_n62);
	nor (gm_n5282, gm_n5281, gm_n71, gm_n45);
	or (gm_n5283, in_12, in_11, in_10, gm_n1900, gm_n49);
	nor (gm_n5284, in_16, gm_n63, in_14, gm_n5283, gm_n81);
	nand (gm_n5285, in_20, in_19, gm_n47, gm_n5284, gm_n71);
	nand (gm_n5286, in_15, gm_n50, in_13, gm_n3628, in_16);
	nor (gm_n5287, gm_n62, in_18, gm_n81, gm_n5286, in_20);
	nand (gm_n5288, gm_n5287, gm_n71);
	and (gm_n5289, gm_n3768, gm_n52, gm_n51);
	nand (gm_n5290, gm_n49, gm_n48, gm_n53, gm_n5289, gm_n50);
	nor (gm_n5291, gm_n81, in_16, gm_n63, gm_n5290, in_18);
	nand (gm_n5292, gm_n71, in_20, in_19, gm_n5291);
	nand (gm_n5293, gm_n50, in_13, gm_n48, gm_n2240, gm_n63);
	nor (gm_n5294, in_18, in_17, in_16, gm_n5293, in_19);
	nand (gm_n5295, gm_n5294, in_21, gm_n45);
	nand (gm_n5296, in_18, gm_n81, in_16, gm_n370, in_19);
	nor (gm_n5297, gm_n5296, gm_n71, gm_n45);
	nand (gm_n5298, in_7, gm_n82, gm_n72, gm_n598, in_8);
	or (gm_n5299, gm_n53, gm_n52, gm_n51, gm_n5298, in_12);
	nor (gm_n5300, in_15, in_14, gm_n49, gm_n5299, in_16);
	nand (gm_n5301, gm_n62, gm_n47, gm_n81, gm_n5300, gm_n45);
	nor (gm_n5302, gm_n5301, gm_n71);
	nand (gm_n5303, gm_n81, in_16, gm_n63, gm_n2272, gm_n47);
	nor (gm_n5304, in_21, gm_n45, in_19, gm_n5303);
	nor (gm_n5305, gm_n1629, gm_n52, gm_n51);
	and (gm_n5306, in_13, gm_n48, in_11, gm_n5305);
	nand (gm_n5307, in_16, gm_n63, in_14, gm_n5306, gm_n81);
	nor (gm_n5308, in_20, gm_n62, gm_n47, gm_n5307, in_21);
	nand (gm_n5309, gm_n48, in_11, gm_n52, gm_n1941, gm_n49);
	nor (gm_n5310, gm_n46, gm_n63, in_14, gm_n5309, gm_n81);
	nand (gm_n5311, in_20, gm_n62, gm_n47, gm_n5310, gm_n71);
	nand (gm_n5312, in_12, gm_n53, gm_n52, gm_n2619, gm_n49);
	nor (gm_n5313, in_16, in_15, in_14, gm_n5312, in_17);
	nand (gm_n5314, gm_n45, gm_n62, gm_n47, gm_n5313, in_21);
	nor (gm_n5315, gm_n3743, gm_n52, gm_n51);
	nand (gm_n5316, in_13, in_12, gm_n53, gm_n5315, gm_n50);
	nor (gm_n5317, gm_n81, in_16, gm_n63, gm_n5316, gm_n47);
	nand (gm_n5318, in_21, in_20, gm_n62, gm_n5317);
	nand (gm_n5319, in_12, in_11, in_10, gm_n889, in_13);
	nor (gm_n5320, in_16, gm_n63, gm_n50, gm_n5319, in_17);
	nand (gm_n5321, in_20, in_19, gm_n47, gm_n5320, gm_n71);
	or (gm_n5322, in_8, in_7, gm_n82, gm_n1429, gm_n51);
	nor (gm_n5323, gm_n48, in_11, gm_n52, gm_n5322, gm_n49);
	nand (gm_n5324, in_16, in_15, gm_n50, gm_n5323, in_17);
	nor (gm_n5325, in_20, in_19, gm_n47, gm_n5324, in_21);
	nand (gm_n5326, in_8, in_7, gm_n82, gm_n1075, gm_n51);
	nor (gm_n5327, gm_n48, in_11, gm_n52, gm_n5326, gm_n49);
	nand (gm_n5328, in_16, gm_n63, gm_n50, gm_n5327, gm_n81);
	nor (gm_n5329, in_20, in_19, in_18, gm_n5328, gm_n71);
	nor (gm_n5330, in_13, gm_n48, in_11, gm_n1884, in_14);
	nand (gm_n5331, gm_n81, in_16, gm_n63, gm_n5330, gm_n47);
	nor (gm_n5332, gm_n71, gm_n45, gm_n62, gm_n5331);
	nor (gm_n5333, in_12, in_11, in_10, gm_n1372, gm_n49);
	nand (gm_n5334, in_16, gm_n63, gm_n50, gm_n5333, gm_n81);
	nor (gm_n5335, in_20, gm_n62, gm_n47, gm_n5334, gm_n71);
	nor (gm_n5336, in_11, gm_n52, in_9, gm_n1439, gm_n48);
	nand (gm_n5337, gm_n63, in_14, gm_n49, gm_n5336, gm_n46);
	nor (gm_n5338, in_19, gm_n47, gm_n81, gm_n5337, gm_n45);
	nand (gm_n5339, gm_n5338, in_21);
	nor (gm_n5340, in_7, in_6, in_5, gm_n483, gm_n64);
	and (gm_n5341, gm_n53, gm_n52, gm_n51, gm_n5340, in_12);
	nand (gm_n5342, in_15, gm_n50, in_13, gm_n5341, in_16);
	nor (gm_n5343, gm_n62, in_18, in_17, gm_n5342, in_20);
	nand (gm_n5344, gm_n5343, in_21);
	nand (gm_n5345, in_12, gm_n53, gm_n52, gm_n1755, in_13);
	nor (gm_n5346, in_16, gm_n63, gm_n50, gm_n5345, gm_n81);
	nand (gm_n5347, in_20, in_19, in_18, gm_n5346, in_21);
	nand (gm_n5348, gm_n63, gm_n50, in_13, gm_n3735, gm_n46);
	nor (gm_n5349, in_19, gm_n47, gm_n81, gm_n5348, in_20);
	nand (gm_n5350, gm_n5349, in_21);
	and (gm_n5351, gm_n52, gm_n51, gm_n64, gm_n1093, in_11);
	and (gm_n5352, gm_n50, in_13, gm_n48, gm_n5351, in_15);
	nand (gm_n5353, gm_n47, gm_n81, gm_n46, gm_n5352, gm_n62);
	nor (gm_n5354, gm_n5353, in_21, in_20);
	and (gm_n5355, in_12, gm_n53, in_10, gm_n4876, gm_n49);
	nand (gm_n5356, in_16, in_15, in_14, gm_n5355, in_17);
	nor (gm_n5357, gm_n45, gm_n62, gm_n47, gm_n5356, in_21);
	and (gm_n5358, in_10, gm_n51, gm_n64, gm_n316);
	and (gm_n5359, gm_n49, in_12, gm_n53, gm_n5358, in_14);
	nand (gm_n5360, gm_n81, in_16, gm_n63, gm_n5359, gm_n47);
	nor (gm_n5361, gm_n71, gm_n45, gm_n62, gm_n5360);
	nand (gm_n5362, gm_n53, gm_n52, in_9, gm_n458);
	nor (gm_n5363, gm_n50, gm_n49, in_12, gm_n5362, gm_n63);
	nand (gm_n5364, in_18, gm_n81, in_16, gm_n5363, gm_n62);
	nor (gm_n5365, gm_n5364, in_21, in_20);
	nand (gm_n5366, gm_n48, in_11, in_10, gm_n1700, in_13);
	nor (gm_n5367, gm_n46, gm_n63, in_14, gm_n5366, in_17);
	nand (gm_n5368, gm_n45, in_19, in_18, gm_n5367, gm_n71);
	nand (gm_n5369, gm_n49, gm_n48, in_11, gm_n4681, in_14);
	nor (gm_n5370, gm_n81, in_16, gm_n63, gm_n5369, gm_n47);
	nand (gm_n5371, gm_n71, gm_n45, in_19, gm_n5370);
	nand (gm_n5372, gm_n45, gm_n62, gm_n47, gm_n2348, in_21);
	and (gm_n5373, gm_n46, gm_n63, in_14, gm_n4076, in_17);
	nand (gm_n5374, gm_n45, in_19, gm_n47, gm_n5373, in_21);
	nor (gm_n5375, gm_n64, gm_n55, gm_n82, gm_n199, gm_n51);
	and (gm_n5376, gm_n48, gm_n53, in_10, gm_n5375, gm_n49);
	nand (gm_n5377, in_16, gm_n63, in_14, gm_n5376, gm_n81);
	nor (gm_n5378, gm_n45, gm_n62, in_18, gm_n5377, gm_n71);
	or (gm_n5379, in_7, gm_n82, gm_n72, gm_n167);
	or (gm_n5380, in_10, gm_n51, in_8, gm_n5379, gm_n53);
	nor (gm_n5381, in_14, in_13, gm_n48, gm_n5380, in_15);
	nand (gm_n5382, in_18, gm_n81, in_16, gm_n5381, gm_n62);
	nor (gm_n5383, gm_n5382, gm_n71, gm_n45);
	nand (gm_n5384, gm_n53, gm_n52, in_9, gm_n2088, gm_n48);
	nor (gm_n5385, in_15, in_14, gm_n49, gm_n5384, gm_n46);
	nand (gm_n5386, gm_n62, gm_n47, gm_n81, gm_n5385, in_20);
	nor (gm_n5387, gm_n5386, in_21);
	or (gm_n5388, in_11, gm_n52, in_9, gm_n2114, gm_n48);
	nor (gm_n5389, gm_n63, gm_n50, in_13, gm_n5388, in_16);
	nand (gm_n5390, gm_n62, in_18, in_17, gm_n5389, in_20);
	nor (gm_n5391, gm_n5390, gm_n71);
	nor (gm_n5392, gm_n53, in_10, in_9, gm_n5263);
	nand (gm_n5393, in_14, in_13, gm_n48, gm_n5392, in_15);
	nor (gm_n5394, in_18, gm_n81, in_16, gm_n5393, gm_n62);
	nand (gm_n5395, gm_n5394, gm_n71, gm_n45);
	nand (gm_n5396, gm_n48, gm_n53, gm_n52, gm_n4072, in_13);
	nor (gm_n5397, in_16, in_15, gm_n50, gm_n5396, gm_n81);
	nand (gm_n5398, gm_n45, gm_n62, gm_n47, gm_n5397, in_21);
	nand (gm_n5399, in_7, gm_n82, in_5, gm_n1126, in_8);
	nor (gm_n5400, gm_n5399, gm_n51);
	nand (gm_n5401, in_12, gm_n53, gm_n52, gm_n5400, in_13);
	nor (gm_n5402, in_16, gm_n63, gm_n50, gm_n5401, gm_n81);
	nand (gm_n5403, in_20, gm_n62, gm_n47, gm_n5402, gm_n71);
	nand (gm_n5404, gm_n48, in_11, in_10, gm_n5400, in_13);
	nor (gm_n5405, gm_n46, in_15, in_14, gm_n5404, in_17);
	nand (gm_n5406, gm_n45, in_19, in_18, gm_n5405, in_21);
	nor (gm_n5407, gm_n63, gm_n50, in_13, gm_n3215, in_16);
	nand (gm_n5408, gm_n62, gm_n47, in_17, gm_n5407, gm_n45);
	nor (gm_n5409, gm_n5408, gm_n71);
	nor (gm_n5410, gm_n53, in_10, in_9, gm_n583, in_12);
	and (gm_n5411, in_15, in_14, in_13, gm_n5410, in_16);
	nand (gm_n5412, in_19, gm_n47, gm_n81, gm_n5411, gm_n45);
	nor (gm_n5413, gm_n5412, gm_n71);
	nand (gm_n5414, gm_n1634, gm_n52, gm_n51);
	nor (gm_n5415, gm_n49, gm_n48, in_11, gm_n5414, in_14);
	nand (gm_n5416, gm_n81, gm_n46, in_15, gm_n5415, gm_n47);
	nor (gm_n5417, in_21, in_20, in_19, gm_n5416);
	or (gm_n5418, in_11, gm_n52, gm_n51, gm_n607);
	nor (gm_n5419, in_14, in_13, in_12, gm_n5418, gm_n63);
	nand (gm_n5420, gm_n47, in_17, gm_n46, gm_n5419, in_19);
	nor (gm_n5421, gm_n5420, in_21, gm_n45);
	nor (gm_n5422, gm_n55, in_6, gm_n72, gm_n867, gm_n64);
	nand (gm_n5423, gm_n5422, gm_n52, gm_n51);
	nor (gm_n5424, in_13, in_12, gm_n53, gm_n5423);
	and (gm_n5425, in_16, gm_n63, gm_n50, gm_n5424, in_17);
	nand (gm_n5426, in_20, in_19, in_18, gm_n5425, gm_n71);
	nand (gm_n5427, in_14, in_13, in_12, gm_n323, in_15);
	nor (gm_n5428, gm_n47, in_17, in_16, gm_n5427, in_19);
	nand (gm_n5429, gm_n5428, in_21, in_20);
	nand (gm_n5430, gm_n48, gm_n53, gm_n52, gm_n1780, in_13);
	nor (gm_n5431, gm_n46, in_15, gm_n50, gm_n5430, in_17);
	nand (gm_n5432, in_20, gm_n62, in_18, gm_n5431, gm_n71);
	and (gm_n5433, gm_n53, gm_n52, in_9, gm_n1302, gm_n48);
	nand (gm_n5434, gm_n63, in_14, in_13, gm_n5433, gm_n46);
	nor (gm_n5435, in_19, in_18, gm_n81, gm_n5434, in_20);
	nand (gm_n5436, gm_n5435, in_21);
	nor (gm_n5437, in_12, gm_n53, gm_n52, gm_n4530, in_13);
	nand (gm_n5438, in_16, gm_n63, gm_n50, gm_n5437, gm_n81);
	nor (gm_n5439, in_20, gm_n62, in_18, gm_n5438, in_21);
	and (gm_n5440, gm_n48, in_11, in_10, gm_n1700, gm_n49);
	nand (gm_n5441, in_16, in_15, gm_n50, gm_n5440, gm_n81);
	nor (gm_n5442, gm_n45, in_19, gm_n47, gm_n5441, in_21);
	and (gm_n5443, in_12, in_11, in_10, gm_n1385, in_13);
	nand (gm_n5444, in_16, gm_n63, gm_n50, gm_n5443, gm_n81);
	nor (gm_n5445, gm_n45, in_19, in_18, gm_n5444, in_21);
	nand (gm_n5446, in_16, gm_n63, gm_n50, gm_n3040, in_17);
	nor (gm_n5447, in_20, in_19, in_18, gm_n5446, in_21);
	or (gm_n5448, in_12, gm_n53, gm_n52, gm_n766, in_13);
	nor (gm_n5449, gm_n46, in_15, gm_n50, gm_n5448, gm_n81);
	nand (gm_n5450, in_20, in_19, in_18, gm_n5449, in_21);
	and (gm_n5451, gm_n3299, in_10, in_9);
	nand (gm_n5452, in_13, in_12, gm_n53, gm_n5451, in_14);
	nor (gm_n5453, gm_n81, in_16, gm_n63, gm_n5452, in_18);
	nand (gm_n5454, gm_n71, gm_n45, in_19, gm_n5453);
	nand (gm_n5455, gm_n50, gm_n49, in_12, gm_n58, in_15);
	nor (gm_n5456, in_18, gm_n81, gm_n46, gm_n5455, in_19);
	nand (gm_n5457, gm_n5456, in_21, gm_n45);
	and (gm_n5458, in_8, gm_n55, in_6, gm_n374, in_9);
	nand (gm_n5459, gm_n48, in_11, in_10, gm_n5458, in_13);
	nor (gm_n5460, gm_n46, in_15, gm_n50, gm_n5459, in_17);
	nand (gm_n5461, gm_n45, gm_n62, gm_n47, gm_n5460, gm_n71);
	nor (gm_n5462, gm_n63, in_14, gm_n49, gm_n1294, gm_n46);
	nand (gm_n5463, in_19, gm_n47, gm_n81, gm_n5462, in_20);
	nor (gm_n5464, gm_n5463, gm_n71);
	nor (gm_n5465, gm_n48, in_11, gm_n52, gm_n1900, gm_n49);
	nand (gm_n5466, in_16, gm_n63, gm_n50, gm_n5465, gm_n81);
	nor (gm_n5467, gm_n45, gm_n62, in_18, gm_n5466, in_21);
	and (gm_n5468, gm_n1550, in_10, in_9);
	and (gm_n5469, gm_n49, in_12, gm_n53, gm_n5468, in_14);
	nand (gm_n5470, gm_n81, gm_n46, gm_n63, gm_n5469, gm_n47);
	nor (gm_n5471, in_21, gm_n45, gm_n62, gm_n5470);
	nor (gm_n5472, gm_n53, in_10, gm_n51, gm_n916, in_12);
	nand (gm_n5473, gm_n5472, in_14, gm_n49);
	or (gm_n5474, gm_n81, gm_n46, gm_n63, gm_n5473, in_18);
	nor (gm_n5475, in_21, in_20, gm_n62, gm_n5474);
	nor (gm_n5476, gm_n53, gm_n52, in_9, gm_n3697, gm_n48);
	nand (gm_n5477, gm_n63, gm_n50, gm_n49, gm_n5476, gm_n46);
	nor (gm_n5478, gm_n62, in_18, gm_n81, gm_n5477, in_20);
	nand (gm_n5479, gm_n5478, gm_n71);
	nand (gm_n5480, gm_n48, in_11, in_10, gm_n1692, in_13);
	nor (gm_n5481, in_16, in_15, gm_n50, gm_n5480, gm_n81);
	nand (gm_n5482, in_20, gm_n62, gm_n47, gm_n5481, gm_n71);
	or (gm_n5483, gm_n49, in_12, in_11, gm_n722, in_14);
	nor (gm_n5484, in_17, gm_n46, in_15, gm_n5483, gm_n47);
	nand (gm_n5485, gm_n71, in_20, gm_n62, gm_n5484);
	nand (gm_n5486, gm_n50, in_13, gm_n48, gm_n4887, gm_n63);
	nor (gm_n5487, gm_n47, gm_n81, in_16, gm_n5486, gm_n62);
	nand (gm_n5488, gm_n5487, in_21, in_20);
	nand (gm_n5489, gm_n53, in_10, gm_n51, gm_n494, in_12);
	nor (gm_n5490, gm_n63, in_14, in_13, gm_n5489, gm_n46);
	nand (gm_n5491, gm_n62, gm_n47, gm_n81, gm_n5490, in_20);
	nor (gm_n5492, gm_n5491, in_21);
	nand (gm_n5493, in_11, gm_n52, gm_n51, gm_n1111, gm_n48);
	nor (gm_n5494, in_15, gm_n50, gm_n49, gm_n5493, in_16);
	nand (gm_n5495, in_19, in_18, gm_n81, gm_n5494, gm_n45);
	nor (gm_n5496, gm_n5495, in_21);
	nor (gm_n5497, gm_n49, in_12, in_11, gm_n2288, gm_n50);
	nand (gm_n5498, in_17, in_16, in_15, gm_n5497, gm_n47);
	nor (gm_n5499, in_21, in_20, in_19, gm_n5498);
	nand (gm_n5500, gm_n62, in_18, gm_n81, gm_n3156, in_20);
	nor (gm_n5501, gm_n5500, in_21);
	nor (gm_n5502, in_11, in_10, in_9, gm_n1709);
	nand (gm_n5503, in_14, in_13, in_12, gm_n5502, gm_n63);
	nor (gm_n5504, gm_n47, in_17, gm_n46, gm_n5503, gm_n62);
	nand (gm_n5505, gm_n5504, in_21, gm_n45);
	nand (gm_n5506, gm_n49, in_12, gm_n53, gm_n579);
	nor (gm_n5507, in_16, in_15, gm_n50, gm_n5506, gm_n81);
	nand (gm_n5508, gm_n45, gm_n62, in_18, gm_n5507, gm_n71);
	and (gm_n5509, gm_n1714, gm_n52, gm_n51);
	nand (gm_n5510, in_13, gm_n48, in_11, gm_n5509, in_14);
	nor (gm_n5511, in_17, in_16, in_15, gm_n5510, in_18);
	nand (gm_n5512, in_21, gm_n45, in_19, gm_n5511);
	nand (gm_n5513, in_14, in_13, in_12, gm_n1470, gm_n63);
	nor (gm_n5514, in_18, gm_n81, gm_n46, gm_n5513, in_19);
	nand (gm_n5515, gm_n5514, gm_n71, gm_n45);
	nor (gm_n5516, in_12, in_11, gm_n52, gm_n1599, in_13);
	nand (gm_n5517, gm_n46, in_15, gm_n50, gm_n5516, in_17);
	nor (gm_n5518, gm_n45, in_19, gm_n47, gm_n5517, in_21);
	nand (gm_n5519, gm_n717, in_9);
	nor (gm_n5520, gm_n48, in_11, gm_n52, gm_n5519, gm_n49);
	nand (gm_n5521, gm_n46, in_15, gm_n50, gm_n5520, in_17);
	nor (gm_n5522, gm_n45, gm_n62, gm_n47, gm_n5521, in_21);
	nor (gm_n5523, in_11, in_10, gm_n51, gm_n1750, in_12);
	and (gm_n5524, gm_n63, in_14, in_13, gm_n5523, in_16);
	nand (gm_n5525, in_19, gm_n47, gm_n81, gm_n5524, in_20);
	nor (gm_n5526, gm_n5525, gm_n71);
	nand (gm_n5527, gm_n64, gm_n55, gm_n82, gm_n374, in_9);
	nor (gm_n5528, in_12, gm_n53, in_10, gm_n5527, in_13);
	nand (gm_n5529, gm_n46, gm_n63, in_14, gm_n5528, in_17);
	nor (gm_n5530, gm_n45, gm_n62, in_18, gm_n5529, gm_n71);
	nor (gm_n5531, gm_n285, in_10, in_9);
	nand (gm_n5532, in_13, in_12, in_11, gm_n5531, gm_n50);
	nor (gm_n5533, in_17, in_16, gm_n63, gm_n5532, gm_n47);
	nand (gm_n5534, gm_n71, gm_n45, gm_n62, gm_n5533);
	nor (gm_n5535, gm_n53, gm_n52, in_9, gm_n247, gm_n48);
	nand (gm_n5536, gm_n63, gm_n50, gm_n49, gm_n5535, gm_n46);
	nor (gm_n5537, gm_n62, in_18, gm_n81, gm_n5536, in_20);
	nand (gm_n5538, gm_n5537, in_21);
	and (gm_n5539, gm_n53, in_10, gm_n51, gm_n3519, in_12);
	nand (gm_n5540, gm_n63, gm_n50, in_13, gm_n5539, gm_n46);
	nor (gm_n5541, in_19, gm_n47, in_17, gm_n5540, in_20);
	nand (gm_n5542, gm_n5541, gm_n71);
	and (gm_n5543, in_16, gm_n63, gm_n50, gm_n1781, gm_n81);
	nand (gm_n5544, gm_n45, in_19, gm_n47, gm_n5543, gm_n71);
	or (gm_n5545, gm_n53, in_10, in_9, gm_n410, gm_n48);
	nor (gm_n5546, in_15, gm_n50, in_13, gm_n5545, gm_n46);
	nand (gm_n5547, in_19, in_18, gm_n81, gm_n5546, gm_n45);
	nor (gm_n5548, gm_n5547, in_21);
	or (gm_n5549, gm_n4153, gm_n51);
	nor (gm_n5550, in_12, in_11, in_10, gm_n5549, gm_n49);
	nand (gm_n5551, gm_n46, gm_n63, gm_n50, gm_n5550, in_17);
	nor (gm_n5552, in_20, gm_n62, gm_n47, gm_n5551, gm_n71);
	nand (gm_n5553, in_11, gm_n52, in_9, gm_n1183, in_12);
	nor (gm_n5554, gm_n63, gm_n50, gm_n49, gm_n5553);
	nand (gm_n5555, gm_n47, in_17, gm_n46, gm_n5554, in_19);
	nor (gm_n5556, gm_n5555, gm_n71, gm_n45);
	nand (gm_n5557, in_17, in_16, gm_n63, gm_n4237, in_18);
	nor (gm_n5558, gm_n71, gm_n45, gm_n62, gm_n5557);
	nand (gm_n5559, in_13, in_12, gm_n53, gm_n3905, gm_n50);
	nor (gm_n5560, gm_n81, in_16, gm_n63, gm_n5559, in_18);
	nand (gm_n5561, gm_n71, gm_n45, gm_n62, gm_n5560);
	and (gm_n5562, gm_n1714, gm_n52, in_9);
	nand (gm_n5563, gm_n49, gm_n48, in_11, gm_n5562, in_14);
	nor (gm_n5564, gm_n81, in_16, in_15, gm_n5563, in_18);
	nand (gm_n5565, gm_n71, gm_n45, in_19, gm_n5564);
	nand (gm_n5566, gm_n49, in_12, gm_n53, gm_n3687, gm_n50);
	nor (gm_n5567, in_17, gm_n46, in_15, gm_n5566, gm_n47);
	nand (gm_n5568, gm_n71, gm_n45, in_19, gm_n5567);
	and (gm_n5569, gm_n53, gm_n52, in_9, gm_n700, gm_n48);
	nand (gm_n5570, gm_n63, gm_n50, gm_n49, gm_n5569, in_16);
	nor (gm_n5571, gm_n62, in_18, in_17, gm_n5570, gm_n45);
	nand (gm_n5572, gm_n5571, gm_n71);
	nor (gm_n5573, in_13, in_12, in_11, gm_n1920, in_14);
	nand (gm_n5574, gm_n81, gm_n46, in_15, gm_n5573, gm_n47);
	nor (gm_n5575, in_21, gm_n45, gm_n62, gm_n5574);
	nand (gm_n5576, gm_n52, in_9, gm_n64, gm_n663, gm_n53);
	nor (gm_n5577, gm_n50, in_13, in_12, gm_n5576, gm_n63);
	nand (gm_n5578, gm_n47, in_17, gm_n46, gm_n5577, gm_n62);
	nor (gm_n5579, gm_n5578, gm_n71, in_20);
	nor (gm_n5580, in_15, gm_n50, gm_n49, gm_n3114, gm_n46);
	nand (gm_n5581, gm_n62, in_18, gm_n81, gm_n5580, gm_n45);
	nor (gm_n5582, gm_n5581, in_21);
	and (gm_n5583, in_14, gm_n49, in_12, gm_n3128, in_15);
	nand (gm_n5584, in_18, gm_n81, gm_n46, gm_n5583, in_19);
	nor (gm_n5585, gm_n5584, in_21, gm_n45);
	or (gm_n5586, in_7, in_6, in_5, gm_n321, in_8);
	nor (gm_n5587, gm_n53, in_10, in_9, gm_n5586);
	nand (gm_n5588, in_14, gm_n49, gm_n48, gm_n5587, in_15);
	nor (gm_n5589, in_18, gm_n81, gm_n46, gm_n5588, gm_n62);
	nand (gm_n5590, gm_n5589, in_21, in_20);
	and (gm_n5591, gm_n3489, gm_n52, gm_n51);
	and (gm_n5592, in_13, in_12, in_11, gm_n5591);
	and (gm_n5593, gm_n46, in_15, in_14, gm_n5592, in_17);
	nand (gm_n5594, in_20, in_19, in_18, gm_n5593, in_21);
	nor (gm_n5595, gm_n53, in_10, in_9, gm_n247);
	nand (gm_n5596, gm_n50, in_13, in_12, gm_n5595, in_15);
	nor (gm_n5597, gm_n47, in_17, gm_n46, gm_n5596, gm_n62);
	nand (gm_n5598, gm_n5597, in_21, gm_n45);
	nor (gm_n5599, gm_n47, in_17, in_16, gm_n1737, gm_n62);
	nand (gm_n5600, gm_n5599, in_21, in_20);
	nor (gm_n5601, gm_n1629, in_10, gm_n51);
	and (gm_n5602, gm_n49, gm_n48, in_11, gm_n5601, gm_n50);
	nand (gm_n5603, in_17, gm_n46, in_15, gm_n5602, gm_n47);
	nor (gm_n5604, gm_n71, gm_n45, gm_n62, gm_n5603);
	or (gm_n5605, in_8, gm_n55, gm_n82, gm_n204, in_9);
	nor (gm_n5606, in_12, in_11, gm_n52, gm_n5605, in_13);
	nand (gm_n5607, gm_n46, gm_n63, in_14, gm_n5606, gm_n81);
	nor (gm_n5608, gm_n45, in_19, gm_n47, gm_n5607, in_21);
	and (gm_n5609, in_13, gm_n48, in_11, gm_n3480, gm_n50);
	nand (gm_n5610, gm_n81, gm_n46, gm_n63, gm_n5609, in_18);
	nor (gm_n5611, gm_n71, gm_n45, in_19, gm_n5610);
	nand (gm_n5612, in_11, gm_n52, in_9, gm_n1788, in_12);
	nor (gm_n5613, in_15, in_14, in_13, gm_n5612, in_16);
	nand (gm_n5614, in_19, gm_n47, in_17, gm_n5613, in_20);
	nor (gm_n5615, gm_n5614, gm_n71);
	and (gm_n5616, gm_n297, in_9);
	nand (gm_n5617, in_12, in_11, in_10, gm_n5616, gm_n49);
	nor (gm_n5618, in_16, gm_n63, in_14, gm_n5617, gm_n81);
	nand (gm_n5619, in_20, in_19, gm_n47, gm_n5618, gm_n71);
	nand (gm_n5620, gm_n64, in_7, gm_n82, gm_n2640, gm_n51);
	or (gm_n5621, in_12, in_11, gm_n52, gm_n5620, gm_n49);
	nor (gm_n5622, in_16, in_15, gm_n50, gm_n5621, gm_n81);
	nand (gm_n5623, in_20, gm_n62, gm_n47, gm_n5622, in_21);
	nand (gm_n5624, gm_n48, gm_n53, in_10, gm_n1080, in_13);
	nor (gm_n5625, gm_n46, in_15, gm_n50, gm_n5624, gm_n81);
	nand (gm_n5626, gm_n45, gm_n62, gm_n47, gm_n5625, gm_n71);
	nand (gm_n5627, gm_n48, in_11, in_10, gm_n1966, gm_n49);
	nor (gm_n5628, gm_n46, in_15, gm_n50, gm_n5627, in_17);
	nand (gm_n5629, in_20, in_19, gm_n47, gm_n5628, gm_n71);
	nand (gm_n5630, in_16, in_15, gm_n50, gm_n2878, gm_n81);
	nor (gm_n5631, gm_n45, in_19, gm_n47, gm_n5630, gm_n71);
	nor (gm_n5632, in_12, gm_n53, gm_n52, gm_n97, in_13);
	nand (gm_n5633, gm_n46, in_15, in_14, gm_n5632, in_17);
	nor (gm_n5634, gm_n45, in_19, gm_n47, gm_n5633, in_21);
	nand (gm_n5635, gm_n46, gm_n63, gm_n50, gm_n2658, in_17);
	nor (gm_n5636, gm_n45, gm_n62, gm_n47, gm_n5635, gm_n71);
	or (gm_n5637, in_10, gm_n51, in_8, gm_n478, in_11);
	nor (gm_n5638, in_14, in_13, in_12, gm_n5637, gm_n63);
	nand (gm_n5639, gm_n47, in_17, in_16, gm_n5638, in_19);
	nor (gm_n5640, gm_n5639, gm_n71, in_20);
	nand (gm_n5641, in_13, gm_n48, in_11, gm_n4515, gm_n50);
	nor (gm_n5642, gm_n81, gm_n46, in_15, gm_n5641, in_18);
	nand (gm_n5643, in_21, gm_n45, in_19, gm_n5642);
	nor (gm_n5644, gm_n2849, in_10, in_9);
	nand (gm_n5645, in_13, in_12, gm_n53, gm_n5644, gm_n50);
	nor (gm_n5646, in_17, in_16, gm_n63, gm_n5645, gm_n47);
	nand (gm_n5647, gm_n71, in_20, gm_n62, gm_n5646);
	nand (gm_n5648, gm_n49, in_12, gm_n53, gm_n1311, in_14);
	nor (gm_n5649, gm_n81, gm_n46, in_15, gm_n5648, in_18);
	nand (gm_n5650, in_21, gm_n45, in_19, gm_n5649);
	and (gm_n5651, in_11, gm_n52, in_9, gm_n2508, in_12);
	nand (gm_n5652, gm_n63, gm_n50, gm_n49, gm_n5651, gm_n46);
	nor (gm_n5653, in_19, in_18, in_17, gm_n5652, in_20);
	nand (gm_n5654, gm_n5653, in_21);
	nor (gm_n5655, in_12, gm_n53, in_10, gm_n3245, in_13);
	nand (gm_n5656, gm_n46, gm_n63, in_14, gm_n5655, gm_n81);
	nor (gm_n5657, gm_n45, gm_n62, in_18, gm_n5656, in_21);
	nor (gm_n5658, gm_n49, in_12, in_11, gm_n622, gm_n50);
	nand (gm_n5659, in_17, in_16, in_15, gm_n5658, gm_n47);
	nor (gm_n5660, in_21, in_20, gm_n62, gm_n5659);
	nor (gm_n5661, gm_n5384, in_13);
	nand (gm_n5662, gm_n46, in_15, in_14, gm_n5661, gm_n81);
	nor (gm_n5663, gm_n45, gm_n62, gm_n47, gm_n5662, in_21);
	nand (gm_n5664, in_11, in_10, gm_n51, gm_n1459, in_12);
	nor (gm_n5665, in_15, gm_n50, gm_n49, gm_n5664, in_16);
	nand (gm_n5666, gm_n62, in_18, in_17, gm_n5665, gm_n45);
	nor (gm_n5667, gm_n5666, gm_n71);
	nor (gm_n5668, in_7, in_6, in_5, gm_n643, gm_n64);
	and (gm_n5669, gm_n5668, gm_n52, gm_n51);
	nand (gm_n5670, gm_n49, in_12, gm_n53, gm_n5669, gm_n50);
	nor (gm_n5671, in_17, gm_n46, gm_n63, gm_n5670, in_18);
	nand (gm_n5672, gm_n71, gm_n45, in_19, gm_n5671);
	nand (gm_n5673, gm_n48, in_11, in_10, gm_n747, in_13);
	nor (gm_n5674, gm_n46, gm_n63, gm_n50, gm_n5673, gm_n81);
	nand (gm_n5675, in_20, gm_n62, gm_n47, gm_n5674, in_21);
	nor (gm_n5676, gm_n64, gm_n55, in_6, gm_n103, in_9);
	nand (gm_n5677, gm_n48, in_11, gm_n52, gm_n5676, in_13);
	nor (gm_n5678, gm_n46, in_15, in_14, gm_n5677, gm_n81);
	nand (gm_n5679, gm_n45, gm_n62, gm_n47, gm_n5678, in_21);
	nand (gm_n5680, in_14, gm_n49, in_12, gm_n4080, in_15);
	nor (gm_n5681, in_18, in_17, gm_n46, gm_n5680, gm_n62);
	nand (gm_n5682, gm_n5681, gm_n71, gm_n45);
	and (gm_n5683, gm_n48, gm_n53, in_10, gm_n2619, in_13);
	nand (gm_n5684, in_16, in_15, gm_n50, gm_n5683, in_17);
	nor (gm_n5685, in_20, gm_n62, in_18, gm_n5684, gm_n71);
	nor (gm_n5686, gm_n63, gm_n50, in_13, gm_n1577, gm_n46);
	nand (gm_n5687, in_19, in_18, gm_n81, gm_n5686, gm_n45);
	nor (gm_n5688, gm_n5687, gm_n71);
	or (gm_n5689, gm_n52, gm_n51, in_8, gm_n907, gm_n53);
	nor (gm_n5690, in_14, gm_n49, in_12, gm_n5689, gm_n63);
	nand (gm_n5691, gm_n47, gm_n81, gm_n46, gm_n5690, gm_n62);
	nor (gm_n5692, gm_n5691, in_21, gm_n45);
	nor (gm_n5693, in_11, in_10, in_9, gm_n5586);
	nand (gm_n5694, in_14, in_13, gm_n48, gm_n5693, gm_n63);
	or (gm_n5695, in_18, in_17, gm_n46, gm_n5694, in_19);
	nor (gm_n5696, gm_n5695, gm_n71, gm_n45);
	nand (gm_n5697, in_12, gm_n53, gm_n52, gm_n1780, in_13);
	nor (gm_n5698, gm_n46, in_15, in_14, gm_n5697, gm_n81);
	nand (gm_n5699, in_20, in_19, gm_n47, gm_n5698, in_21);
	nand (gm_n5700, in_12, in_11, in_10, gm_n2641, in_13);
	nor (gm_n5701, in_16, gm_n63, gm_n50, gm_n5700, in_17);
	nand (gm_n5702, in_20, gm_n62, gm_n47, gm_n5701, in_21);
	nand (gm_n5703, gm_n5702, gm_n5699);
	nor (gm_n5704, gm_n5692, gm_n5688, gm_n5685, gm_n5703, gm_n5696);
	nand (gm_n5705, gm_n5679, gm_n5675, gm_n5672, gm_n5704, gm_n5682);
	nor (gm_n5706, gm_n5663, gm_n5660, gm_n5657, gm_n5705, gm_n5667);
	nand (gm_n5707, gm_n5650, gm_n5647, gm_n5643, gm_n5706, gm_n5654);
	nor (gm_n5708, gm_n5636, gm_n5634, gm_n5631, gm_n5707, gm_n5640);
	nand (gm_n5709, gm_n5626, gm_n5623, gm_n5619, gm_n5708, gm_n5629);
	nor (gm_n5710, gm_n5611, gm_n5608, gm_n5604, gm_n5709, gm_n5615);
	nand (gm_n5711, gm_n5598, gm_n5594, gm_n5590, gm_n5710, gm_n5600);
	nor (gm_n5712, gm_n5582, gm_n5579, gm_n5575, gm_n5711, gm_n5585);
	nand (gm_n5713, gm_n5568, gm_n5565, gm_n5561, gm_n5712, gm_n5572);
	nor (gm_n5714, gm_n5556, gm_n5552, gm_n5548, gm_n5713, gm_n5558);
	nand (gm_n5715, gm_n5542, gm_n5538, gm_n5534, gm_n5714, gm_n5544);
	nor (gm_n5716, gm_n5526, gm_n5522, gm_n5518, gm_n5715, gm_n5530);
	nand (gm_n5717, gm_n5512, gm_n5508, gm_n5505, gm_n5716, gm_n5515);
	nor (gm_n5718, gm_n5499, gm_n5496, gm_n5492, gm_n5717, gm_n5501);
	nand (gm_n5719, gm_n5485, gm_n5482, gm_n5479, gm_n5718, gm_n5488);
	nor (gm_n5720, gm_n5471, gm_n5467, gm_n5464, gm_n5719, gm_n5475);
	nand (gm_n5721, gm_n5457, gm_n5454, gm_n5450, gm_n5720, gm_n5461);
	nor (gm_n5722, gm_n5445, gm_n5442, gm_n5439, gm_n5721, gm_n5447);
	nand (gm_n5723, gm_n5432, gm_n5429, gm_n5426, gm_n5722, gm_n5436);
	nor (gm_n5724, gm_n5417, gm_n5413, gm_n5409, gm_n5723, gm_n5421);
	nand (gm_n5725, gm_n5403, gm_n5398, gm_n5395, gm_n5724, gm_n5406);
	nor (gm_n5726, gm_n5387, gm_n5383, gm_n5378, gm_n5725, gm_n5391);
	nand (gm_n5727, gm_n5372, gm_n5371, gm_n5368, gm_n5726, gm_n5374);
	nor (gm_n5728, gm_n5361, gm_n5357, gm_n5354, gm_n5727, gm_n5365);
	nand (gm_n5729, gm_n5347, gm_n5344, gm_n5339, gm_n5728, gm_n5350);
	nor (gm_n5730, gm_n5332, gm_n5329, gm_n5325, gm_n5729, gm_n5335);
	nand (gm_n5731, gm_n5318, gm_n5314, gm_n5311, gm_n5730, gm_n5321);
	nor (gm_n5732, gm_n5304, gm_n5302, gm_n5297, gm_n5731, gm_n5308);
	nand (gm_n5733, gm_n5292, gm_n5288, gm_n5285, gm_n5732, gm_n5295);
	nor (gm_n5734, gm_n5278, gm_n5275, gm_n5271, gm_n5733, gm_n5282);
	nand (gm_n5735, gm_n5262, gm_n5259, gm_n5256, gm_n5734, gm_n5267);
	nor (gm_n5736, gm_n5247, gm_n5244, gm_n5241, gm_n5735, gm_n5251);
	nand (gm_n5737, gm_n5235, gm_n5232, gm_n5228, gm_n5736, gm_n5238);
	nor (gm_n5738, gm_n5221, gm_n5218, gm_n5216, gm_n5737, gm_n5224);
	nand (gm_n5739, gm_n5209, gm_n5205, gm_n5201, gm_n5738, gm_n5213);
	nor (out_8, gm_n5193, gm_n5189, gm_n5184, gm_n5739, gm_n5197);
	nand (gm_n5741, gm_n53, in_10, gm_n51, gm_n1057, in_12);
	nor (gm_n5742, gm_n63, in_14, in_13, gm_n5741, in_16);
	nand (gm_n5743, gm_n62, in_18, in_17, gm_n5742, gm_n45);
	nor (gm_n5744, gm_n5743, in_21);
	nand (gm_n5745, in_13, gm_n48, gm_n53, gm_n5531, gm_n50);
	nor (gm_n5746, in_17, gm_n46, in_15, gm_n5745, gm_n47);
	nand (gm_n5747, gm_n71, gm_n45, gm_n62, gm_n5746);
	and (gm_n5748, gm_n48, in_11, gm_n52, gm_n400, gm_n49);
	and (gm_n5749, in_16, in_15, gm_n50, gm_n5748, gm_n81);
	nand (gm_n5750, in_20, in_19, in_18, gm_n5749, gm_n71);
	nor (gm_n5751, in_17, in_16, gm_n63, gm_n3982, gm_n47);
	nand (gm_n5752, gm_n71, gm_n45, gm_n62, gm_n5751);
	nand (gm_n5753, in_12, gm_n53, in_10, gm_n1932, gm_n49);
	nor (gm_n5754, in_16, gm_n63, in_14, gm_n5753, in_17);
	nand (gm_n5755, in_20, gm_n62, in_18, gm_n5754, in_21);
	nor (gm_n5756, gm_n53, gm_n52, in_9, gm_n649);
	and (gm_n5757, in_14, gm_n49, gm_n48, gm_n5756, in_15);
	nand (gm_n5758, gm_n47, in_17, in_16, gm_n5757, gm_n62);
	nor (gm_n5759, gm_n5758, in_21, in_20);
	nand (gm_n5760, gm_n291, in_10, in_9);
	nor (gm_n5761, gm_n49, gm_n48, gm_n53, gm_n5760, gm_n50);
	nand (gm_n5762, in_17, gm_n46, in_15, gm_n5761, in_18);
	nor (gm_n5763, gm_n71, gm_n45, in_19, gm_n5762);
	nor (gm_n5764, in_11, in_10, gm_n51, gm_n2419, in_12);
	and (gm_n5765, in_15, gm_n50, in_13, gm_n5764, in_16);
	nand (gm_n5766, in_19, gm_n47, in_17, gm_n5765, gm_n45);
	nor (gm_n5767, gm_n5766, gm_n71);
	nand (gm_n5768, in_8, gm_n55, gm_n82, gm_n2640, gm_n51);
	nor (gm_n5769, in_12, in_11, gm_n52, gm_n5768, gm_n49);
	nand (gm_n5770, gm_n46, in_15, in_14, gm_n5769, gm_n81);
	nor (gm_n5771, in_20, in_19, in_18, gm_n5770, in_21);
	nor (gm_n5772, gm_n53, in_10, in_9, gm_n3428);
	nand (gm_n5773, gm_n50, in_13, gm_n48, gm_n5772, gm_n63);
	nor (gm_n5774, gm_n47, gm_n81, in_16, gm_n5773, gm_n62);
	nand (gm_n5775, gm_n5774, in_21, gm_n45);
	nor (gm_n5776, in_11, in_10, in_9, gm_n183);
	nand (gm_n5777, in_14, in_13, in_12, gm_n5776, gm_n63);
	nor (gm_n5778, gm_n47, in_17, gm_n46, gm_n5777, gm_n62);
	nand (gm_n5779, gm_n5778, in_21, in_20);
	and (gm_n5780, gm_n53, in_10, in_9, gm_n1339, gm_n48);
	nand (gm_n5781, in_15, gm_n50, in_13, gm_n5780, in_16);
	nor (gm_n5782, in_19, in_18, gm_n81, gm_n5781, gm_n45);
	nand (gm_n5783, gm_n5782, gm_n71);
	nor (gm_n5784, gm_n51, in_8, in_7, gm_n588, in_10);
	nand (gm_n5785, gm_n49, gm_n48, gm_n53, gm_n5784, gm_n50);
	nor (gm_n5786, in_17, in_16, in_15, gm_n5785, in_18);
	nand (gm_n5787, gm_n71, gm_n45, gm_n62, gm_n5786);
	and (gm_n5788, gm_n55, gm_n82, gm_n72, gm_n284);
	nand (gm_n5789, in_10, gm_n51, gm_n64, gm_n5788, in_11);
	nor (gm_n5790, gm_n50, gm_n49, gm_n48, gm_n5789, gm_n63);
	nand (gm_n5791, in_18, gm_n81, gm_n46, gm_n5790, gm_n62);
	nor (gm_n5792, gm_n5791, in_21, in_20);
	nor (gm_n5793, gm_n64, gm_n55, gm_n82, gm_n96, gm_n51);
	and (gm_n5794, gm_n48, in_11, gm_n52, gm_n5793, in_13);
	nand (gm_n5795, gm_n46, gm_n63, in_14, gm_n5794, in_17);
	nor (gm_n5796, in_20, in_19, in_18, gm_n5795, gm_n71);
	nor (gm_n5797, gm_n50, in_13, in_12, gm_n5689, in_15);
	nand (gm_n5798, gm_n47, in_17, in_16, gm_n5797, gm_n62);
	nor (gm_n5799, gm_n5798, gm_n71, in_20);
	nor (gm_n5800, in_13, in_12, in_11, gm_n1916, gm_n50);
	nand (gm_n5801, gm_n81, gm_n46, in_15, gm_n5800, in_18);
	nor (gm_n5802, in_21, in_20, in_19, gm_n5801);
	nor (gm_n5803, in_11, in_10, in_9, gm_n3557, gm_n48);
	nand (gm_n5804, gm_n63, in_14, gm_n49, gm_n5803, in_16);
	nor (gm_n5805, gm_n62, in_18, gm_n81, gm_n5804, in_20);
	nand (gm_n5806, gm_n5805, in_21);
	nand (gm_n5807, gm_n48, in_11, in_10, gm_n1755, gm_n49);
	nor (gm_n5808, gm_n46, in_15, gm_n50, gm_n5807, in_17);
	nand (gm_n5809, gm_n45, in_19, in_18, gm_n5808, in_21);
	nand (gm_n5810, in_13, gm_n48, gm_n53, gm_n3712);
	nor (gm_n5811, in_16, in_15, gm_n50, gm_n5810, in_17);
	nand (gm_n5812, gm_n45, in_19, gm_n47, gm_n5811, gm_n71);
	nand (gm_n5813, in_14, in_13, gm_n48, gm_n3471, in_15);
	nor (gm_n5814, in_18, in_17, gm_n46, gm_n5813, in_19);
	nand (gm_n5815, gm_n5814, gm_n71, in_20);
	or (gm_n5816, gm_n51, in_8, gm_n55, gm_n525, in_10);
	nor (gm_n5817, in_13, gm_n48, in_11, gm_n5816, in_14);
	nand (gm_n5818, gm_n81, in_16, in_15, gm_n5817, in_18);
	nor (gm_n5819, gm_n71, gm_n45, gm_n62, gm_n5818);
	nand (gm_n5820, gm_n47, in_17, in_16, gm_n127, in_19);
	nor (gm_n5821, gm_n5820, gm_n71, gm_n45);
	and (gm_n5822, in_8, gm_n55, gm_n82, gm_n757, gm_n51);
	and (gm_n5823, in_12, gm_n53, in_10, gm_n5822, gm_n49);
	nand (gm_n5824, in_16, gm_n63, in_14, gm_n5823, in_17);
	nor (gm_n5825, in_20, in_19, in_18, gm_n5824, gm_n71);
	nand (gm_n5826, in_11, in_10, in_9, gm_n1222);
	nor (gm_n5827, in_14, gm_n49, gm_n48, gm_n5826, in_15);
	nand (gm_n5828, in_18, in_17, gm_n46, gm_n5827, in_19);
	nor (gm_n5829, gm_n5828, gm_n71, gm_n45);
	and (gm_n5830, gm_n46, in_15, gm_n50, gm_n2936, gm_n81);
	nand (gm_n5831, gm_n45, in_19, in_18, gm_n5830, in_21);
	nor (gm_n5832, in_17, gm_n46, gm_n63, gm_n952, gm_n47);
	nand (gm_n5833, gm_n71, gm_n45, gm_n62, gm_n5832);
	nor (gm_n5834, gm_n2926, in_10, gm_n51);
	nand (gm_n5835, in_13, in_12, in_11, gm_n5834, in_14);
	nor (gm_n5836, gm_n81, in_16, gm_n63, gm_n5835, in_18);
	nand (gm_n5837, in_21, gm_n45, gm_n62, gm_n5836);
	and (gm_n5838, in_10, gm_n51, in_8, gm_n57);
	nand (gm_n5839, in_13, in_12, gm_n53, gm_n5838, in_14);
	nor (gm_n5840, in_17, in_16, in_15, gm_n5839, gm_n47);
	nand (gm_n5841, in_21, gm_n45, in_19, gm_n5840);
	and (gm_n5842, gm_n3904, in_9);
	and (gm_n5843, gm_n48, in_11, in_10, gm_n5842, in_13);
	nand (gm_n5844, in_16, gm_n63, gm_n50, gm_n5843, gm_n81);
	nor (gm_n5845, gm_n45, in_19, gm_n47, gm_n5844, in_21);
	nor (gm_n5846, gm_n48, gm_n53, gm_n52, gm_n531, in_13);
	nand (gm_n5847, in_16, gm_n63, in_14, gm_n5846, in_17);
	nor (gm_n5848, in_20, in_19, in_18, gm_n5847, gm_n71);
	nor (gm_n5849, in_13, in_12, in_11, gm_n3300, in_14);
	nand (gm_n5850, in_17, in_16, in_15, gm_n5849, in_18);
	nor (gm_n5851, in_21, gm_n45, in_19, gm_n5850);
	and (gm_n5852, gm_n48, in_11, gm_n52, gm_n1671, in_13);
	nand (gm_n5853, in_16, gm_n63, in_14, gm_n5852, in_17);
	nor (gm_n5854, in_20, in_19, in_18, gm_n5853, gm_n71);
	nand (gm_n5855, in_13, gm_n48, in_11, gm_n85, in_14);
	nor (gm_n5856, in_17, in_16, in_15, gm_n5855, gm_n47);
	nand (gm_n5857, in_21, in_20, gm_n62, gm_n5856);
	and (gm_n5858, in_9, gm_n64, in_7, gm_n151, in_10);
	nand (gm_n5859, in_13, in_12, in_11, gm_n5858, in_14);
	nor (gm_n5860, in_17, in_16, gm_n63, gm_n5859, in_18);
	nand (gm_n5861, gm_n71, gm_n45, gm_n62, gm_n5860);
	nand (gm_n5862, in_12, in_11, gm_n52, gm_n2097, gm_n49);
	nor (gm_n5863, in_16, gm_n63, in_14, gm_n5862, in_17);
	nand (gm_n5864, in_20, gm_n62, in_18, gm_n5863, in_21);
	nor (gm_n5865, in_11, gm_n52, gm_n51, gm_n2610, gm_n48);
	nand (gm_n5866, in_15, in_14, gm_n49, gm_n5865, gm_n46);
	nor (gm_n5867, gm_n62, in_18, gm_n81, gm_n5866, gm_n45);
	nand (gm_n5868, gm_n5867, gm_n71);
	nand (gm_n5869, in_16, in_15, gm_n50, gm_n401, gm_n81);
	nor (gm_n5870, gm_n45, gm_n62, in_18, gm_n5869, in_21);
	and (gm_n5871, gm_n48, in_11, in_10, gm_n1975, gm_n49);
	nand (gm_n5872, gm_n46, in_15, in_14, gm_n5871, in_17);
	nor (gm_n5873, in_20, gm_n62, in_18, gm_n5872, gm_n71);
	nor (gm_n5874, in_14, gm_n49, gm_n48, gm_n4943, in_15);
	nand (gm_n5875, in_18, in_17, gm_n46, gm_n5874, gm_n62);
	nor (gm_n5876, gm_n5875, gm_n71, gm_n45);
	nand (gm_n5877, gm_n52, gm_n51, in_8, gm_n384);
	nor (gm_n5878, gm_n49, gm_n48, gm_n53, gm_n5877, in_14);
	nand (gm_n5879, in_17, gm_n46, gm_n63, gm_n5878, in_18);
	nor (gm_n5880, in_21, in_20, gm_n62, gm_n5879);
	nor (gm_n5881, gm_n5298, in_10, gm_n51);
	nand (gm_n5882, in_13, in_12, in_11, gm_n5881, in_14);
	nor (gm_n5883, in_17, gm_n46, gm_n63, gm_n5882, in_18);
	nand (gm_n5884, gm_n71, in_20, gm_n62, gm_n5883);
	nand (gm_n5885, gm_n48, in_11, gm_n52, gm_n1719, gm_n49);
	nor (gm_n5886, in_16, gm_n63, in_14, gm_n5885, in_17);
	nand (gm_n5887, gm_n45, in_19, in_18, gm_n5886, gm_n71);
	nand (gm_n5888, in_7, gm_n82, gm_n72, gm_n252, gm_n64);
	nor (gm_n5889, in_11, gm_n52, in_9, gm_n5888, in_12);
	nand (gm_n5890, in_15, in_14, gm_n49, gm_n5889, in_16);
	nor (gm_n5891, gm_n62, in_18, in_17, gm_n5890, in_20);
	nand (gm_n5892, gm_n5891, in_21);
	nor (gm_n5893, in_8, gm_n55, gm_n82, gm_n1429, in_9);
	nand (gm_n5894, in_12, gm_n53, gm_n52, gm_n5893, gm_n49);
	nor (gm_n5895, gm_n46, gm_n63, gm_n50, gm_n5894, gm_n81);
	nand (gm_n5896, in_20, gm_n62, in_18, gm_n5895, gm_n71);
	nor (gm_n5897, in_15, in_14, gm_n49, gm_n5194, in_16);
	nand (gm_n5898, in_19, gm_n47, gm_n81, gm_n5897, gm_n45);
	nor (gm_n5899, gm_n5898, in_21);
	and (gm_n5900, in_12, gm_n53, gm_n52, gm_n1671, in_13);
	nand (gm_n5901, gm_n46, gm_n63, gm_n50, gm_n5900, in_17);
	nor (gm_n5902, gm_n45, in_19, gm_n47, gm_n5901, in_21);
	nor (gm_n5903, in_12, gm_n53, in_10, gm_n2645, in_13);
	nand (gm_n5904, in_16, gm_n63, in_14, gm_n5903, gm_n81);
	nor (gm_n5905, gm_n45, in_19, in_18, gm_n5904, in_21);
	nand (gm_n5906, gm_n51, in_8, in_7, gm_n136);
	nor (gm_n5907, gm_n48, gm_n53, gm_n52, gm_n5906, in_13);
	nand (gm_n5908, gm_n46, gm_n63, gm_n50, gm_n5907, gm_n81);
	nor (gm_n5909, in_20, in_19, gm_n47, gm_n5908, in_21);
	nand (gm_n5910, gm_n50, in_13, in_12, gm_n4196, gm_n63);
	nor (gm_n5911, in_18, in_17, in_16, gm_n5910, gm_n62);
	nand (gm_n5912, gm_n5911, gm_n71, gm_n45);
	nor (gm_n5913, in_11, in_10, in_9, gm_n3697, gm_n48);
	nand (gm_n5914, in_15, in_14, gm_n49, gm_n5913, gm_n46);
	nor (gm_n5915, gm_n62, gm_n47, gm_n81, gm_n5914, gm_n45);
	nand (gm_n5916, gm_n5915, in_21);
	nor (gm_n5917, gm_n52, in_9, gm_n64, gm_n4514, gm_n53);
	nand (gm_n5918, gm_n50, in_13, in_12, gm_n5917, in_15);
	nor (gm_n5919, gm_n47, gm_n81, in_16, gm_n5918, gm_n62);
	nand (gm_n5920, gm_n5919, in_21, in_20);
	nand (gm_n5921, gm_n49, gm_n48, in_11, gm_n5468, gm_n50);
	nor (gm_n5922, gm_n81, gm_n46, gm_n63, gm_n5921, gm_n47);
	nand (gm_n5923, in_21, gm_n45, gm_n62, gm_n5922);
	nor (gm_n5924, in_11, gm_n52, in_9, gm_n3198);
	and (gm_n5925, in_14, gm_n49, in_12, gm_n5924, in_15);
	nand (gm_n5926, gm_n47, gm_n81, gm_n46, gm_n5925, in_19);
	nor (gm_n5927, gm_n5926, gm_n71, in_20);
	and (gm_n5928, gm_n2653, gm_n52, gm_n51);
	and (gm_n5929, gm_n49, gm_n48, in_11, gm_n5928, gm_n50);
	nand (gm_n5930, in_17, in_16, gm_n63, gm_n5929, in_18);
	nor (gm_n5931, gm_n71, in_20, gm_n62, gm_n5930);
	nor (gm_n5932, gm_n3198, gm_n52, gm_n51);
	and (gm_n5933, in_13, gm_n48, in_11, gm_n5932, gm_n50);
	nand (gm_n5934, gm_n81, in_16, gm_n63, gm_n5933, in_18);
	nor (gm_n5935, gm_n71, gm_n45, in_19, gm_n5934);
	and (gm_n5936, in_12, gm_n53, gm_n52, gm_n3069, gm_n49);
	nand (gm_n5937, gm_n46, in_15, gm_n50, gm_n5936, gm_n81);
	nor (gm_n5938, in_20, gm_n62, in_18, gm_n5937, in_21);
	nand (gm_n5939, in_15, in_14, in_13, gm_n2398, gm_n46);
	nor (gm_n5940, gm_n62, in_18, gm_n81, gm_n5939, in_20);
	nand (gm_n5941, gm_n5940, in_21);
	and (gm_n5942, gm_n46, in_15, in_14, gm_n386, gm_n81);
	nand (gm_n5943, gm_n45, gm_n62, gm_n47, gm_n5942, in_21);
	nor (gm_n5944, in_11, in_10, in_9, gm_n410, in_12);
	nand (gm_n5945, in_15, gm_n50, in_13, gm_n5944, in_16);
	nor (gm_n5946, in_19, in_18, in_17, gm_n5945, gm_n45);
	nand (gm_n5947, gm_n5946, gm_n71);
	nor (gm_n5948, gm_n53, in_10, in_9, gm_n2275, gm_n48);
	nand (gm_n5949, in_15, in_14, in_13, gm_n5948, in_16);
	nor (gm_n5950, gm_n62, gm_n47, in_17, gm_n5949, in_20);
	nand (gm_n5951, gm_n5950, gm_n71);
	or (gm_n5952, in_11, in_10, in_9, gm_n873, gm_n48);
	nor (gm_n5953, in_15, in_14, in_13, gm_n5952, in_16);
	nand (gm_n5954, in_19, in_18, in_17, gm_n5953, in_20);
	nor (gm_n5955, gm_n5954, in_21);
	nor (gm_n5956, in_13, in_12, gm_n53, gm_n4891, in_14);
	nand (gm_n5957, gm_n81, gm_n46, in_15, gm_n5956, in_18);
	nor (gm_n5958, in_21, gm_n45, in_19, gm_n5957);
	or (gm_n5959, in_11, in_10, gm_n51, gm_n4562, gm_n48);
	nor (gm_n5960, in_15, in_14, gm_n49, gm_n5959, in_16);
	nand (gm_n5961, gm_n62, gm_n47, in_17, gm_n5960, gm_n45);
	nor (gm_n5962, gm_n5961, in_21);
	and (gm_n5963, gm_n49, gm_n48, in_11, gm_n436, gm_n50);
	nand (gm_n5964, gm_n81, in_16, in_15, gm_n5963, in_18);
	nor (gm_n5965, gm_n71, in_20, in_19, gm_n5964);
	or (gm_n5966, gm_n1970, gm_n52, in_9);
	or (gm_n5967, in_13, gm_n48, gm_n53, gm_n5966, in_14);
	nor (gm_n5968, in_17, gm_n46, in_15, gm_n5967, gm_n47);
	nand (gm_n5969, in_21, in_20, gm_n62, gm_n5968);
	nor (gm_n5970, gm_n53, in_10, in_9, gm_n90, in_12);
	nand (gm_n5971, gm_n63, gm_n50, gm_n49, gm_n5970, gm_n46);
	nor (gm_n5972, in_19, in_18, in_17, gm_n5971, gm_n45);
	nand (gm_n5973, gm_n5972, in_21);
	nand (gm_n5974, gm_n49, gm_n48, gm_n53, gm_n4640, gm_n50);
	nor (gm_n5975, gm_n81, gm_n46, gm_n63, gm_n5974, gm_n47);
	nand (gm_n5976, gm_n71, gm_n45, in_19, gm_n5975);
	nor (gm_n5977, gm_n51, gm_n64, in_7, gm_n525, in_10);
	nand (gm_n5978, in_13, in_12, gm_n53, gm_n5977, gm_n50);
	nor (gm_n5979, in_17, gm_n46, in_15, gm_n5978, in_18);
	nand (gm_n5980, gm_n71, in_20, in_19, gm_n5979);
	nand (gm_n5981, in_9, gm_n64, gm_n55, gm_n151, in_10);
	nor (gm_n5982, gm_n49, gm_n48, gm_n53, gm_n5981, gm_n50);
	nand (gm_n5983, in_17, in_16, in_15, gm_n5982, in_18);
	nor (gm_n5984, in_21, in_20, in_19, gm_n5983);
	nand (gm_n5985, gm_n46, gm_n63, in_14, gm_n4502, gm_n81);
	nor (gm_n5986, gm_n45, in_19, gm_n47, gm_n5985, in_21);
	nand (gm_n5987, in_12, in_11, in_10, gm_n3941, in_13);
	or (gm_n5988, in_16, in_15, in_14, gm_n5987, gm_n81);
	nor (gm_n5989, in_20, gm_n62, in_18, gm_n5988, in_21);
	and (gm_n5990, gm_n63, gm_n50, gm_n49, gm_n1534, gm_n46);
	nand (gm_n5991, gm_n62, gm_n47, gm_n81, gm_n5990, in_20);
	nor (gm_n5992, gm_n5991, in_21);
	nor (gm_n5993, in_11, gm_n52, in_9, gm_n322);
	nand (gm_n5994, gm_n50, in_13, in_12, gm_n5993, in_15);
	nor (gm_n5995, in_18, gm_n81, gm_n46, gm_n5994, gm_n62);
	nand (gm_n5996, gm_n5995, gm_n71, in_20);
	nand (gm_n5997, in_12, gm_n53, in_10, gm_n3443, in_13);
	nor (gm_n5998, in_16, gm_n63, in_14, gm_n5997, in_17);
	nand (gm_n5999, gm_n45, gm_n62, in_18, gm_n5998, in_21);
	nand (gm_n6000, in_12, gm_n53, gm_n52, gm_n1692, in_13);
	nor (gm_n6001, gm_n46, in_15, gm_n50, gm_n6000, gm_n81);
	nand (gm_n6002, in_20, in_19, gm_n47, gm_n6001, in_21);
	nor (gm_n6003, in_17, in_16, in_15, gm_n1998, in_18);
	nand (gm_n6004, gm_n71, gm_n45, in_19, gm_n6003);
	nor (gm_n6005, gm_n1040, gm_n49);
	nand (gm_n6006, gm_n46, gm_n63, gm_n50, gm_n6005, in_17);
	nor (gm_n6007, gm_n45, gm_n62, in_18, gm_n6006, in_21);
	nor (gm_n6008, in_12, gm_n53, gm_n52, gm_n3773, in_13);
	nand (gm_n6009, in_16, gm_n63, gm_n50, gm_n6008, gm_n81);
	nor (gm_n6010, in_20, gm_n62, gm_n47, gm_n6009, in_21);
	and (gm_n6011, gm_n49, gm_n48, gm_n53, gm_n3170, in_14);
	nand (gm_n6012, gm_n81, gm_n46, gm_n63, gm_n6011, in_18);
	nor (gm_n6013, gm_n71, gm_n45, in_19, gm_n6012);
	nor (gm_n6014, gm_n53, in_10, in_9, gm_n2397, in_12);
	nand (gm_n6015, gm_n6014, gm_n49);
	or (gm_n6016, gm_n46, in_15, in_14, gm_n6015, in_17);
	nor (gm_n6017, in_20, in_19, gm_n47, gm_n6016, gm_n71);
	and (gm_n6018, in_16, gm_n63, in_14, gm_n1653, in_17);
	nand (gm_n6019, gm_n45, gm_n62, gm_n47, gm_n6018, in_21);
	nand (gm_n6020, gm_n63, gm_n50, in_13, gm_n2903, in_16);
	nor (gm_n6021, gm_n62, in_18, in_17, gm_n6020, gm_n45);
	nand (gm_n6022, gm_n6021, gm_n71);
	or (gm_n6023, gm_n48, in_11, gm_n52, gm_n1744, in_13);
	nor (gm_n6024, gm_n46, gm_n63, gm_n50, gm_n6023, gm_n81);
	nand (gm_n6025, gm_n45, in_19, in_18, gm_n6024, in_21);
	nand (gm_n6026, in_14, gm_n49, gm_n48, gm_n5924, in_15);
	nor (gm_n6027, in_18, gm_n81, in_16, gm_n6026, gm_n62);
	nand (gm_n6028, gm_n6027, gm_n71, gm_n45);
	and (gm_n6029, in_13, in_12, gm_n53, gm_n2828, gm_n50);
	nand (gm_n6030, gm_n81, gm_n46, gm_n63, gm_n6029, in_18);
	nor (gm_n6031, in_21, in_20, in_19, gm_n6030);
	nand (gm_n6032, gm_n64, in_7, in_6, gm_n379, in_9);
	nor (gm_n6033, in_12, gm_n53, gm_n52, gm_n6032, in_13);
	nand (gm_n6034, in_16, gm_n63, in_14, gm_n6033, gm_n81);
	nor (gm_n6035, gm_n45, gm_n62, gm_n47, gm_n6034, gm_n71);
	nor (gm_n6036, in_13, gm_n48, gm_n53, gm_n4325, gm_n50);
	nand (gm_n6037, in_17, gm_n46, in_15, gm_n6036, in_18);
	nor (gm_n6038, gm_n71, gm_n45, gm_n62, gm_n6037);
	and (gm_n6039, in_12, in_11, gm_n52, gm_n1332, in_13);
	nand (gm_n6040, in_16, in_15, in_14, gm_n6039, gm_n81);
	nor (gm_n6041, in_20, gm_n62, in_18, gm_n6040, gm_n71);
	nand (gm_n6042, gm_n48, in_11, gm_n52, gm_n3909, in_13);
	nor (gm_n6043, gm_n46, in_15, gm_n50, gm_n6042, in_17);
	nand (gm_n6044, in_20, gm_n62, in_18, gm_n6043, in_21);
	nand (gm_n6045, in_12, in_11, in_10, gm_n2056, in_13);
	nor (gm_n6046, gm_n46, in_15, gm_n50, gm_n6045, gm_n81);
	nand (gm_n6047, gm_n45, gm_n62, gm_n47, gm_n6046, gm_n71);
	nor (gm_n6048, gm_n53, gm_n52, in_9, gm_n3340);
	nand (gm_n6049, gm_n50, in_13, in_12, gm_n6048, gm_n63);
	nor (gm_n6050, in_18, in_17, gm_n46, gm_n6049, in_19);
	nand (gm_n6051, gm_n6050, in_21, in_20);
	nor (gm_n6052, in_8, in_7, gm_n82, gm_n161, gm_n51);
	nand (gm_n6053, in_12, in_11, gm_n52, gm_n6052, in_13);
	nor (gm_n6054, gm_n46, in_15, gm_n50, gm_n6053, gm_n81);
	nand (gm_n6055, in_20, in_19, gm_n47, gm_n6054, in_21);
	nand (gm_n6056, gm_n64, gm_n55, gm_n82, gm_n1075, gm_n51);
	nor (gm_n6057, gm_n48, gm_n53, gm_n52, gm_n6056, in_13);
	nand (gm_n6058, gm_n46, gm_n63, gm_n50, gm_n6057, gm_n81);
	nor (gm_n6059, in_20, gm_n62, in_18, gm_n6058, gm_n71);
	nor (gm_n6060, gm_n48, in_11, in_10, gm_n5030, gm_n49);
	nand (gm_n6061, gm_n46, in_15, gm_n50, gm_n6060, gm_n81);
	nor (gm_n6062, gm_n45, gm_n62, in_18, gm_n6061, in_21);
	nor (gm_n6063, in_12, gm_n53, gm_n52, gm_n5030, gm_n49);
	nand (gm_n6064, gm_n46, gm_n63, in_14, gm_n6063, in_17);
	nor (gm_n6065, gm_n45, in_19, in_18, gm_n6064, gm_n71);
	nor (gm_n6066, gm_n49, gm_n48, in_11, gm_n4398, in_14);
	nand (gm_n6067, gm_n81, gm_n46, gm_n63, gm_n6066, gm_n47);
	nor (gm_n6068, in_21, gm_n45, in_19, gm_n6067);
	nor (gm_n6069, gm_n53, gm_n52, in_9, gm_n1831);
	nand (gm_n6070, gm_n50, gm_n49, in_12, gm_n6069, in_15);
	nor (gm_n6071, in_18, gm_n81, in_16, gm_n6070, in_19);
	nand (gm_n6072, gm_n6071, gm_n71, in_20);
	nand (gm_n6073, gm_n48, gm_n53, gm_n52, gm_n2334, gm_n49);
	nor (gm_n6074, in_16, gm_n63, gm_n50, gm_n6073, in_17);
	nand (gm_n6075, in_20, in_19, in_18, gm_n6074, gm_n71);
	and (gm_n6076, in_10, in_9, in_8, gm_n338);
	nand (gm_n6077, in_13, gm_n48, gm_n53, gm_n6076, in_14);
	nor (gm_n6078, gm_n81, gm_n46, in_15, gm_n6077, gm_n47);
	nand (gm_n6079, gm_n71, gm_n45, in_19, gm_n6078);
	nor (gm_n6080, gm_n52, gm_n51, in_8, gm_n478, in_11);
	and (gm_n6081, gm_n6080, in_13, gm_n48);
	and (gm_n6082, gm_n46, in_15, in_14, gm_n6081, in_17);
	nand (gm_n6083, gm_n45, in_19, in_18, gm_n6082, gm_n71);
	nor (gm_n6084, in_12, gm_n53, gm_n52, gm_n264, in_13);
	nand (gm_n6085, in_16, gm_n63, in_14, gm_n6084, gm_n81);
	nor (gm_n6086, gm_n45, gm_n62, in_18, gm_n6085, gm_n71);
	and (gm_n6087, in_13, gm_n48, gm_n53, gm_n3035, in_14);
	nand (gm_n6088, in_17, in_16, gm_n63, gm_n6087, in_18);
	nor (gm_n6089, gm_n71, gm_n45, in_19, gm_n6088);
	nor (gm_n6090, gm_n50, in_13, in_12, gm_n5789, in_15);
	nand (gm_n6091, in_18, gm_n81, gm_n46, gm_n6090, in_19);
	nor (gm_n6092, gm_n6091, in_21, in_20);
	or (gm_n6093, gm_n53, in_10, gm_n51, gm_n2823, in_12);
	nor (gm_n6094, gm_n63, in_14, gm_n49, gm_n6093, gm_n46);
	nand (gm_n6095, gm_n62, in_18, in_17, gm_n6094, gm_n45);
	nor (gm_n6096, gm_n6095, gm_n71);
	nor (gm_n6097, gm_n53, gm_n52, gm_n51, gm_n1831, in_12);
	nand (gm_n6098, in_15, in_14, in_13, gm_n6097, gm_n46);
	nor (gm_n6099, in_19, in_18, gm_n81, gm_n6098, in_20);
	nand (gm_n6100, gm_n6099, in_21);
	nor (gm_n6101, in_11, in_10, gm_n51, gm_n2397, gm_n48);
	nand (gm_n6102, in_15, gm_n50, gm_n49, gm_n6101, gm_n46);
	nor (gm_n6103, in_19, in_18, in_17, gm_n6102, gm_n45);
	nand (gm_n6104, gm_n6103, gm_n71);
	and (gm_n6105, gm_n1550, gm_n52, in_9);
	nand (gm_n6106, gm_n49, gm_n48, in_11, gm_n6105, in_14);
	nor (gm_n6107, gm_n81, in_16, in_15, gm_n6106, in_18);
	nand (gm_n6108, gm_n71, gm_n45, gm_n62, gm_n6107);
	and (gm_n6109, gm_n46, gm_n63, gm_n50, gm_n3901, gm_n81);
	nand (gm_n6110, in_20, gm_n62, in_18, gm_n6109, gm_n71);
	nor (gm_n6111, gm_n48, gm_n53, gm_n52, gm_n1076, in_13);
	nand (gm_n6112, in_16, in_15, in_14, gm_n6111, in_17);
	nor (gm_n6113, in_20, in_19, gm_n47, gm_n6112, in_21);
	nor (gm_n6114, gm_n49, gm_n48, gm_n53, gm_n2589, in_14);
	nand (gm_n6115, gm_n81, in_16, in_15, gm_n6114, in_18);
	nor (gm_n6116, in_21, gm_n45, gm_n62, gm_n6115);
	and (gm_n6117, gm_n48, gm_n53, gm_n52, gm_n1440, gm_n49);
	nand (gm_n6118, in_16, gm_n63, gm_n50, gm_n6117, in_17);
	nor (gm_n6119, in_20, in_19, in_18, gm_n6118, gm_n71);
	nand (gm_n6120, gm_n52, in_9, gm_n64, gm_n838, gm_n53);
	nor (gm_n6121, in_14, gm_n49, in_12, gm_n6120, gm_n63);
	nand (gm_n6122, gm_n47, gm_n81, gm_n46, gm_n6121, in_19);
	nor (gm_n6123, gm_n6122, gm_n71, in_20);
	and (gm_n6124, gm_n1274, gm_n52, in_9);
	nand (gm_n6125, gm_n49, gm_n48, gm_n53, gm_n6124, in_14);
	nor (gm_n6126, in_17, gm_n46, gm_n63, gm_n6125, in_18);
	nand (gm_n6127, in_21, in_20, gm_n62, gm_n6126);
	nor (gm_n6128, in_17, in_16, gm_n63, gm_n1998, gm_n47);
	nand (gm_n6129, in_21, gm_n45, gm_n62, gm_n6128);
	nand (gm_n6130, in_12, in_11, gm_n52, gm_n5842, gm_n49);
	nor (gm_n6131, gm_n46, gm_n63, in_14, gm_n6130, gm_n81);
	nand (gm_n6132, in_20, in_19, gm_n47, gm_n6131, gm_n71);
	nor (gm_n6133, in_16, gm_n63, gm_n50, gm_n5236, in_17);
	nand (gm_n6134, gm_n45, in_19, gm_n47, gm_n6133, in_21);
	nand (gm_n6135, gm_n52, gm_n51, gm_n64, gm_n302);
	nor (gm_n6136, in_13, in_12, in_11, gm_n6135);
	nand (gm_n6137, gm_n46, in_15, in_14, gm_n6136, gm_n81);
	nor (gm_n6138, gm_n45, in_19, in_18, gm_n6137, gm_n71);
	and (gm_n6139, gm_n64, gm_n55, gm_n82, gm_n379, in_9);
	and (gm_n6140, gm_n48, in_11, gm_n52, gm_n6139, gm_n49);
	nand (gm_n6141, gm_n46, in_15, gm_n50, gm_n6140, in_17);
	nor (gm_n6142, gm_n45, in_19, in_18, gm_n6141, gm_n71);
	nor (gm_n6143, in_10, gm_n51, in_8, gm_n390, in_11);
	nand (gm_n6144, gm_n6143, in_13, gm_n48);
	or (gm_n6145, in_16, in_15, gm_n50, gm_n6144, gm_n81);
	nor (gm_n6146, gm_n45, in_19, gm_n47, gm_n6145, gm_n71);
	nand (gm_n6147, gm_n1002, gm_n51);
	nor (gm_n6148, in_12, in_11, gm_n52, gm_n6147, gm_n49);
	nand (gm_n6149, gm_n46, in_15, gm_n50, gm_n6148, gm_n81);
	nor (gm_n6150, gm_n45, gm_n62, gm_n47, gm_n6149, gm_n71);
	nor (gm_n6151, in_10, in_9, in_8, gm_n5180, in_11);
	nand (gm_n6152, gm_n50, gm_n49, in_12, gm_n6151, in_15);
	nor (gm_n6153, in_18, in_17, in_16, gm_n6152, in_19);
	nand (gm_n6154, gm_n6153, in_21, in_20);
	nand (gm_n6155, in_7, gm_n82, in_5, gm_n519, gm_n64);
	nor (gm_n6156, gm_n53, gm_n52, in_9, gm_n6155);
	nand (gm_n6157, gm_n50, gm_n49, in_12, gm_n6156, in_15);
	nor (gm_n6158, gm_n47, in_17, gm_n46, gm_n6157, gm_n62);
	nand (gm_n6159, gm_n6158, gm_n71, gm_n45);
	nor (gm_n6160, gm_n53, in_10, in_9, gm_n3146, in_12);
	nand (gm_n6161, in_15, in_14, gm_n49, gm_n6160, gm_n46);
	nor (gm_n6162, in_19, gm_n47, in_17, gm_n6161, in_20);
	nand (gm_n6163, gm_n6162, gm_n71);
	and (gm_n6164, gm_n53, gm_n52, in_9, gm_n1183, gm_n48);
	and (gm_n6165, gm_n6164, gm_n50, in_13);
	and (gm_n6166, gm_n81, gm_n46, in_15, gm_n6165, in_18);
	nand (gm_n6167, in_21, gm_n45, in_19, gm_n6166);
	nand (gm_n6168, in_11, gm_n52, gm_n51, gm_n792, gm_n48);
	nor (gm_n6169, gm_n63, gm_n50, gm_n49, gm_n6168);
	nand (gm_n6170, gm_n47, gm_n81, gm_n46, gm_n6169, gm_n62);
	nor (gm_n6171, gm_n6170, in_21, in_20);
	nor (gm_n6172, in_15, gm_n50, gm_n49, gm_n4306, gm_n46);
	nand (gm_n6173, gm_n62, in_18, in_17, gm_n6172, in_20);
	nor (gm_n6174, gm_n6173, in_21);
	nor (gm_n6175, in_14, in_13, gm_n48, gm_n3328, in_15);
	nand (gm_n6176, gm_n47, in_17, gm_n46, gm_n6175, in_19);
	nor (gm_n6177, gm_n6176, in_21, in_20);
	nor (gm_n6178, gm_n48, gm_n53, gm_n52, gm_n5549, gm_n49);
	nand (gm_n6179, gm_n46, in_15, gm_n50, gm_n6178, in_17);
	nor (gm_n6180, gm_n45, gm_n62, gm_n47, gm_n6179, in_21);
	nand (gm_n6181, gm_n49, gm_n48, in_11, gm_n1107, gm_n50);
	nor (gm_n6182, in_17, gm_n46, gm_n63, gm_n6181, gm_n47);
	nand (gm_n6183, in_21, in_20, gm_n62, gm_n6182);
	and (gm_n6184, gm_n52, gm_n51, in_8, gm_n691, in_11);
	nand (gm_n6185, in_14, gm_n49, gm_n48, gm_n6184, gm_n63);
	nor (gm_n6186, gm_n47, gm_n81, gm_n46, gm_n6185, in_19);
	nand (gm_n6187, gm_n6186, in_21, in_20);
	or (gm_n6188, in_12, gm_n53, gm_n52, gm_n2355, gm_n49);
	nor (gm_n6189, in_16, gm_n63, gm_n50, gm_n6188, in_17);
	nand (gm_n6190, in_20, in_19, in_18, gm_n6189, gm_n71);
	nor (gm_n6191, in_16, in_15, in_14, gm_n5700, gm_n81);
	nand (gm_n6192, in_20, gm_n62, in_18, gm_n6191, gm_n71);
	or (gm_n6193, gm_n64, in_7, gm_n82, gm_n96, in_9);
	nor (gm_n6194, gm_n48, gm_n53, gm_n52, gm_n6193, in_13);
	nand (gm_n6195, gm_n46, gm_n63, in_14, gm_n6194, in_17);
	nor (gm_n6196, gm_n45, in_19, gm_n47, gm_n6195, in_21);
	nand (gm_n6197, gm_n53, gm_n52, gm_n51, gm_n194, gm_n48);
	nor (gm_n6198, gm_n63, gm_n50, in_13, gm_n6197, gm_n46);
	nand (gm_n6199, gm_n62, in_18, in_17, gm_n6198, in_20);
	nor (gm_n6200, gm_n6199, in_21);
	nor (gm_n6201, gm_n50, gm_n49, gm_n48, gm_n3644, in_15);
	nand (gm_n6202, in_18, gm_n81, gm_n46, gm_n6201, in_19);
	nor (gm_n6203, gm_n6202, in_21, gm_n45);
	or (gm_n6204, gm_n64, in_7, in_6, gm_n161, gm_n51);
	nor (gm_n6205, in_12, in_11, gm_n52, gm_n6204, in_13);
	nand (gm_n6206, gm_n46, gm_n63, gm_n50, gm_n6205, in_17);
	nor (gm_n6207, in_20, gm_n62, gm_n47, gm_n6206, gm_n71);
	nor (gm_n6208, gm_n51, in_8, in_7, gm_n84, gm_n52);
	nand (gm_n6209, gm_n49, in_12, gm_n53, gm_n6208, gm_n50);
	nor (gm_n6210, gm_n81, in_16, in_15, gm_n6209, in_18);
	nand (gm_n6211, in_21, in_20, in_19, gm_n6210);
	or (gm_n6212, in_12, in_11, in_10, gm_n2043, gm_n49);
	nor (gm_n6213, in_16, in_15, gm_n50, gm_n6212, gm_n81);
	nand (gm_n6214, in_20, gm_n62, in_18, gm_n6213, in_21);
	nor (gm_n6215, in_16, in_15, in_14, gm_n904, gm_n81);
	nand (gm_n6216, in_20, gm_n62, gm_n47, gm_n6215, gm_n71);
	nor (gm_n6217, in_8, in_7, in_6, gm_n530, in_9);
	nand (gm_n6218, gm_n48, in_11, gm_n52, gm_n6217, gm_n49);
	nor (gm_n6219, gm_n46, in_15, in_14, gm_n6218, in_17);
	nand (gm_n6220, in_20, gm_n62, in_18, gm_n6219, gm_n71);
	nand (gm_n6221, gm_n53, gm_n52, in_9, gm_n668);
	nor (gm_n6222, in_14, gm_n49, in_12, gm_n6221);
	nand (gm_n6223, in_17, in_16, in_15, gm_n6222, gm_n47);
	nor (gm_n6224, gm_n71, gm_n45, in_19, gm_n6223);
	nor (gm_n6225, gm_n49, gm_n48, in_11, gm_n1953, in_14);
	nand (gm_n6226, gm_n81, in_16, gm_n63, gm_n6225, in_18);
	nor (gm_n6227, in_21, in_20, gm_n62, gm_n6226);
	nand (gm_n6228, in_17, gm_n46, gm_n63, gm_n6165, gm_n47);
	nor (gm_n6229, in_21, in_20, in_19, gm_n6228);
	and (gm_n6230, in_12, gm_n53, gm_n52, gm_n375, in_13);
	nand (gm_n6231, gm_n46, in_15, in_14, gm_n6230, gm_n81);
	nor (gm_n6232, gm_n45, gm_n62, in_18, gm_n6231, gm_n71);
	nand (gm_n6233, gm_n49, gm_n48, in_11, gm_n3615, in_14);
	nor (gm_n6234, gm_n81, in_16, in_15, gm_n6233, gm_n47);
	nand (gm_n6235, in_21, gm_n45, in_19, gm_n6234);
	and (gm_n6236, gm_n53, gm_n52, gm_n51, gm_n3856);
	nand (gm_n6237, in_14, in_13, in_12, gm_n6236, gm_n63);
	nor (gm_n6238, gm_n47, in_17, in_16, gm_n6237, in_19);
	nand (gm_n6239, gm_n6238, gm_n71, gm_n45);
	nor (gm_n6240, in_11, gm_n52, in_9, gm_n1434);
	nand (gm_n6241, in_14, in_13, in_12, gm_n6240, gm_n63);
	nor (gm_n6242, gm_n47, gm_n81, gm_n46, gm_n6241, gm_n62);
	nand (gm_n6243, gm_n6242, in_21, gm_n45);
	nand (gm_n6244, gm_n50, in_13, gm_n48, gm_n1122, gm_n63);
	nor (gm_n6245, gm_n47, gm_n81, in_16, gm_n6244, in_19);
	nand (gm_n6246, gm_n6245, gm_n71, in_20);
	nand (gm_n6247, in_12, in_11, gm_n52, gm_n3744, in_13);
	nor (gm_n6248, gm_n46, in_15, gm_n50, gm_n6247, in_17);
	nand (gm_n6249, in_20, in_19, gm_n47, gm_n6248, in_21);
	nand (gm_n6250, gm_n6243, gm_n6239, gm_n6235, gm_n6249, gm_n6246);
	nor (gm_n6251, gm_n6229, gm_n6227, gm_n6224, gm_n6250, gm_n6232);
	nand (gm_n6252, gm_n6216, gm_n6214, gm_n6211, gm_n6251, gm_n6220);
	nor (gm_n6253, gm_n6203, gm_n6200, gm_n6196, gm_n6252, gm_n6207);
	nand (gm_n6254, gm_n6190, gm_n6187, gm_n6183, gm_n6253, gm_n6192);
	nor (gm_n6255, gm_n6177, gm_n6174, gm_n6171, gm_n6254, gm_n6180);
	nand (gm_n6256, gm_n6163, gm_n6159, gm_n6154, gm_n6255, gm_n6167);
	nor (gm_n6257, gm_n6146, gm_n6142, gm_n6138, gm_n6256, gm_n6150);
	nand (gm_n6258, gm_n6132, gm_n6129, gm_n6127, gm_n6257, gm_n6134);
	nor (gm_n6259, gm_n6119, gm_n6116, gm_n6113, gm_n6258, gm_n6123);
	nand (gm_n6260, gm_n6108, gm_n6104, gm_n6100, gm_n6259, gm_n6110);
	nor (gm_n6261, gm_n6092, gm_n6089, gm_n6086, gm_n6260, gm_n6096);
	nand (gm_n6262, gm_n6079, gm_n6075, gm_n6072, gm_n6261, gm_n6083);
	nor (gm_n6263, gm_n6065, gm_n6062, gm_n6059, gm_n6262, gm_n6068);
	nand (gm_n6264, gm_n6051, gm_n6047, gm_n6044, gm_n6263, gm_n6055);
	nor (gm_n6265, gm_n6038, gm_n6035, gm_n6031, gm_n6264, gm_n6041);
	nand (gm_n6266, gm_n6025, gm_n6022, gm_n6019, gm_n6265, gm_n6028);
	nor (gm_n6267, gm_n6013, gm_n6010, gm_n6007, gm_n6266, gm_n6017);
	nand (gm_n6268, gm_n6002, gm_n5999, gm_n5996, gm_n6267, gm_n6004);
	nor (gm_n6269, gm_n5989, gm_n5986, gm_n5984, gm_n6268, gm_n5992);
	nand (gm_n6270, gm_n5976, gm_n5973, gm_n5969, gm_n6269, gm_n5980);
	nor (gm_n6271, gm_n5962, gm_n5958, gm_n5955, gm_n6270, gm_n5965);
	nand (gm_n6272, gm_n5947, gm_n5943, gm_n5941, gm_n6271, gm_n5951);
	nor (gm_n6273, gm_n5935, gm_n5931, gm_n5927, gm_n6272, gm_n5938);
	nand (gm_n6274, gm_n5920, gm_n5916, gm_n5912, gm_n6273, gm_n5923);
	nor (gm_n6275, gm_n5905, gm_n5902, gm_n5899, gm_n6274, gm_n5909);
	nand (gm_n6276, gm_n5892, gm_n5887, gm_n5884, gm_n6275, gm_n5896);
	nor (gm_n6277, gm_n5876, gm_n5873, gm_n5870, gm_n6276, gm_n5880);
	nand (gm_n6278, gm_n5864, gm_n5861, gm_n5857, gm_n6277, gm_n5868);
	nor (gm_n6279, gm_n5851, gm_n5848, gm_n5845, gm_n6278, gm_n5854);
	nand (gm_n6280, gm_n5837, gm_n5833, gm_n5831, gm_n6279, gm_n5841);
	nor (gm_n6281, gm_n5825, gm_n5821, gm_n5819, gm_n6280, gm_n5829);
	nand (gm_n6282, gm_n5812, gm_n5809, gm_n5806, gm_n6281, gm_n5815);
	nor (gm_n6283, gm_n5799, gm_n5796, gm_n5792, gm_n6282, gm_n5802);
	nand (gm_n6284, gm_n5783, gm_n5779, gm_n5775, gm_n6283, gm_n5787);
	nor (gm_n6285, gm_n5767, gm_n5763, gm_n5759, gm_n6284, gm_n5771);
	nand (gm_n6286, gm_n5752, gm_n5750, gm_n5747, gm_n6285, gm_n5755);
	nor (out_9, gm_n6286, gm_n5744);
	and (gm_n6288, gm_n50, gm_n49, gm_n48, gm_n4485, in_15);
	nand (gm_n6289, gm_n47, in_17, gm_n46, gm_n6288, gm_n62);
	nor (gm_n6290, gm_n6289, gm_n71, gm_n45);
	nand (gm_n6291, in_13, in_12, gm_n53, gm_n5932, in_14);
	nor (gm_n6292, gm_n81, gm_n46, in_15, gm_n6291, gm_n47);
	nand (gm_n6293, in_21, gm_n45, in_19, gm_n6292);
	nor (gm_n6294, gm_n51, in_8, in_7, gm_n843);
	nand (gm_n6295, in_12, gm_n53, gm_n52, gm_n6294, gm_n49);
	nor (gm_n6296, gm_n46, in_15, gm_n50, gm_n6295, in_17);
	nand (gm_n6297, gm_n45, gm_n62, in_18, gm_n6296, in_21);
	nand (gm_n6298, in_13, in_12, gm_n53, gm_n137, gm_n50);
	nor (gm_n6299, in_17, gm_n46, gm_n63, gm_n6298, in_18);
	nand (gm_n6300, in_21, gm_n45, gm_n62, gm_n6299);
	nor (gm_n6301, in_9, in_8, gm_n55, gm_n223, gm_n52);
	nand (gm_n6302, gm_n49, gm_n48, in_11, gm_n6301, in_14);
	nor (gm_n6303, in_17, gm_n46, gm_n63, gm_n6302, in_18);
	nand (gm_n6304, gm_n71, gm_n45, in_19, gm_n6303);
	nand (gm_n6305, gm_n1583, in_10, in_9);
	nor (gm_n6306, in_13, gm_n48, gm_n53, gm_n6305, gm_n50);
	nand (gm_n6307, gm_n81, gm_n46, gm_n63, gm_n6306, gm_n47);
	nor (gm_n6308, gm_n71, in_20, in_19, gm_n6307);
	or (gm_n6309, gm_n390, in_9, in_8);
	nor (gm_n6310, gm_n48, gm_n53, gm_n52, gm_n6309, gm_n49);
	nand (gm_n6311, in_16, in_15, in_14, gm_n6310, in_17);
	nor (gm_n6312, gm_n45, gm_n62, gm_n47, gm_n6311, in_21);
	and (gm_n6313, gm_n3451, in_10, gm_n51);
	and (gm_n6314, in_13, in_12, in_11, gm_n6313, in_14);
	nand (gm_n6315, gm_n81, gm_n46, in_15, gm_n6314, gm_n47);
	nor (gm_n6316, in_21, gm_n45, in_19, gm_n6315);
	nand (gm_n6317, in_10, gm_n51, in_8, gm_n1608, in_11);
	nor (gm_n6318, in_14, in_13, in_12, gm_n6317, in_15);
	nand (gm_n6319, gm_n47, in_17, in_16, gm_n6318, in_19);
	nor (gm_n6320, gm_n6319, gm_n71, in_20);
	nand (gm_n6321, in_12, gm_n53, gm_n52, gm_n2877, in_13);
	nor (gm_n6322, in_16, in_15, in_14, gm_n6321, gm_n81);
	nand (gm_n6323, in_20, in_19, gm_n47, gm_n6322, in_21);
	nand (gm_n6324, gm_n50, gm_n49, in_12, gm_n3210, gm_n63);
	nor (gm_n6325, gm_n47, gm_n81, in_16, gm_n6324, in_19);
	nand (gm_n6326, gm_n6325, gm_n71, in_20);
	nor (gm_n6327, in_9, in_8, gm_n55, gm_n553, in_10);
	nand (gm_n6328, in_13, gm_n48, in_11, gm_n6327, in_14);
	nor (gm_n6329, in_17, gm_n46, in_15, gm_n6328, in_18);
	nand (gm_n6330, gm_n71, in_20, gm_n62, gm_n6329);
	nor (gm_n6331, gm_n3174, gm_n51, in_8);
	nand (gm_n6332, gm_n48, gm_n53, in_10, gm_n6331, gm_n49);
	nor (gm_n6333, gm_n46, in_15, gm_n50, gm_n6332, in_17);
	nand (gm_n6334, gm_n45, in_19, in_18, gm_n6333, in_21);
	and (gm_n6335, gm_n48, gm_n53, gm_n52, gm_n5893, in_13);
	nand (gm_n6336, gm_n46, in_15, gm_n50, gm_n6335, gm_n81);
	nor (gm_n6337, in_20, gm_n62, in_18, gm_n6336, gm_n71);
	nand (gm_n6338, in_11, gm_n52, in_9, gm_n1057, in_12);
	nor (gm_n6339, gm_n6338, gm_n49);
	nand (gm_n6340, gm_n46, in_15, in_14, gm_n6339, gm_n81);
	nor (gm_n6341, in_20, gm_n62, gm_n47, gm_n6340, gm_n71);
	and (gm_n6342, in_8, in_7, in_6, gm_n2640, gm_n51);
	and (gm_n6343, gm_n48, gm_n53, gm_n52, gm_n6342, in_13);
	nand (gm_n6344, gm_n46, gm_n63, in_14, gm_n6343, gm_n81);
	nor (gm_n6345, gm_n45, in_19, in_18, gm_n6344, in_21);
	nand (gm_n6346, gm_n46, gm_n63, in_14, gm_n6230, in_17);
	nor (gm_n6347, gm_n45, gm_n62, in_18, gm_n6346, in_21);
	and (gm_n6348, gm_n53, gm_n52, gm_n51, gm_n232, in_12);
	nand (gm_n6349, in_15, gm_n50, gm_n49, gm_n6348, in_16);
	nor (gm_n6350, gm_n62, gm_n47, in_17, gm_n6349, in_20);
	nand (gm_n6351, gm_n6350, gm_n71);
	nand (gm_n6352, in_15, gm_n50, gm_n49, gm_n674, gm_n46);
	nor (gm_n6353, gm_n62, gm_n47, in_17, gm_n6352, gm_n45);
	nand (gm_n6354, gm_n6353, in_21);
	and (gm_n6355, gm_n53, in_10, gm_n51, gm_n1683);
	nand (gm_n6356, gm_n50, gm_n49, gm_n48, gm_n6355, in_15);
	nor (gm_n6357, gm_n47, gm_n81, in_16, gm_n6356, in_19);
	nand (gm_n6358, gm_n6357, in_21, gm_n45);
	nand (gm_n6359, in_12, gm_n53, in_10, gm_n1675, gm_n49);
	nor (gm_n6360, gm_n46, in_15, gm_n50, gm_n6359, in_17);
	nand (gm_n6361, in_20, in_19, gm_n47, gm_n6360, gm_n71);
	nand (gm_n6362, in_9, in_8, in_7, gm_n151, gm_n52);
	nor (gm_n6363, gm_n49, in_12, in_11, gm_n6362, in_14);
	nand (gm_n6364, gm_n81, gm_n46, gm_n63, gm_n6363, in_18);
	nor (gm_n6365, in_21, in_20, in_19, gm_n6364);
	nor (gm_n6366, gm_n48, in_11, gm_n52, gm_n4169, in_13);
	nand (gm_n6367, gm_n46, gm_n63, in_14, gm_n6366, in_17);
	nor (gm_n6368, gm_n45, gm_n62, in_18, gm_n6367, in_21);
	or (gm_n6369, in_16, gm_n63, gm_n50, gm_n2044, in_17);
	nor (gm_n6370, in_20, in_19, in_18, gm_n6369, gm_n71);
	and (gm_n6371, in_13, gm_n48, gm_n53, gm_n6105, gm_n50);
	nand (gm_n6372, in_17, in_16, gm_n63, gm_n6371, in_18);
	nor (gm_n6373, in_21, gm_n45, in_19, gm_n6372);
	nor (gm_n6374, gm_n53, in_10, in_9, gm_n774, in_12);
	nand (gm_n6375, gm_n63, gm_n50, gm_n49, gm_n6374, gm_n46);
	nor (gm_n6376, gm_n62, in_18, in_17, gm_n6375, in_20);
	nand (gm_n6377, gm_n6376, gm_n71);
	nor (gm_n6378, gm_n53, in_10, gm_n51, gm_n1052, gm_n48);
	nand (gm_n6379, in_15, gm_n50, gm_n49, gm_n6378, gm_n46);
	nor (gm_n6380, in_19, gm_n47, gm_n81, gm_n6379, in_20);
	nand (gm_n6381, gm_n6380, gm_n71);
	nand (gm_n6382, in_12, gm_n53, gm_n52, gm_n1759, gm_n49);
	nor (gm_n6383, in_16, in_15, in_14, gm_n6382, gm_n81);
	nand (gm_n6384, gm_n45, gm_n62, gm_n47, gm_n6383, in_21);
	nand (gm_n6385, gm_n63, gm_n50, gm_n49, gm_n5944, in_16);
	nor (gm_n6386, in_19, gm_n47, in_17, gm_n6385, in_20);
	nand (gm_n6387, gm_n6386, gm_n71);
	nor (gm_n6388, in_12, in_11, gm_n52, gm_n4362, gm_n49);
	nand (gm_n6389, in_16, in_15, gm_n50, gm_n6388, in_17);
	nor (gm_n6390, in_20, gm_n62, in_18, gm_n6389, gm_n71);
	nor (gm_n6391, in_12, in_11, gm_n52, gm_n5030, in_13);
	nand (gm_n6392, gm_n46, in_15, gm_n50, gm_n6391, gm_n81);
	nor (gm_n6393, gm_n45, in_19, gm_n47, gm_n6392, gm_n71);
	nor (gm_n6394, gm_n63, in_14, in_13, gm_n3501, gm_n46);
	nand (gm_n6395, gm_n62, in_18, in_17, gm_n6394, gm_n45);
	nor (gm_n6396, gm_n6395, in_21);
	nand (gm_n6397, gm_n1044, gm_n52, in_9);
	nor (gm_n6398, gm_n49, in_12, gm_n53, gm_n6397, gm_n50);
	nand (gm_n6399, gm_n81, in_16, gm_n63, gm_n6398, gm_n47);
	nor (gm_n6400, in_21, gm_n45, in_19, gm_n6399);
	nor (gm_n6401, gm_n3484, in_10, in_9);
	nand (gm_n6402, gm_n49, in_12, gm_n53, gm_n6401, in_14);
	nor (gm_n6403, in_17, gm_n46, in_15, gm_n6402, in_18);
	nand (gm_n6404, in_21, in_20, in_19, gm_n6403);
	and (gm_n6405, gm_n316, in_9, gm_n64);
	nand (gm_n6406, in_12, gm_n53, in_10, gm_n6405, gm_n49);
	nor (gm_n6407, in_16, in_15, gm_n50, gm_n6406, in_17);
	nand (gm_n6408, in_20, in_19, in_18, gm_n6407, gm_n71);
	nor (gm_n6409, gm_n53, in_10, gm_n51, gm_n440);
	nand (gm_n6410, gm_n50, gm_n49, gm_n48, gm_n6409, in_15);
	nor (gm_n6411, in_18, gm_n81, in_16, gm_n6410, in_19);
	nand (gm_n6412, gm_n6411, gm_n71, gm_n45);
	nand (gm_n6413, gm_n63, in_14, gm_n49, gm_n3880, gm_n46);
	nor (gm_n6414, in_19, gm_n47, gm_n81, gm_n6413, gm_n45);
	nand (gm_n6415, gm_n6414, in_21);
	nor (gm_n6416, gm_n48, gm_n53, in_10, gm_n1599, gm_n49);
	nand (gm_n6417, in_16, in_15, gm_n50, gm_n6416, in_17);
	nor (gm_n6418, gm_n45, gm_n62, gm_n47, gm_n6417, gm_n71);
	and (gm_n6419, gm_n48, gm_n53, gm_n52, gm_n2877, gm_n49);
	nand (gm_n6420, gm_n46, gm_n63, in_14, gm_n6419, in_17);
	nor (gm_n6421, in_20, in_19, gm_n47, gm_n6420, in_21);
	nand (gm_n6422, in_11, gm_n52, gm_n51, gm_n1583, gm_n48);
	nor (gm_n6423, gm_n63, in_14, gm_n49, gm_n6422, gm_n46);
	nand (gm_n6424, in_19, in_18, in_17, gm_n6423, gm_n45);
	nor (gm_n6425, gm_n6424, in_21);
	and (gm_n6426, in_11, gm_n52, in_9, gm_n5340, gm_n48);
	and (gm_n6427, in_15, in_14, gm_n49, gm_n6426, in_16);
	nand (gm_n6428, in_19, gm_n47, gm_n81, gm_n6427, gm_n45);
	nor (gm_n6429, gm_n6428, gm_n71);
	and (gm_n6430, in_8, gm_n55, in_6, gm_n2640, in_9);
	nand (gm_n6431, gm_n48, gm_n53, gm_n52, gm_n6430, gm_n49);
	nor (gm_n6432, gm_n46, gm_n63, in_14, gm_n6431, gm_n81);
	nand (gm_n6433, gm_n45, in_19, in_18, gm_n6432, in_21);
	or (gm_n6434, gm_n48, in_11, gm_n52, gm_n6032, in_13);
	nor (gm_n6435, gm_n46, in_15, gm_n50, gm_n6434, gm_n81);
	nand (gm_n6436, in_20, in_19, in_18, gm_n6435, gm_n71);
	and (gm_n6437, gm_n47, gm_n81, gm_n46, gm_n4559, gm_n62);
	nand (gm_n6438, gm_n6437, gm_n71, gm_n45);
	nand (gm_n6439, gm_n63, gm_n50, gm_n49, gm_n4784, in_16);
	nor (gm_n6440, gm_n62, in_18, gm_n81, gm_n6439, gm_n45);
	nand (gm_n6441, gm_n6440, in_21);
	and (gm_n6442, gm_n49, in_12, gm_n53, gm_n3320, gm_n50);
	nand (gm_n6443, in_17, gm_n46, in_15, gm_n6442, in_18);
	nor (gm_n6444, gm_n71, gm_n45, in_19, gm_n6443);
	and (gm_n6445, gm_n49, gm_n48, in_11, gm_n4688, in_14);
	nand (gm_n6446, in_17, gm_n46, in_15, gm_n6445, gm_n47);
	nor (gm_n6447, in_21, gm_n45, gm_n62, gm_n6446);
	nor (gm_n6448, in_12, in_11, in_10, gm_n162, in_13);
	nand (gm_n6449, gm_n46, gm_n63, gm_n50, gm_n6448, in_17);
	nor (gm_n6450, gm_n45, in_19, in_18, gm_n6449, gm_n71);
	nand (gm_n6451, gm_n2699, in_9);
	nor (gm_n6452, gm_n48, gm_n53, in_10, gm_n6451, in_13);
	nand (gm_n6453, gm_n46, gm_n63, in_14, gm_n6452, gm_n81);
	nor (gm_n6454, gm_n45, gm_n62, gm_n47, gm_n6453, gm_n71);
	nand (gm_n6455, in_12, in_11, in_10, gm_n4329, in_13);
	nor (gm_n6456, in_16, in_15, gm_n50, gm_n6455, in_17);
	nand (gm_n6457, gm_n45, in_19, gm_n47, gm_n6456, gm_n71);
	nand (gm_n6458, gm_n50, in_13, in_12, gm_n1937, in_15);
	nor (gm_n6459, in_18, gm_n81, in_16, gm_n6458, gm_n62);
	nand (gm_n6460, gm_n6459, in_21, gm_n45);
	nand (gm_n6461, in_14, in_13, in_12, gm_n4377, gm_n63);
	nor (gm_n6462, gm_n47, in_17, in_16, gm_n6461, gm_n62);
	nand (gm_n6463, gm_n6462, gm_n71, gm_n45);
	nand (gm_n6464, gm_n50, in_13, in_12, gm_n908, in_15);
	nor (gm_n6465, gm_n47, gm_n81, in_16, gm_n6464, gm_n62);
	nand (gm_n6466, gm_n6465, in_21, gm_n45);
	nand (gm_n6467, gm_n53, gm_n52, in_9, gm_n3086, gm_n48);
	nor (gm_n6468, in_15, in_14, in_13, gm_n6467, gm_n46);
	nand (gm_n6469, in_19, in_18, in_17, gm_n6468, in_20);
	nor (gm_n6470, gm_n6469, gm_n71);
	nand (gm_n6471, in_11, gm_n52, in_9, gm_n484, in_12);
	nor (gm_n6472, gm_n6471, gm_n49);
	nand (gm_n6473, gm_n46, in_15, in_14, gm_n6472, gm_n81);
	nor (gm_n6474, in_20, gm_n62, in_18, gm_n6473, in_21);
	or (gm_n6475, in_8, in_7, in_6, gm_n1429, gm_n51);
	nor (gm_n6476, in_12, in_11, gm_n52, gm_n6475, gm_n49);
	nand (gm_n6477, gm_n46, in_15, in_14, gm_n6476, gm_n81);
	nor (gm_n6478, gm_n45, in_19, gm_n47, gm_n6477, in_21);
	or (gm_n6479, in_7, gm_n82, in_5, gm_n124, in_8);
	nor (gm_n6480, in_11, in_10, in_9, gm_n6479, in_12);
	nand (gm_n6481, gm_n63, in_14, in_13, gm_n6480, in_16);
	or (gm_n6482, in_19, gm_n47, in_17, gm_n6481, in_20);
	nor (gm_n6483, gm_n6482, gm_n71);
	nand (gm_n6484, in_15, gm_n50, gm_n49, gm_n5248, gm_n46);
	nor (gm_n6485, gm_n62, gm_n47, gm_n81, gm_n6484, in_20);
	nand (gm_n6486, gm_n6485, in_21);
	nor (gm_n6487, gm_n53, gm_n52, gm_n51, gm_n4489, gm_n48);
	nand (gm_n6488, gm_n63, gm_n50, in_13, gm_n6487, gm_n46);
	nor (gm_n6489, in_19, in_18, gm_n81, gm_n6488, gm_n45);
	nand (gm_n6490, gm_n6489, in_21);
	nand (gm_n6491, gm_n48, in_11, gm_n52, gm_n1932, in_13);
	nor (gm_n6492, gm_n46, in_15, in_14, gm_n6491, gm_n81);
	nand (gm_n6493, in_20, in_19, gm_n47, gm_n6492, in_21);
	nor (gm_n6494, gm_n46, gm_n63, gm_n50, gm_n4158, gm_n81);
	nand (gm_n6495, in_20, gm_n62, gm_n47, gm_n6494, in_21);
	nor (gm_n6496, in_11, in_10, gm_n51, gm_n955, in_12);
	and (gm_n6497, gm_n63, in_14, in_13, gm_n6496, gm_n46);
	nand (gm_n6498, gm_n62, gm_n47, gm_n81, gm_n6497, gm_n45);
	nor (gm_n6499, gm_n6498, in_21);
	nor (gm_n6500, gm_n55, gm_n82, gm_n72, gm_n130, gm_n64);
	nand (gm_n6501, in_11, in_10, gm_n51, gm_n6500, in_12);
	nor (gm_n6502, in_15, gm_n50, gm_n49, gm_n6501, in_16);
	nand (gm_n6503, gm_n62, in_18, in_17, gm_n6502, gm_n45);
	nor (gm_n6504, gm_n6503, in_21);
	nor (gm_n6505, in_12, gm_n53, gm_n52, gm_n1617, gm_n49);
	nand (gm_n6506, gm_n46, in_15, gm_n50, gm_n6505, in_17);
	nor (gm_n6507, in_20, in_19, gm_n47, gm_n6506, gm_n71);
	nand (gm_n6508, gm_n53, gm_n52, gm_n51, gm_n4723, gm_n48);
	nor (gm_n6509, gm_n63, gm_n50, in_13, gm_n6508, gm_n46);
	nand (gm_n6510, in_19, gm_n47, gm_n81, gm_n6509, gm_n45);
	nor (gm_n6511, gm_n6510, in_21);
	nor (gm_n6512, in_17, in_16, in_15, gm_n3074, in_18);
	nand (gm_n6513, gm_n71, in_20, in_19, gm_n6512);
	and (gm_n6514, gm_n53, in_10, gm_n51, gm_n4042, in_12);
	nand (gm_n6515, in_15, in_14, gm_n49, gm_n6514, in_16);
	nor (gm_n6516, gm_n62, gm_n47, gm_n81, gm_n6515, in_20);
	nand (gm_n6517, gm_n6516, gm_n71);
	or (gm_n6518, gm_n64, gm_n55, gm_n82, gm_n199, in_9);
	or (gm_n6519, in_12, gm_n53, in_10, gm_n6518, gm_n49);
	nor (gm_n6520, gm_n46, in_15, in_14, gm_n6519, in_17);
	nand (gm_n6521, in_20, gm_n62, in_18, gm_n6520, in_21);
	or (gm_n6522, gm_n63, gm_n50, gm_n49, gm_n515, gm_n46);
	nor (gm_n6523, gm_n62, in_18, in_17, gm_n6522, in_20);
	nand (gm_n6524, gm_n6523, gm_n71);
	and (gm_n6525, gm_n2034, in_9);
	and (gm_n6526, gm_n48, in_11, in_10, gm_n6525, in_13);
	nand (gm_n6527, in_16, in_15, gm_n50, gm_n6526, gm_n81);
	nor (gm_n6528, in_20, gm_n62, in_18, gm_n6527, in_21);
	nor (gm_n6529, gm_n48, gm_n53, gm_n52, gm_n411, gm_n49);
	nand (gm_n6530, gm_n46, gm_n63, in_14, gm_n6529, gm_n81);
	nor (gm_n6531, gm_n45, in_19, gm_n47, gm_n6530, gm_n71);
	nand (gm_n6532, in_11, gm_n52, in_9, gm_n1563, gm_n48);
	nor (gm_n6533, in_15, gm_n50, in_13, gm_n6532, in_16);
	nand (gm_n6534, gm_n62, in_18, in_17, gm_n6533, in_20);
	nor (gm_n6535, gm_n6534, in_21);
	nor (gm_n6536, gm_n50, gm_n49, gm_n48, gm_n4494, in_15);
	nand (gm_n6537, gm_n47, gm_n81, gm_n46, gm_n6536, gm_n62);
	nor (gm_n6538, gm_n6537, in_21, in_20);
	nor (gm_n6539, gm_n64, in_7, gm_n82, gm_n103, in_9);
	nand (gm_n6540, gm_n48, in_11, gm_n52, gm_n6539, gm_n49);
	nor (gm_n6541, in_16, in_15, gm_n50, gm_n6540, gm_n81);
	nand (gm_n6542, in_20, in_19, gm_n47, gm_n6541, gm_n71);
	nand (gm_n6543, in_13, in_12, in_11, gm_n3189, gm_n50);
	nor (gm_n6544, gm_n81, in_16, gm_n63, gm_n6543, in_18);
	nand (gm_n6545, gm_n71, gm_n45, gm_n62, gm_n6544);
	nand (gm_n6546, gm_n48, gm_n53, gm_n52, gm_n1688, in_13);
	nor (gm_n6547, in_16, in_15, in_14, gm_n6546, gm_n81);
	nand (gm_n6548, gm_n45, gm_n62, gm_n47, gm_n6547, gm_n71);
	and (gm_n6549, in_7, gm_n82, gm_n72, gm_n209, in_8);
	and (gm_n6550, gm_n53, in_10, in_9, gm_n6549);
	nand (gm_n6551, in_14, in_13, in_12, gm_n6550, in_15);
	nor (gm_n6552, gm_n47, gm_n81, in_16, gm_n6551, gm_n62);
	nand (gm_n6553, gm_n6552, gm_n71, in_20);
	nor (gm_n6554, gm_n49, gm_n48, in_11, gm_n464, gm_n50);
	nand (gm_n6555, gm_n81, in_16, gm_n63, gm_n6554, in_18);
	nor (gm_n6556, in_21, in_20, in_19, gm_n6555);
	and (gm_n6557, in_14, in_13, in_12, gm_n2371, in_15);
	nand (gm_n6558, in_18, gm_n81, gm_n46, gm_n6557, in_19);
	nor (gm_n6559, gm_n6558, in_21, in_20);
	nand (gm_n6560, in_11, in_10, in_9, gm_n509, gm_n48);
	nor (gm_n6561, gm_n63, in_14, in_13, gm_n6560, gm_n46);
	nand (gm_n6562, gm_n62, gm_n47, gm_n81, gm_n6561, gm_n45);
	nor (gm_n6563, gm_n6562, gm_n71);
	and (gm_n6564, gm_n53, gm_n52, gm_n51, gm_n3299);
	and (gm_n6565, in_14, in_13, in_12, gm_n6564, in_15);
	nand (gm_n6566, gm_n47, in_17, gm_n46, gm_n6565, in_19);
	nor (gm_n6567, gm_n6566, in_21, gm_n45);
	and (gm_n6568, gm_n3804, in_10, gm_n51);
	nand (gm_n6569, in_13, in_12, gm_n53, gm_n6568, gm_n50);
	nor (gm_n6570, gm_n81, in_16, gm_n63, gm_n6569, gm_n47);
	nand (gm_n6571, in_21, gm_n45, in_19, gm_n6570);
	nor (gm_n6572, gm_n2559, gm_n51);
	nand (gm_n6573, gm_n48, gm_n53, gm_n52, gm_n6572, in_13);
	nor (gm_n6574, in_16, gm_n63, in_14, gm_n6573, in_17);
	nand (gm_n6575, in_20, in_19, gm_n47, gm_n6574, gm_n71);
	nor (gm_n6576, gm_n916, gm_n52, gm_n51);
	nand (gm_n6577, gm_n49, gm_n48, gm_n53, gm_n6576, in_14);
	nor (gm_n6578, in_17, in_16, in_15, gm_n6577, in_18);
	nand (gm_n6579, gm_n71, gm_n45, gm_n62, gm_n6578);
	nand (gm_n6580, gm_n48, in_11, in_10, gm_n2555, gm_n49);
	nor (gm_n6581, in_16, in_15, in_14, gm_n6580, in_17);
	nand (gm_n6582, in_20, gm_n62, in_18, gm_n6581, gm_n71);
	and (gm_n6583, gm_n3183, in_9);
	and (gm_n6584, gm_n48, gm_n53, in_10, gm_n6583, in_13);
	nand (gm_n6585, in_16, in_15, gm_n50, gm_n6584, in_17);
	nor (gm_n6586, gm_n45, in_19, gm_n47, gm_n6585, in_21);
	nor (gm_n6587, gm_n48, gm_n53, gm_n52, gm_n1117, in_13);
	nand (gm_n6588, gm_n46, gm_n63, gm_n50, gm_n6587, in_17);
	nor (gm_n6589, in_20, gm_n62, in_18, gm_n6588, in_21);
	nand (gm_n6590, in_18, gm_n81, in_16, gm_n6169, in_19);
	nor (gm_n6591, gm_n6590, gm_n71, gm_n45);
	nand (gm_n6592, gm_n53, in_10, in_9, gm_n1895);
	nor (gm_n6593, gm_n50, in_13, in_12, gm_n6592, in_15);
	nand (gm_n6594, in_18, gm_n81, in_16, gm_n6593, in_19);
	nor (gm_n6595, gm_n6594, in_21, gm_n45);
	nand (gm_n6596, gm_n50, in_13, in_12, gm_n4999, in_15);
	nor (gm_n6597, in_18, gm_n81, in_16, gm_n6596, in_19);
	nand (gm_n6598, gm_n6597, gm_n71, in_20);
	nand (gm_n6599, gm_n48, in_11, gm_n52, gm_n3309, in_13);
	nor (gm_n6600, in_16, in_15, gm_n50, gm_n6599, gm_n81);
	nand (gm_n6601, gm_n45, in_19, in_18, gm_n6600, in_21);
	nand (gm_n6602, in_14, gm_n49, gm_n48, gm_n469, in_15);
	nor (gm_n6603, gm_n47, in_17, in_16, gm_n6602, in_19);
	nand (gm_n6604, gm_n6603, in_21, gm_n45);
	nand (gm_n6605, in_9, in_8, in_7, gm_n1007, gm_n52);
	or (gm_n6606, in_13, gm_n48, in_11, gm_n6605);
	nor (gm_n6607, in_16, gm_n63, in_14, gm_n6606, gm_n81);
	nand (gm_n6608, in_20, in_19, gm_n47, gm_n6607, gm_n71);
	nand (gm_n6609, gm_n52, in_9, gm_n64, gm_n838);
	nor (gm_n6610, in_13, in_12, gm_n53, gm_n6609, in_14);
	nand (gm_n6611, gm_n81, in_16, in_15, gm_n6610, in_18);
	nor (gm_n6612, in_21, gm_n45, gm_n62, gm_n6611);
	nand (gm_n6613, in_11, gm_n52, gm_n51, gm_n1279, in_12);
	nor (gm_n6614, in_15, in_14, gm_n49, gm_n6613, gm_n46);
	nand (gm_n6615, in_19, gm_n47, gm_n81, gm_n6614, gm_n45);
	nor (gm_n6616, gm_n6615, in_21);
	nand (gm_n6617, in_11, gm_n52, in_9, gm_n593, gm_n48);
	nor (gm_n6618, gm_n63, gm_n50, gm_n49, gm_n6617, in_16);
	nand (gm_n6619, in_19, gm_n47, in_17, gm_n6618, in_20);
	nor (gm_n6620, gm_n6619, gm_n71);
	nand (gm_n6621, gm_n52, gm_n51, gm_n64, gm_n5788);
	nor (gm_n6622, in_13, in_12, in_11, gm_n6621);
	nand (gm_n6623, in_16, in_15, gm_n50, gm_n6622, in_17);
	nor (gm_n6624, in_20, in_19, gm_n47, gm_n6623, gm_n71);
	nand (gm_n6625, gm_n48, gm_n53, in_10, gm_n1966, in_13);
	nor (gm_n6626, in_16, in_15, in_14, gm_n6625, in_17);
	nand (gm_n6627, gm_n45, in_19, gm_n47, gm_n6626, gm_n71);
	nand (gm_n6628, gm_n49, gm_n48, gm_n53, gm_n3253, in_14);
	nor (gm_n6629, in_17, gm_n46, in_15, gm_n6628, gm_n47);
	nand (gm_n6630, in_21, gm_n45, gm_n62, gm_n6629);
	nand (gm_n6631, in_14, gm_n49, in_12, gm_n4315, gm_n63);
	nor (gm_n6632, in_18, in_17, in_16, gm_n6631, in_19);
	nand (gm_n6633, gm_n6632, gm_n71, gm_n45);
	nand (gm_n6634, gm_n50, gm_n49, gm_n48, gm_n6564, in_15);
	nor (gm_n6635, in_18, in_17, gm_n46, gm_n6634, in_19);
	nand (gm_n6636, gm_n6635, gm_n71, in_20);
	nor (gm_n6637, gm_n48, gm_n53, in_10, gm_n1430, in_13);
	nand (gm_n6638, in_16, in_15, in_14, gm_n6637, gm_n81);
	nor (gm_n6639, gm_n45, in_19, in_18, gm_n6638, in_21);
	nor (gm_n6640, gm_n50, gm_n49, in_12, gm_n2832, gm_n63);
	nand (gm_n6641, gm_n47, in_17, in_16, gm_n6640, in_19);
	nor (gm_n6642, gm_n6641, in_21, in_20);
	nor (gm_n6643, gm_n55, gm_n82, gm_n72, gm_n130, in_8);
	nand (gm_n6644, gm_n6643, gm_n52, gm_n51);
	nor (gm_n6645, gm_n49, gm_n48, gm_n53, gm_n6644, in_14);
	nand (gm_n6646, gm_n81, gm_n46, gm_n63, gm_n6645, gm_n47);
	nor (gm_n6647, gm_n71, in_20, gm_n62, gm_n6646);
	nor (gm_n6648, gm_n50, gm_n49, in_12, gm_n1348, in_15);
	nand (gm_n6649, in_18, in_17, gm_n46, gm_n6648, gm_n62);
	nor (gm_n6650, gm_n6649, in_21, gm_n45);
	nand (gm_n6651, gm_n48, gm_n53, gm_n52, gm_n3562, gm_n49);
	nor (gm_n6652, in_16, gm_n63, gm_n50, gm_n6651, gm_n81);
	nand (gm_n6653, in_20, in_19, in_18, gm_n6652, gm_n71);
	nand (gm_n6654, gm_n48, in_11, gm_n52, gm_n2555, gm_n49);
	nor (gm_n6655, in_16, gm_n63, in_14, gm_n6654, in_17);
	nand (gm_n6656, in_20, gm_n62, in_18, gm_n6655, gm_n71);
	nor (gm_n6657, in_9, in_8, gm_n55, gm_n1256, in_10);
	nand (gm_n6658, gm_n49, gm_n48, gm_n53, gm_n6657, in_14);
	nor (gm_n6659, in_17, in_16, in_15, gm_n6658, in_18);
	nand (gm_n6660, in_21, gm_n45, gm_n62, gm_n6659);
	nand (gm_n6661, in_12, gm_n53, in_10, gm_n3354, gm_n49);
	nor (gm_n6662, in_16, gm_n63, in_14, gm_n6661, in_17);
	nand (gm_n6663, in_20, gm_n62, gm_n47, gm_n6662, in_21);
	nand (gm_n6664, in_11, gm_n52, in_9, gm_n1952, in_12);
	nor (gm_n6665, in_15, in_14, in_13, gm_n6664, in_16);
	nand (gm_n6666, in_19, gm_n47, gm_n81, gm_n6665, gm_n45);
	nor (gm_n6667, gm_n6666, gm_n71);
	nor (gm_n6668, in_8, in_7, in_6, gm_n141, in_9);
	and (gm_n6669, gm_n48, in_11, gm_n52, gm_n6668, gm_n49);
	nand (gm_n6670, in_16, gm_n63, gm_n50, gm_n6669, gm_n81);
	nor (gm_n6671, gm_n45, gm_n62, in_18, gm_n6670, gm_n71);
	or (gm_n6672, in_8, in_7, in_6, gm_n96, gm_n51);
	nor (gm_n6673, gm_n48, gm_n53, gm_n52, gm_n6672, in_13);
	nand (gm_n6674, gm_n46, gm_n63, in_14, gm_n6673, gm_n81);
	nor (gm_n6675, gm_n45, in_19, gm_n47, gm_n6674, gm_n71);
	and (gm_n6676, gm_n50, gm_n49, gm_n48, gm_n4298, in_15);
	nand (gm_n6677, gm_n47, in_17, gm_n46, gm_n6676, in_19);
	nor (gm_n6678, gm_n6677, gm_n71, gm_n45);
	and (gm_n6679, gm_n53, gm_n52, in_9, gm_n1156, gm_n48);
	nand (gm_n6680, gm_n63, in_14, in_13, gm_n6679, gm_n46);
	nor (gm_n6681, in_19, gm_n47, gm_n81, gm_n6680, gm_n45);
	nand (gm_n6682, gm_n6681, in_21);
	and (gm_n6683, in_11, in_10, gm_n51, gm_n1634, in_12);
	nand (gm_n6684, gm_n63, gm_n50, gm_n49, gm_n6683, in_16);
	nor (gm_n6685, gm_n62, in_18, gm_n81, gm_n6684, gm_n45);
	nand (gm_n6686, gm_n6685, in_21);
	nand (gm_n6687, in_14, gm_n49, in_12, gm_n2437, gm_n63);
	nor (gm_n6688, in_18, gm_n81, in_16, gm_n6687, in_19);
	nand (gm_n6689, gm_n6688, gm_n71, in_20);
	nand (gm_n6690, gm_n49, in_12, gm_n53, gm_n1542, gm_n50);
	nor (gm_n6691, in_17, in_16, in_15, gm_n6690, in_18);
	nand (gm_n6692, gm_n71, gm_n45, gm_n62, gm_n6691);
	nand (gm_n6693, gm_n53, gm_n52, in_9, gm_n5668, gm_n48);
	nor (gm_n6694, in_15, gm_n50, gm_n49, gm_n6693, in_16);
	nand (gm_n6695, gm_n62, in_18, in_17, gm_n6694, in_20);
	nor (gm_n6696, gm_n6695, gm_n71);
	and (gm_n6697, in_12, in_11, in_10, gm_n3748, gm_n49);
	nand (gm_n6698, gm_n46, in_15, gm_n50, gm_n6697, gm_n81);
	nor (gm_n6699, in_20, in_19, gm_n47, gm_n6698, gm_n71);
	nand (gm_n6700, in_17, in_16, gm_n63, gm_n631, gm_n47);
	nor (gm_n6701, in_21, gm_n45, in_19, gm_n6700);
	nand (gm_n6702, gm_n242, in_10, gm_n51);
	nor (gm_n6703, gm_n49, in_12, in_11, gm_n6702, in_14);
	nand (gm_n6704, gm_n81, in_16, gm_n63, gm_n6703, in_18);
	nor (gm_n6705, gm_n71, gm_n45, gm_n62, gm_n6704);
	nor (gm_n6706, in_11, gm_n52, gm_n51, gm_n333, gm_n48);
	nand (gm_n6707, gm_n63, gm_n50, gm_n49, gm_n6706, gm_n46);
	nor (gm_n6708, in_19, gm_n47, gm_n81, gm_n6707, in_20);
	nand (gm_n6709, gm_n6708, in_21);
	nor (gm_n6710, gm_n53, in_10, gm_n51, gm_n2902, in_12);
	nand (gm_n6711, gm_n63, gm_n50, gm_n49, gm_n6710, in_16);
	nor (gm_n6712, gm_n62, in_18, in_17, gm_n6711, in_20);
	nand (gm_n6713, gm_n6712, gm_n71);
	nor (gm_n6714, gm_n64, gm_n55, in_6, gm_n156, gm_n51);
	nand (gm_n6715, in_12, in_11, in_10, gm_n6714, gm_n49);
	nor (gm_n6716, in_16, gm_n63, in_14, gm_n6715, gm_n81);
	nand (gm_n6717, gm_n45, in_19, in_18, gm_n6716, gm_n71);
	nor (gm_n6718, in_10, in_9, in_8, gm_n907, gm_n53);
	nand (gm_n6719, in_14, in_13, in_12, gm_n6718, in_15);
	nor (gm_n6720, in_18, gm_n81, in_16, gm_n6719, in_19);
	nand (gm_n6721, gm_n6720, gm_n71, in_20);
	and (gm_n6722, in_14, gm_n49, in_12, gm_n3633, in_15);
	nand (gm_n6723, in_18, in_17, gm_n46, gm_n6722, gm_n62);
	nor (gm_n6724, gm_n6723, in_21, in_20);
	or (gm_n6725, in_10, gm_n51, in_8, gm_n853, gm_n53);
	nor (gm_n6726, gm_n50, in_13, gm_n48, gm_n6725, gm_n63);
	nand (gm_n6727, in_18, gm_n81, in_16, gm_n6726, in_19);
	nor (gm_n6728, gm_n6727, gm_n71, in_20);
	and (gm_n6729, in_15, gm_n50, gm_n49, gm_n917, in_16);
	nand (gm_n6730, in_19, in_18, in_17, gm_n6729, in_20);
	nor (gm_n6731, gm_n6730, in_21);
	nor (gm_n6732, in_10, in_9, gm_n64, gm_n907);
	and (gm_n6733, gm_n49, in_12, gm_n53, gm_n6732, in_14);
	nand (gm_n6734, gm_n81, gm_n46, gm_n63, gm_n6733, in_18);
	nor (gm_n6735, in_21, in_20, gm_n62, gm_n6734);
	nand (gm_n6736, gm_n961, in_13, gm_n48);
	nor (gm_n6737, in_16, in_15, in_14, gm_n6736, gm_n81);
	nand (gm_n6738, gm_n45, in_19, gm_n47, gm_n6737, gm_n71);
	nand (gm_n6739, in_12, in_11, gm_n52, gm_n1808, gm_n49);
	nor (gm_n6740, gm_n46, in_15, gm_n50, gm_n6739, in_17);
	nand (gm_n6741, gm_n45, gm_n62, gm_n47, gm_n6740, in_21);
	nor (gm_n6742, gm_n3949, gm_n51);
	nand (gm_n6743, gm_n48, gm_n53, in_10, gm_n6742, in_13);
	nor (gm_n6744, in_16, gm_n63, gm_n50, gm_n6743, gm_n81);
	nand (gm_n6745, gm_n45, gm_n62, in_18, gm_n6744, gm_n71);
	nor (gm_n6746, gm_n53, gm_n52, gm_n51, gm_n571, in_12);
	nand (gm_n6747, gm_n63, in_14, gm_n49, gm_n6746, gm_n46);
	nor (gm_n6748, in_19, gm_n47, in_17, gm_n6747, in_20);
	nand (gm_n6749, gm_n6748, gm_n71);
	or (gm_n6750, in_11, in_10, in_9, gm_n3428, gm_n48);
	nor (gm_n6751, in_15, gm_n50, gm_n49, gm_n6750, gm_n46);
	nand (gm_n6752, in_19, in_18, in_17, gm_n6751, in_20);
	nor (gm_n6753, gm_n6752, in_21);
	nor (gm_n6754, gm_n48, gm_n53, in_10, gm_n2931, gm_n49);
	nand (gm_n6755, in_16, in_15, gm_n50, gm_n6754, in_17);
	nor (gm_n6756, gm_n45, gm_n62, in_18, gm_n6755, in_21);
	and (gm_n6757, gm_n48, gm_n53, gm_n52, gm_n2956, in_13);
	nand (gm_n6758, gm_n46, gm_n63, in_14, gm_n6757, gm_n81);
	nor (gm_n6759, gm_n45, gm_n62, in_18, gm_n6758, gm_n71);
	nand (gm_n6760, in_8, in_7, in_6, gm_n757, in_9);
	nor (gm_n6761, in_12, gm_n53, gm_n52, gm_n6760, gm_n49);
	nand (gm_n6762, gm_n46, in_15, in_14, gm_n6761, gm_n81);
	nor (gm_n6763, gm_n45, gm_n62, in_18, gm_n6762, gm_n71);
	and (gm_n6764, in_11, gm_n52, gm_n51, gm_n458, in_12);
	nand (gm_n6765, in_15, gm_n50, in_13, gm_n6764, gm_n46);
	nor (gm_n6766, gm_n62, gm_n47, in_17, gm_n6765, gm_n45);
	nand (gm_n6767, gm_n6766, in_21);
	or (gm_n6768, gm_n64, in_7, in_6, gm_n156, in_9);
	nor (gm_n6769, gm_n6768, gm_n52);
	nand (gm_n6770, gm_n49, in_12, gm_n53, gm_n6769, gm_n50);
	nor (gm_n6771, gm_n81, gm_n46, in_15, gm_n6770, gm_n47);
	nand (gm_n6772, in_21, in_20, in_19, gm_n6771);
	nor (gm_n6773, in_9, gm_n64, gm_n55, gm_n525, in_10);
	nand (gm_n6774, in_13, in_12, gm_n53, gm_n6773, gm_n50);
	nor (gm_n6775, gm_n81, gm_n46, gm_n63, gm_n6774, gm_n47);
	nand (gm_n6776, gm_n71, gm_n45, in_19, gm_n6775);
	nor (gm_n6777, gm_n53, in_10, in_9, gm_n2546, in_12);
	nand (gm_n6778, in_15, in_14, in_13, gm_n6777, in_16);
	nor (gm_n6779, in_19, gm_n47, gm_n81, gm_n6778, gm_n45);
	nand (gm_n6780, gm_n6779, in_21);
	or (gm_n6781, gm_n53, in_10, in_9, gm_n2564, in_12);
	nor (gm_n6782, gm_n63, gm_n50, in_13, gm_n6781, gm_n46);
	nand (gm_n6783, in_19, gm_n47, gm_n81, gm_n6782, in_20);
	nor (gm_n6784, gm_n6783, gm_n71);
	nand (gm_n6785, gm_n53, in_10, in_9, gm_n644, gm_n48);
	nor (gm_n6786, gm_n63, in_14, in_13, gm_n6785, in_16);
	nand (gm_n6787, gm_n62, in_18, gm_n81, gm_n6786, gm_n45);
	nor (gm_n6788, gm_n6787, in_21);
	nor (gm_n6789, in_11, in_10, gm_n51, gm_n1127, in_12);
	and (gm_n6790, in_15, in_14, in_13, gm_n6789, in_16);
	nand (gm_n6791, in_19, gm_n47, in_17, gm_n6790, gm_n45);
	nor (gm_n6792, gm_n6791, in_21);
	nand (gm_n6793, gm_n53, gm_n52, gm_n51, gm_n1044, gm_n48);
	nor (gm_n6794, in_15, gm_n50, in_13, gm_n6793, gm_n46);
	nand (gm_n6795, gm_n62, in_18, gm_n81, gm_n6794, gm_n45);
	nor (gm_n6796, gm_n6795, gm_n71);
	nand (gm_n6797, gm_n48, in_11, in_10, gm_n5793, gm_n49);
	nor (gm_n6798, gm_n46, in_15, in_14, gm_n6797, gm_n81);
	nand (gm_n6799, in_20, gm_n62, gm_n47, gm_n6798, gm_n71);
	and (gm_n6800, gm_n4200, gm_n52, in_9);
	nand (gm_n6801, gm_n49, gm_n48, gm_n53, gm_n6800, gm_n50);
	nor (gm_n6802, gm_n81, gm_n46, gm_n63, gm_n6801, gm_n47);
	nand (gm_n6803, gm_n71, in_20, in_19, gm_n6802);
	nor (gm_n6804, in_11, gm_n52, gm_n51, gm_n6155, in_12);
	nand (gm_n6805, in_15, gm_n50, in_13, gm_n6804, in_16);
	nor (gm_n6806, gm_n62, in_18, in_17, gm_n6805, gm_n45);
	nand (gm_n6807, gm_n6806, in_21);
	and (gm_n6808, in_11, in_10, gm_n51, gm_n997, gm_n48);
	nand (gm_n6809, gm_n63, gm_n50, in_13, gm_n6808, gm_n46);
	nor (gm_n6810, gm_n62, gm_n47, gm_n81, gm_n6809, gm_n45);
	nand (gm_n6811, gm_n6810, gm_n71);
	nand (gm_n6812, in_12, in_11, in_10, gm_n562, in_13);
	nor (gm_n6813, in_16, in_15, gm_n50, gm_n6812, in_17);
	nand (gm_n6814, in_20, in_19, in_18, gm_n6813, in_21);
	nand (gm_n6815, gm_n6807, gm_n6803, gm_n6799, gm_n6814, gm_n6811);
	nor (gm_n6816, gm_n6792, gm_n6788, gm_n6784, gm_n6815, gm_n6796);
	nand (gm_n6817, gm_n6776, gm_n6772, gm_n6767, gm_n6816, gm_n6780);
	nor (gm_n6818, gm_n6759, gm_n6756, gm_n6753, gm_n6817, gm_n6763);
	nand (gm_n6819, gm_n6745, gm_n6741, gm_n6738, gm_n6818, gm_n6749);
	nor (gm_n6820, gm_n6731, gm_n6728, gm_n6724, gm_n6819, gm_n6735);
	nand (gm_n6821, gm_n6717, gm_n6713, gm_n6709, gm_n6820, gm_n6721);
	nor (gm_n6822, gm_n6701, gm_n6699, gm_n6696, gm_n6821, gm_n6705);
	nand (gm_n6823, gm_n6689, gm_n6686, gm_n6682, gm_n6822, gm_n6692);
	nor (gm_n6824, gm_n6675, gm_n6671, gm_n6667, gm_n6823, gm_n6678);
	nand (gm_n6825, gm_n6660, gm_n6656, gm_n6653, gm_n6824, gm_n6663);
	nor (gm_n6826, gm_n6647, gm_n6642, gm_n6639, gm_n6825, gm_n6650);
	nand (gm_n6827, gm_n6633, gm_n6630, gm_n6627, gm_n6826, gm_n6636);
	nor (gm_n6828, gm_n6620, gm_n6616, gm_n6612, gm_n6827, gm_n6624);
	nand (gm_n6829, gm_n6604, gm_n6601, gm_n6598, gm_n6828, gm_n6608);
	nor (gm_n6830, gm_n6591, gm_n6589, gm_n6586, gm_n6829, gm_n6595);
	nand (gm_n6831, gm_n6579, gm_n6575, gm_n6571, gm_n6830, gm_n6582);
	nor (gm_n6832, gm_n6563, gm_n6559, gm_n6556, gm_n6831, gm_n6567);
	nand (gm_n6833, gm_n6548, gm_n6545, gm_n6542, gm_n6832, gm_n6553);
	nor (gm_n6834, gm_n6535, gm_n6531, gm_n6528, gm_n6833, gm_n6538);
	nand (gm_n6835, gm_n6521, gm_n6517, gm_n6513, gm_n6834, gm_n6524);
	nor (gm_n6836, gm_n6507, gm_n6504, gm_n6499, gm_n6835, gm_n6511);
	nand (gm_n6837, gm_n6493, gm_n6490, gm_n6486, gm_n6836, gm_n6495);
	nor (gm_n6838, gm_n6478, gm_n6474, gm_n6470, gm_n6837, gm_n6483);
	nand (gm_n6839, gm_n6463, gm_n6460, gm_n6457, gm_n6838, gm_n6466);
	nor (gm_n6840, gm_n6450, gm_n6447, gm_n6444, gm_n6839, gm_n6454);
	nand (gm_n6841, gm_n6438, gm_n6436, gm_n6433, gm_n6840, gm_n6441);
	nor (gm_n6842, gm_n6425, gm_n6421, gm_n6418, gm_n6841, gm_n6429);
	nand (gm_n6843, gm_n6412, gm_n6408, gm_n6404, gm_n6842, gm_n6415);
	nor (gm_n6844, gm_n6396, gm_n6393, gm_n6390, gm_n6843, gm_n6400);
	nand (gm_n6845, gm_n6384, gm_n6381, gm_n6377, gm_n6844, gm_n6387);
	nor (gm_n6846, gm_n6370, gm_n6368, gm_n6365, gm_n6845, gm_n6373);
	nand (gm_n6847, gm_n6358, gm_n6354, gm_n6351, gm_n6846, gm_n6361);
	nor (gm_n6848, gm_n6345, gm_n6341, gm_n6337, gm_n6847, gm_n6347);
	nand (gm_n6849, gm_n6330, gm_n6326, gm_n6323, gm_n6848, gm_n6334);
	nor (gm_n6850, gm_n6316, gm_n6312, gm_n6308, gm_n6849, gm_n6320);
	nand (gm_n6851, gm_n6300, gm_n6297, gm_n6293, gm_n6850, gm_n6304);
	nor (out_10, gm_n6851, gm_n6290);
	and (gm_n6853, gm_n2254, gm_n52, in_9);
	and (gm_n6854, in_13, gm_n48, gm_n53, gm_n6853, gm_n50);
	nand (gm_n6855, in_17, in_16, gm_n63, gm_n6854, in_18);
	nor (gm_n6856, gm_n71, gm_n45, gm_n62, gm_n6855);
	nor (gm_n6857, gm_n5252, in_9);
	nand (gm_n6858, gm_n48, in_11, in_10, gm_n6857, in_13);
	nor (gm_n6859, in_16, in_15, in_14, gm_n6858, in_17);
	nand (gm_n6860, gm_n45, gm_n62, gm_n47, gm_n6859, gm_n71);
	nor (gm_n6861, gm_n53, gm_n52, in_9, gm_n955, gm_n48);
	nand (gm_n6862, gm_n63, in_14, in_13, gm_n6861, in_16);
	nor (gm_n6863, gm_n62, in_18, in_17, gm_n6862, in_20);
	nand (gm_n6864, gm_n6863, in_21);
	nor (gm_n6865, gm_n53, in_10, gm_n51, gm_n1709, gm_n48);
	nand (gm_n6866, in_15, in_14, gm_n49, gm_n6865, gm_n46);
	nor (gm_n6867, in_19, in_18, in_17, gm_n6866, in_20);
	nand (gm_n6868, gm_n6867, gm_n71);
	nand (gm_n6869, in_12, in_11, in_10, gm_n4968, gm_n49);
	nor (gm_n6870, in_16, gm_n63, gm_n50, gm_n6869, in_17);
	nand (gm_n6871, in_20, in_19, gm_n47, gm_n6870, gm_n71);
	nand (gm_n6872, in_11, in_10, gm_n51, gm_n2034, gm_n48);
	nor (gm_n6873, gm_n63, in_14, in_13, gm_n6872, gm_n46);
	nand (gm_n6874, in_19, gm_n47, in_17, gm_n6873, gm_n45);
	nor (gm_n6875, gm_n6874, gm_n71);
	nand (gm_n6876, in_16, gm_n63, gm_n50, gm_n4307, gm_n81);
	nor (gm_n6877, in_20, in_19, in_18, gm_n6876, gm_n71);
	and (gm_n6878, in_12, gm_n53, gm_n52, gm_n6539, gm_n49);
	nand (gm_n6879, in_16, in_15, gm_n50, gm_n6878, gm_n81);
	nor (gm_n6880, in_20, in_19, gm_n47, gm_n6879, gm_n71);
	or (gm_n6881, in_16, gm_n63, in_14, gm_n2090, in_17);
	nor (gm_n6882, gm_n45, in_19, in_18, gm_n6881, in_21);
	nor (gm_n6883, gm_n5298, in_9);
	nand (gm_n6884, gm_n48, in_11, in_10, gm_n6883, gm_n49);
	nor (gm_n6885, in_16, in_15, in_14, gm_n6884, gm_n81);
	nand (gm_n6886, in_20, gm_n62, gm_n47, gm_n6885, in_21);
	nand (gm_n6887, in_12, gm_n53, in_10, gm_n3060, in_13);
	nor (gm_n6888, in_16, gm_n63, in_14, gm_n6887, gm_n81);
	nand (gm_n6889, gm_n45, gm_n62, in_18, gm_n6888, gm_n71);
	nor (gm_n6890, in_10, in_9, gm_n64, gm_n4079, in_11);
	nand (gm_n6891, gm_n50, gm_n49, in_12, gm_n6890, in_15);
	nor (gm_n6892, in_18, in_17, in_16, gm_n6891, in_19);
	nand (gm_n6893, gm_n6892, in_21, gm_n45);
	nand (gm_n6894, in_12, gm_n53, gm_n52, gm_n6742, gm_n49);
	nor (gm_n6895, in_16, gm_n63, gm_n50, gm_n6894, gm_n81);
	nand (gm_n6896, in_20, in_19, in_18, gm_n6895, in_21);
	nand (gm_n6897, gm_n64, in_7, in_6, gm_n638, gm_n51);
	nor (gm_n6898, in_12, in_11, gm_n52, gm_n6897, gm_n49);
	nand (gm_n6899, gm_n46, in_15, in_14, gm_n6898, in_17);
	nor (gm_n6900, in_20, in_19, in_18, gm_n6899, gm_n71);
	nand (gm_n6901, gm_n53, in_10, in_9, gm_n1874, in_12);
	nor (gm_n6902, in_15, gm_n50, in_13, gm_n6901, gm_n46);
	nand (gm_n6903, gm_n62, in_18, gm_n81, gm_n6902, in_20);
	nor (gm_n6904, gm_n6903, gm_n71);
	and (gm_n6905, gm_n1134, in_9);
	and (gm_n6906, in_12, gm_n53, gm_n52, gm_n6905, gm_n49);
	nand (gm_n6907, gm_n46, in_15, in_14, gm_n6906, in_17);
	nor (gm_n6908, in_20, in_19, in_18, gm_n6907, gm_n71);
	nand (gm_n6909, in_10, in_9, in_8, gm_n57, in_11);
	nor (gm_n6910, in_14, gm_n49, in_12, gm_n6909, gm_n63);
	nand (gm_n6911, gm_n47, in_17, gm_n46, gm_n6910, in_19);
	nor (gm_n6912, gm_n6911, gm_n71, in_20);
	nor (gm_n6913, gm_n52, gm_n51, gm_n64, gm_n907, gm_n53);
	nand (gm_n6914, gm_n50, gm_n49, gm_n48, gm_n6913, in_15);
	nor (gm_n6915, in_18, in_17, in_16, gm_n6914, gm_n62);
	nand (gm_n6916, gm_n6915, gm_n71, in_20);
	or (gm_n6917, in_11, gm_n52, gm_n51, gm_n686);
	or (gm_n6918, gm_n50, in_13, in_12, gm_n6917, in_15);
	nor (gm_n6919, gm_n47, gm_n81, gm_n46, gm_n6918, in_19);
	nand (gm_n6920, gm_n6919, gm_n71, in_20);
	or (gm_n6921, gm_n50, in_13, gm_n48, gm_n6221, gm_n63);
	nor (gm_n6922, in_18, gm_n81, in_16, gm_n6921, in_19);
	nand (gm_n6923, gm_n6922, gm_n71, in_20);
	and (gm_n6924, gm_n46, in_15, gm_n50, gm_n5306, in_17);
	nand (gm_n6925, in_20, gm_n62, gm_n47, gm_n6924, in_21);
	nand (gm_n6926, gm_n46, in_15, in_14, gm_n5078, in_17);
	nor (gm_n6927, in_20, in_19, in_18, gm_n6926, in_21);
	nor (gm_n6928, in_12, gm_n53, gm_n52, gm_n1280, gm_n49);
	nand (gm_n6929, in_16, gm_n63, in_14, gm_n6928, gm_n81);
	nor (gm_n6930, in_20, in_19, in_18, gm_n6929, gm_n71);
	and (gm_n6931, in_14, in_13, gm_n48, gm_n3547, gm_n63);
	nand (gm_n6932, in_18, gm_n81, in_16, gm_n6931, gm_n62);
	nor (gm_n6933, gm_n6932, gm_n71, gm_n45);
	and (gm_n6934, in_12, in_11, in_10, gm_n1719, in_13);
	nand (gm_n6935, in_16, gm_n63, gm_n50, gm_n6934, gm_n81);
	nor (gm_n6936, gm_n45, gm_n62, gm_n47, gm_n6935, gm_n71);
	or (gm_n6937, gm_n48, in_11, in_10, gm_n5268, in_13);
	nor (gm_n6938, gm_n46, gm_n63, in_14, gm_n6937, gm_n81);
	nand (gm_n6939, gm_n45, in_19, in_18, gm_n6938, in_21);
	nand (gm_n6940, in_12, gm_n53, in_10, gm_n3354, in_13);
	nor (gm_n6941, gm_n46, in_15, gm_n50, gm_n6940, in_17);
	nand (gm_n6942, in_20, in_19, gm_n47, gm_n6941, in_21);
	and (gm_n6943, in_11, in_10, in_9, gm_n2513);
	nand (gm_n6944, in_14, in_13, in_12, gm_n6943, in_15);
	nor (gm_n6945, gm_n47, in_17, in_16, gm_n6944, in_19);
	nand (gm_n6946, gm_n6945, in_21, gm_n45);
	nand (gm_n6947, gm_n48, gm_n53, gm_n52, gm_n2685, gm_n49);
	nor (gm_n6948, in_16, in_15, gm_n50, gm_n6947, gm_n81);
	nand (gm_n6949, gm_n45, gm_n62, in_18, gm_n6948, gm_n71);
	nor (gm_n6950, gm_n3884, in_10, in_9);
	and (gm_n6951, gm_n49, in_12, gm_n53, gm_n6950, in_14);
	nand (gm_n6952, gm_n81, gm_n46, gm_n63, gm_n6951, gm_n47);
	nor (gm_n6953, gm_n71, in_20, in_19, gm_n6952);
	nand (gm_n6954, in_11, gm_n52, in_9, gm_n4050, in_12);
	nor (gm_n6955, gm_n63, in_14, gm_n49, gm_n6954, in_16);
	nand (gm_n6956, in_19, in_18, in_17, gm_n6955, in_20);
	nor (gm_n6957, gm_n6956, in_21);
	nand (gm_n6958, gm_n48, gm_n53, in_10, gm_n1700, in_13);
	or (gm_n6959, gm_n46, in_15, gm_n50, gm_n6958, gm_n81);
	nor (gm_n6960, gm_n45, in_19, gm_n47, gm_n6959, gm_n71);
	nor (gm_n6961, gm_n53, gm_n52, in_9, gm_n1879);
	and (gm_n6962, in_14, in_13, gm_n48, gm_n6961, in_15);
	nand (gm_n6963, in_18, in_17, in_16, gm_n6962, gm_n62);
	nor (gm_n6964, gm_n6963, in_21, in_20);
	and (gm_n6965, gm_n53, gm_n52, gm_n51, gm_n1874, gm_n48);
	nand (gm_n6966, in_15, in_14, in_13, gm_n6965, gm_n46);
	nor (gm_n6967, in_19, gm_n47, in_17, gm_n6966, in_20);
	nand (gm_n6968, gm_n6967, in_21);
	or (gm_n6969, gm_n48, gm_n53, in_10, gm_n2327, in_13);
	nor (gm_n6970, in_16, in_15, in_14, gm_n6969, in_17);
	nand (gm_n6971, gm_n45, in_19, gm_n47, gm_n6970, in_21);
	nand (gm_n6972, in_14, gm_n49, in_12, gm_n4619, in_15);
	nor (gm_n6973, in_18, gm_n81, gm_n46, gm_n6972, in_19);
	nand (gm_n6974, gm_n6973, in_21, gm_n45);
	nor (gm_n6975, gm_n2275, gm_n52, in_9);
	nand (gm_n6976, in_13, gm_n48, gm_n53, gm_n6975, gm_n50);
	nor (gm_n6977, in_17, in_16, gm_n63, gm_n6976, gm_n47);
	nand (gm_n6978, in_21, gm_n45, in_19, gm_n6977);
	and (gm_n6979, in_15, gm_n50, gm_n49, gm_n3752, gm_n46);
	nand (gm_n6980, gm_n62, gm_n47, gm_n81, gm_n6979, in_20);
	nor (gm_n6981, gm_n6980, gm_n71);
	nor (gm_n6982, in_12, in_11, gm_n52, gm_n2597, gm_n49);
	nand (gm_n6983, in_16, in_15, in_14, gm_n6982, in_17);
	nor (gm_n6984, in_20, in_19, gm_n47, gm_n6983, gm_n71);
	nor (gm_n6985, in_12, in_11, in_10, gm_n3508, in_13);
	nand (gm_n6986, gm_n46, gm_n63, in_14, gm_n6985, in_17);
	nor (gm_n6987, in_20, gm_n62, gm_n47, gm_n6986, gm_n71);
	nand (gm_n6988, gm_n53, in_10, gm_n51, gm_n1222, gm_n48);
	nor (gm_n6989, gm_n63, gm_n50, gm_n49, gm_n6988, in_16);
	nand (gm_n6990, in_19, gm_n47, gm_n81, gm_n6989, gm_n45);
	nor (gm_n6991, gm_n6990, in_21);
	nor (gm_n6992, gm_n53, in_10, in_9, gm_n6155, gm_n48);
	nand (gm_n6993, in_15, gm_n50, in_13, gm_n6992, in_16);
	nor (gm_n6994, in_19, gm_n47, in_17, gm_n6993, in_20);
	nand (gm_n6995, gm_n6994, gm_n71);
	and (gm_n6996, gm_n53, in_10, gm_n51, gm_n4273, in_12);
	nand (gm_n6997, in_15, in_14, gm_n49, gm_n6996, in_16);
	nor (gm_n6998, in_19, gm_n47, gm_n81, gm_n6997, gm_n45);
	nand (gm_n6999, gm_n6998, in_21);
	nor (gm_n7000, gm_n53, in_10, gm_n51, gm_n2266, in_12);
	nand (gm_n7001, gm_n63, gm_n50, in_13, gm_n7000, gm_n46);
	nor (gm_n7002, in_19, gm_n47, gm_n81, gm_n7001, gm_n45);
	nand (gm_n7003, gm_n7002, gm_n71);
	nand (gm_n7004, in_13, gm_n48, gm_n53, gm_n2244, in_14);
	nor (gm_n7005, in_17, in_16, in_15, gm_n7004, in_18);
	nand (gm_n7006, gm_n71, in_20, gm_n62, gm_n7005);
	nand (gm_n7007, gm_n53, in_10, gm_n51, gm_n458, gm_n48);
	nor (gm_n7008, in_15, gm_n50, in_13, gm_n7007, in_16);
	nand (gm_n7009, in_19, in_18, gm_n81, gm_n7008, gm_n45);
	nor (gm_n7010, gm_n7009, in_21);
	nand (gm_n7011, in_11, in_10, gm_n51, gm_n3214, gm_n48);
	nor (gm_n7012, gm_n63, in_14, in_13, gm_n7011, gm_n46);
	nand (gm_n7013, gm_n62, in_18, gm_n81, gm_n7012, in_20);
	nor (gm_n7014, gm_n7013, gm_n71);
	or (gm_n7015, in_16, gm_n63, in_14, gm_n5987, gm_n81);
	nor (gm_n7016, in_20, gm_n62, in_18, gm_n7015, gm_n71);
	and (gm_n7017, in_12, in_11, in_10, gm_n589, gm_n49);
	nand (gm_n7018, gm_n46, gm_n63, in_14, gm_n7017, in_17);
	nor (gm_n7019, gm_n45, gm_n62, gm_n47, gm_n7018, gm_n71);
	nand (gm_n7020, gm_n63, gm_n50, in_13, gm_n3199, in_16);
	nor (gm_n7021, in_19, in_18, gm_n81, gm_n7020, in_20);
	nand (gm_n7022, gm_n7021, in_21);
	and (gm_n7023, gm_n1895, gm_n52, in_9);
	nand (gm_n7024, gm_n49, in_12, in_11, gm_n7023, gm_n50);
	nor (gm_n7025, gm_n81, in_16, gm_n63, gm_n7024, gm_n47);
	nand (gm_n7026, gm_n71, in_20, in_19, gm_n7025);
	nand (gm_n7027, gm_n48, gm_n53, in_10, gm_n1307, in_13);
	nor (gm_n7028, gm_n46, gm_n63, in_14, gm_n7027, in_17);
	nand (gm_n7029, in_20, in_19, in_18, gm_n7028, gm_n71);
	nand (gm_n7030, gm_n50, in_13, in_12, gm_n6355, in_15);
	nor (gm_n7031, gm_n47, gm_n81, in_16, gm_n7030, gm_n62);
	nand (gm_n7032, gm_n7031, gm_n71, gm_n45);
	nand (gm_n7033, in_11, gm_n52, gm_n51, gm_n4723, in_12);
	nor (gm_n7034, gm_n63, in_14, gm_n49, gm_n7033, in_16);
	nand (gm_n7035, in_19, in_18, gm_n81, gm_n7034, in_20);
	nor (gm_n7036, gm_n7035, gm_n71);
	nor (gm_n7037, gm_n48, in_11, in_10, gm_n4097, in_13);
	nand (gm_n7038, gm_n46, in_15, gm_n50, gm_n7037, gm_n81);
	nor (gm_n7039, in_20, gm_n62, gm_n47, gm_n7038, gm_n71);
	nand (gm_n7040, gm_n53, in_10, in_9, gm_n1279, in_12);
	nor (gm_n7041, in_15, gm_n50, gm_n49, gm_n7040, gm_n46);
	nand (gm_n7042, gm_n62, gm_n47, in_17, gm_n7041, in_20);
	nor (gm_n7043, gm_n7042, gm_n71);
	and (gm_n7044, in_11, in_10, in_9, gm_n3856, in_12);
	and (gm_n7045, gm_n63, in_14, in_13, gm_n7044, gm_n46);
	nand (gm_n7046, gm_n62, in_18, in_17, gm_n7045, gm_n45);
	nor (gm_n7047, gm_n7046, in_21);
	nor (gm_n7048, gm_n1735, gm_n51);
	nand (gm_n7049, gm_n48, gm_n53, gm_n52, gm_n7048, in_13);
	nor (gm_n7050, gm_n46, in_15, gm_n50, gm_n7049, gm_n81);
	nand (gm_n7051, in_20, in_19, gm_n47, gm_n7050, in_21);
	nand (gm_n7052, gm_n48, gm_n53, in_10, gm_n3553, gm_n49);
	nor (gm_n7053, gm_n46, gm_n63, gm_n50, gm_n7052, in_17);
	nand (gm_n7054, in_20, gm_n62, in_18, gm_n7053, gm_n71);
	nor (gm_n7055, gm_n55, in_6, in_5, gm_n643, gm_n64);
	and (gm_n7056, in_11, gm_n52, gm_n51, gm_n7055, in_12);
	nand (gm_n7057, gm_n63, gm_n50, gm_n49, gm_n7056, gm_n46);
	nor (gm_n7058, in_19, in_18, in_17, gm_n7057, in_20);
	nand (gm_n7059, gm_n7058, gm_n71);
	and (gm_n7060, in_11, gm_n52, gm_n51, gm_n484);
	nand (gm_n7061, in_14, gm_n49, gm_n48, gm_n7060, gm_n63);
	nor (gm_n7062, in_18, gm_n81, in_16, gm_n7061, in_19);
	nand (gm_n7063, gm_n7062, gm_n71, gm_n45);
	and (gm_n7064, in_11, gm_n52, in_9, gm_n4119, in_12);
	and (gm_n7065, gm_n63, gm_n50, in_13, gm_n7064, in_16);
	nand (gm_n7066, in_19, gm_n47, gm_n81, gm_n7065, in_20);
	nor (gm_n7067, gm_n7066, in_21);
	or (gm_n7068, in_8, in_7, in_6, gm_n119, gm_n51);
	nor (gm_n7069, in_12, gm_n53, in_10, gm_n7068, gm_n49);
	nand (gm_n7070, gm_n46, gm_n63, gm_n50, gm_n7069, in_17);
	nor (gm_n7071, gm_n45, in_19, gm_n47, gm_n7070, in_21);
	nand (gm_n7072, in_8, gm_n55, in_6, gm_n638, gm_n51);
	nor (gm_n7073, gm_n48, in_11, gm_n52, gm_n7072, in_13);
	nand (gm_n7074, gm_n46, in_15, in_14, gm_n7073, gm_n81);
	nor (gm_n7075, gm_n45, in_19, gm_n47, gm_n7074, in_21);
	nor (gm_n7076, gm_n48, in_11, in_10, gm_n4715, in_13);
	nand (gm_n7077, in_16, in_15, in_14, gm_n7076, in_17);
	nor (gm_n7078, in_20, gm_n62, gm_n47, gm_n7077, gm_n71);
	nand (gm_n7079, gm_n63, gm_n50, gm_n49, gm_n645, gm_n46);
	nor (gm_n7080, gm_n62, in_18, in_17, gm_n7079, in_20);
	nand (gm_n7081, gm_n7080, gm_n71);
	nand (gm_n7082, gm_n48, in_11, in_10, gm_n7048, gm_n49);
	nor (gm_n7083, in_16, in_15, in_14, gm_n7082, in_17);
	nand (gm_n7084, in_20, gm_n62, in_18, gm_n7083, gm_n71);
	nand (gm_n7085, gm_n63, in_14, gm_n49, gm_n5523);
	nor (gm_n7086, in_18, in_17, in_16, gm_n7085, gm_n62);
	nand (gm_n7087, gm_n7086, in_21, gm_n45);
	nor (gm_n7088, gm_n253, in_9);
	nand (gm_n7089, gm_n48, gm_n53, in_10, gm_n7088, gm_n49);
	nor (gm_n7090, gm_n46, in_15, gm_n50, gm_n7089, in_17);
	nand (gm_n7091, in_20, in_19, in_18, gm_n7090, in_21);
	nand (gm_n7092, gm_n51, in_8, gm_n55, gm_n136);
	nor (gm_n7093, gm_n48, in_11, gm_n52, gm_n7092, gm_n49);
	nand (gm_n7094, gm_n46, gm_n63, in_14, gm_n7093, gm_n81);
	nor (gm_n7095, gm_n45, in_19, in_18, gm_n7094, in_21);
	or (gm_n7096, gm_n5399, in_10, in_9);
	nor (gm_n7097, gm_n49, in_12, in_11, gm_n7096, gm_n50);
	nand (gm_n7098, gm_n81, in_16, in_15, gm_n7097, gm_n47);
	nor (gm_n7099, gm_n71, gm_n45, in_19, gm_n7098);
	nor (gm_n7100, gm_n48, gm_n53, in_10, gm_n6147, gm_n49);
	nand (gm_n7101, gm_n46, in_15, in_14, gm_n7100, gm_n81);
	nor (gm_n7102, gm_n45, in_19, gm_n47, gm_n7101, gm_n71);
	nor (gm_n7103, gm_n1481, in_10, gm_n51);
	and (gm_n7104, gm_n49, gm_n48, in_11, gm_n7103, in_14);
	nand (gm_n7105, gm_n81, in_16, in_15, gm_n7104, in_18);
	nor (gm_n7106, gm_n71, gm_n45, in_19, gm_n7105);
	and (gm_n7107, in_11, in_10, in_9, gm_n189);
	nand (gm_n7108, in_14, in_13, in_12, gm_n7107, gm_n63);
	nor (gm_n7109, gm_n47, in_17, gm_n46, gm_n7108, gm_n62);
	nand (gm_n7110, gm_n7109, gm_n71, in_20);
	and (gm_n7111, in_11, in_10, gm_n51, gm_n1339);
	nand (gm_n7112, gm_n50, gm_n49, gm_n48, gm_n7111, in_15);
	nor (gm_n7113, gm_n47, gm_n81, in_16, gm_n7112, in_19);
	nand (gm_n7114, gm_n7113, in_21, in_20);
	nor (gm_n7115, in_8, gm_n55, in_6, gm_n530, in_9);
	nand (gm_n7116, gm_n48, gm_n53, in_10, gm_n7115, gm_n49);
	nor (gm_n7117, in_16, in_15, gm_n50, gm_n7116, gm_n81);
	nand (gm_n7118, gm_n45, gm_n62, gm_n47, gm_n7117, in_21);
	nand (gm_n7119, in_12, in_11, gm_n52, gm_n5822, in_13);
	nor (gm_n7120, in_16, gm_n63, gm_n50, gm_n7119, in_17);
	nand (gm_n7121, in_20, in_19, gm_n47, gm_n7120, gm_n71);
	nand (gm_n7122, gm_n52, gm_n51, in_8, gm_n838, in_11);
	nor (gm_n7123, in_14, in_13, gm_n48, gm_n7122, gm_n63);
	nand (gm_n7124, gm_n47, in_17, in_16, gm_n7123, gm_n62);
	nor (gm_n7125, gm_n7124, in_21, gm_n45);
	nand (gm_n7126, in_11, in_10, gm_n51, gm_n2181, gm_n48);
	nor (gm_n7127, in_15, gm_n50, gm_n49, gm_n7126, gm_n46);
	nand (gm_n7128, in_19, gm_n47, gm_n81, gm_n7127, in_20);
	nor (gm_n7129, gm_n7128, gm_n71);
	nand (gm_n7130, gm_n53, gm_n52, gm_n51, gm_n2047, gm_n48);
	nor (gm_n7131, gm_n63, gm_n50, in_13, gm_n7130, gm_n46);
	nand (gm_n7132, gm_n62, gm_n47, in_17, gm_n7131, in_20);
	nor (gm_n7133, gm_n7132, in_21);
	and (gm_n7134, gm_n1603, in_9);
	and (gm_n7135, gm_n48, in_11, gm_n52, gm_n7134, gm_n49);
	nand (gm_n7136, gm_n46, in_15, gm_n50, gm_n7135, gm_n81);
	nor (gm_n7137, gm_n45, gm_n62, in_18, gm_n7136, gm_n71);
	and (gm_n7138, in_11, gm_n52, gm_n51, gm_n612, in_12);
	nand (gm_n7139, in_15, in_14, gm_n49, gm_n7138, in_16);
	nor (gm_n7140, in_19, in_18, gm_n81, gm_n7139, gm_n45);
	nand (gm_n7141, gm_n7140, gm_n71);
	nand (gm_n7142, in_13, in_12, gm_n53, gm_n3528, gm_n50);
	nor (gm_n7143, in_17, in_16, gm_n63, gm_n7142, in_18);
	nand (gm_n7144, in_21, gm_n45, gm_n62, gm_n7143);
	nand (gm_n7145, gm_n48, in_11, gm_n52, gm_n968, gm_n49);
	nor (gm_n7146, in_16, gm_n63, in_14, gm_n7145, gm_n81);
	nand (gm_n7147, gm_n45, gm_n62, gm_n47, gm_n7146, gm_n71);
	nor (gm_n7148, in_16, gm_n63, in_14, gm_n5810, in_17);
	nand (gm_n7149, in_20, gm_n62, in_18, gm_n7148, in_21);
	or (gm_n7150, in_11, gm_n52, gm_n51, gm_n3542, gm_n48);
	nor (gm_n7151, in_15, gm_n50, in_13, gm_n7150, in_16);
	nand (gm_n7152, in_19, in_18, gm_n81, gm_n7151, in_20);
	nor (gm_n7153, gm_n7152, gm_n71);
	or (gm_n7154, in_8, gm_n55, in_6, gm_n103, in_9);
	nor (gm_n7155, in_12, gm_n53, gm_n52, gm_n7154, gm_n49);
	nand (gm_n7156, gm_n46, gm_n63, gm_n50, gm_n7155, gm_n81);
	nor (gm_n7157, gm_n45, gm_n62, in_18, gm_n7156, in_21);
	and (gm_n7158, gm_n49, gm_n48, gm_n53, gm_n4741, in_14);
	nand (gm_n7159, in_17, in_16, gm_n63, gm_n7158, gm_n47);
	nor (gm_n7160, gm_n71, gm_n45, gm_n62, gm_n7159);
	and (gm_n7161, gm_n49, in_12, gm_n53, gm_n5834, gm_n50);
	nand (gm_n7162, gm_n81, gm_n46, in_15, gm_n7161, gm_n47);
	nor (gm_n7163, in_21, gm_n45, in_19, gm_n7162);
	nand (gm_n7164, gm_n48, in_11, gm_n52, gm_n696, gm_n49);
	nor (gm_n7165, gm_n46, in_15, gm_n50, gm_n7164, gm_n81);
	nand (gm_n7166, gm_n45, gm_n62, in_18, gm_n7165, gm_n71);
	nand (gm_n7167, gm_n49, gm_n48, in_11, gm_n5669, gm_n50);
	nor (gm_n7168, gm_n81, in_16, gm_n63, gm_n7167, gm_n47);
	nand (gm_n7169, gm_n71, gm_n45, in_19, gm_n7168);
	nor (gm_n7170, in_16, in_15, gm_n50, gm_n6606, in_17);
	nand (gm_n7171, in_20, in_19, gm_n47, gm_n7170, in_21);
	nor (gm_n7172, gm_n3475, gm_n51);
	nand (gm_n7173, gm_n48, gm_n53, gm_n52, gm_n7172, in_13);
	nor (gm_n7174, gm_n46, in_15, in_14, gm_n7173, gm_n81);
	nand (gm_n7175, gm_n45, in_19, in_18, gm_n7174, gm_n71);
	and (gm_n7176, in_9, in_8, gm_n55, gm_n504);
	and (gm_n7177, gm_n48, gm_n53, in_10, gm_n7176, in_13);
	nand (gm_n7178, in_16, gm_n63, in_14, gm_n7177, in_17);
	nor (gm_n7179, in_20, in_19, in_18, gm_n7178, in_21);
	nand (gm_n7180, gm_n46, in_15, in_14, gm_n6230, in_17);
	nor (gm_n7181, gm_n45, gm_n62, gm_n47, gm_n7180, in_21);
	nand (gm_n7182, gm_n53, in_10, gm_n51, gm_n2472, gm_n48);
	nor (gm_n7183, in_15, gm_n50, gm_n49, gm_n7182, gm_n46);
	nand (gm_n7184, gm_n62, in_18, in_17, gm_n7183, gm_n45);
	nor (gm_n7185, gm_n7184, gm_n71);
	nor (gm_n7186, gm_n64, gm_n55, gm_n82, gm_n204, gm_n51);
	and (gm_n7187, gm_n48, gm_n53, in_10, gm_n7186, in_13);
	nand (gm_n7188, in_16, gm_n63, gm_n50, gm_n7187, gm_n81);
	nor (gm_n7189, gm_n45, in_19, gm_n47, gm_n7188, in_21);
	nand (gm_n7190, gm_n48, in_11, gm_n52, gm_n7088, in_13);
	nor (gm_n7191, gm_n46, in_15, in_14, gm_n7190, in_17);
	nand (gm_n7192, in_20, gm_n62, gm_n47, gm_n7191, gm_n71);
	nor (gm_n7193, gm_n1533, in_10, in_9);
	nand (gm_n7194, gm_n49, in_12, gm_n53, gm_n7193, gm_n50);
	nor (gm_n7195, in_17, gm_n46, in_15, gm_n7194, in_18);
	nand (gm_n7196, gm_n71, in_20, gm_n62, gm_n7195);
	nand (gm_n7197, gm_n48, in_11, gm_n52, gm_n6525, in_13);
	nor (gm_n7198, in_16, in_15, in_14, gm_n7197, in_17);
	nand (gm_n7199, gm_n45, in_19, in_18, gm_n7198, gm_n71);
	nand (gm_n7200, in_12, gm_n53, gm_n52, gm_n146, gm_n49);
	nor (gm_n7201, gm_n46, gm_n63, in_14, gm_n7200, gm_n81);
	nand (gm_n7202, gm_n45, gm_n62, gm_n47, gm_n7201, gm_n71);
	and (gm_n7203, gm_n48, in_11, in_10, gm_n3909, gm_n49);
	nand (gm_n7204, gm_n46, in_15, in_14, gm_n7203, in_17);
	nor (gm_n7205, gm_n45, in_19, gm_n47, gm_n7204, in_21);
	nand (gm_n7206, gm_n1293, in_10, gm_n51);
	nor (gm_n7207, gm_n49, gm_n48, in_11, gm_n7206, gm_n50);
	nand (gm_n7208, gm_n81, gm_n46, in_15, gm_n7207, gm_n47);
	nor (gm_n7209, gm_n71, in_20, in_19, gm_n7208);
	nand (gm_n7210, gm_n53, in_10, gm_n51, gm_n76, in_12);
	nor (gm_n7211, in_15, gm_n50, gm_n49, gm_n7210, gm_n46);
	nand (gm_n7212, in_19, gm_n47, gm_n81, gm_n7211, gm_n45);
	nor (gm_n7213, gm_n7212, in_21);
	nor (gm_n7214, in_21, gm_n45, gm_n62, gm_n424);
	nand (gm_n7215, in_15, gm_n50, gm_n49, gm_n4065, gm_n46);
	nor (gm_n7216, in_19, gm_n47, gm_n81, gm_n7215, gm_n45);
	nand (gm_n7217, gm_n7216, gm_n71);
	nand (gm_n7218, gm_n49, gm_n48, gm_n53, gm_n539, gm_n50);
	nor (gm_n7219, gm_n81, gm_n46, gm_n63, gm_n7218, gm_n47);
	nand (gm_n7220, in_21, in_20, gm_n62, gm_n7219);
	nand (gm_n7221, gm_n48, gm_n53, gm_n52, gm_n4127, in_13);
	nor (gm_n7222, in_16, gm_n63, gm_n50, gm_n7221, in_17);
	nand (gm_n7223, gm_n45, gm_n62, in_18, gm_n7222, in_21);
	and (gm_n7224, in_13, in_12, in_11, gm_n2218);
	and (gm_n7225, gm_n46, gm_n63, in_14, gm_n7224, gm_n81);
	nand (gm_n7226, gm_n45, in_19, gm_n47, gm_n7225, in_21);
	or (gm_n7227, gm_n64, gm_n55, gm_n82, gm_n204, in_9);
	nor (gm_n7228, in_12, gm_n53, gm_n52, gm_n7227, gm_n49);
	nand (gm_n7229, gm_n46, gm_n63, in_14, gm_n7228, in_17);
	nor (gm_n7230, gm_n45, in_19, in_18, gm_n7229, gm_n71);
	and (gm_n7231, gm_n2014, gm_n51);
	and (gm_n7232, in_12, in_11, gm_n52, gm_n7231, gm_n49);
	nand (gm_n7233, gm_n46, in_15, in_14, gm_n7232, in_17);
	nor (gm_n7234, in_20, in_19, gm_n47, gm_n7233, gm_n71);
	or (gm_n7235, in_8, in_7, gm_n82, gm_n141, gm_n51);
	nor (gm_n7236, in_12, in_11, in_10, gm_n7235, gm_n49);
	nand (gm_n7237, gm_n46, gm_n63, gm_n50, gm_n7236, gm_n81);
	nor (gm_n7238, gm_n45, in_19, in_18, gm_n7237, gm_n71);
	nand (gm_n7239, in_11, gm_n52, gm_n51, gm_n210, gm_n48);
	nor (gm_n7240, gm_n63, in_14, gm_n49, gm_n7239, in_16);
	nand (gm_n7241, gm_n62, gm_n47, gm_n81, gm_n7240, in_20);
	nor (gm_n7242, gm_n7241, in_21);
	nand (gm_n7243, gm_n49, in_12, gm_n53, gm_n743, in_14);
	nor (gm_n7244, in_17, gm_n46, gm_n63, gm_n7243, in_18);
	nand (gm_n7245, in_21, in_20, gm_n62, gm_n7244);
	and (gm_n7246, gm_n53, gm_n52, gm_n51, gm_n3519);
	nand (gm_n7247, gm_n50, gm_n49, gm_n48, gm_n7246, in_15);
	nor (gm_n7248, gm_n47, gm_n81, in_16, gm_n7247, gm_n62);
	nand (gm_n7249, gm_n7248, in_21, in_20);
	nor (gm_n7250, gm_n51, gm_n64, gm_n55, gm_n588, gm_n52);
	nand (gm_n7251, gm_n49, gm_n48, gm_n53, gm_n7250, gm_n50);
	nor (gm_n7252, in_17, gm_n46, in_15, gm_n7251, gm_n47);
	nand (gm_n7253, in_21, gm_n45, gm_n62, gm_n7252);
	nand (gm_n7254, in_12, in_11, in_10, gm_n5676, gm_n49);
	nor (gm_n7255, in_16, gm_n63, gm_n50, gm_n7254, gm_n81);
	nand (gm_n7256, gm_n45, gm_n62, in_18, gm_n7255, in_21);
	and (gm_n7257, gm_n48, in_11, in_10, gm_n4984, in_13);
	nand (gm_n7258, gm_n46, in_15, gm_n50, gm_n7257, gm_n81);
	nor (gm_n7259, in_20, gm_n62, in_18, gm_n7258, gm_n71);
	nor (gm_n7260, in_12, in_11, in_10, gm_n5620, gm_n49);
	nand (gm_n7261, gm_n46, in_15, in_14, gm_n7260, gm_n81);
	nor (gm_n7262, in_20, gm_n62, in_18, gm_n7261, gm_n71);
	nand (gm_n7263, in_11, gm_n52, gm_n51, gm_n3086, in_12);
	nor (gm_n7264, gm_n63, in_14, gm_n49, gm_n7263, in_16);
	nand (gm_n7265, gm_n62, in_18, in_17, gm_n7264, gm_n45);
	nor (gm_n7266, gm_n7265, in_21);
	and (gm_n7267, in_13, in_12, in_11, gm_n1542, in_14);
	nand (gm_n7268, in_17, in_16, in_15, gm_n7267, gm_n47);
	nor (gm_n7269, in_21, gm_n45, gm_n62, gm_n7268);
	nor (gm_n7270, in_10, gm_n51, in_8, gm_n5379, in_11);
	nand (gm_n7271, gm_n50, in_13, gm_n48, gm_n7270, gm_n63);
	nor (gm_n7272, gm_n47, in_17, in_16, gm_n7271, gm_n62);
	nand (gm_n7273, gm_n7272, gm_n71, in_20);
	nand (gm_n7274, gm_n48, gm_n53, in_10, gm_n1201, in_13);
	nor (gm_n7275, in_16, in_15, gm_n50, gm_n7274, gm_n81);
	nand (gm_n7276, in_20, gm_n62, gm_n47, gm_n7275, gm_n71);
	nand (gm_n7277, gm_n48, gm_n53, in_10, gm_n2819, gm_n49);
	nor (gm_n7278, gm_n46, gm_n63, in_14, gm_n7277, gm_n81);
	nand (gm_n7279, in_20, gm_n62, gm_n47, gm_n7278, in_21);
	nand (gm_n7280, in_12, in_11, gm_n52, gm_n1941, gm_n49);
	nor (gm_n7281, gm_n46, gm_n63, in_14, gm_n7280, in_17);
	nand (gm_n7282, in_20, in_19, gm_n47, gm_n7281, in_21);
	nor (gm_n7283, gm_n48, gm_n53, gm_n52, gm_n4381, in_13);
	nand (gm_n7284, gm_n46, gm_n63, in_14, gm_n7283, in_17);
	nor (gm_n7285, in_20, in_19, gm_n47, gm_n7284, in_21);
	nor (gm_n7286, gm_n48, gm_n53, in_10, gm_n1723, gm_n49);
	nand (gm_n7287, gm_n46, gm_n63, gm_n50, gm_n7286, in_17);
	nor (gm_n7288, in_20, in_19, in_18, gm_n7287, in_21);
	nor (gm_n7289, in_12, in_11, gm_n52, gm_n4696, in_13);
	nand (gm_n7290, gm_n46, gm_n63, in_14, gm_n7289, gm_n81);
	nor (gm_n7291, in_20, in_19, in_18, gm_n7290, in_21);
	nand (gm_n7292, in_11, gm_n52, in_9, gm_n2432, gm_n48);
	nor (gm_n7293, in_15, in_14, in_13, gm_n7292, in_16);
	nand (gm_n7294, in_19, gm_n47, in_17, gm_n7293, gm_n45);
	nor (gm_n7295, gm_n7294, gm_n71);
	nand (gm_n7296, in_13, gm_n48, in_11, gm_n844, in_14);
	nor (gm_n7297, gm_n81, in_16, gm_n63, gm_n7296, gm_n47);
	nand (gm_n7298, gm_n71, in_20, gm_n62, gm_n7297);
	nand (gm_n7299, gm_n49, in_12, gm_n53, gm_n2214, in_14);
	nor (gm_n7300, gm_n81, in_16, in_15, gm_n7299, in_18);
	nand (gm_n7301, in_21, in_20, gm_n62, gm_n7300);
	nand (gm_n7302, in_15, gm_n50, gm_n49, gm_n5410, gm_n46);
	nor (gm_n7303, in_19, gm_n47, gm_n81, gm_n7302, in_20);
	nand (gm_n7304, gm_n7303, in_21);
	nor (gm_n7305, gm_n514, in_9);
	nand (gm_n7306, in_12, gm_n53, gm_n52, gm_n7305, in_13);
	nor (gm_n7307, gm_n46, gm_n63, in_14, gm_n7306, gm_n81);
	nand (gm_n7308, in_20, in_19, in_18, gm_n7307, gm_n71);
	nand (gm_n7309, in_11, in_10, in_9, gm_n1142);
	nor (gm_n7310, in_14, gm_n49, gm_n48, gm_n7309, in_15);
	nand (gm_n7311, in_18, in_17, gm_n46, gm_n7310, in_19);
	nor (gm_n7312, gm_n7311, gm_n71, in_20);
	nor (gm_n7313, gm_n49, in_12, in_11, gm_n1031, in_14);
	nand (gm_n7314, gm_n81, in_16, gm_n63, gm_n7313, in_18);
	nor (gm_n7315, gm_n71, in_20, gm_n62, gm_n7314);
	nor (gm_n7316, gm_n63, gm_n50, in_13, gm_n4929, gm_n46);
	nand (gm_n7317, in_19, in_18, in_17, gm_n7316, gm_n45);
	nor (gm_n7318, gm_n7317, gm_n71);
	nand (gm_n7319, gm_n51, gm_n64, gm_n55, gm_n136, gm_n52);
	nor (gm_n7320, in_13, in_12, gm_n53, gm_n7319, gm_n50);
	nand (gm_n7321, gm_n81, gm_n46, in_15, gm_n7320, gm_n47);
	nor (gm_n7322, gm_n71, in_20, in_19, gm_n7321);
	nand (gm_n7323, in_14, in_13, gm_n48, gm_n5917, gm_n63);
	nor (gm_n7324, gm_n47, in_17, in_16, gm_n7323, gm_n62);
	nand (gm_n7325, gm_n7324, gm_n71, gm_n45);
	nor (gm_n7326, gm_n53, in_10, gm_n51, gm_n183, gm_n48);
	nand (gm_n7327, gm_n63, gm_n50, in_13, gm_n7326, gm_n46);
	nor (gm_n7328, in_19, gm_n47, in_17, gm_n7327, in_20);
	nand (gm_n7329, gm_n7328, gm_n71);
	or (gm_n7330, gm_n45, gm_n62, in_18, gm_n3766, in_21);
	nand (gm_n7331, gm_n50, gm_n49, gm_n48, gm_n5502, in_15);
	nor (gm_n7332, gm_n47, in_17, gm_n46, gm_n7331, in_19);
	nand (gm_n7333, gm_n7332, in_21, in_20);
	nand (gm_n7334, gm_n53, gm_n52, gm_n51, gm_n3904, in_12);
	nor (gm_n7335, in_15, in_14, in_13, gm_n7334, gm_n46);
	nand (gm_n7336, in_19, gm_n47, in_17, gm_n7335, gm_n45);
	nor (gm_n7337, gm_n7336, in_21);
	nor (gm_n7338, gm_n50, in_13, gm_n48, gm_n5418, in_15);
	nand (gm_n7339, in_18, gm_n81, gm_n46, gm_n7338, gm_n62);
	nor (gm_n7340, gm_n7339, in_21, in_20);
	nor (gm_n7341, gm_n49, gm_n48, in_11, gm_n169, gm_n50);
	nand (gm_n7342, in_17, gm_n46, gm_n63, gm_n7341, gm_n47);
	nor (gm_n7343, in_21, in_20, gm_n62, gm_n7342);
	nor (gm_n7344, gm_n48, in_11, in_10, gm_n1398, in_13);
	nand (gm_n7345, in_16, in_15, gm_n50, gm_n7344, gm_n81);
	nor (gm_n7346, in_20, in_19, gm_n47, gm_n7345, gm_n71);
	nand (gm_n7347, in_12, gm_n53, in_10, gm_n4127, gm_n49);
	nor (gm_n7348, in_16, in_15, in_14, gm_n7347, in_17);
	nand (gm_n7349, gm_n45, in_19, gm_n47, gm_n7348, gm_n71);
	nor (gm_n7350, in_17, in_16, in_15, gm_n5473, in_18);
	nand (gm_n7351, in_21, gm_n45, in_19, gm_n7350);
	nand (gm_n7352, gm_n48, gm_n53, gm_n52, gm_n6583, in_13);
	nor (gm_n7353, gm_n46, gm_n63, gm_n50, gm_n7352, in_17);
	nand (gm_n7354, in_20, in_19, in_18, gm_n7353, in_21);
	nand (gm_n7355, in_12, gm_n53, in_10, gm_n3909, in_13);
	nor (gm_n7356, gm_n46, gm_n63, gm_n50, gm_n7355, in_17);
	nand (gm_n7357, in_20, in_19, in_18, gm_n7356, in_21);
	nor (gm_n7358, in_11, gm_n52, gm_n51, gm_n738);
	nand (gm_n7359, gm_n50, in_13, in_12, gm_n7358, in_15);
	nor (gm_n7360, in_18, in_17, in_16, gm_n7359, gm_n62);
	nand (gm_n7361, gm_n7360, gm_n71, in_20);
	nand (gm_n7362, gm_n7354, gm_n7351, gm_n7349, gm_n7361, gm_n7357);
	nor (gm_n7363, gm_n7343, gm_n7340, gm_n7337, gm_n7362, gm_n7346);
	nand (gm_n7364, gm_n7330, gm_n7329, gm_n7325, gm_n7363, gm_n7333);
	nor (gm_n7365, gm_n7318, gm_n7315, gm_n7312, gm_n7364, gm_n7322);
	nand (gm_n7366, gm_n7304, gm_n7301, gm_n7298, gm_n7365, gm_n7308);
	nor (gm_n7367, gm_n7291, gm_n7288, gm_n7285, gm_n7366, gm_n7295);
	nand (gm_n7368, gm_n7279, gm_n7276, gm_n7273, gm_n7367, gm_n7282);
	nor (gm_n7369, gm_n7266, gm_n7262, gm_n7259, gm_n7368, gm_n7269);
	nand (gm_n7370, gm_n7253, gm_n7249, gm_n7245, gm_n7369, gm_n7256);
	nor (gm_n7371, gm_n7238, gm_n7234, gm_n7230, gm_n7370, gm_n7242);
	nand (gm_n7372, gm_n7223, gm_n7220, gm_n7217, gm_n7371, gm_n7226);
	nor (gm_n7373, gm_n7213, gm_n7209, gm_n7205, gm_n7372, gm_n7214);
	nand (gm_n7374, gm_n7199, gm_n7196, gm_n7192, gm_n7373, gm_n7202);
	nor (gm_n7375, gm_n7185, gm_n7181, gm_n7179, gm_n7374, gm_n7189);
	nand (gm_n7376, gm_n7171, gm_n7169, gm_n7166, gm_n7375, gm_n7175);
	nor (gm_n7377, gm_n7160, gm_n7157, gm_n7153, gm_n7376, gm_n7163);
	nand (gm_n7378, gm_n7147, gm_n7144, gm_n7141, gm_n7377, gm_n7149);
	nor (gm_n7379, gm_n7133, gm_n7129, gm_n7125, gm_n7378, gm_n7137);
	nand (gm_n7380, gm_n7118, gm_n7114, gm_n7110, gm_n7379, gm_n7121);
	nor (gm_n7381, gm_n7102, gm_n7099, gm_n7095, gm_n7380, gm_n7106);
	nand (gm_n7382, gm_n7087, gm_n7084, gm_n7081, gm_n7381, gm_n7091);
	nor (gm_n7383, gm_n7075, gm_n7071, gm_n7067, gm_n7382, gm_n7078);
	nand (gm_n7384, gm_n7059, gm_n7054, gm_n7051, gm_n7383, gm_n7063);
	nor (gm_n7385, gm_n7043, gm_n7039, gm_n7036, gm_n7384, gm_n7047);
	nand (gm_n7386, gm_n7029, gm_n7026, gm_n7022, gm_n7385, gm_n7032);
	nor (gm_n7387, gm_n7016, gm_n7014, gm_n7010, gm_n7386, gm_n7019);
	nand (gm_n7388, gm_n7003, gm_n6999, gm_n6995, gm_n7387, gm_n7006);
	nor (gm_n7389, gm_n6987, gm_n6984, gm_n6981, gm_n7388, gm_n6991);
	nand (gm_n7390, gm_n6974, gm_n6971, gm_n6968, gm_n7389, gm_n6978);
	nor (gm_n7391, gm_n6960, gm_n6957, gm_n6953, gm_n7390, gm_n6964);
	nand (gm_n7392, gm_n6946, gm_n6942, gm_n6939, gm_n7391, gm_n6949);
	nor (gm_n7393, gm_n6933, gm_n6930, gm_n6927, gm_n7392, gm_n6936);
	nand (gm_n7394, gm_n6923, gm_n6920, gm_n6916, gm_n7393, gm_n6925);
	nor (gm_n7395, gm_n6908, gm_n6904, gm_n6900, gm_n7394, gm_n6912);
	nand (gm_n7396, gm_n6893, gm_n6889, gm_n6886, gm_n7395, gm_n6896);
	nor (gm_n7397, gm_n6880, gm_n6877, gm_n6875, gm_n7396, gm_n6882);
	nand (gm_n7398, gm_n6868, gm_n6864, gm_n6860, gm_n7397, gm_n6871);
	nor (out_11, gm_n7398, gm_n6856);
	nand (gm_n7400, in_9, in_8, gm_n55, gm_n136);
	nor (gm_n7401, gm_n48, in_11, in_10, gm_n7400, gm_n49);
	nand (gm_n7402, gm_n46, in_15, in_14, gm_n7401, gm_n81);
	nor (gm_n7403, gm_n45, gm_n62, in_18, gm_n7402, in_21);
	nand (gm_n7404, gm_n48, in_11, gm_n52, gm_n1975, gm_n49);
	nor (gm_n7405, gm_n46, gm_n63, gm_n50, gm_n7404, gm_n81);
	nand (gm_n7406, gm_n45, in_19, gm_n47, gm_n7405, gm_n71);
	nand (gm_n7407, in_13, in_12, gm_n53, gm_n5562, in_14);
	nor (gm_n7408, in_17, in_16, in_15, gm_n7407, in_18);
	nand (gm_n7409, in_21, gm_n45, gm_n62, gm_n7408);
	nand (gm_n7410, in_12, gm_n53, in_10, gm_n617, gm_n49);
	nor (gm_n7411, gm_n46, in_15, in_14, gm_n7410, in_17);
	nand (gm_n7412, in_20, in_19, gm_n47, gm_n7411, in_21);
	nand (gm_n7413, in_14, gm_n49, gm_n48, gm_n5279, gm_n63);
	nor (gm_n7414, in_18, in_17, in_16, gm_n7413, in_19);
	nand (gm_n7415, gm_n7414, gm_n71, in_20);
	nand (gm_n7416, in_16, gm_n63, gm_n50, gm_n2007, in_17);
	nor (gm_n7417, gm_n45, in_19, in_18, gm_n7416, gm_n71);
	or (gm_n7418, in_11, gm_n52, gm_n51, gm_n1481, in_12);
	nor (gm_n7419, gm_n63, gm_n50, in_13, gm_n7418, in_16);
	nand (gm_n7420, in_19, gm_n47, gm_n81, gm_n7419, gm_n45);
	nor (gm_n7421, gm_n7420, in_21);
	nor (gm_n7422, in_12, gm_n53, in_10, gm_n2743, gm_n49);
	nand (gm_n7423, gm_n46, in_15, gm_n50, gm_n7422, gm_n81);
	nor (gm_n7424, gm_n45, in_19, gm_n47, gm_n7423, in_21);
	nor (gm_n7425, gm_n686, in_10, gm_n51);
	and (gm_n7426, gm_n49, in_12, gm_n53, gm_n7425, in_14);
	nand (gm_n7427, in_17, gm_n46, gm_n63, gm_n7426, in_18);
	nor (gm_n7428, gm_n71, in_20, in_19, gm_n7427);
	nand (gm_n7429, in_12, gm_n53, in_10, gm_n2760, in_13);
	nor (gm_n7430, in_16, gm_n63, gm_n50, gm_n7429, in_17);
	nand (gm_n7431, gm_n45, in_19, in_18, gm_n7430, in_21);
	nand (gm_n7432, in_13, in_12, in_11, gm_n5451, gm_n50);
	nor (gm_n7433, in_17, in_16, in_15, gm_n7432, in_18);
	nand (gm_n7434, in_21, gm_n45, gm_n62, gm_n7433);
	nor (gm_n7435, gm_n46, gm_n63, in_14, gm_n4912, in_17);
	nand (gm_n7436, gm_n45, gm_n62, in_18, gm_n7435, gm_n71);
	nand (gm_n7437, in_12, in_11, in_10, gm_n1982, gm_n49);
	nor (gm_n7438, gm_n46, gm_n63, in_14, gm_n7437, in_17);
	nand (gm_n7439, in_20, gm_n62, gm_n47, gm_n7438, in_21);
	nor (gm_n7440, in_12, in_11, gm_n52, gm_n6032, in_13);
	nand (gm_n7441, gm_n46, gm_n63, gm_n50, gm_n7440, gm_n81);
	nor (gm_n7442, gm_n45, gm_n62, in_18, gm_n7441, in_21);
	nor (gm_n7443, gm_n48, gm_n53, in_10, gm_n1824, in_13);
	nand (gm_n7444, gm_n46, gm_n63, in_14, gm_n7443, gm_n81);
	nor (gm_n7445, gm_n45, gm_n62, gm_n47, gm_n7444, in_21);
	and (gm_n7446, gm_n48, gm_n53, in_10, gm_n3562, in_13);
	nand (gm_n7447, gm_n46, gm_n63, in_14, gm_n7446, gm_n81);
	nor (gm_n7448, gm_n45, gm_n62, gm_n47, gm_n7447, in_21);
	nand (gm_n7449, gm_n46, in_15, in_14, gm_n2572, in_17);
	nor (gm_n7450, in_20, gm_n62, gm_n47, gm_n7449, in_21);
	and (gm_n7451, gm_n46, in_15, gm_n50, gm_n4316, in_17);
	nand (gm_n7452, gm_n45, gm_n62, gm_n47, gm_n7451, gm_n71);
	nand (gm_n7453, in_14, gm_n49, gm_n48, gm_n5776, in_15);
	nor (gm_n7454, gm_n47, in_17, in_16, gm_n7453, gm_n62);
	nand (gm_n7455, gm_n7454, in_21, in_20);
	nand (gm_n7456, gm_n48, gm_n53, in_10, gm_n1808, in_13);
	nor (gm_n7457, gm_n46, gm_n63, in_14, gm_n7456, gm_n81);
	nand (gm_n7458, in_20, in_19, in_18, gm_n7457, in_21);
	nor (gm_n7459, gm_n53, gm_n52, in_9, gm_n2266);
	nand (gm_n7460, in_14, gm_n49, in_12, gm_n7459, gm_n63);
	nor (gm_n7461, in_18, in_17, in_16, gm_n7460, in_19);
	nand (gm_n7462, gm_n7461, in_21, gm_n45);
	nand (gm_n7463, gm_n46, in_15, in_14, gm_n1938, gm_n81);
	nor (gm_n7464, in_20, in_19, in_18, gm_n7463, gm_n71);
	nor (gm_n7465, gm_n48, gm_n53, gm_n52, gm_n5906, gm_n49);
	nand (gm_n7466, in_16, gm_n63, in_14, gm_n7465, in_17);
	nor (gm_n7467, gm_n45, in_19, gm_n47, gm_n7466, gm_n71);
	and (gm_n7468, in_13, in_12, in_11, gm_n5838, gm_n50);
	nand (gm_n7469, in_17, in_16, in_15, gm_n7468, gm_n47);
	nor (gm_n7470, gm_n71, gm_n45, in_19, gm_n7469);
	and (gm_n7471, gm_n49, gm_n48, in_11, gm_n4794, gm_n50);
	nand (gm_n7472, in_17, in_16, gm_n63, gm_n7471, in_18);
	nor (gm_n7473, in_21, in_20, in_19, gm_n7472);
	or (gm_n7474, in_13, in_12, gm_n53, gm_n938, in_14);
	nor (gm_n7475, in_17, in_16, in_15, gm_n7474, gm_n47);
	nand (gm_n7476, in_21, gm_n45, gm_n62, gm_n7475);
	and (gm_n7477, gm_n52, in_9, in_8, gm_n2708, gm_n53);
	nand (gm_n7478, in_14, gm_n49, in_12, gm_n7477, gm_n63);
	nor (gm_n7479, gm_n47, gm_n81, in_16, gm_n7478, in_19);
	nand (gm_n7480, gm_n7479, gm_n71, in_20);
	nand (gm_n7481, in_15, in_14, gm_n49, gm_n7064, in_16);
	nor (gm_n7482, in_19, in_18, in_17, gm_n7481, gm_n45);
	nand (gm_n7483, gm_n7482, in_21);
	and (gm_n7484, gm_n53, gm_n52, gm_n51, gm_n2194, gm_n48);
	nand (gm_n7485, gm_n63, gm_n50, in_13, gm_n7484, gm_n46);
	nor (gm_n7486, in_19, in_18, gm_n81, gm_n7485, in_20);
	nand (gm_n7487, gm_n7486, in_21);
	nand (gm_n7488, in_11, in_10, gm_n51, gm_n2088, in_12);
	nor (gm_n7489, in_15, in_14, gm_n49, gm_n7488, in_16);
	nand (gm_n7490, gm_n62, gm_n47, gm_n81, gm_n7489, gm_n45);
	nor (gm_n7491, gm_n7490, gm_n71);
	nand (gm_n7492, in_11, gm_n52, gm_n51, gm_n2088, in_12);
	nor (gm_n7493, in_15, in_14, in_13, gm_n7492, gm_n46);
	nand (gm_n7494, gm_n62, in_18, in_17, gm_n7493, gm_n45);
	nor (gm_n7495, gm_n7494, gm_n71);
	nor (gm_n7496, gm_n3826, gm_n49, gm_n48);
	nand (gm_n7497, gm_n46, in_15, gm_n50, gm_n7496, gm_n81);
	nor (gm_n7498, in_20, in_19, in_18, gm_n7497, gm_n71);
	or (gm_n7499, gm_n53, gm_n52, gm_n51, gm_n5263, in_12);
	nor (gm_n7500, in_15, in_14, in_13, gm_n7499, in_16);
	nand (gm_n7501, gm_n62, gm_n47, in_17, gm_n7500, in_20);
	nor (gm_n7502, gm_n7501, in_21);
	nand (gm_n7503, gm_n48, in_11, in_10, gm_n1688, in_13);
	nor (gm_n7504, in_16, gm_n63, in_14, gm_n7503, gm_n81);
	nand (gm_n7505, gm_n45, gm_n62, gm_n47, gm_n7504, gm_n71);
	nor (gm_n7506, in_10, gm_n51, in_8, gm_n3821);
	nand (gm_n7507, in_13, gm_n48, in_11, gm_n7506, gm_n50);
	nor (gm_n7508, gm_n81, gm_n46, in_15, gm_n7507, gm_n47);
	nand (gm_n7509, gm_n71, in_20, in_19, gm_n7508);
	nor (gm_n7510, in_9, gm_n64, in_7, gm_n463, in_10);
	nand (gm_n7511, gm_n49, in_12, gm_n53, gm_n7510, gm_n50);
	nor (gm_n7512, gm_n81, in_16, gm_n63, gm_n7511, in_18);
	nand (gm_n7513, gm_n71, in_20, gm_n62, gm_n7512);
	nor (gm_n7514, gm_n53, in_10, gm_n51, gm_n2445);
	nand (gm_n7515, in_14, gm_n49, in_12, gm_n7514, in_15);
	nor (gm_n7516, in_18, in_17, gm_n46, gm_n7515, in_19);
	nand (gm_n7517, gm_n7516, gm_n71, in_20);
	or (gm_n7518, in_16, gm_n63, in_14, gm_n1841, in_17);
	nor (gm_n7519, in_20, gm_n62, in_18, gm_n7518, gm_n71);
	nand (gm_n7520, gm_n929, gm_n52, gm_n51);
	nor (gm_n7521, gm_n49, gm_n48, gm_n53, gm_n7520, in_14);
	nand (gm_n7522, gm_n81, gm_n46, gm_n63, gm_n7521, gm_n47);
	nor (gm_n7523, gm_n71, gm_n45, in_19, gm_n7522);
	and (gm_n7524, gm_n53, gm_n52, gm_n51, gm_n1222);
	and (gm_n7525, in_14, in_13, gm_n48, gm_n7524, in_15);
	nand (gm_n7526, gm_n47, in_17, gm_n46, gm_n7525, in_19);
	nor (gm_n7527, gm_n7526, in_21, in_20);
	and (gm_n7528, in_15, in_14, gm_n49, gm_n1705, in_16);
	nand (gm_n7529, gm_n62, in_18, in_17, gm_n7528, gm_n45);
	nor (gm_n7530, gm_n7529, gm_n71);
	or (gm_n7531, in_12, in_11, in_10, gm_n6897, in_13);
	nor (gm_n7532, gm_n46, gm_n63, gm_n50, gm_n7531, in_17);
	nand (gm_n7533, gm_n45, in_19, in_18, gm_n7532, gm_n71);
	nor (gm_n7534, gm_n53, in_10, gm_n51, gm_n607, gm_n48);
	nand (gm_n7535, in_15, gm_n50, in_13, gm_n7534, in_16);
	nor (gm_n7536, gm_n62, in_18, in_17, gm_n7535, in_20);
	nand (gm_n7537, gm_n7536, gm_n71);
	nand (gm_n7538, in_14, in_13, in_12, gm_n7111, gm_n63);
	nor (gm_n7539, gm_n47, gm_n81, gm_n46, gm_n7538, gm_n62);
	nand (gm_n7540, gm_n7539, gm_n71, gm_n45);
	nand (gm_n7541, in_13, gm_n48, gm_n53, gm_n1776, in_14);
	nor (gm_n7542, gm_n81, gm_n46, gm_n63, gm_n7541, gm_n47);
	nand (gm_n7543, in_21, gm_n45, in_19, gm_n7542);
	nor (gm_n7544, gm_n48, gm_n53, in_10, gm_n639, in_13);
	nand (gm_n7545, in_16, in_15, gm_n50, gm_n7544, in_17);
	nor (gm_n7546, gm_n45, in_19, in_18, gm_n7545, in_21);
	and (gm_n7547, gm_n49, in_12, in_11, gm_n5784, in_14);
	nand (gm_n7548, in_17, gm_n46, in_15, gm_n7547, gm_n47);
	nor (gm_n7549, gm_n71, in_20, in_19, gm_n7548);
	nor (gm_n7550, in_14, in_13, gm_n48, gm_n5060, gm_n63);
	nand (gm_n7551, in_18, gm_n81, gm_n46, gm_n7550, gm_n62);
	nor (gm_n7552, gm_n7551, gm_n71, in_20);
	nor (gm_n7553, in_14, in_13, gm_n48, gm_n2504, gm_n63);
	nand (gm_n7554, gm_n47, gm_n81, gm_n46, gm_n7553, gm_n62);
	nor (gm_n7555, gm_n7554, gm_n71, gm_n45);
	nor (gm_n7556, gm_n81, in_16, in_15, gm_n1539, in_18);
	nand (gm_n7557, in_21, in_20, in_19, gm_n7556);
	nand (gm_n7558, gm_n49, gm_n48, in_11, gm_n1584, gm_n50);
	nor (gm_n7559, in_17, in_16, in_15, gm_n7558, in_18);
	nand (gm_n7560, in_21, in_20, gm_n62, gm_n7559);
	or (gm_n7561, gm_n48, gm_n53, gm_n52, gm_n3773, in_13);
	nor (gm_n7562, in_16, gm_n63, in_14, gm_n7561, gm_n81);
	nand (gm_n7563, gm_n45, in_19, in_18, gm_n7562, in_21);
	and (gm_n7564, in_10, gm_n51, gm_n64, gm_n302, gm_n53);
	and (gm_n7565, gm_n50, gm_n49, gm_n48, gm_n7564, in_15);
	and (gm_n7566, gm_n47, gm_n81, in_16, gm_n7565, in_19);
	nand (gm_n7567, gm_n7566, gm_n71, in_20);
	nor (gm_n7568, gm_n53, gm_n52, gm_n51, gm_n4314, gm_n48);
	nand (gm_n7569, gm_n7568, gm_n50, gm_n49);
	or (gm_n7570, gm_n81, gm_n46, in_15, gm_n7569, in_18);
	nor (gm_n7571, gm_n71, gm_n45, gm_n62, gm_n7570);
	or (gm_n7572, in_9, gm_n64, gm_n55, gm_n259, in_10);
	nor (gm_n7573, gm_n49, in_12, in_11, gm_n7572, gm_n50);
	nand (gm_n7574, gm_n81, in_16, in_15, gm_n7573, in_18);
	nor (gm_n7575, gm_n71, gm_n45, gm_n62, gm_n7574);
	nor (gm_n7576, in_14, gm_n49, in_12, gm_n4258, gm_n63);
	nand (gm_n7577, in_18, gm_n81, in_16, gm_n7576, in_19);
	nor (gm_n7578, gm_n7577, in_21, gm_n45);
	and (gm_n7579, gm_n929, in_10, gm_n51);
	and (gm_n7580, gm_n49, gm_n48, in_11, gm_n7579, in_14);
	nand (gm_n7581, gm_n81, in_16, in_15, gm_n7580, in_18);
	nor (gm_n7582, in_21, gm_n45, in_19, gm_n7581);
	nand (gm_n7583, in_14, in_13, in_12, gm_n7524, in_15);
	nor (gm_n7584, gm_n47, gm_n81, gm_n46, gm_n7583, gm_n62);
	nand (gm_n7585, gm_n7584, in_21, in_20);
	nand (gm_n7586, in_12, in_11, gm_n52, gm_n3309, in_13);
	nor (gm_n7587, in_16, in_15, in_14, gm_n7586, in_17);
	nand (gm_n7588, gm_n45, in_19, gm_n47, gm_n7587, gm_n71);
	nand (gm_n7589, in_12, gm_n53, gm_n52, gm_n4911, in_13);
	nor (gm_n7590, gm_n46, in_15, in_14, gm_n7589, in_17);
	nand (gm_n7591, gm_n45, in_19, in_18, gm_n7590, in_21);
	nand (gm_n7592, gm_n48, in_11, gm_n52, gm_n589, gm_n49);
	nor (gm_n7593, in_16, gm_n63, in_14, gm_n7592, in_17);
	nand (gm_n7594, in_20, gm_n62, in_18, gm_n7593, in_21);
	nor (gm_n7595, in_15, gm_n50, in_13, gm_n1880, in_16);
	nand (gm_n7596, gm_n62, in_18, in_17, gm_n7595, gm_n45);
	nor (gm_n7597, gm_n7596, in_21);
	nand (gm_n7598, in_16, gm_n63, gm_n50, gm_n4644, gm_n81);
	nor (gm_n7599, in_20, gm_n62, gm_n47, gm_n7598, in_21);
	nor (gm_n7600, in_12, gm_n53, in_10, gm_n1398, gm_n49);
	nand (gm_n7601, in_16, in_15, gm_n50, gm_n7600, gm_n81);
	nor (gm_n7602, gm_n45, in_19, gm_n47, gm_n7601, gm_n71);
	nand (gm_n7603, in_17, in_16, in_15, gm_n516, gm_n47);
	nor (gm_n7604, in_21, in_20, gm_n62, gm_n7603);
	nand (gm_n7605, in_12, gm_n53, in_10, gm_n2819, in_13);
	nor (gm_n7606, in_16, gm_n63, gm_n50, gm_n7605, in_17);
	nand (gm_n7607, gm_n45, in_19, in_18, gm_n7606, gm_n71);
	nand (gm_n7608, gm_n48, in_11, gm_n52, gm_n200, in_13);
	nor (gm_n7609, gm_n46, gm_n63, in_14, gm_n7608, gm_n81);
	nand (gm_n7610, in_20, in_19, gm_n47, gm_n7609, gm_n71);
	and (gm_n7611, gm_n1380, in_10, gm_n51);
	nand (gm_n7612, gm_n49, in_12, gm_n53, gm_n7611, in_14);
	nor (gm_n7613, gm_n81, gm_n46, gm_n63, gm_n7612, in_18);
	nand (gm_n7614, in_21, gm_n45, gm_n62, gm_n7613);
	and (gm_n7615, gm_n53, gm_n52, in_9, gm_n1788, gm_n48);
	nand (gm_n7616, gm_n63, in_14, in_13, gm_n7615, gm_n46);
	nor (gm_n7617, gm_n62, gm_n47, in_17, gm_n7616, gm_n45);
	nand (gm_n7618, gm_n7617, gm_n71);
	nand (gm_n7619, in_11, gm_n52, gm_n51, gm_n1704);
	nor (gm_n7620, gm_n50, in_13, gm_n48, gm_n7619, in_15);
	nand (gm_n7621, in_18, in_17, gm_n46, gm_n7620, in_19);
	nor (gm_n7622, gm_n7621, in_21, in_20);
	nor (gm_n7623, gm_n50, in_13, in_12, gm_n4748, gm_n63);
	nand (gm_n7624, in_18, gm_n81, in_16, gm_n7623, gm_n62);
	nor (gm_n7625, gm_n7624, in_21, in_20);
	nor (gm_n7626, in_11, in_10, in_9, gm_n453);
	and (gm_n7627, in_14, in_13, in_12, gm_n7626, in_15);
	nand (gm_n7628, in_18, gm_n81, gm_n46, gm_n7627, gm_n62);
	nor (gm_n7629, gm_n7628, gm_n71, in_20);
	nand (gm_n7630, in_11, gm_n52, in_9, gm_n1360, in_12);
	nor (gm_n7631, in_15, in_14, gm_n49, gm_n7630, in_16);
	nand (gm_n7632, in_19, gm_n47, gm_n81, gm_n7631, gm_n45);
	nor (gm_n7633, gm_n7632, gm_n71);
	nor (gm_n7634, gm_n53, gm_n52, gm_n51, gm_n1763, gm_n48);
	nand (gm_n7635, in_15, in_14, in_13, gm_n7634, gm_n46);
	nor (gm_n7636, gm_n62, gm_n47, in_17, gm_n7635, in_20);
	nand (gm_n7637, gm_n7636, in_21);
	nand (gm_n7638, in_12, in_11, gm_n52, gm_n654, in_13);
	nor (gm_n7639, in_16, in_15, gm_n50, gm_n7638, in_17);
	nand (gm_n7640, gm_n45, in_19, gm_n47, gm_n7639, gm_n71);
	nand (gm_n7641, gm_n48, in_11, gm_n52, gm_n5616, gm_n49);
	nor (gm_n7642, gm_n46, gm_n63, gm_n50, gm_n7641, gm_n81);
	nand (gm_n7643, in_20, gm_n62, in_18, gm_n7642, gm_n71);
	or (gm_n7644, in_12, gm_n53, in_10, gm_n1824, gm_n49);
	nor (gm_n7645, in_16, gm_n63, in_14, gm_n7644, gm_n81);
	nand (gm_n7646, in_20, in_19, gm_n47, gm_n7645, gm_n71);
	nor (gm_n7647, gm_n49, gm_n48, gm_n53, gm_n938);
	nand (gm_n7648, in_16, gm_n63, in_14, gm_n7647, gm_n81);
	nor (gm_n7649, gm_n45, in_19, in_18, gm_n7648, gm_n71);
	or (gm_n7650, in_9, in_8, in_7, gm_n588, gm_n52);
	nor (gm_n7651, in_13, in_12, gm_n53, gm_n7650, gm_n50);
	nand (gm_n7652, in_17, gm_n46, in_15, gm_n7651, gm_n47);
	nor (gm_n7653, gm_n71, in_20, in_19, gm_n7652);
	and (gm_n7654, in_21, in_20, gm_n62, gm_n953);
	nor (gm_n7655, in_13, in_12, gm_n53, gm_n6621, gm_n50);
	nand (gm_n7656, gm_n81, in_16, in_15, gm_n7655, in_18);
	nor (gm_n7657, in_21, gm_n45, gm_n62, gm_n7656);
	nand (gm_n7658, gm_n48, gm_n53, in_10, gm_n1840, gm_n49);
	nor (gm_n7659, in_16, gm_n63, gm_n50, gm_n7658, gm_n81);
	nand (gm_n7660, in_20, gm_n62, in_18, gm_n7659, in_21);
	nor (gm_n7661, gm_n3697, in_10, gm_n51);
	nand (gm_n7662, in_13, gm_n48, gm_n53, gm_n7661, in_14);
	nor (gm_n7663, gm_n81, gm_n46, gm_n63, gm_n7662, gm_n47);
	nand (gm_n7664, in_21, gm_n45, gm_n62, gm_n7663);
	nor (gm_n7665, gm_n46, gm_n63, in_14, gm_n3045, gm_n81);
	nand (gm_n7666, in_20, gm_n62, gm_n47, gm_n7665, gm_n71);
	nand (gm_n7667, in_12, in_11, in_10, gm_n589, in_13);
	nor (gm_n7668, in_16, gm_n63, in_14, gm_n7667, gm_n81);
	nand (gm_n7669, gm_n45, gm_n62, in_18, gm_n7668, gm_n71);
	nand (gm_n7670, in_11, in_10, in_9, gm_n4042, in_12);
	nor (gm_n7671, in_15, gm_n50, in_13, gm_n7670, in_16);
	nand (gm_n7672, in_19, in_18, gm_n81, gm_n7671, gm_n45);
	nor (gm_n7673, gm_n7672, gm_n71);
	and (gm_n7674, in_12, in_11, in_10, gm_n980, gm_n49);
	nand (gm_n7675, in_16, in_15, in_14, gm_n7674, gm_n81);
	nor (gm_n7676, in_20, in_19, gm_n47, gm_n7675, gm_n71);
	or (gm_n7677, in_9, in_8, gm_n55, gm_n463, gm_n52);
	nor (gm_n7678, in_13, gm_n48, in_11, gm_n7677, gm_n50);
	nand (gm_n7679, gm_n81, gm_n46, in_15, gm_n7678, gm_n47);
	nor (gm_n7680, gm_n71, gm_n45, in_19, gm_n7679);
	nand (gm_n7681, gm_n52, gm_n51, gm_n64, gm_n1088, in_11);
	nor (gm_n7682, gm_n7681, gm_n49, gm_n48);
	nand (gm_n7683, in_16, in_15, in_14, gm_n7682, in_17);
	nor (gm_n7684, gm_n45, in_19, gm_n47, gm_n7683, gm_n71);
	or (gm_n7685, in_12, gm_n53, in_10, gm_n3924, gm_n49);
	nor (gm_n7686, in_16, in_15, in_14, gm_n7685, in_17);
	nand (gm_n7687, in_20, gm_n62, gm_n47, gm_n7686, in_21);
	and (gm_n7688, gm_n53, in_10, gm_n51, gm_n210, gm_n48);
	nand (gm_n7689, gm_n63, in_14, gm_n49, gm_n7688, gm_n46);
	nor (gm_n7690, gm_n62, in_18, in_17, gm_n7689, gm_n45);
	nand (gm_n7691, gm_n7690, in_21);
	nand (gm_n7692, gm_n49, in_12, gm_n53, gm_n7506, in_14);
	nor (gm_n7693, gm_n81, gm_n46, gm_n63, gm_n7692, gm_n47);
	nand (gm_n7694, in_21, gm_n45, in_19, gm_n7693);
	nor (gm_n7695, gm_n1533, gm_n52, gm_n51);
	nand (gm_n7696, gm_n49, in_12, gm_n53, gm_n7695, in_14);
	nor (gm_n7697, in_17, gm_n46, gm_n63, gm_n7696, in_18);
	nand (gm_n7698, gm_n71, in_20, in_19, gm_n7697);
	nor (gm_n7699, gm_n50, in_13, gm_n48, gm_n869, in_15);
	nand (gm_n7700, gm_n47, in_17, in_16, gm_n7699, gm_n62);
	nor (gm_n7701, gm_n7700, in_21, gm_n45);
	nand (gm_n7702, in_8, in_7, gm_n82, gm_n379, gm_n51);
	nor (gm_n7703, gm_n48, in_11, in_10, gm_n7702, gm_n49);
	nand (gm_n7704, gm_n46, in_15, gm_n50, gm_n7703, in_17);
	nor (gm_n7705, in_20, gm_n62, in_18, gm_n7704, in_21);
	nand (gm_n7706, in_16, gm_n63, in_14, gm_n4320, gm_n81);
	nor (gm_n7707, gm_n45, in_19, gm_n47, gm_n7706, in_21);
	nand (gm_n7708, gm_n53, in_10, in_9, gm_n2254, gm_n48);
	nor (gm_n7709, in_15, in_14, in_13, gm_n7708, in_16);
	nand (gm_n7710, gm_n62, gm_n47, in_17, gm_n7709, in_20);
	nor (gm_n7711, gm_n7710, gm_n71);
	nand (gm_n7712, in_12, gm_n53, in_10, gm_n2182, in_13);
	nor (gm_n7713, in_16, in_15, gm_n50, gm_n7712, in_17);
	nand (gm_n7714, gm_n45, in_19, gm_n47, gm_n7713, gm_n71);
	and (gm_n7715, in_11, in_10, in_9, gm_n1360, in_12);
	nand (gm_n7716, gm_n63, in_14, gm_n49, gm_n7715, gm_n46);
	nor (gm_n7717, in_19, gm_n47, in_17, gm_n7716, gm_n45);
	nand (gm_n7718, gm_n7717, gm_n71);
	and (gm_n7719, in_12, gm_n53, gm_n52, gm_n2672, in_13);
	and (gm_n7720, gm_n46, gm_n63, gm_n50, gm_n7719, gm_n81);
	nand (gm_n7721, gm_n45, in_19, gm_n47, gm_n7720, in_21);
	nand (gm_n7722, in_13, gm_n48, gm_n53, gm_n2499, gm_n50);
	nor (gm_n7723, in_17, in_16, in_15, gm_n7722, in_18);
	nand (gm_n7724, gm_n71, in_20, in_19, gm_n7723);
	nand (gm_n7725, in_11, gm_n52, in_9, gm_n1192, gm_n48);
	nor (gm_n7726, gm_n63, in_14, in_13, gm_n7725, in_16);
	nand (gm_n7727, gm_n62, in_18, in_17, gm_n7726, gm_n45);
	nor (gm_n7728, gm_n7727, in_21);
	and (gm_n7729, gm_n53, gm_n52, in_9, gm_n3768);
	and (gm_n7730, gm_n50, gm_n49, gm_n48, gm_n7729, in_15);
	nand (gm_n7731, gm_n47, in_17, in_16, gm_n7730, gm_n62);
	nor (gm_n7732, gm_n7731, in_21, in_20);
	and (gm_n7733, in_12, gm_n53, in_10, gm_n2890, in_13);
	nand (gm_n7734, gm_n46, gm_n63, gm_n50, gm_n7733, in_17);
	nor (gm_n7735, gm_n45, gm_n62, gm_n47, gm_n7734, gm_n71);
	nor (gm_n7736, gm_n48, gm_n53, gm_n52, gm_n5268, gm_n49);
	nand (gm_n7737, gm_n46, gm_n63, gm_n50, gm_n7736, gm_n81);
	nor (gm_n7738, gm_n45, gm_n62, gm_n47, gm_n7737, gm_n71);
	nor (gm_n7739, gm_n53, gm_n52, in_9, gm_n4489, gm_n48);
	nand (gm_n7740, gm_n63, gm_n50, in_13, gm_n7739, in_16);
	nor (gm_n7741, gm_n62, gm_n47, in_17, gm_n7740, gm_n45);
	nand (gm_n7742, gm_n7741, in_21);
	nand (gm_n7743, gm_n48, gm_n53, gm_n52, gm_n1861, in_13);
	nor (gm_n7744, gm_n46, gm_n63, gm_n50, gm_n7743, in_17);
	nand (gm_n7745, gm_n45, gm_n62, in_18, gm_n7744, in_21);
	nor (gm_n7746, gm_n52, in_9, in_8, gm_n907, gm_n53);
	nand (gm_n7747, in_14, gm_n49, in_12, gm_n7746, gm_n63);
	nor (gm_n7748, in_18, gm_n81, in_16, gm_n7747, gm_n62);
	nand (gm_n7749, gm_n7748, gm_n71, in_20);
	nand (gm_n7750, in_13, gm_n48, in_11, gm_n1257, in_14);
	nor (gm_n7751, gm_n81, in_16, gm_n63, gm_n7750, gm_n47);
	nand (gm_n7752, in_21, gm_n45, gm_n62, gm_n7751);
	nor (gm_n7753, gm_n50, gm_n49, gm_n48, gm_n6592, in_15);
	nand (gm_n7754, gm_n47, in_17, gm_n46, gm_n7753, in_19);
	nor (gm_n7755, gm_n7754, in_21, in_20);
	or (gm_n7756, in_11, gm_n52, gm_n51, gm_n2902, in_12);
	nor (gm_n7757, gm_n63, gm_n50, in_13, gm_n7756, in_16);
	nand (gm_n7758, gm_n62, in_18, gm_n81, gm_n7757, gm_n45);
	nor (gm_n7759, gm_n7758, gm_n71);
	nand (gm_n7760, gm_n46, gm_n63, in_14, gm_n5061, gm_n81);
	nor (gm_n7761, in_20, gm_n62, in_18, gm_n7760, in_21);
	nor (gm_n7762, gm_n48, in_11, gm_n52, gm_n6451, in_13);
	nand (gm_n7763, gm_n46, gm_n63, gm_n50, gm_n7762, in_17);
	nor (gm_n7764, gm_n45, in_19, gm_n47, gm_n7763, in_21);
	nor (gm_n7765, gm_n3077, gm_n51, gm_n64);
	nand (gm_n7766, in_12, in_11, in_10, gm_n7765, gm_n49);
	nor (gm_n7767, in_16, gm_n63, gm_n50, gm_n7766, in_17);
	nand (gm_n7768, gm_n45, gm_n62, in_18, gm_n7767, gm_n71);
	nand (gm_n7769, in_14, gm_n49, in_12, gm_n5693, in_15);
	nor (gm_n7770, in_18, gm_n81, in_16, gm_n7769, gm_n62);
	nand (gm_n7771, gm_n7770, gm_n71, gm_n45);
	and (gm_n7772, in_16, gm_n63, in_14, gm_n4522, gm_n81);
	nand (gm_n7773, in_20, in_19, gm_n47, gm_n7772, in_21);
	nor (gm_n7774, in_11, in_10, gm_n51, gm_n873, gm_n48);
	nand (gm_n7775, in_15, in_14, in_13, gm_n7774, in_16);
	nor (gm_n7776, gm_n62, gm_n47, gm_n81, gm_n7775, in_20);
	nand (gm_n7777, gm_n7776, in_21);
	nand (gm_n7778, gm_n53, in_10, in_9, gm_n1192, gm_n48);
	nor (gm_n7779, in_15, gm_n50, in_13, gm_n7778, gm_n46);
	nand (gm_n7780, gm_n62, in_18, in_17, gm_n7779, in_20);
	nor (gm_n7781, gm_n7780, in_21);
	and (gm_n7782, gm_n48, gm_n53, in_10, gm_n6572, gm_n49);
	nand (gm_n7783, gm_n46, gm_n63, in_14, gm_n7782, in_17);
	nor (gm_n7784, in_20, gm_n62, gm_n47, gm_n7783, gm_n71);
	nor (gm_n7785, in_12, in_11, in_10, gm_n7068, in_13);
	nand (gm_n7786, in_16, in_15, in_14, gm_n7785, in_17);
	nor (gm_n7787, gm_n45, gm_n62, gm_n47, gm_n7786, gm_n71);
	and (gm_n7788, gm_n6500, gm_n52, in_9);
	and (gm_n7789, in_13, gm_n48, in_11, gm_n7788, in_14);
	nand (gm_n7790, in_17, gm_n46, gm_n63, gm_n7789, gm_n47);
	nor (gm_n7791, in_21, in_20, in_19, gm_n7790);
	nor (gm_n7792, gm_n48, gm_n53, gm_n52, gm_n7072, gm_n49);
	and (gm_n7793, gm_n46, gm_n63, gm_n50, gm_n7792, in_17);
	nand (gm_n7794, in_20, gm_n62, gm_n47, gm_n7793, gm_n71);
	nand (gm_n7795, gm_n50, in_13, gm_n48, gm_n572, in_15);
	nor (gm_n7796, in_18, in_17, in_16, gm_n7795, gm_n62);
	nand (gm_n7797, gm_n7796, gm_n71, gm_n45);
	nand (gm_n7798, gm_n49, gm_n48, gm_n53, gm_n2203, gm_n50);
	nor (gm_n7799, gm_n81, gm_n46, in_15, gm_n7798, gm_n47);
	nand (gm_n7800, in_21, gm_n45, gm_n62, gm_n7799);
	nand (gm_n7801, in_12, gm_n53, gm_n52, gm_n3039, gm_n49);
	nor (gm_n7802, gm_n46, in_15, in_14, gm_n7801, in_17);
	nand (gm_n7803, in_20, gm_n62, in_18, gm_n7802, gm_n71);
	nor (gm_n7804, gm_n50, gm_n49, gm_n48, gm_n3341, in_15);
	nand (gm_n7805, in_18, gm_n81, gm_n46, gm_n7804, gm_n62);
	nor (gm_n7806, gm_n7805, in_21, in_20);
	and (gm_n7807, in_14, in_13, gm_n48, gm_n406, in_15);
	nand (gm_n7808, gm_n47, in_17, in_16, gm_n7807, in_19);
	nor (gm_n7809, gm_n7808, in_21, in_20);
	nor (gm_n7810, in_13, gm_n48, in_11, gm_n6644, in_14);
	nand (gm_n7811, gm_n81, gm_n46, gm_n63, gm_n7810, in_18);
	nor (gm_n7812, gm_n71, in_20, gm_n62, gm_n7811);
	and (gm_n7813, in_11, gm_n52, gm_n51, gm_n232, gm_n48);
	and (gm_n7814, gm_n63, gm_n50, gm_n49, gm_n7813, in_16);
	nand (gm_n7815, in_19, in_18, gm_n81, gm_n7814, gm_n45);
	nor (gm_n7816, gm_n7815, in_21);
	and (gm_n7817, in_12, in_11, gm_n52, gm_n6405, gm_n49);
	and (gm_n7818, gm_n46, gm_n63, gm_n50, gm_n7817, in_17);
	nand (gm_n7819, in_20, gm_n62, gm_n47, gm_n7818, gm_n71);
	nand (gm_n7820, in_12, in_11, gm_n52, gm_n311, gm_n49);
	nor (gm_n7821, gm_n46, gm_n63, in_14, gm_n7820, in_17);
	nand (gm_n7822, gm_n45, gm_n62, in_18, gm_n7821, gm_n71);
	or (gm_n7823, in_9, gm_n64, gm_n55, gm_n588, in_10);
	nor (gm_n7824, gm_n49, gm_n48, in_11, gm_n7823, in_14);
	and (gm_n7825, in_17, in_16, in_15, gm_n7824, in_18);
	nand (gm_n7826, in_21, gm_n45, gm_n62, gm_n7825);
	nor (gm_n7827, in_17, gm_n46, gm_n63, gm_n5978, in_18);
	nand (gm_n7828, gm_n71, gm_n45, in_19, gm_n7827);
	nor (gm_n7829, gm_n50, gm_n49, in_12, gm_n3584, gm_n63);
	nand (gm_n7830, in_18, in_17, gm_n46, gm_n7829, in_19);
	nor (gm_n7831, gm_n7830, gm_n71, in_20);
	nor (gm_n7832, in_13, in_12, gm_n53, gm_n5052, in_14);
	nand (gm_n7833, gm_n81, in_16, in_15, gm_n7832, gm_n47);
	nor (gm_n7834, in_21, gm_n45, gm_n62, gm_n7833);
	nor (gm_n7835, gm_n48, gm_n53, in_10, gm_n7227, gm_n49);
	nand (gm_n7836, gm_n46, gm_n63, gm_n50, gm_n7835, gm_n81);
	nor (gm_n7837, in_20, gm_n62, gm_n47, gm_n7836, in_21);
	nor (gm_n7838, gm_n50, gm_n49, in_12, gm_n1193, in_15);
	nand (gm_n7839, gm_n47, gm_n81, in_16, gm_n7838, in_19);
	nor (gm_n7840, gm_n7839, in_21, in_20);
	nand (gm_n7841, gm_n49, in_12, in_11, gm_n505, in_14);
	nor (gm_n7842, gm_n81, in_16, in_15, gm_n7841, gm_n47);
	nand (gm_n7843, gm_n71, in_20, gm_n62, gm_n7842);
	nor (gm_n7844, in_17, in_16, gm_n63, gm_n7569, in_18);
	nand (gm_n7845, in_21, gm_n45, gm_n62, gm_n7844);
	nor (gm_n7846, in_11, in_10, in_9, gm_n2914, in_12);
	nand (gm_n7847, in_15, gm_n50, in_13, gm_n7846, gm_n46);
	nor (gm_n7848, in_19, in_18, gm_n81, gm_n7847, gm_n45);
	nand (gm_n7849, gm_n7848, gm_n71);
	nand (gm_n7850, in_15, gm_n50, in_13, gm_n5071, gm_n46);
	nor (gm_n7851, in_19, in_18, gm_n81, gm_n7850, in_20);
	nand (gm_n7852, gm_n7851, in_21);
	nand (gm_n7853, gm_n7055, in_9);
	nor (gm_n7854, in_12, in_11, in_10, gm_n7853, in_13);
	nand (gm_n7855, in_16, gm_n63, in_14, gm_n7854, in_17);
	nor (gm_n7856, gm_n45, in_19, in_18, gm_n7855, in_21);
	nor (gm_n7857, gm_n53, in_10, gm_n51, gm_n2849);
	and (gm_n7858, in_14, in_13, in_12, gm_n7857, gm_n63);
	nand (gm_n7859, gm_n47, gm_n81, gm_n46, gm_n7858, in_19);
	nor (gm_n7860, gm_n7859, gm_n71, gm_n45);
	nand (gm_n7861, gm_n53, in_10, in_9, gm_n997, in_12);
	nor (gm_n7862, in_15, gm_n50, gm_n49, gm_n7861, in_16);
	nand (gm_n7863, gm_n62, gm_n47, gm_n81, gm_n7862, gm_n45);
	nor (gm_n7864, gm_n7863, gm_n71);
	nand (gm_n7865, in_11, in_10, gm_n51, gm_n848, gm_n48);
	nor (gm_n7866, in_15, in_14, gm_n49, gm_n7865, in_16);
	nand (gm_n7867, in_19, in_18, gm_n81, gm_n7866, in_20);
	nor (gm_n7868, gm_n7867, gm_n71);
	nand (gm_n7869, gm_n63, gm_n50, gm_n49, gm_n6496, in_16);
	nor (gm_n7870, gm_n62, in_18, gm_n81, gm_n7869, in_20);
	nand (gm_n7871, gm_n7870, gm_n71);
	nor (gm_n7872, in_11, gm_n52, gm_n51, gm_n322, in_12);
	nand (gm_n7873, gm_n63, gm_n50, gm_n49, gm_n7872, gm_n46);
	nor (gm_n7874, gm_n62, in_18, gm_n81, gm_n7873, gm_n45);
	nand (gm_n7875, gm_n7874, in_21);
	nand (gm_n7876, gm_n48, gm_n53, gm_n52, gm_n3659, gm_n49);
	nor (gm_n7877, in_16, gm_n63, in_14, gm_n7876, in_17);
	nand (gm_n7878, in_20, gm_n62, in_18, gm_n7877, in_21);
	and (gm_n7879, in_11, gm_n52, in_9, gm_n3043, gm_n48);
	nand (gm_n7880, gm_n63, in_14, gm_n49, gm_n7879, gm_n46);
	nor (gm_n7881, in_19, in_18, gm_n81, gm_n7880, gm_n45);
	nand (gm_n7882, gm_n7881, gm_n71);
	nor (gm_n7883, gm_n51, in_8, in_7, gm_n588, gm_n52);
	nand (gm_n7884, gm_n49, gm_n48, in_11, gm_n7883, in_14);
	nor (gm_n7885, gm_n81, gm_n46, gm_n63, gm_n7884, gm_n47);
	nand (gm_n7886, in_21, in_20, gm_n62, gm_n7885);
	nand (gm_n7887, gm_n7878, gm_n7875, gm_n7871, gm_n7886, gm_n7882);
	nor (gm_n7888, gm_n7864, gm_n7860, gm_n7856, gm_n7887, gm_n7868);
	nand (gm_n7889, gm_n7849, gm_n7845, gm_n7843, gm_n7888, gm_n7852);
	nor (gm_n7890, gm_n7837, gm_n7834, gm_n7831, gm_n7889, gm_n7840);
	nand (gm_n7891, gm_n7826, gm_n7822, gm_n7819, gm_n7890, gm_n7828);
	nor (gm_n7892, gm_n7812, gm_n7809, gm_n7806, gm_n7891, gm_n7816);
	nand (gm_n7893, gm_n7800, gm_n7797, gm_n7794, gm_n7892, gm_n7803);
	nor (gm_n7894, gm_n7787, gm_n7784, gm_n7781, gm_n7893, gm_n7791);
	nand (gm_n7895, gm_n7773, gm_n7771, gm_n7768, gm_n7894, gm_n7777);
	nor (gm_n7896, gm_n7761, gm_n7759, gm_n7755, gm_n7895, gm_n7764);
	nand (gm_n7897, gm_n7749, gm_n7745, gm_n7742, gm_n7896, gm_n7752);
	nor (gm_n7898, gm_n7735, gm_n7732, gm_n7728, gm_n7897, gm_n7738);
	nand (gm_n7899, gm_n7721, gm_n7718, gm_n7714, gm_n7898, gm_n7724);
	nor (gm_n7900, gm_n7707, gm_n7705, gm_n7701, gm_n7899, gm_n7711);
	nand (gm_n7901, gm_n7694, gm_n7691, gm_n7687, gm_n7900, gm_n7698);
	nor (gm_n7902, gm_n7680, gm_n7676, gm_n7673, gm_n7901, gm_n7684);
	nand (gm_n7903, gm_n7666, gm_n7664, gm_n7660, gm_n7902, gm_n7669);
	nor (gm_n7904, gm_n7654, gm_n7653, gm_n7649, gm_n7903, gm_n7657);
	nand (gm_n7905, gm_n7643, gm_n7640, gm_n7637, gm_n7904, gm_n7646);
	nor (gm_n7906, gm_n7629, gm_n7625, gm_n7622, gm_n7905, gm_n7633);
	nand (gm_n7907, gm_n7614, gm_n7610, gm_n7607, gm_n7906, gm_n7618);
	nor (gm_n7908, gm_n7602, gm_n7599, gm_n7597, gm_n7907, gm_n7604);
	nand (gm_n7909, gm_n7591, gm_n7588, gm_n7585, gm_n7908, gm_n7594);
	nor (gm_n7910, gm_n7578, gm_n7575, gm_n7571, gm_n7909, gm_n7582);
	nand (gm_n7911, gm_n7563, gm_n7560, gm_n7557, gm_n7910, gm_n7567);
	nor (gm_n7912, gm_n7552, gm_n7549, gm_n7546, gm_n7911, gm_n7555);
	nand (gm_n7913, gm_n7540, gm_n7537, gm_n7533, gm_n7912, gm_n7543);
	nor (gm_n7914, gm_n7527, gm_n7523, gm_n7519, gm_n7913, gm_n7530);
	nand (gm_n7915, gm_n7513, gm_n7509, gm_n7505, gm_n7914, gm_n7517);
	nor (gm_n7916, gm_n7498, gm_n7495, gm_n7491, gm_n7915, gm_n7502);
	nand (gm_n7917, gm_n7483, gm_n7480, gm_n7476, gm_n7916, gm_n7487);
	nor (gm_n7918, gm_n7470, gm_n7467, gm_n7464, gm_n7917, gm_n7473);
	nand (gm_n7919, gm_n7458, gm_n7455, gm_n7452, gm_n7918, gm_n7462);
	nor (gm_n7920, gm_n7448, gm_n7445, gm_n7442, gm_n7919, gm_n7450);
	nand (gm_n7921, gm_n7436, gm_n7434, gm_n7431, gm_n7920, gm_n7439);
	nor (gm_n7922, gm_n7424, gm_n7421, gm_n7417, gm_n7921, gm_n7428);
	nand (gm_n7923, gm_n7412, gm_n7409, gm_n7406, gm_n7922, gm_n7415);
	nor (out_12, gm_n7923, gm_n7403);
	and (gm_n7925, gm_n52, gm_n51, gm_n64, gm_n921, in_11);
	and (gm_n7926, in_14, in_13, gm_n48, gm_n7925, in_15);
	nand (gm_n7927, gm_n47, in_17, in_16, gm_n7926, in_19);
	nor (gm_n7928, gm_n7927, gm_n71, gm_n45);
	and (gm_n7929, gm_n53, gm_n52, gm_n51, gm_n566, gm_n48);
	nand (gm_n7930, in_15, gm_n50, in_13, gm_n7929, gm_n46);
	nor (gm_n7931, gm_n62, gm_n47, in_17, gm_n7930, gm_n45);
	nand (gm_n7932, gm_n7931, in_21);
	nand (gm_n7933, in_14, in_13, gm_n48, gm_n2267, in_15);
	nor (gm_n7934, gm_n47, gm_n81, gm_n46, gm_n7933, in_19);
	nand (gm_n7935, gm_n7934, in_21, gm_n45);
	nand (gm_n7936, in_12, gm_n53, in_10, gm_n5822, in_13);
	nor (gm_n7937, gm_n46, in_15, in_14, gm_n7936, gm_n81);
	nand (gm_n7938, in_20, gm_n62, gm_n47, gm_n7937, in_21);
	and (gm_n7939, in_9, gm_n64, gm_n55, gm_n404, gm_n52);
	nand (gm_n7940, in_13, in_12, gm_n53, gm_n7939, gm_n50);
	nor (gm_n7941, in_17, in_16, in_15, gm_n7940, in_18);
	nand (gm_n7942, in_21, in_20, in_19, gm_n7941);
	nor (gm_n7943, gm_n63, gm_n50, gm_n49, gm_n6197, gm_n46);
	nand (gm_n7944, in_19, in_18, in_17, gm_n7943, gm_n45);
	nor (gm_n7945, gm_n7944, in_21);
	nand (gm_n7946, gm_n52, gm_n51, gm_n64, gm_n2708, in_11);
	nor (gm_n7947, gm_n50, in_13, gm_n48, gm_n7946, gm_n63);
	nand (gm_n7948, in_18, in_17, gm_n46, gm_n7947, gm_n62);
	nor (gm_n7949, gm_n7948, gm_n71, in_20);
	nor (gm_n7950, in_13, in_12, gm_n53, gm_n3494);
	nand (gm_n7951, in_16, in_15, gm_n50, gm_n7950, in_17);
	nor (gm_n7952, gm_n45, in_19, gm_n47, gm_n7951, gm_n71);
	nand (gm_n7953, in_11, in_10, in_9, gm_n1952);
	nor (gm_n7954, in_14, in_13, in_12, gm_n7953, in_15);
	nand (gm_n7955, in_18, in_17, in_16, gm_n7954, in_19);
	nor (gm_n7956, gm_n7955, gm_n71, in_20);
	nand (gm_n7957, in_13, in_12, gm_n53, gm_n3687, gm_n50);
	nor (gm_n7958, in_17, in_16, gm_n63, gm_n7957, in_18);
	nand (gm_n7959, gm_n71, in_20, in_19, gm_n7958);
	nand (gm_n7960, in_13, gm_n48, in_11, gm_n2218, in_14);
	nor (gm_n7961, gm_n81, in_16, gm_n63, gm_n7960, gm_n47);
	nand (gm_n7962, in_21, in_20, gm_n62, gm_n7961);
	nand (gm_n7963, gm_n50, in_13, gm_n48, gm_n6048, in_15);
	nor (gm_n7964, gm_n47, gm_n81, in_16, gm_n7963, gm_n62);
	nand (gm_n7965, gm_n7964, gm_n71, in_20);
	nor (gm_n7966, gm_n53, in_10, in_9, gm_n3198, in_12);
	nand (gm_n7967, in_15, in_14, gm_n49, gm_n7966, in_16);
	nor (gm_n7968, in_19, in_18, in_17, gm_n7967, gm_n45);
	nand (gm_n7969, gm_n7968, gm_n71);
	and (gm_n7970, gm_n48, in_11, in_10, gm_n5822, in_13);
	nand (gm_n7971, gm_n46, gm_n63, in_14, gm_n7970, in_17);
	nor (gm_n7972, in_20, in_19, gm_n47, gm_n7971, in_21);
	nand (gm_n7973, gm_n46, gm_n63, in_14, gm_n6005, gm_n81);
	nor (gm_n7974, in_20, gm_n62, gm_n47, gm_n7973, in_21);
	nor (gm_n7975, gm_n48, in_11, gm_n52, gm_n3764, gm_n49);
	nand (gm_n7976, in_16, in_15, in_14, gm_n7975, in_17);
	nor (gm_n7977, in_20, in_19, in_18, gm_n7976, in_21);
	nor (gm_n7978, gm_n63, in_14, gm_n49, gm_n5120, gm_n46);
	nand (gm_n7979, gm_n62, in_18, in_17, gm_n7978, gm_n45);
	nor (gm_n7980, gm_n7979, gm_n71);
	nand (gm_n7981, gm_n48, gm_n53, in_10, gm_n6668, gm_n49);
	nor (gm_n7982, in_16, gm_n63, gm_n50, gm_n7981, in_17);
	nand (gm_n7983, gm_n45, in_19, in_18, gm_n7982, gm_n71);
	nor (gm_n7984, gm_n6479, gm_n51);
	nand (gm_n7985, gm_n48, in_11, in_10, gm_n7984, in_13);
	nor (gm_n7986, in_16, in_15, in_14, gm_n7985, gm_n81);
	nand (gm_n7987, gm_n45, in_19, gm_n47, gm_n7986, in_21);
	nand (gm_n7988, in_12, gm_n53, gm_n52, gm_n2522, gm_n49);
	nor (gm_n7989, gm_n46, gm_n63, gm_n50, gm_n7988, gm_n81);
	nand (gm_n7990, in_20, in_19, gm_n47, gm_n7989, in_21);
	and (gm_n7991, gm_n4484, gm_n52, in_9);
	nand (gm_n7992, in_13, gm_n48, gm_n53, gm_n7991, gm_n50);
	nor (gm_n7993, in_17, in_16, gm_n63, gm_n7992, gm_n47);
	nand (gm_n7994, gm_n71, gm_n45, in_19, gm_n7993);
	and (gm_n7995, in_12, in_11, in_10, gm_n3287, in_13);
	nand (gm_n7996, gm_n46, gm_n63, in_14, gm_n7995, in_17);
	nor (gm_n7997, gm_n45, in_19, gm_n47, gm_n7996, gm_n71);
	nand (gm_n7998, in_11, in_10, in_9, gm_n76);
	nor (gm_n7999, gm_n50, in_13, gm_n48, gm_n7998, gm_n63);
	nand (gm_n8000, in_18, in_17, gm_n46, gm_n7999, in_19);
	nor (gm_n8001, gm_n8000, in_21, in_20);
	or (gm_n8002, in_11, in_10, in_9, gm_n1970, in_12);
	nor (gm_n8003, in_15, in_14, in_13, gm_n8002, in_16);
	nand (gm_n8004, in_19, in_18, gm_n81, gm_n8003, in_20);
	nor (gm_n8005, gm_n8004, in_21);
	and (gm_n8006, in_12, gm_n53, in_10, gm_n339, in_13);
	nand (gm_n8007, in_16, gm_n63, in_14, gm_n8006, in_17);
	nor (gm_n8008, gm_n45, gm_n62, in_18, gm_n8007, in_21);
	or (gm_n8009, in_12, in_11, gm_n52, gm_n7154, in_13);
	nor (gm_n8010, gm_n46, gm_n63, gm_n50, gm_n8009, gm_n81);
	nand (gm_n8011, gm_n45, gm_n62, gm_n47, gm_n8010, gm_n71);
	nor (gm_n8012, gm_n2546, gm_n52, in_9);
	nand (gm_n8013, gm_n49, gm_n48, gm_n53, gm_n8012, gm_n50);
	nor (gm_n8014, in_17, gm_n46, in_15, gm_n8013, gm_n47);
	nand (gm_n8015, gm_n71, in_20, in_19, gm_n8014);
	nor (gm_n8016, gm_n53, gm_n52, gm_n51, gm_n2005, in_12);
	nand (gm_n8017, gm_n63, gm_n50, gm_n49, gm_n8016, gm_n46);
	nor (gm_n8018, gm_n62, in_18, gm_n81, gm_n8017, in_20);
	nand (gm_n8019, gm_n8018, gm_n71);
	nand (gm_n8020, in_12, in_11, in_10, gm_n968, in_13);
	nor (gm_n8021, in_16, in_15, gm_n50, gm_n8020, gm_n81);
	nand (gm_n8022, in_20, gm_n62, in_18, gm_n8021, gm_n71);
	nand (gm_n8023, gm_n81, gm_n46, gm_n63, gm_n2869, gm_n47);
	nor (gm_n8024, in_21, gm_n45, gm_n62, gm_n8023);
	and (gm_n8025, gm_n48, gm_n53, in_10, gm_n912, in_13);
	nand (gm_n8026, in_16, gm_n63, gm_n50, gm_n8025, in_17);
	nor (gm_n8027, in_20, gm_n62, gm_n47, gm_n8026, in_21);
	nand (gm_n8028, in_10, gm_n51, in_8, gm_n302, gm_n53);
	nor (gm_n8029, in_14, in_13, in_12, gm_n8028, in_15);
	nand (gm_n8030, in_18, gm_n81, gm_n46, gm_n8029, in_19);
	nor (gm_n8031, gm_n8030, in_21, gm_n45);
	and (gm_n8032, gm_n49, in_12, in_11, gm_n6769, gm_n50);
	nand (gm_n8033, gm_n81, gm_n46, gm_n63, gm_n8032, gm_n47);
	nor (gm_n8034, gm_n71, gm_n45, in_19, gm_n8033);
	nand (gm_n8035, gm_n50, in_13, gm_n48, gm_n3048, gm_n63);
	nor (gm_n8036, in_18, gm_n81, gm_n46, gm_n8035, gm_n62);
	nand (gm_n8037, gm_n8036, in_21, gm_n45);
	nor (gm_n8038, gm_n2885, in_9);
	nand (gm_n8039, gm_n48, in_11, gm_n52, gm_n8038, gm_n49);
	nor (gm_n8040, in_16, gm_n63, gm_n50, gm_n8039, in_17);
	nand (gm_n8041, gm_n45, in_19, gm_n47, gm_n8040, gm_n71);
	or (gm_n8042, in_13, gm_n48, gm_n53, gm_n1908, in_14);
	nor (gm_n8043, in_17, gm_n46, in_15, gm_n8042, gm_n47);
	nand (gm_n8044, in_21, in_20, gm_n62, gm_n8043);
	nand (gm_n8045, in_12, gm_n53, gm_n52, gm_n3909, gm_n49);
	nor (gm_n8046, in_16, in_15, in_14, gm_n8045, gm_n81);
	nand (gm_n8047, in_20, in_19, in_18, gm_n8046, gm_n71);
	or (gm_n8048, gm_n53, in_10, gm_n51, gm_n955, gm_n48);
	nor (gm_n8049, gm_n63, in_14, gm_n49, gm_n8048, gm_n46);
	nand (gm_n8050, gm_n62, in_18, gm_n81, gm_n8049, in_20);
	nor (gm_n8051, gm_n8050, in_21);
	or (gm_n8052, gm_n53, gm_n52, gm_n51, gm_n1474, in_12);
	nor (gm_n8053, in_15, in_14, gm_n49, gm_n8052, in_16);
	nand (gm_n8054, in_19, in_18, in_17, gm_n8053, gm_n45);
	nor (gm_n8055, gm_n8054, gm_n71);
	nor (gm_n8056, in_12, in_11, in_10, gm_n4294, in_13);
	nand (gm_n8057, in_16, in_15, gm_n50, gm_n8056, in_17);
	nor (gm_n8058, in_20, in_19, gm_n47, gm_n8057, in_21);
	or (gm_n8059, in_11, gm_n52, in_9, gm_n2119, gm_n48);
	nor (gm_n8060, in_15, in_14, gm_n49, gm_n8059, gm_n46);
	nand (gm_n8061, gm_n62, gm_n47, gm_n81, gm_n8060, in_20);
	nor (gm_n8062, gm_n8061, in_21);
	and (gm_n8063, in_7, gm_n82, gm_n72, gm_n420, in_8);
	and (gm_n8064, gm_n53, in_10, in_9, gm_n8063);
	nand (gm_n8065, in_14, in_13, in_12, gm_n8064, gm_n63);
	nor (gm_n8066, gm_n47, in_17, in_16, gm_n8065, gm_n62);
	nand (gm_n8067, gm_n8066, in_21, gm_n45);
	nand (gm_n8068, gm_n48, gm_n53, in_10, gm_n3562, gm_n49);
	nor (gm_n8069, gm_n46, in_15, gm_n50, gm_n8068, gm_n81);
	nand (gm_n8070, in_20, in_19, in_18, gm_n8069, gm_n71);
	and (gm_n8071, gm_n189, gm_n52, in_9);
	nand (gm_n8072, gm_n49, in_12, gm_n53, gm_n8071, gm_n50);
	nor (gm_n8073, in_17, gm_n46, in_15, gm_n8072, gm_n47);
	nand (gm_n8074, gm_n71, in_20, in_19, gm_n8073);
	and (gm_n8075, in_16, gm_n63, gm_n50, gm_n7719, in_17);
	nand (gm_n8076, gm_n45, gm_n62, in_18, gm_n8075, in_21);
	nand (gm_n8077, in_16, in_15, in_14, gm_n4279, gm_n81);
	nor (gm_n8078, gm_n45, in_19, in_18, gm_n8077, in_21);
	nand (gm_n8079, in_17, gm_n46, gm_n63, gm_n2669, in_18);
	nor (gm_n8080, gm_n71, in_20, in_19, gm_n8079);
	or (gm_n8081, gm_n46, gm_n63, in_14, gm_n4537, gm_n81);
	nor (gm_n8082, gm_n45, gm_n62, in_18, gm_n8081, in_21);
	nand (gm_n8083, gm_n46, in_15, gm_n50, gm_n6472, gm_n81);
	nor (gm_n8084, gm_n45, gm_n62, in_18, gm_n8083, gm_n71);
	or (gm_n8085, in_12, in_11, in_10, gm_n5030, gm_n49);
	nor (gm_n8086, in_16, gm_n63, gm_n50, gm_n8085, in_17);
	nand (gm_n8087, in_20, in_19, in_18, gm_n8086, in_21);
	nor (gm_n8088, in_11, gm_n52, in_9, gm_n395, in_12);
	nand (gm_n8089, gm_n63, gm_n50, in_13, gm_n8088, in_16);
	nor (gm_n8090, gm_n62, gm_n47, gm_n81, gm_n8089, gm_n45);
	nand (gm_n8091, gm_n8090, in_21);
	or (gm_n8092, in_13, in_12, in_11, gm_n5052, in_14);
	nor (gm_n8093, in_17, gm_n46, in_15, gm_n8092, gm_n47);
	nand (gm_n8094, gm_n71, in_20, in_19, gm_n8093);
	or (gm_n8095, gm_n53, in_10, in_9, gm_n440);
	or (gm_n8096, gm_n50, gm_n49, in_12, gm_n8095, in_15);
	nor (gm_n8097, gm_n47, gm_n81, in_16, gm_n8096, gm_n62);
	nand (gm_n8098, gm_n8097, in_21, gm_n45);
	nand (gm_n8099, gm_n81, gm_n46, gm_n63, gm_n7824, gm_n47);
	nor (gm_n8100, gm_n71, in_20, gm_n62, gm_n8099);
	nand (gm_n8101, in_11, gm_n52, gm_n51, gm_n2234, gm_n48);
	nor (gm_n8102, in_15, in_14, gm_n49, gm_n8101, in_16);
	nand (gm_n8103, gm_n62, in_18, gm_n81, gm_n8102, in_20);
	nor (gm_n8104, gm_n8103, gm_n71);
	nor (gm_n8105, gm_n520, in_10, gm_n51);
	and (gm_n8106, in_13, gm_n48, gm_n53, gm_n8105, gm_n50);
	nand (gm_n8107, gm_n81, gm_n46, gm_n63, gm_n8106, in_18);
	nor (gm_n8108, gm_n71, gm_n45, gm_n62, gm_n8107);
	nand (gm_n8109, gm_n53, in_10, gm_n51, gm_n1339, gm_n48);
	nor (gm_n8110, gm_n63, in_14, gm_n49, gm_n8109, gm_n46);
	nand (gm_n8111, gm_n62, gm_n47, gm_n81, gm_n8110, in_20);
	nor (gm_n8112, gm_n8111, in_21);
	or (gm_n8113, gm_n53, in_10, in_9, gm_n2345);
	nor (gm_n8114, in_14, gm_n49, gm_n48, gm_n8113, gm_n63);
	and (gm_n8115, in_18, gm_n81, in_16, gm_n8114, gm_n62);
	nand (gm_n8116, gm_n8115, in_21, gm_n45);
	nand (gm_n8117, in_12, gm_n53, gm_n52, gm_n2877, gm_n49);
	nor (gm_n8118, in_16, in_15, gm_n50, gm_n8117, gm_n81);
	nand (gm_n8119, in_20, gm_n62, in_18, gm_n8118, in_21);
	and (gm_n8120, gm_n46, in_15, gm_n50, gm_n5661, in_17);
	nand (gm_n8121, in_20, gm_n62, in_18, gm_n8120, gm_n71);
	or (gm_n8122, in_7, in_6, in_5, gm_n124, gm_n64);
	nor (gm_n8123, in_11, gm_n52, in_9, gm_n8122);
	nand (gm_n8124, in_14, gm_n49, in_12, gm_n8123, in_15);
	nor (gm_n8125, gm_n47, gm_n81, in_16, gm_n8124, in_19);
	nand (gm_n8126, gm_n8125, in_21, in_20);
	nor (gm_n8127, gm_n48, gm_n53, gm_n52, gm_n7853, in_13);
	nand (gm_n8128, in_16, gm_n63, in_14, gm_n8127, gm_n81);
	nor (gm_n8129, in_20, gm_n62, in_18, gm_n8128, gm_n71);
	nor (gm_n8130, in_12, in_11, in_10, gm_n1824, in_13);
	nand (gm_n8131, gm_n46, gm_n63, in_14, gm_n8130, in_17);
	nor (gm_n8132, gm_n45, in_19, gm_n47, gm_n8131, in_21);
	nand (gm_n8133, in_18, in_17, in_16, gm_n5554, in_19);
	nor (gm_n8134, gm_n8133, in_21, gm_n45);
	nor (gm_n8135, in_12, gm_n53, in_10, gm_n347, gm_n49);
	nand (gm_n8136, gm_n46, gm_n63, in_14, gm_n8135, gm_n81);
	nor (gm_n8137, in_20, gm_n62, gm_n47, gm_n8136, gm_n71);
	and (gm_n8138, gm_n53, in_10, gm_n51, gm_n1563);
	nand (gm_n8139, gm_n50, gm_n49, in_12, gm_n8138, gm_n63);
	nor (gm_n8140, in_18, gm_n81, in_16, gm_n8139, gm_n62);
	nand (gm_n8141, gm_n8140, gm_n71, in_20);
	nand (gm_n8142, in_12, in_11, in_10, gm_n6052, gm_n49);
	nor (gm_n8143, gm_n46, in_15, gm_n50, gm_n8142, in_17);
	nand (gm_n8144, in_20, gm_n62, in_18, gm_n8143, gm_n71);
	nand (gm_n8145, gm_n48, gm_n53, gm_n52, gm_n4950, in_13);
	nor (gm_n8146, in_16, gm_n63, in_14, gm_n8145, gm_n81);
	nand (gm_n8147, gm_n45, gm_n62, gm_n47, gm_n8146, in_21);
	nor (gm_n8148, in_11, gm_n52, in_9, gm_n1533, gm_n48);
	nand (gm_n8149, in_15, gm_n50, gm_n49, gm_n8148, gm_n46);
	nor (gm_n8150, in_19, gm_n47, in_17, gm_n8149, gm_n45);
	nand (gm_n8151, gm_n8150, in_21);
	nand (gm_n8152, gm_n51, in_8, in_7, gm_n504, gm_n52);
	nor (gm_n8153, in_13, gm_n48, gm_n53, gm_n8152, in_14);
	nand (gm_n8154, gm_n81, in_16, in_15, gm_n8153, in_18);
	nor (gm_n8155, gm_n71, gm_n45, in_19, gm_n8154);
	nand (gm_n8156, gm_n46, in_15, in_14, gm_n7950, gm_n81);
	nor (gm_n8157, gm_n45, gm_n62, gm_n47, gm_n8156, in_21);
	or (gm_n8158, in_17, in_16, in_15, gm_n3351, gm_n47);
	nor (gm_n8159, gm_n71, gm_n45, in_19, gm_n8158);
	and (gm_n8160, gm_n3316, in_13, gm_n48);
	nand (gm_n8161, in_16, gm_n63, in_14, gm_n8160, in_17);
	nor (gm_n8162, gm_n45, gm_n62, gm_n47, gm_n8161, in_21);
	nor (gm_n8163, gm_n64, in_7, gm_n82, gm_n96, gm_n51);
	nand (gm_n8164, in_12, gm_n53, in_10, gm_n8163, in_13);
	nor (gm_n8165, gm_n46, in_15, gm_n50, gm_n8164, in_17);
	nand (gm_n8166, gm_n45, in_19, gm_n47, gm_n8165, in_21);
	nor (gm_n8167, in_9, in_8, in_7, gm_n279, gm_n52);
	nand (gm_n8168, gm_n49, gm_n48, in_11, gm_n8167, gm_n50);
	nor (gm_n8169, gm_n81, in_16, gm_n63, gm_n8168, gm_n47);
	nand (gm_n8170, in_21, in_20, gm_n62, gm_n8169);
	nand (gm_n8171, in_12, gm_n53, gm_n52, gm_n2641, gm_n49);
	nor (gm_n8172, in_16, in_15, gm_n50, gm_n8171, gm_n81);
	nand (gm_n8173, in_20, in_19, in_18, gm_n8172, gm_n71);
	nor (gm_n8174, in_11, in_10, gm_n51, gm_n1393, in_12);
	nand (gm_n8175, gm_n63, in_14, in_13, gm_n8174, in_16);
	nor (gm_n8176, in_19, in_18, gm_n81, gm_n8175, in_20);
	nand (gm_n8177, gm_n8176, in_21);
	or (gm_n8178, in_16, in_15, gm_n50, gm_n4965, gm_n81);
	nor (gm_n8179, in_20, in_19, gm_n47, gm_n8178, in_21);
	nand (gm_n8180, in_10, in_9, in_8, gm_n691, in_11);
	nor (gm_n8181, gm_n50, gm_n49, gm_n48, gm_n8180, in_15);
	nand (gm_n8182, gm_n47, in_17, gm_n46, gm_n8181, gm_n62);
	nor (gm_n8183, gm_n8182, in_21, in_20);
	nor (gm_n8184, in_12, gm_n53, gm_n52, gm_n2280, in_13);
	nand (gm_n8185, gm_n46, in_15, gm_n50, gm_n8184, gm_n81);
	nor (gm_n8186, in_20, in_19, gm_n47, gm_n8185, gm_n71);
	nand (gm_n8187, gm_n53, in_10, gm_n51, gm_n4618, gm_n48);
	nor (gm_n8188, gm_n63, gm_n50, in_13, gm_n8187, gm_n46);
	nand (gm_n8189, gm_n62, gm_n47, in_17, gm_n8188, in_20);
	nor (gm_n8190, gm_n8189, in_21);
	nand (gm_n8191, in_12, in_11, in_10, gm_n1759, gm_n49);
	nor (gm_n8192, in_16, gm_n63, gm_n50, gm_n8191, gm_n81);
	nand (gm_n8193, in_20, in_19, in_18, gm_n8192, gm_n71);
	and (gm_n8194, gm_n4723, in_9);
	nand (gm_n8195, gm_n48, in_11, gm_n52, gm_n8194, in_13);
	nor (gm_n8196, in_16, in_15, in_14, gm_n8195, in_17);
	nand (gm_n8197, in_20, gm_n62, in_18, gm_n8196, in_21);
	nor (gm_n8198, gm_n48, gm_n53, gm_n52, gm_n1723, in_13);
	and (gm_n8199, in_16, in_15, gm_n50, gm_n8198, gm_n81);
	nand (gm_n8200, gm_n45, in_19, gm_n47, gm_n8199, in_21);
	or (gm_n8201, gm_n48, gm_n53, gm_n52, gm_n264, in_13);
	nor (gm_n8202, in_16, in_15, gm_n50, gm_n8201, gm_n81);
	nand (gm_n8203, gm_n45, gm_n62, gm_n47, gm_n8202, gm_n71);
	nor (gm_n8204, gm_n48, gm_n53, in_10, gm_n6518, in_13);
	nand (gm_n8205, in_16, in_15, gm_n50, gm_n8204, in_17);
	nor (gm_n8206, in_20, gm_n62, gm_n47, gm_n8205, in_21);
	nand (gm_n8207, in_16, gm_n63, in_14, gm_n4881, gm_n81);
	nor (gm_n8208, in_20, gm_n62, gm_n47, gm_n8207, in_21);
	and (gm_n8209, gm_n63, in_14, gm_n49, gm_n7634, gm_n46);
	nand (gm_n8210, gm_n62, in_18, in_17, gm_n8209, in_20);
	nor (gm_n8211, gm_n8210, in_21);
	and (gm_n8212, in_12, in_11, gm_n52, gm_n2729, in_13);
	nand (gm_n8213, in_16, gm_n63, gm_n50, gm_n8212, gm_n81);
	nor (gm_n8214, gm_n45, in_19, gm_n47, gm_n8213, in_21);
	nand (gm_n8215, gm_n3845, gm_n49);
	nor (gm_n8216, gm_n46, gm_n63, in_14, gm_n8215, gm_n81);
	nand (gm_n8217, gm_n45, in_19, in_18, gm_n8216, gm_n71);
	nand (gm_n8218, gm_n50, in_13, in_12, gm_n3577, in_15);
	nor (gm_n8219, gm_n47, gm_n81, gm_n46, gm_n8218, gm_n62);
	nand (gm_n8220, gm_n8219, gm_n71, gm_n45);
	nand (gm_n8221, gm_n49, gm_n48, in_11, gm_n3262, gm_n50);
	nor (gm_n8222, gm_n81, in_16, gm_n63, gm_n8221, gm_n47);
	nand (gm_n8223, in_21, in_20, in_19, gm_n8222);
	nand (gm_n8224, in_7, in_6, gm_n72, gm_n327, in_8);
	nor (gm_n8225, gm_n53, in_10, gm_n51, gm_n8224, in_12);
	nand (gm_n8226, in_15, gm_n50, gm_n49, gm_n8225, in_16);
	nor (gm_n8227, gm_n62, in_18, gm_n81, gm_n8226, gm_n45);
	nand (gm_n8228, gm_n8227, in_21);
	nor (gm_n8229, gm_n48, in_11, in_10, gm_n5768, gm_n49);
	nand (gm_n8230, in_16, in_15, in_14, gm_n8229, gm_n81);
	nor (gm_n8231, gm_n45, in_19, in_18, gm_n8230, gm_n71);
	nor (gm_n8232, in_11, in_10, gm_n51, gm_n328, gm_n48);
	and (gm_n8233, in_15, in_14, gm_n49, gm_n8232, gm_n46);
	nand (gm_n8234, in_19, in_18, gm_n81, gm_n8233, in_20);
	nor (gm_n8235, gm_n8234, gm_n71);
	nand (gm_n8236, in_16, in_15, in_14, gm_n6622, in_17);
	nor (gm_n8237, gm_n45, gm_n62, in_18, gm_n8236, in_21);
	nand (gm_n8238, in_16, in_15, gm_n50, gm_n1249, in_17);
	nor (gm_n8239, in_20, in_19, gm_n47, gm_n8238, in_21);
	nand (gm_n8240, in_14, gm_n49, in_12, gm_n4051, in_15);
	nor (gm_n8241, gm_n47, in_17, in_16, gm_n8240, in_19);
	nand (gm_n8242, gm_n8241, gm_n71, gm_n45);
	nor (gm_n8243, in_9, gm_n64, in_7, gm_n588, gm_n52);
	nand (gm_n8244, gm_n49, gm_n48, in_11, gm_n8243, gm_n50);
	nor (gm_n8245, gm_n81, gm_n46, in_15, gm_n8244, in_18);
	nand (gm_n8246, in_21, gm_n45, in_19, gm_n8245);
	or (gm_n8247, gm_n48, gm_n53, gm_n52, gm_n4692, in_13);
	nor (gm_n8248, gm_n46, gm_n63, gm_n50, gm_n8247, in_17);
	nand (gm_n8249, in_20, gm_n62, in_18, gm_n8248, in_21);
	or (gm_n8250, in_13, in_12, gm_n53, gm_n4432, gm_n50);
	nor (gm_n8251, in_17, gm_n46, in_15, gm_n8250, gm_n47);
	nand (gm_n8252, in_21, in_20, in_19, gm_n8251);
	nor (gm_n8253, gm_n49, in_12, in_11, gm_n859, in_14);
	nand (gm_n8254, gm_n81, in_16, in_15, gm_n8253, gm_n47);
	nor (gm_n8255, gm_n71, in_20, in_19, gm_n8254);
	nor (gm_n8256, in_8, gm_n55, gm_n82, gm_n141, gm_n51);
	and (gm_n8257, gm_n48, gm_n53, gm_n52, gm_n8256, in_13);
	nand (gm_n8258, gm_n46, gm_n63, in_14, gm_n8257, gm_n81);
	nor (gm_n8259, in_20, in_19, gm_n47, gm_n8258, in_21);
	or (gm_n8260, in_11, gm_n52, in_9, gm_n6155, in_12);
	nor (gm_n8261, in_15, in_14, gm_n49, gm_n8260, gm_n46);
	nand (gm_n8262, gm_n62, gm_n47, in_17, gm_n8261, in_20);
	nor (gm_n8263, gm_n8262, gm_n71);
	nor (gm_n8264, gm_n50, in_13, gm_n48, gm_n2998, gm_n63);
	nand (gm_n8265, gm_n47, gm_n81, in_16, gm_n8264, gm_n62);
	nor (gm_n8266, gm_n8265, in_21, in_20);
	nand (gm_n8267, gm_n48, gm_n53, in_10, gm_n2415, gm_n49);
	nor (gm_n8268, in_16, gm_n63, gm_n50, gm_n8267, in_17);
	nand (gm_n8269, in_20, gm_n62, in_18, gm_n8268, in_21);
	or (gm_n8270, in_12, gm_n53, gm_n52, gm_n1174, gm_n49);
	nor (gm_n8271, in_16, in_15, gm_n50, gm_n8270, gm_n81);
	nand (gm_n8272, in_20, gm_n62, gm_n47, gm_n8271, in_21);
	nand (gm_n8273, in_12, in_11, in_10, gm_n7231, in_13);
	nor (gm_n8274, gm_n46, in_15, gm_n50, gm_n8273, gm_n81);
	nand (gm_n8275, gm_n45, in_19, gm_n47, gm_n8274, gm_n71);
	or (gm_n8276, gm_n583, in_10, gm_n51);
	nor (gm_n8277, gm_n49, in_12, in_11, gm_n8276);
	and (gm_n8278, gm_n46, in_15, in_14, gm_n8277, gm_n81);
	nand (gm_n8279, gm_n45, gm_n62, in_18, gm_n8278, gm_n71);
	nand (gm_n8280, in_11, gm_n52, in_9, gm_n1634, in_12);
	nor (gm_n8281, gm_n63, gm_n50, in_13, gm_n8280, gm_n46);
	nand (gm_n8282, in_19, in_18, gm_n81, gm_n8281, in_20);
	nor (gm_n8283, gm_n8282, in_21);
	and (gm_n8284, gm_n50, gm_n49, gm_n48, gm_n4936, in_15);
	nand (gm_n8285, gm_n47, gm_n81, gm_n46, gm_n8284, in_19);
	nor (gm_n8286, gm_n8285, in_21, in_20);
	nor (gm_n8287, gm_n49, in_12, in_11, gm_n2006, in_14);
	nand (gm_n8288, in_17, gm_n46, gm_n63, gm_n8287, gm_n47);
	nor (gm_n8289, gm_n71, gm_n45, in_19, gm_n8288);
	nor (gm_n8290, gm_n52, gm_n51, in_8, gm_n390, in_11);
	and (gm_n8291, gm_n50, gm_n49, in_12, gm_n8290, gm_n63);
	nand (gm_n8292, in_18, gm_n81, gm_n46, gm_n8291, in_19);
	nor (gm_n8293, gm_n8292, in_21, gm_n45);
	or (gm_n8294, gm_n63, gm_n50, gm_n49, gm_n734, gm_n46);
	nor (gm_n8295, gm_n62, gm_n47, gm_n81, gm_n8294, gm_n45);
	nand (gm_n8296, gm_n8295, in_21);
	nand (gm_n8297, gm_n48, gm_n53, in_10, gm_n280, in_13);
	nor (gm_n8298, gm_n46, in_15, gm_n50, gm_n8297, gm_n81);
	nand (gm_n8299, in_20, in_19, gm_n47, gm_n8298, gm_n71);
	nor (gm_n8300, gm_n46, in_15, gm_n50, gm_n4940, gm_n81);
	nand (gm_n8301, in_20, in_19, gm_n47, gm_n8300, gm_n71);
	nand (gm_n8302, in_12, in_11, gm_n52, gm_n5375, gm_n49);
	nor (gm_n8303, gm_n46, in_15, in_14, gm_n8302, in_17);
	nand (gm_n8304, in_20, gm_n62, in_18, gm_n8303, in_21);
	nor (gm_n8305, gm_n48, in_11, in_10, gm_n1252, gm_n49);
	nand (gm_n8306, gm_n46, in_15, in_14, gm_n8305, gm_n81);
	nor (gm_n8307, gm_n45, in_19, in_18, gm_n8306, gm_n71);
	and (gm_n8308, gm_n48, in_11, gm_n52, gm_n1941, in_13);
	nand (gm_n8309, gm_n46, gm_n63, in_14, gm_n8308, gm_n81);
	nor (gm_n8310, in_20, gm_n62, gm_n47, gm_n8309, gm_n71);
	nor (gm_n8311, gm_n2559, in_10, in_9);
	and (gm_n8312, in_13, in_12, gm_n53, gm_n8311, in_14);
	nand (gm_n8313, in_17, gm_n46, gm_n63, gm_n8312, in_18);
	nor (gm_n8314, gm_n71, gm_n45, in_19, gm_n8313);
	nand (gm_n8315, gm_n52, gm_n51, gm_n64, gm_n338, gm_n53);
	nor (gm_n8316, in_14, in_13, in_12, gm_n8315, in_15);
	nand (gm_n8317, in_18, in_17, in_16, gm_n8316, gm_n62);
	nor (gm_n8318, gm_n8317, in_21, gm_n45);
	or (gm_n8319, in_12, gm_n53, in_10, gm_n1617, in_13);
	nor (gm_n8320, gm_n46, in_15, in_14, gm_n8319, gm_n81);
	nand (gm_n8321, gm_n45, gm_n62, in_18, gm_n8320, gm_n71);
	nand (gm_n8322, gm_n48, gm_n53, in_10, gm_n4072, in_13);
	nor (gm_n8323, gm_n46, in_15, gm_n50, gm_n8322, in_17);
	nand (gm_n8324, gm_n45, gm_n62, in_18, gm_n8323, gm_n71);
	nand (gm_n8325, in_12, in_11, gm_n52, gm_n6139, gm_n49);
	nor (gm_n8326, in_16, gm_n63, gm_n50, gm_n8325, gm_n81);
	nand (gm_n8327, in_20, in_19, in_18, gm_n8326, gm_n71);
	and (gm_n8328, gm_n7107, gm_n49, gm_n48);
	and (gm_n8329, gm_n46, in_15, in_14, gm_n8328, in_17);
	nand (gm_n8330, gm_n45, in_19, gm_n47, gm_n8329, gm_n71);
	nor (gm_n8331, in_12, in_11, in_10, gm_n7068, gm_n49);
	nand (gm_n8332, in_16, gm_n63, gm_n50, gm_n8331, gm_n81);
	nor (gm_n8333, in_20, in_19, gm_n47, gm_n8332, in_21);
	nand (gm_n8334, gm_n53, in_10, gm_n51, gm_n297, gm_n48);
	nor (gm_n8335, gm_n63, gm_n50, in_13, gm_n8334, gm_n46);
	nand (gm_n8336, gm_n62, in_18, in_17, gm_n8335, gm_n45);
	nor (gm_n8337, gm_n8336, in_21);
	nand (gm_n8338, in_11, in_10, in_9, gm_n3519, gm_n48);
	nor (gm_n8339, gm_n63, gm_n50, in_13, gm_n8338, gm_n46);
	nand (gm_n8340, gm_n62, gm_n47, in_17, gm_n8339, gm_n45);
	nor (gm_n8341, gm_n8340, gm_n71);
	nand (gm_n8342, in_11, in_10, in_9, gm_n3086, gm_n48);
	nor (gm_n8343, in_15, gm_n50, gm_n49, gm_n8342, in_16);
	nand (gm_n8344, in_19, gm_n47, gm_n81, gm_n8343, gm_n45);
	nor (gm_n8345, gm_n8344, gm_n71);
	nor (gm_n8346, gm_n46, in_15, gm_n50, gm_n1466, in_17);
	nand (gm_n8347, gm_n45, gm_n62, gm_n47, gm_n8346, in_21);
	nand (gm_n8348, in_12, gm_n53, in_10, gm_n2749, gm_n49);
	nor (gm_n8349, in_16, gm_n63, gm_n50, gm_n8348, in_17);
	nand (gm_n8350, gm_n45, in_19, in_18, gm_n8349, gm_n71);
	nor (gm_n8351, gm_n53, in_10, gm_n51, gm_n368, gm_n48);
	nand (gm_n8352, in_15, gm_n50, gm_n49, gm_n8351, in_16);
	nor (gm_n8353, gm_n62, gm_n47, gm_n81, gm_n8352, in_20);
	nand (gm_n8354, gm_n8353, gm_n71);
	nor (gm_n8355, in_11, in_10, gm_n51, gm_n2564, gm_n48);
	nand (gm_n8356, in_15, gm_n50, in_13, gm_n8355, in_16);
	nor (gm_n8357, gm_n62, in_18, in_17, gm_n8356, in_20);
	nand (gm_n8358, gm_n8357, in_21);
	nor (gm_n8359, in_12, in_11, gm_n52, gm_n5620, in_13);
	nand (gm_n8360, in_16, gm_n63, gm_n50, gm_n8359, in_17);
	nor (gm_n8361, gm_n45, in_19, gm_n47, gm_n8360, in_21);
	nor (gm_n8362, gm_n49, gm_n48, gm_n53, gm_n4351, in_14);
	nand (gm_n8363, gm_n81, gm_n46, in_15, gm_n8362, in_18);
	nor (gm_n8364, in_21, in_20, gm_n62, gm_n8363);
	nor (gm_n8365, gm_n63, in_14, gm_n49, gm_n2689, in_16);
	nand (gm_n8366, in_19, gm_n47, gm_n81, gm_n8365, in_20);
	nor (gm_n8367, gm_n8366, gm_n71);
	or (gm_n8368, gm_n64, in_7, gm_n82, gm_n119, gm_n51);
	nor (gm_n8369, in_12, gm_n53, gm_n52, gm_n8368, in_13);
	nand (gm_n8370, in_16, in_15, in_14, gm_n8369, in_17);
	nor (gm_n8371, gm_n45, gm_n62, in_18, gm_n8370, gm_n71);
	nand (gm_n8372, gm_n48, gm_n53, in_10, gm_n2729, in_13);
	nor (gm_n8373, gm_n46, gm_n63, in_14, gm_n8372, gm_n81);
	nand (gm_n8374, in_20, in_19, in_18, gm_n8373, gm_n71);
	nor (gm_n8375, gm_n53, gm_n52, gm_n51, gm_n4562, gm_n48);
	nand (gm_n8376, gm_n63, gm_n50, gm_n49, gm_n8375, in_16);
	nor (gm_n8377, in_19, in_18, in_17, gm_n8376, gm_n45);
	nand (gm_n8378, gm_n8377, in_21);
	nand (gm_n8379, gm_n50, gm_n49, in_12, gm_n6961, in_15);
	nor (gm_n8380, gm_n47, gm_n81, gm_n46, gm_n8379, gm_n62);
	nand (gm_n8381, gm_n8380, in_21, in_20);
	or (gm_n8382, in_13, in_12, gm_n53, gm_n1920, gm_n50);
	nor (gm_n8383, gm_n81, in_16, gm_n63, gm_n8382, in_18);
	nand (gm_n8384, in_21, gm_n45, gm_n62, gm_n8383);
	or (gm_n8385, in_11, gm_n52, gm_n51, gm_n2077, in_12);
	nor (gm_n8386, in_15, gm_n50, gm_n49, gm_n8385, gm_n46);
	nand (gm_n8387, in_19, gm_n47, gm_n81, gm_n8386, in_20);
	nor (gm_n8388, gm_n8387, in_21);
	nand (gm_n8389, gm_n46, gm_n63, gm_n50, gm_n6081, gm_n81);
	nor (gm_n8390, in_20, gm_n62, in_18, gm_n8389, in_21);
	nor (gm_n8391, gm_n48, gm_n53, in_10, gm_n2623, in_13);
	nand (gm_n8392, in_16, in_15, gm_n50, gm_n8391, in_17);
	nor (gm_n8393, in_20, in_19, in_18, gm_n8392, in_21);
	nor (gm_n8394, gm_n49, in_12, in_11, gm_n2225, gm_n50);
	nand (gm_n8395, gm_n81, in_16, in_15, gm_n8394, in_18);
	nor (gm_n8396, gm_n71, gm_n45, gm_n62, gm_n8395);
	and (gm_n8397, in_11, gm_n52, in_9, gm_n1142, gm_n48);
	nand (gm_n8398, in_15, in_14, gm_n49, gm_n8397, in_16);
	nor (gm_n8399, in_19, gm_n47, in_17, gm_n8398, in_20);
	nand (gm_n8400, gm_n8399, in_21);
	nor (gm_n8401, in_11, gm_n52, gm_n51, gm_n2836, in_12);
	nand (gm_n8402, in_15, in_14, gm_n49, gm_n8401, in_16);
	nor (gm_n8403, in_19, in_18, in_17, gm_n8402, in_20);
	nand (gm_n8404, gm_n8403, gm_n71);
	nor (gm_n8405, gm_n53, gm_n52, gm_n51, gm_n1879, gm_n48);
	nand (gm_n8406, gm_n63, gm_n50, gm_n49, gm_n8405, gm_n46);
	nor (gm_n8407, in_19, in_18, in_17, gm_n8406, gm_n45);
	nand (gm_n8408, gm_n8407, in_21);
	and (gm_n8409, gm_n52, in_9, in_8, gm_n431, gm_n53);
	nand (gm_n8410, gm_n50, in_13, gm_n48, gm_n8409, gm_n63);
	nor (gm_n8411, in_18, gm_n81, gm_n46, gm_n8410, in_19);
	nand (gm_n8412, gm_n8411, in_21, gm_n45);
	nand (gm_n8413, gm_n50, in_13, gm_n48, gm_n7857, in_15);
	nor (gm_n8414, in_18, in_17, in_16, gm_n8413, gm_n62);
	nand (gm_n8415, gm_n8414, gm_n71, in_20);
	nand (gm_n8416, gm_n8408, gm_n8404, gm_n8400, gm_n8415, gm_n8412);
	nor (gm_n8417, gm_n8393, gm_n8390, gm_n8388, gm_n8416, gm_n8396);
	nand (gm_n8418, gm_n8381, gm_n8378, gm_n8374, gm_n8417, gm_n8384);
	nor (gm_n8419, gm_n8367, gm_n8364, gm_n8361, gm_n8418, gm_n8371);
	nand (gm_n8420, gm_n8354, gm_n8350, gm_n8347, gm_n8419, gm_n8358);
	nor (gm_n8421, gm_n8341, gm_n8337, gm_n8333, gm_n8420, gm_n8345);
	nand (gm_n8422, gm_n8327, gm_n8324, gm_n8321, gm_n8421, gm_n8330);
	nor (gm_n8423, gm_n8314, gm_n8310, gm_n8307, gm_n8422, gm_n8318);
	nand (gm_n8424, gm_n8301, gm_n8299, gm_n8296, gm_n8423, gm_n8304);
	nor (gm_n8425, gm_n8289, gm_n8286, gm_n8283, gm_n8424, gm_n8293);
	nand (gm_n8426, gm_n8275, gm_n8272, gm_n8269, gm_n8425, gm_n8279);
	nor (gm_n8427, gm_n8263, gm_n8259, gm_n8255, gm_n8426, gm_n8266);
	nand (gm_n8428, gm_n8249, gm_n8246, gm_n8242, gm_n8427, gm_n8252);
	nor (gm_n8429, gm_n8237, gm_n8235, gm_n8231, gm_n8428, gm_n8239);
	nand (gm_n8430, gm_n8223, gm_n8220, gm_n8217, gm_n8429, gm_n8228);
	nor (gm_n8431, gm_n8211, gm_n8208, gm_n8206, gm_n8430, gm_n8214);
	nand (gm_n8432, gm_n8200, gm_n8197, gm_n8193, gm_n8431, gm_n8203);
	nor (gm_n8433, gm_n8186, gm_n8183, gm_n8179, gm_n8432, gm_n8190);
	nand (gm_n8434, gm_n8173, gm_n8170, gm_n8166, gm_n8433, gm_n8177);
	nor (gm_n8435, gm_n8159, gm_n8157, gm_n8155, gm_n8434, gm_n8162);
	nand (gm_n8436, gm_n8147, gm_n8144, gm_n8141, gm_n8435, gm_n8151);
	nor (gm_n8437, gm_n8134, gm_n8132, gm_n8129, gm_n8436, gm_n8137);
	nand (gm_n8438, gm_n8121, gm_n8119, gm_n8116, gm_n8437, gm_n8126);
	nor (gm_n8439, gm_n8108, gm_n8104, gm_n8100, gm_n8438, gm_n8112);
	nand (gm_n8440, gm_n8094, gm_n8091, gm_n8087, gm_n8439, gm_n8098);
	nor (gm_n8441, gm_n8082, gm_n8080, gm_n8078, gm_n8440, gm_n8084);
	nand (gm_n8442, gm_n8074, gm_n8070, gm_n8067, gm_n8441, gm_n8076);
	nor (gm_n8443, gm_n8058, gm_n8055, gm_n8051, gm_n8442, gm_n8062);
	nand (gm_n8444, gm_n8044, gm_n8041, gm_n8037, gm_n8443, gm_n8047);
	nor (gm_n8445, gm_n8031, gm_n8027, gm_n8024, gm_n8444, gm_n8034);
	nand (gm_n8446, gm_n8019, gm_n8015, gm_n8011, gm_n8445, gm_n8022);
	nor (gm_n8447, gm_n8005, gm_n8001, gm_n7997, gm_n8446, gm_n8008);
	nand (gm_n8448, gm_n7990, gm_n7987, gm_n7983, gm_n8447, gm_n7994);
	nor (gm_n8449, gm_n7977, gm_n7974, gm_n7972, gm_n8448, gm_n7980);
	nand (gm_n8450, gm_n7965, gm_n7962, gm_n7959, gm_n8449, gm_n7969);
	nor (gm_n8451, gm_n7952, gm_n7949, gm_n7945, gm_n8450, gm_n7956);
	nand (gm_n8452, gm_n7938, gm_n7935, gm_n7932, gm_n8451, gm_n7942);
	nor (out_13, gm_n8452, gm_n7928);
	nor (gm_n8454, gm_n48, in_11, gm_n52, gm_n4104, gm_n49);
	nand (gm_n8455, in_16, in_15, gm_n50, gm_n8454, in_17);
	nor (gm_n8456, gm_n45, gm_n62, in_18, gm_n8455, in_21);
	nor (gm_n8457, in_16, gm_n63, gm_n50, gm_n7644, gm_n81);
	nand (gm_n8458, in_20, in_19, gm_n47, gm_n8457, gm_n71);
	nand (gm_n8459, gm_n49, in_12, in_11, gm_n436, gm_n50);
	nor (gm_n8460, gm_n81, in_16, in_15, gm_n8459, gm_n47);
	nand (gm_n8461, gm_n71, in_20, in_19, gm_n8460);
	nand (gm_n8462, in_12, gm_n53, gm_n52, gm_n2284, gm_n49);
	nor (gm_n8463, gm_n46, in_15, gm_n50, gm_n8462, in_17);
	nand (gm_n8464, in_20, gm_n62, in_18, gm_n8463, in_21);
	nand (gm_n8465, in_14, gm_n49, in_12, gm_n2019, gm_n63);
	nor (gm_n8466, in_18, in_17, gm_n46, gm_n8465, in_19);
	nand (gm_n8467, gm_n8466, gm_n71, gm_n45);
	nand (gm_n8468, in_16, gm_n63, gm_n50, gm_n8198, in_17);
	nor (gm_n8469, in_20, gm_n62, in_18, gm_n8468, in_21);
	and (gm_n8470, gm_n48, in_11, in_10, gm_n912, in_13);
	nand (gm_n8471, in_16, in_15, in_14, gm_n8470, in_17);
	nor (gm_n8472, gm_n45, in_19, in_18, gm_n8471, gm_n71);
	nand (gm_n8473, gm_n53, in_10, in_9, gm_n3214, gm_n48);
	nor (gm_n8474, gm_n63, in_14, in_13, gm_n8473, in_16);
	nand (gm_n8475, in_19, gm_n47, gm_n81, gm_n8474, gm_n45);
	nor (gm_n8476, gm_n8475, in_21);
	and (gm_n8477, gm_n50, in_13, in_12, gm_n2654, in_15);
	nand (gm_n8478, gm_n47, in_17, in_16, gm_n8477, in_19);
	nor (gm_n8479, gm_n8478, in_21, in_20);
	nand (gm_n8480, gm_n48, gm_n53, gm_n52, gm_n946, gm_n49);
	nor (gm_n8481, in_16, gm_n63, in_14, gm_n8480, gm_n81);
	nand (gm_n8482, in_20, gm_n62, in_18, gm_n8481, in_21);
	nand (gm_n8483, gm_n63, gm_n50, in_13, gm_n7813, gm_n46);
	nor (gm_n8484, gm_n62, in_18, in_17, gm_n8483, gm_n45);
	nand (gm_n8485, gm_n8484, gm_n71);
	and (gm_n8486, in_18, in_17, gm_n46, gm_n3093, in_19);
	nand (gm_n8487, gm_n8486, in_21, gm_n45);
	nand (gm_n8488, in_13, in_12, in_11, gm_n4922, in_14);
	nor (gm_n8489, gm_n81, in_16, gm_n63, gm_n8488, gm_n47);
	nand (gm_n8490, in_21, gm_n45, in_19, gm_n8489);
	nand (gm_n8491, in_10, gm_n51, in_8, gm_n1088, gm_n53);
	nor (gm_n8492, gm_n50, gm_n49, gm_n48, gm_n8491, in_15);
	nand (gm_n8493, in_18, gm_n81, in_16, gm_n8492, gm_n62);
	nor (gm_n8494, gm_n8493, in_21, in_20);
	nor (gm_n8495, gm_n53, gm_n52, in_9, gm_n1434);
	and (gm_n8496, in_14, gm_n49, in_12, gm_n8495, gm_n63);
	nand (gm_n8497, gm_n47, in_17, gm_n46, gm_n8496, in_19);
	nor (gm_n8498, gm_n8497, in_21, gm_n45);
	and (gm_n8499, in_12, gm_n53, gm_n52, gm_n3354, gm_n49);
	nand (gm_n8500, gm_n46, in_15, in_14, gm_n8499, in_17);
	nor (gm_n8501, in_20, gm_n62, gm_n47, gm_n8500, gm_n71);
	nor (gm_n8502, in_12, gm_n53, gm_n52, gm_n758, gm_n49);
	nand (gm_n8503, gm_n46, in_15, in_14, gm_n8502, gm_n81);
	nor (gm_n8504, gm_n45, gm_n62, in_18, gm_n8503, gm_n71);
	nor (gm_n8505, in_8, gm_n55, gm_n82, gm_n103, gm_n51);
	nand (gm_n8506, gm_n48, in_11, in_10, gm_n8505, gm_n49);
	nor (gm_n8507, in_16, gm_n63, gm_n50, gm_n8506, gm_n81);
	nand (gm_n8508, in_20, gm_n62, in_18, gm_n8507, gm_n71);
	nand (gm_n8509, in_13, in_12, in_11, gm_n3708, in_14);
	nor (gm_n8510, gm_n81, in_16, gm_n63, gm_n8509, in_18);
	nand (gm_n8511, in_21, in_20, gm_n62, gm_n8510);
	nand (gm_n8512, gm_n53, gm_n52, in_9, gm_n3091, in_12);
	nor (gm_n8513, gm_n8512, in_13);
	and (gm_n8514, gm_n46, gm_n63, in_14, gm_n8513, gm_n81);
	nand (gm_n8515, gm_n45, in_19, in_18, gm_n8514, in_21);
	nor (gm_n8516, in_11, in_10, in_9, gm_n774);
	nand (gm_n8517, in_14, gm_n49, in_12, gm_n8516, gm_n63);
	nor (gm_n8518, in_18, in_17, gm_n46, gm_n8517, gm_n62);
	nand (gm_n8519, gm_n8518, in_21, gm_n45);
	nor (gm_n8520, gm_n48, in_11, in_10, gm_n8368, in_13);
	nand (gm_n8521, in_16, in_15, in_14, gm_n8520, gm_n81);
	nor (gm_n8522, in_20, gm_n62, gm_n47, gm_n8521, in_21);
	and (gm_n8523, in_12, in_11, gm_n52, gm_n6331, gm_n49);
	nand (gm_n8524, in_16, in_15, in_14, gm_n8523, in_17);
	nor (gm_n8525, gm_n45, gm_n62, in_18, gm_n8524, gm_n71);
	and (gm_n8526, in_13, in_12, in_11, gm_n7193, in_14);
	nand (gm_n8527, in_17, gm_n46, in_15, gm_n8526, gm_n47);
	nor (gm_n8528, in_21, in_20, gm_n62, gm_n8527);
	and (gm_n8529, in_12, in_11, in_10, gm_n2284, in_13);
	nand (gm_n8530, gm_n46, gm_n63, gm_n50, gm_n8529, gm_n81);
	nor (gm_n8531, gm_n45, gm_n62, in_18, gm_n8530, gm_n71);
	and (gm_n8532, gm_n47, gm_n81, gm_n46, gm_n1149, in_19);
	nand (gm_n8533, gm_n8532, gm_n71, in_20);
	nand (gm_n8534, gm_n49, gm_n48, in_11, gm_n1652, in_14);
	nor (gm_n8535, in_17, in_16, gm_n63, gm_n8534, gm_n47);
	nand (gm_n8536, gm_n71, gm_n45, gm_n62, gm_n8535);
	and (gm_n8537, gm_n53, gm_n52, in_9, gm_n1936);
	nand (gm_n8538, in_14, in_13, in_12, gm_n8537, in_15);
	nor (gm_n8539, gm_n47, gm_n81, in_16, gm_n8538, gm_n62);
	nand (gm_n8540, gm_n8539, gm_n71, gm_n45);
	and (gm_n8541, in_16, in_15, in_14, gm_n7682, gm_n81);
	nand (gm_n8542, in_20, in_19, gm_n47, gm_n8541, in_21);
	nand (gm_n8543, in_11, in_10, in_9, gm_n1302, gm_n48);
	nor (gm_n8544, gm_n63, gm_n50, in_13, gm_n8543, gm_n46);
	nand (gm_n8545, in_19, gm_n47, gm_n81, gm_n8544, in_20);
	nor (gm_n8546, gm_n8545, gm_n71);
	nand (gm_n8547, in_11, gm_n52, in_9, gm_n4388, in_12);
	nor (gm_n8548, in_15, gm_n50, in_13, gm_n8547, in_16);
	nand (gm_n8549, gm_n62, in_18, in_17, gm_n8548, in_20);
	nor (gm_n8550, gm_n8549, gm_n71);
	and (gm_n8551, in_12, in_11, gm_n52, gm_n4072, in_13);
	nand (gm_n8552, gm_n46, in_15, in_14, gm_n8551, gm_n81);
	nor (gm_n8553, in_20, in_19, in_18, gm_n8552, gm_n71);
	nand (gm_n8554, gm_n46, in_15, gm_n50, gm_n670, in_17);
	nor (gm_n8555, gm_n45, in_19, in_18, gm_n8554, gm_n71);
	nand (gm_n8556, in_12, gm_n53, in_10, gm_n343, in_13);
	nor (gm_n8557, in_16, gm_n63, gm_n50, gm_n8556, in_17);
	nand (gm_n8558, gm_n45, in_19, gm_n47, gm_n8557, gm_n71);
	nand (gm_n8559, in_15, gm_n50, gm_n49, gm_n4436, in_16);
	nor (gm_n8560, gm_n62, in_18, gm_n81, gm_n8559, gm_n45);
	nand (gm_n8561, gm_n8560, gm_n71);
	nor (gm_n8562, gm_n53, gm_n52, in_9, gm_n8122, in_12);
	nand (gm_n8563, in_15, gm_n50, in_13, gm_n8562, in_16);
	nor (gm_n8564, gm_n62, in_18, in_17, gm_n8563, gm_n45);
	nand (gm_n8565, gm_n8564, gm_n71);
	nor (gm_n8566, gm_n53, gm_n52, in_9, gm_n2926, gm_n48);
	nand (gm_n8567, in_15, in_14, in_13, gm_n8566, gm_n46);
	nor (gm_n8568, in_19, gm_n47, in_17, gm_n8567, in_20);
	nand (gm_n8569, gm_n8568, gm_n71);
	nor (gm_n8570, gm_n783, gm_n51);
	and (gm_n8571, gm_n48, in_11, gm_n52, gm_n8570, gm_n49);
	nand (gm_n8572, in_16, gm_n63, gm_n50, gm_n8571, gm_n81);
	nor (gm_n8573, gm_n45, in_19, in_18, gm_n8572, gm_n71);
	and (gm_n8574, in_12, gm_n53, gm_n52, gm_n2097, gm_n49);
	nand (gm_n8575, gm_n46, gm_n63, gm_n50, gm_n8574, in_17);
	nor (gm_n8576, in_20, gm_n62, gm_n47, gm_n8575, gm_n71);
	and (gm_n8577, in_12, in_11, gm_n52, gm_n7115, in_13);
	nand (gm_n8578, in_16, in_15, gm_n50, gm_n8577, in_17);
	nor (gm_n8579, in_20, gm_n62, gm_n47, gm_n8578, gm_n71);
	nor (gm_n8580, gm_n48, gm_n53, in_10, gm_n2355, in_13);
	nand (gm_n8581, in_16, gm_n63, in_14, gm_n8580, in_17);
	nor (gm_n8582, in_20, gm_n62, gm_n47, gm_n8581, in_21);
	nor (gm_n8583, gm_n53, gm_n52, gm_n51, gm_n3557, gm_n48);
	nand (gm_n8584, gm_n63, gm_n50, in_13, gm_n8583, in_16);
	nor (gm_n8585, gm_n62, gm_n47, in_17, gm_n8584, gm_n45);
	nand (gm_n8586, gm_n8585, in_21);
	nand (gm_n8587, in_13, gm_n48, gm_n53, gm_n4027, gm_n50);
	nor (gm_n8588, in_17, gm_n46, gm_n63, gm_n8587, in_18);
	nand (gm_n8589, in_21, gm_n45, in_19, gm_n8588);
	nand (gm_n8590, in_14, gm_n49, in_12, gm_n3295, gm_n63);
	nor (gm_n8591, in_18, gm_n81, gm_n46, gm_n8590, in_19);
	nand (gm_n8592, gm_n8591, gm_n71, in_20);
	or (gm_n8593, gm_n48, in_11, gm_n52, gm_n2841, in_13);
	nor (gm_n8594, gm_n46, gm_n63, gm_n50, gm_n8593, gm_n81);
	nand (gm_n8595, in_20, in_19, in_18, gm_n8594, gm_n71);
	nor (gm_n8596, gm_n48, in_11, in_10, gm_n639, gm_n49);
	nand (gm_n8597, in_16, gm_n63, gm_n50, gm_n8596, in_17);
	nor (gm_n8598, in_20, in_19, in_18, gm_n8597, in_21);
	and (gm_n8599, in_14, in_13, gm_n48, gm_n6240, gm_n63);
	nand (gm_n8600, gm_n47, gm_n81, in_16, gm_n8599, in_19);
	nor (gm_n8601, gm_n8600, gm_n71, in_20);
	nand (gm_n8602, gm_n53, gm_n52, in_9, gm_n1147, gm_n48);
	nor (gm_n8603, in_15, gm_n50, in_13, gm_n8602, in_16);
	nand (gm_n8604, in_19, in_18, in_17, gm_n8603, gm_n45);
	nor (gm_n8605, gm_n8604, in_21);
	nand (gm_n8606, gm_n53, gm_n52, in_9, gm_n1339, gm_n48);
	nor (gm_n8607, in_15, in_14, gm_n49, gm_n8606, in_16);
	nand (gm_n8608, gm_n62, gm_n47, in_17, gm_n8607, in_20);
	nor (gm_n8609, gm_n8608, gm_n71);
	nor (gm_n8610, gm_n51, gm_n64, gm_n55, gm_n1256, gm_n52);
	nand (gm_n8611, gm_n49, in_12, gm_n53, gm_n8610, in_14);
	nor (gm_n8612, in_17, in_16, in_15, gm_n8611, gm_n47);
	nand (gm_n8613, gm_n71, in_20, gm_n62, gm_n8612);
	nand (gm_n8614, gm_n49, in_12, in_11, gm_n5133, in_14);
	nor (gm_n8615, gm_n81, gm_n46, in_15, gm_n8614, gm_n47);
	nand (gm_n8616, in_21, in_20, in_19, gm_n8615);
	or (gm_n8617, in_12, gm_n53, in_10, gm_n104, in_13);
	nor (gm_n8618, in_16, in_15, gm_n50, gm_n8617, gm_n81);
	nand (gm_n8619, in_20, gm_n62, gm_n47, gm_n8618, gm_n71);
	and (gm_n8620, gm_n46, in_15, gm_n50, gm_n4144, gm_n81);
	nand (gm_n8621, gm_n45, in_19, gm_n47, gm_n8620, in_21);
	nand (gm_n8622, in_11, gm_n52, gm_n51, gm_n1339, in_12);
	nor (gm_n8623, gm_n63, in_14, gm_n49, gm_n8622, in_16);
	nand (gm_n8624, gm_n62, gm_n47, gm_n81, gm_n8623, in_20);
	nor (gm_n8625, gm_n8624, in_21);
	and (gm_n8626, gm_n63, gm_n50, gm_n49, gm_n7739, in_16);
	nand (gm_n8627, in_19, gm_n47, gm_n81, gm_n8626, in_20);
	nor (gm_n8628, gm_n8627, in_21);
	nor (gm_n8629, in_8, in_7, gm_n82, gm_n530, in_9);
	and (gm_n8630, gm_n48, gm_n53, in_10, gm_n8629, in_13);
	nand (gm_n8631, in_16, in_15, in_14, gm_n8630, gm_n81);
	nor (gm_n8632, in_20, in_19, gm_n47, gm_n8631, in_21);
	nand (gm_n8633, gm_n53, gm_n52, in_9, gm_n4388);
	nor (gm_n8634, gm_n50, gm_n49, gm_n48, gm_n8633, gm_n63);
	nand (gm_n8635, gm_n47, gm_n81, in_16, gm_n8634, in_19);
	nor (gm_n8636, gm_n8635, gm_n71, gm_n45);
	and (gm_n8637, gm_n53, gm_n52, in_9, gm_n3451);
	nand (gm_n8638, in_14, gm_n49, gm_n48, gm_n8637, in_15);
	nor (gm_n8639, gm_n47, in_17, gm_n46, gm_n8638, gm_n62);
	nand (gm_n8640, gm_n8639, in_21, gm_n45);
	nor (gm_n8641, gm_n52, gm_n51, in_8, gm_n2239, gm_n53);
	nand (gm_n8642, gm_n50, gm_n49, in_12, gm_n8641, gm_n63);
	nor (gm_n8643, gm_n47, gm_n81, gm_n46, gm_n8642, gm_n62);
	nand (gm_n8644, gm_n8643, in_21, gm_n45);
	nand (gm_n8645, in_13, gm_n48, in_11, gm_n5133, gm_n50);
	nor (gm_n8646, gm_n81, gm_n46, gm_n63, gm_n8645, in_18);
	nand (gm_n8647, in_21, gm_n45, in_19, gm_n8646);
	nand (gm_n8648, gm_n49, gm_n48, gm_n53, gm_n4872, in_14);
	nor (gm_n8649, in_17, in_16, gm_n63, gm_n8648, gm_n47);
	nand (gm_n8650, in_21, gm_n45, gm_n62, gm_n8649);
	nor (gm_n8651, in_11, gm_n52, in_9, gm_n5586);
	and (gm_n8652, gm_n50, in_13, in_12, gm_n8651, in_15);
	nand (gm_n8653, gm_n47, in_17, in_16, gm_n8652, in_19);
	nor (gm_n8654, gm_n8653, in_21, in_20);
	nor (gm_n8655, in_14, gm_n49, in_12, gm_n8633, in_15);
	nand (gm_n8656, gm_n47, gm_n81, in_16, gm_n8655, gm_n62);
	nor (gm_n8657, gm_n8656, in_21, gm_n45);
	and (gm_n8658, in_13, gm_n48, gm_n53, gm_n5003, in_14);
	nand (gm_n8659, gm_n81, gm_n46, gm_n63, gm_n8658, gm_n47);
	nor (gm_n8660, in_21, in_20, gm_n62, gm_n8659);
	and (gm_n8661, in_13, gm_n48, in_11, gm_n1958, gm_n50);
	nand (gm_n8662, gm_n81, gm_n46, gm_n63, gm_n8661, in_18);
	nor (gm_n8663, gm_n71, in_20, in_19, gm_n8662);
	and (gm_n8664, gm_n48, in_11, gm_n52, gm_n4418, in_13);
	and (gm_n8665, gm_n46, in_15, in_14, gm_n8664, in_17);
	nand (gm_n8666, gm_n45, gm_n62, in_18, gm_n8665, gm_n71);
	nand (gm_n8667, gm_n49, gm_n48, gm_n53, gm_n137, gm_n50);
	nor (gm_n8668, in_17, gm_n46, in_15, gm_n8667, in_18);
	nand (gm_n8669, gm_n71, gm_n45, gm_n62, gm_n8668);
	nand (gm_n8670, gm_n50, gm_n49, in_12, gm_n7925, in_15);
	nor (gm_n8671, gm_n47, gm_n81, in_16, gm_n8670, in_19);
	nand (gm_n8672, gm_n8671, gm_n71, gm_n45);
	nand (gm_n8673, in_15, in_14, in_13, gm_n5476, gm_n46);
	nor (gm_n8674, gm_n62, gm_n47, in_17, gm_n8673, gm_n45);
	nand (gm_n8675, gm_n8674, gm_n71);
	nor (gm_n8676, gm_n1750, gm_n52, in_9);
	and (gm_n8677, in_13, gm_n48, in_11, gm_n8676, in_14);
	nand (gm_n8678, in_17, gm_n46, in_15, gm_n8677, in_18);
	nor (gm_n8679, in_21, in_20, gm_n62, gm_n8678);
	and (gm_n8680, gm_n50, gm_n49, in_12, gm_n5587, gm_n63);
	nand (gm_n8681, gm_n47, in_17, in_16, gm_n8680, gm_n62);
	nor (gm_n8682, gm_n8681, gm_n71, in_20);
	nor (gm_n8683, gm_n55, in_6, gm_n72, gm_n124, in_8);
	nand (gm_n8684, gm_n53, in_10, in_9, gm_n8683, in_12);
	nor (gm_n8685, in_15, gm_n50, in_13, gm_n8684, in_16);
	nand (gm_n8686, gm_n62, in_18, gm_n81, gm_n8685, in_20);
	nor (gm_n8687, gm_n8686, in_21);
	nor (gm_n8688, gm_n48, gm_n53, in_10, gm_n2052, gm_n49);
	nand (gm_n8689, in_16, gm_n63, in_14, gm_n8688, gm_n81);
	nor (gm_n8690, gm_n45, gm_n62, gm_n47, gm_n8689, in_21);
	and (gm_n8691, gm_n53, in_10, gm_n51, gm_n5422, in_12);
	nand (gm_n8692, in_15, in_14, gm_n49, gm_n8691, in_16);
	nor (gm_n8693, gm_n62, in_18, in_17, gm_n8692, in_20);
	nand (gm_n8694, gm_n8693, gm_n71);
	nor (gm_n8695, gm_n51, gm_n64, in_7, gm_n259, in_10);
	nand (gm_n8696, gm_n49, in_12, in_11, gm_n8695, gm_n50);
	nor (gm_n8697, in_17, gm_n46, gm_n63, gm_n8696, in_18);
	nand (gm_n8698, in_21, gm_n45, in_19, gm_n8697);
	nand (gm_n8699, in_14, gm_n49, gm_n48, gm_n4802, gm_n63);
	nor (gm_n8700, gm_n47, in_17, in_16, gm_n8699, gm_n62);
	nand (gm_n8701, gm_n8700, in_21, gm_n45);
	nor (gm_n8702, in_10, in_9, in_8, gm_n468, in_11);
	nand (gm_n8703, in_14, gm_n49, gm_n48, gm_n8702, gm_n63);
	nor (gm_n8704, gm_n47, in_17, in_16, gm_n8703, in_19);
	nand (gm_n8705, gm_n8704, gm_n71, in_20);
	nand (gm_n8706, in_17, gm_n46, gm_n63, gm_n5042, in_18);
	nor (gm_n8707, gm_n71, in_20, in_19, gm_n8706);
	or (gm_n8708, gm_n53, gm_n52, gm_n51, gm_n2546, gm_n48);
	nor (gm_n8709, gm_n8708, gm_n50, in_13);
	nand (gm_n8710, in_17, gm_n46, in_15, gm_n8709, in_18);
	nor (gm_n8711, gm_n71, in_20, gm_n62, gm_n8710);
	nand (gm_n8712, in_16, in_15, gm_n50, gm_n3495, gm_n81);
	nor (gm_n8713, gm_n45, in_19, in_18, gm_n8712, in_21);
	nor (gm_n8714, gm_n48, in_11, gm_n52, gm_n4262, gm_n49);
	nand (gm_n8715, in_16, in_15, gm_n50, gm_n8714, gm_n81);
	nor (gm_n8716, in_20, gm_n62, in_18, gm_n8715, in_21);
	nand (gm_n8717, gm_n48, gm_n53, in_10, gm_n2235, in_13);
	nor (gm_n8718, in_16, in_15, in_14, gm_n8717, gm_n81);
	nand (gm_n8719, in_20, gm_n62, gm_n47, gm_n8718, gm_n71);
	nand (gm_n8720, in_13, in_12, gm_n53, gm_n224, gm_n50);
	nor (gm_n8721, gm_n81, in_16, in_15, gm_n8720, in_18);
	nand (gm_n8722, gm_n71, gm_n45, in_19, gm_n8721);
	nand (gm_n8723, gm_n48, in_11, gm_n52, gm_n7176, gm_n49);
	nor (gm_n8724, gm_n46, gm_n63, in_14, gm_n8723, gm_n81);
	nand (gm_n8725, gm_n45, in_19, in_18, gm_n8724, gm_n71);
	nand (gm_n8726, gm_n48, in_11, in_10, gm_n2890, in_13);
	nor (gm_n8727, gm_n46, in_15, in_14, gm_n8726, in_17);
	nand (gm_n8728, in_20, in_19, in_18, gm_n8727, in_21);
	and (gm_n8729, gm_n48, gm_n53, in_10, gm_n2760, gm_n49);
	nand (gm_n8730, in_16, gm_n63, gm_n50, gm_n8729, gm_n81);
	nor (gm_n8731, gm_n45, gm_n62, gm_n47, gm_n8730, in_21);
	nor (gm_n8732, in_11, in_10, gm_n51, gm_n3257);
	and (gm_n8733, gm_n50, in_13, in_12, gm_n8732, gm_n63);
	nand (gm_n8734, in_18, in_17, gm_n46, gm_n8733, gm_n62);
	nor (gm_n8735, gm_n8734, in_21, in_20);
	and (gm_n8736, gm_n6679, gm_n50, gm_n49);
	nand (gm_n8737, gm_n81, gm_n46, in_15, gm_n8736, in_18);
	nor (gm_n8738, in_21, gm_n45, in_19, gm_n8737);
	and (gm_n8739, in_14, gm_n49, gm_n48, gm_n6943, in_15);
	nand (gm_n8740, gm_n47, gm_n81, gm_n46, gm_n8739, gm_n62);
	nor (gm_n8741, gm_n8740, gm_n71, in_20);
	or (gm_n8742, gm_n48, gm_n53, gm_n52, gm_n7227, in_13);
	nor (gm_n8743, in_16, in_15, gm_n50, gm_n8742, gm_n81);
	nand (gm_n8744, gm_n45, in_19, gm_n47, gm_n8743, gm_n71);
	nand (gm_n8745, gm_n48, in_11, in_10, gm_n268, gm_n49);
	nor (gm_n8746, in_16, gm_n63, gm_n50, gm_n8745, in_17);
	nand (gm_n8747, gm_n45, gm_n62, in_18, gm_n8746, in_21);
	nand (gm_n8748, gm_n63, gm_n50, gm_n49, gm_n1248, in_16);
	nor (gm_n8749, in_19, gm_n47, gm_n81, gm_n8748, gm_n45);
	nand (gm_n8750, gm_n8749, gm_n71);
	nand (gm_n8751, gm_n48, gm_n53, gm_n52, gm_n617, gm_n49);
	nor (gm_n8752, in_16, in_15, in_14, gm_n8751, gm_n81);
	nand (gm_n8753, gm_n45, in_19, gm_n47, gm_n8752, gm_n71);
	and (gm_n8754, in_14, gm_n49, in_12, gm_n6409, in_15);
	nand (gm_n8755, gm_n47, gm_n81, in_16, gm_n8754, gm_n62);
	nor (gm_n8756, gm_n8755, in_21, in_20);
	nor (gm_n8757, in_12, in_11, gm_n52, gm_n7092, in_13);
	nand (gm_n8758, gm_n46, gm_n63, gm_n50, gm_n8757, gm_n81);
	nor (gm_n8759, in_20, in_19, gm_n47, gm_n8758, gm_n71);
	nor (gm_n8760, in_13, in_12, in_11, gm_n1024, gm_n50);
	nand (gm_n8761, gm_n81, in_16, in_15, gm_n8760, gm_n47);
	nor (gm_n8762, in_21, in_20, gm_n62, gm_n8761);
	and (gm_n8763, gm_n49, gm_n48, gm_n53, gm_n3916, in_14);
	nand (gm_n8764, gm_n81, gm_n46, in_15, gm_n8763, gm_n47);
	nor (gm_n8765, gm_n71, in_20, in_19, gm_n8764);
	nor (gm_n8766, in_16, gm_n63, in_14, gm_n5506, gm_n81);
	nand (gm_n8767, gm_n45, in_19, in_18, gm_n8766, gm_n71);
	nor (gm_n8768, gm_n46, gm_n63, in_14, gm_n8068, in_17);
	nand (gm_n8769, gm_n45, in_19, in_18, gm_n8768, in_21);
	nand (gm_n8770, in_14, gm_n49, gm_n48, gm_n2420, gm_n63);
	nor (gm_n8771, in_18, in_17, in_16, gm_n8770, gm_n62);
	nand (gm_n8772, gm_n8771, gm_n71, in_20);
	nand (gm_n8773, gm_n49, gm_n48, gm_n53, gm_n3480, gm_n50);
	nor (gm_n8774, in_17, in_16, gm_n63, gm_n8773, gm_n47);
	nand (gm_n8775, gm_n71, in_20, in_19, gm_n8774);
	nand (gm_n8776, in_11, in_10, gm_n51, gm_n3768, in_12);
	nor (gm_n8777, gm_n63, gm_n50, gm_n49, gm_n8776, in_16);
	nand (gm_n8778, in_19, in_18, gm_n81, gm_n8777, in_20);
	nor (gm_n8779, gm_n8778, in_21);
	and (gm_n8780, in_12, in_11, in_10, gm_n146, gm_n49);
	nand (gm_n8781, gm_n46, in_15, in_14, gm_n8780, in_17);
	nor (gm_n8782, gm_n45, gm_n62, gm_n47, gm_n8781, in_21);
	and (gm_n8783, gm_n48, gm_n53, in_10, gm_n747, in_13);
	nand (gm_n8784, in_16, in_15, gm_n50, gm_n8783, gm_n81);
	nor (gm_n8785, in_20, gm_n62, gm_n47, gm_n8784, gm_n71);
	and (gm_n8786, gm_n51, in_8, in_7, gm_n404);
	and (gm_n8787, in_12, in_11, in_10, gm_n8786, gm_n49);
	nand (gm_n8788, in_16, gm_n63, gm_n50, gm_n8787, gm_n81);
	nor (gm_n8789, gm_n45, gm_n62, gm_n47, gm_n8788, gm_n71);
	nand (gm_n8790, gm_n55, gm_n82, gm_n72, gm_n209, gm_n64);
	nor (gm_n8791, gm_n53, gm_n52, gm_n51, gm_n8790, in_12);
	nand (gm_n8792, gm_n63, gm_n50, in_13, gm_n8791, gm_n46);
	nor (gm_n8793, gm_n62, gm_n47, in_17, gm_n8792, in_20);
	nand (gm_n8794, gm_n8793, gm_n71);
	nor (gm_n8795, in_16, in_15, gm_n50, gm_n6130, in_17);
	nand (gm_n8796, in_20, in_19, in_18, gm_n8795, in_21);
	nand (gm_n8797, in_12, gm_n53, gm_n52, gm_n3268, in_13);
	nor (gm_n8798, in_16, gm_n63, gm_n50, gm_n8797, gm_n81);
	nand (gm_n8799, in_20, in_19, in_18, gm_n8798, gm_n71);
	nand (gm_n8800, gm_n48, in_11, gm_n52, gm_n2819, in_13);
	nor (gm_n8801, gm_n46, gm_n63, in_14, gm_n8800, gm_n81);
	nand (gm_n8802, gm_n45, in_19, gm_n47, gm_n8801, in_21);
	and (gm_n8803, in_13, in_12, in_11, gm_n8610, in_14);
	nand (gm_n8804, in_17, gm_n46, in_15, gm_n8803, in_18);
	nor (gm_n8805, gm_n71, gm_n45, in_19, gm_n8804);
	and (gm_n8806, in_15, in_14, in_13, gm_n1635, gm_n46);
	nand (gm_n8807, gm_n62, in_18, gm_n81, gm_n8806, in_20);
	nor (gm_n8808, gm_n8807, in_21);
	nor (gm_n8809, in_10, in_9, gm_n64, gm_n853);
	and (gm_n8810, gm_n49, in_12, gm_n53, gm_n8809, in_14);
	nand (gm_n8811, gm_n81, in_16, gm_n63, gm_n8810, in_18);
	nor (gm_n8812, in_21, in_20, in_19, gm_n8811);
	and (gm_n8813, in_14, in_13, gm_n48, gm_n2366, gm_n63);
	nand (gm_n8814, in_18, in_17, in_16, gm_n8813, in_19);
	nor (gm_n8815, gm_n8814, in_21, gm_n45);
	nand (gm_n8816, in_12, gm_n53, gm_n52, gm_n7186, in_13);
	nor (gm_n8817, in_16, in_15, in_14, gm_n8816, in_17);
	nand (gm_n8818, in_20, in_19, gm_n47, gm_n8817, gm_n71);
	nand (gm_n8819, in_12, gm_n53, gm_n52, gm_n1982, gm_n49);
	nor (gm_n8820, in_16, gm_n63, gm_n50, gm_n8819, gm_n81);
	nand (gm_n8821, gm_n45, in_19, gm_n47, gm_n8820, gm_n71);
	nand (gm_n8822, in_12, gm_n53, in_10, gm_n2067, gm_n49);
	nor (gm_n8823, in_16, gm_n63, gm_n50, gm_n8822, gm_n81);
	nand (gm_n8824, in_20, in_19, gm_n47, gm_n8823, in_21);
	nand (gm_n8825, gm_n50, in_13, gm_n48, gm_n1223, gm_n63);
	nor (gm_n8826, gm_n47, in_17, in_16, gm_n8825, gm_n62);
	nand (gm_n8827, gm_n8826, gm_n71, gm_n45);
	nor (gm_n8828, gm_n50, gm_n49, in_12, gm_n5826, gm_n63);
	nand (gm_n8829, gm_n47, gm_n81, in_16, gm_n8828, gm_n62);
	nor (gm_n8830, gm_n8829, gm_n71, in_20);
	and (gm_n8831, gm_n48, in_11, in_10, gm_n2685, gm_n49);
	nand (gm_n8832, in_16, in_15, gm_n50, gm_n8831, gm_n81);
	nor (gm_n8833, gm_n45, gm_n62, gm_n47, gm_n8832, gm_n71);
	nand (gm_n8834, in_16, in_15, gm_n50, gm_n3111, gm_n81);
	nor (gm_n8835, gm_n45, in_19, in_18, gm_n8834, in_21);
	nand (gm_n8836, gm_n52, in_9, in_8, gm_n338, gm_n53);
	nor (gm_n8837, in_14, gm_n49, gm_n48, gm_n8836, in_15);
	nand (gm_n8838, in_18, in_17, in_16, gm_n8837, in_19);
	nor (gm_n8839, gm_n8838, gm_n71, in_20);
	nor (gm_n8840, in_18, gm_n81, in_16, gm_n3486, in_19);
	nand (gm_n8841, gm_n8840, in_21, in_20);
	nand (gm_n8842, gm_n48, in_11, gm_n52, gm_n268, gm_n49);
	nor (gm_n8843, gm_n46, gm_n63, in_14, gm_n8842, in_17);
	nand (gm_n8844, in_20, in_19, in_18, gm_n8843, in_21);
	nand (gm_n8845, in_14, gm_n49, gm_n48, gm_n549, in_15);
	nor (gm_n8846, in_18, gm_n81, in_16, gm_n8845, gm_n62);
	nand (gm_n8847, gm_n8846, in_21, gm_n45);
	nand (gm_n8848, gm_n49, gm_n48, in_11, gm_n594, in_14);
	nor (gm_n8849, in_17, in_16, in_15, gm_n8848, in_18);
	nand (gm_n8850, in_21, gm_n45, in_19, gm_n8849);
	and (gm_n8851, gm_n50, in_13, gm_n48, gm_n3456, gm_n63);
	nand (gm_n8852, in_18, gm_n81, in_16, gm_n8851, gm_n62);
	nor (gm_n8853, gm_n8852, gm_n71, in_20);
	and (gm_n8854, gm_n51, gm_n64, gm_n55, gm_n66, gm_n52);
	and (gm_n8855, gm_n49, in_12, gm_n53, gm_n8854, in_14);
	nand (gm_n8856, gm_n81, in_16, in_15, gm_n8855, in_18);
	nor (gm_n8857, in_21, in_20, gm_n62, gm_n8856);
	and (gm_n8858, in_12, gm_n53, in_10, gm_n2729, in_13);
	nand (gm_n8859, gm_n46, gm_n63, in_14, gm_n8858, gm_n81);
	nor (gm_n8860, gm_n45, gm_n62, in_18, gm_n8859, in_21);
	and (gm_n8861, gm_n50, in_13, gm_n48, gm_n5210, in_15);
	nand (gm_n8862, in_18, gm_n81, gm_n46, gm_n8861, gm_n62);
	nor (gm_n8863, gm_n8862, gm_n71, in_20);
	nand (gm_n8864, in_13, in_12, gm_n53, gm_n2120, gm_n50);
	nor (gm_n8865, gm_n81, gm_n46, in_15, gm_n8864, gm_n47);
	nand (gm_n8866, gm_n71, in_20, gm_n62, gm_n8865);
	nand (gm_n8867, in_14, in_13, in_12, gm_n2538, gm_n63);
	nor (gm_n8868, gm_n47, gm_n81, gm_n46, gm_n8867, in_19);
	nand (gm_n8869, gm_n8868, gm_n71, in_20);
	nor (gm_n8870, gm_n2503, gm_n52, gm_n51);
	nand (gm_n8871, gm_n49, gm_n48, in_11, gm_n8870, gm_n50);
	nor (gm_n8872, in_17, in_16, gm_n63, gm_n8871, gm_n47);
	nand (gm_n8873, gm_n71, gm_n45, gm_n62, gm_n8872);
	nand (gm_n8874, in_14, gm_n49, gm_n48, gm_n1188, in_15);
	nor (gm_n8875, gm_n47, in_17, gm_n46, gm_n8874, gm_n62);
	nand (gm_n8876, gm_n8875, in_21, gm_n45);
	or (gm_n8877, gm_n53, in_10, gm_n51, gm_n8790, gm_n48);
	nor (gm_n8878, gm_n8877, in_14, in_13);
	nand (gm_n8879, gm_n81, gm_n46, in_15, gm_n8878, in_18);
	nor (gm_n8880, gm_n71, gm_n45, gm_n62, gm_n8879);
	and (gm_n8881, gm_n5185, gm_n52, gm_n51);
	and (gm_n8882, in_13, in_12, in_11, gm_n8881, in_14);
	nand (gm_n8883, in_17, gm_n46, gm_n63, gm_n8882, in_18);
	nor (gm_n8884, in_21, in_20, gm_n62, gm_n8883);
	nor (gm_n8885, in_12, gm_n53, in_10, gm_n6056, in_13);
	nand (gm_n8886, gm_n46, in_15, gm_n50, gm_n8885, in_17);
	nor (gm_n8887, gm_n45, gm_n62, gm_n47, gm_n8886, in_21);
	nor (gm_n8888, gm_n48, gm_n53, in_10, gm_n5605, in_13);
	nand (gm_n8889, in_16, in_15, in_14, gm_n8888, in_17);
	nor (gm_n8890, in_20, gm_n62, gm_n47, gm_n8889, in_21);
	nand (gm_n8891, gm_n48, in_11, gm_n52, gm_n5138, gm_n49);
	nor (gm_n8892, in_16, gm_n63, gm_n50, gm_n8891, gm_n81);
	nand (gm_n8893, in_20, in_19, gm_n47, gm_n8892, gm_n71);
	nor (gm_n8894, gm_n46, in_15, gm_n50, gm_n6015, gm_n81);
	nand (gm_n8895, in_20, in_19, gm_n47, gm_n8894, gm_n71);
	nand (gm_n8896, gm_n53, in_10, gm_n51, gm_n2229, in_12);
	or (gm_n8897, gm_n63, in_14, gm_n49, gm_n8896, gm_n46);
	nor (gm_n8898, gm_n62, in_18, in_17, gm_n8897, gm_n45);
	nand (gm_n8899, gm_n8898, gm_n71);
	nand (gm_n8900, in_12, in_11, gm_n52, gm_n3039, in_13);
	nor (gm_n8901, gm_n46, gm_n63, gm_n50, gm_n8900, in_17);
	nand (gm_n8902, gm_n45, gm_n62, gm_n47, gm_n8901, gm_n71);
	nand (gm_n8903, in_11, in_10, in_9, gm_n1147, gm_n48);
	nor (gm_n8904, in_15, gm_n50, gm_n49, gm_n8903, in_16);
	nand (gm_n8905, gm_n62, in_18, gm_n81, gm_n8904, gm_n45);
	nor (gm_n8906, gm_n8905, in_21);
	nor (gm_n8907, in_15, gm_n50, in_13, gm_n2994, in_16);
	nand (gm_n8908, in_19, in_18, gm_n81, gm_n8907, gm_n45);
	nor (gm_n8909, gm_n8908, gm_n71);
	and (gm_n8910, gm_n48, gm_n53, in_10, gm_n2984, in_13);
	nand (gm_n8911, in_16, in_15, in_14, gm_n8910, gm_n81);
	nor (gm_n8912, gm_n45, gm_n62, gm_n47, gm_n8911, in_21);
	nor (gm_n8913, in_12, gm_n53, gm_n52, gm_n1744, gm_n49);
	nand (gm_n8914, gm_n46, in_15, in_14, gm_n8913, gm_n81);
	nor (gm_n8915, gm_n45, gm_n62, in_18, gm_n8914, in_21);
	nor (gm_n8916, gm_n62, in_18, gm_n81, gm_n522, gm_n45);
	nand (gm_n8917, gm_n8916, in_21);
	nand (gm_n8918, in_13, gm_n48, in_11, gm_n6568, gm_n50);
	nor (gm_n8919, gm_n81, gm_n46, gm_n63, gm_n8918, in_18);
	nand (gm_n8920, gm_n71, gm_n45, in_19, gm_n8919);
	nand (gm_n8921, gm_n50, gm_n49, in_12, gm_n3078, in_15);
	nor (gm_n8922, gm_n47, in_17, gm_n46, gm_n8921, in_19);
	nand (gm_n8923, gm_n8922, in_21, in_20);
	and (gm_n8924, in_11, gm_n52, gm_n51, gm_n3183, in_12);
	nand (gm_n8925, gm_n63, in_14, gm_n49, gm_n8924, in_16);
	nor (gm_n8926, gm_n62, gm_n47, gm_n81, gm_n8925, gm_n45);
	nand (gm_n8927, gm_n8926, gm_n71);
	nor (gm_n8928, in_10, in_9, gm_n64, gm_n390, gm_n53);
	nand (gm_n8929, in_14, in_13, gm_n48, gm_n8928, in_15);
	nor (gm_n8930, in_18, in_17, in_16, gm_n8929, in_19);
	nand (gm_n8931, gm_n8930, in_21, gm_n45);
	nand (gm_n8932, gm_n8923, gm_n8920, gm_n8917, gm_n8931, gm_n8927);
	nor (gm_n8933, gm_n8912, gm_n8909, gm_n8906, gm_n8932, gm_n8915);
	nand (gm_n8934, gm_n8899, gm_n8895, gm_n8893, gm_n8933, gm_n8902);
	nor (gm_n8935, gm_n8887, gm_n8884, gm_n8880, gm_n8934, gm_n8890);
	nand (gm_n8936, gm_n8873, gm_n8869, gm_n8866, gm_n8935, gm_n8876);
	nor (gm_n8937, gm_n8860, gm_n8857, gm_n8853, gm_n8936, gm_n8863);
	nand (gm_n8938, gm_n8847, gm_n8844, gm_n8841, gm_n8937, gm_n8850);
	nor (gm_n8939, gm_n8835, gm_n8833, gm_n8830, gm_n8938, gm_n8839);
	nand (gm_n8940, gm_n8824, gm_n8821, gm_n8818, gm_n8939, gm_n8827);
	nor (gm_n8941, gm_n8812, gm_n8808, gm_n8805, gm_n8940, gm_n8815);
	nand (gm_n8942, gm_n8799, gm_n8796, gm_n8794, gm_n8941, gm_n8802);
	nor (gm_n8943, gm_n8785, gm_n8782, gm_n8779, gm_n8942, gm_n8789);
	nand (gm_n8944, gm_n8772, gm_n8769, gm_n8767, gm_n8943, gm_n8775);
	nor (gm_n8945, gm_n8762, gm_n8759, gm_n8756, gm_n8944, gm_n8765);
	nand (gm_n8946, gm_n8750, gm_n8747, gm_n8744, gm_n8945, gm_n8753);
	nor (gm_n8947, gm_n8738, gm_n8735, gm_n8731, gm_n8946, gm_n8741);
	nand (gm_n8948, gm_n8725, gm_n8722, gm_n8719, gm_n8947, gm_n8728);
	nor (gm_n8949, gm_n8713, gm_n8711, gm_n8707, gm_n8948, gm_n8716);
	nand (gm_n8950, gm_n8701, gm_n8698, gm_n8694, gm_n8949, gm_n8705);
	nor (gm_n8951, gm_n8687, gm_n8682, gm_n8679, gm_n8950, gm_n8690);
	nand (gm_n8952, gm_n8672, gm_n8669, gm_n8666, gm_n8951, gm_n8675);
	nor (gm_n8953, gm_n8660, gm_n8657, gm_n8654, gm_n8952, gm_n8663);
	nand (gm_n8954, gm_n8647, gm_n8644, gm_n8640, gm_n8953, gm_n8650);
	nor (gm_n8955, gm_n8632, gm_n8628, gm_n8625, gm_n8954, gm_n8636);
	nand (gm_n8956, gm_n8619, gm_n8616, gm_n8613, gm_n8955, gm_n8621);
	nor (gm_n8957, gm_n8605, gm_n8601, gm_n8598, gm_n8956, gm_n8609);
	nand (gm_n8958, gm_n8592, gm_n8589, gm_n8586, gm_n8957, gm_n8595);
	nor (gm_n8959, gm_n8579, gm_n8576, gm_n8573, gm_n8958, gm_n8582);
	nand (gm_n8960, gm_n8565, gm_n8561, gm_n8558, gm_n8959, gm_n8569);
	nor (gm_n8961, gm_n8553, gm_n8550, gm_n8546, gm_n8960, gm_n8555);
	nand (gm_n8962, gm_n8540, gm_n8536, gm_n8533, gm_n8961, gm_n8542);
	nor (gm_n8963, gm_n8528, gm_n8525, gm_n8522, gm_n8962, gm_n8531);
	nand (gm_n8964, gm_n8515, gm_n8511, gm_n8508, gm_n8963, gm_n8519);
	nor (gm_n8965, gm_n8501, gm_n8498, gm_n8494, gm_n8964, gm_n8504);
	nand (gm_n8966, gm_n8487, gm_n8485, gm_n8482, gm_n8965, gm_n8490);
	nor (gm_n8967, gm_n8476, gm_n8472, gm_n8469, gm_n8966, gm_n8479);
	nand (gm_n8968, gm_n8464, gm_n8461, gm_n8458, gm_n8967, gm_n8467);
	nor (out_14, gm_n8968, gm_n8456);
	nor (gm_n8970, in_12, in_11, in_10, gm_n233, in_13);
	nand (gm_n8971, in_16, in_15, in_14, gm_n8970, in_17);
	nor (gm_n8972, in_20, gm_n62, in_18, gm_n8971, gm_n71);
	nand (gm_n8973, gm_n50, in_13, gm_n48, gm_n8495, in_15);
	nor (gm_n8974, gm_n47, in_17, in_16, gm_n8973, in_19);
	nand (gm_n8975, gm_n8974, gm_n71, in_20);
	nor (gm_n8976, in_10, in_9, gm_n64, gm_n468, in_11);
	and (gm_n8977, gm_n50, in_13, in_12, gm_n8976, gm_n63);
	and (gm_n8978, in_18, gm_n81, in_16, gm_n8977, in_19);
	nand (gm_n8979, gm_n8978, in_21, gm_n45);
	nand (gm_n8980, gm_n63, gm_n50, gm_n49, gm_n6861, gm_n46);
	nor (gm_n8981, in_19, gm_n47, gm_n81, gm_n8980, in_20);
	nand (gm_n8982, gm_n8981, in_21);
	nand (gm_n8983, in_15, in_14, gm_n49, gm_n4868, gm_n46);
	nor (gm_n8984, in_19, gm_n47, in_17, gm_n8983, gm_n45);
	nand (gm_n8985, gm_n8984, in_21);
	and (gm_n8986, gm_n50, gm_n49, gm_n48, gm_n3044, in_15);
	nand (gm_n8987, gm_n47, in_17, in_16, gm_n8986, gm_n62);
	nor (gm_n8988, gm_n8987, gm_n71, gm_n45);
	nand (gm_n8989, in_16, in_15, in_14, gm_n8831, in_17);
	nor (gm_n8990, in_20, in_19, gm_n47, gm_n8989, in_21);
	and (gm_n8991, gm_n48, gm_n53, gm_n52, gm_n1719, gm_n49);
	nand (gm_n8992, gm_n46, in_15, gm_n50, gm_n8991, gm_n81);
	nor (gm_n8993, in_20, in_19, in_18, gm_n8992, in_21);
	nand (gm_n8994, in_11, gm_n52, in_9, gm_n1178);
	nor (gm_n8995, gm_n50, gm_n49, gm_n48, gm_n8994, in_15);
	nand (gm_n8996, gm_n47, gm_n81, in_16, gm_n8995, in_19);
	nor (gm_n8997, gm_n8996, gm_n71, in_20);
	nor (gm_n8998, gm_n52, gm_n51, in_8, gm_n5379, in_11);
	nand (gm_n8999, in_14, in_13, in_12, gm_n8998, in_15);
	nor (gm_n9000, in_18, in_17, in_16, gm_n8999, in_19);
	nand (gm_n9001, gm_n9000, gm_n71, gm_n45);
	nand (gm_n9002, gm_n63, gm_n50, in_13, gm_n7879, gm_n46);
	nor (gm_n9003, gm_n62, in_18, gm_n81, gm_n9002, gm_n45);
	nand (gm_n9004, gm_n9003, in_21);
	nand (gm_n9005, in_13, gm_n48, in_11, gm_n6800, gm_n50);
	nor (gm_n9006, in_17, in_16, gm_n63, gm_n9005, in_18);
	nand (gm_n9007, gm_n71, in_20, in_19, gm_n9006);
	nor (gm_n9008, gm_n53, in_10, in_9, gm_n2902);
	nand (gm_n9009, gm_n50, in_13, gm_n48, gm_n9008, in_15);
	nor (gm_n9010, in_18, in_17, in_16, gm_n9009, gm_n62);
	nand (gm_n9011, gm_n9010, gm_n71, in_20);
	nand (gm_n9012, in_17, gm_n46, in_15, gm_n1817, in_18);
	nor (gm_n9013, gm_n71, in_20, in_19, gm_n9012);
	nor (gm_n9014, gm_n48, in_11, in_10, gm_n3515, gm_n49);
	nand (gm_n9015, gm_n46, gm_n63, gm_n50, gm_n9014, gm_n81);
	nor (gm_n9016, gm_n45, gm_n62, in_18, gm_n9015, gm_n71);
	and (gm_n9017, in_12, in_11, in_10, gm_n311, gm_n49);
	nand (gm_n9018, in_16, gm_n63, gm_n50, gm_n9017, gm_n81);
	nor (gm_n9019, gm_n45, gm_n62, in_18, gm_n9018, gm_n71);
	nand (gm_n9020, in_11, gm_n52, in_9, gm_n4273, gm_n48);
	nor (gm_n9021, in_15, in_14, gm_n49, gm_n9020, in_16);
	nand (gm_n9022, gm_n62, in_18, gm_n81, gm_n9021, gm_n45);
	nor (gm_n9023, gm_n9022, in_21);
	nand (gm_n9024, gm_n49, gm_n48, in_11, gm_n3543, gm_n50);
	nor (gm_n9025, in_17, in_16, gm_n63, gm_n9024, in_18);
	nand (gm_n9026, gm_n71, in_20, in_19, gm_n9025);
	nand (gm_n9027, gm_n49, gm_n48, in_11, gm_n1257, in_14);
	nor (gm_n9028, in_17, in_16, in_15, gm_n9027, gm_n47);
	nand (gm_n9029, gm_n71, in_20, in_19, gm_n9028);
	nor (gm_n9030, gm_n53, in_10, gm_n51, gm_n4562, in_12);
	nand (gm_n9031, gm_n63, gm_n50, gm_n49, gm_n9030, in_16);
	nor (gm_n9032, in_19, in_18, in_17, gm_n9031, in_20);
	nand (gm_n9033, gm_n9032, in_21);
	nand (gm_n9034, in_12, in_11, in_10, gm_n692, gm_n49);
	nor (gm_n9035, gm_n46, gm_n63, gm_n50, gm_n9034, in_17);
	nand (gm_n9036, gm_n45, in_19, in_18, gm_n9035, gm_n71);
	and (gm_n9037, in_14, in_13, in_12, gm_n8637, in_15);
	nand (gm_n9038, in_18, gm_n81, gm_n46, gm_n9037, gm_n62);
	nor (gm_n9039, gm_n9038, in_21, in_20);
	nor (gm_n9040, gm_n49, gm_n48, gm_n53, gm_n1179, in_14);
	nand (gm_n9041, in_17, gm_n46, in_15, gm_n9040, gm_n47);
	nor (gm_n9042, gm_n71, gm_n45, gm_n62, gm_n9041);
	nor (gm_n9043, gm_n2503, in_10, in_9);
	and (gm_n9044, gm_n49, gm_n48, gm_n53, gm_n9043, gm_n50);
	nand (gm_n9045, gm_n81, gm_n46, in_15, gm_n9044, in_18);
	nor (gm_n9046, in_21, in_20, in_19, gm_n9045);
	nor (gm_n9047, gm_n48, gm_n53, in_10, gm_n104, in_13);
	nand (gm_n9048, in_16, in_15, in_14, gm_n9047, gm_n81);
	nor (gm_n9049, gm_n45, gm_n62, in_18, gm_n9048, in_21);
	nand (gm_n9050, in_14, in_13, gm_n48, gm_n7626, gm_n63);
	nor (gm_n9051, in_18, in_17, gm_n46, gm_n9050, in_19);
	nand (gm_n9052, gm_n9051, gm_n71, gm_n45);
	nor (gm_n9053, gm_n46, gm_n63, gm_n50, gm_n5283, in_17);
	nand (gm_n9054, in_20, gm_n62, gm_n47, gm_n9053, in_21);
	nand (gm_n9055, in_12, gm_n53, in_10, gm_n5375, gm_n49);
	nor (gm_n9056, in_16, gm_n63, gm_n50, gm_n9055, gm_n81);
	nand (gm_n9057, gm_n45, gm_n62, gm_n47, gm_n9056, in_21);
	nand (gm_n9058, in_12, gm_n53, gm_n52, gm_n1413, in_13);
	nor (gm_n9059, in_16, gm_n63, gm_n50, gm_n9058, gm_n81);
	nand (gm_n9060, in_20, in_19, in_18, gm_n9059, in_21);
	nand (gm_n9061, gm_n53, in_10, in_9, gm_n902, in_12);
	nor (gm_n9062, in_15, gm_n50, gm_n49, gm_n9061, in_16);
	nand (gm_n9063, gm_n62, gm_n47, gm_n81, gm_n9062, gm_n45);
	nor (gm_n9064, gm_n9063, in_21);
	nor (gm_n9065, in_12, gm_n53, in_10, gm_n2043, in_13);
	nand (gm_n9066, in_16, gm_n63, in_14, gm_n9065, in_17);
	nor (gm_n9067, gm_n45, in_19, in_18, gm_n9066, gm_n71);
	and (gm_n9068, in_12, gm_n53, gm_n52, gm_n3727, in_13);
	nand (gm_n9069, gm_n46, gm_n63, in_14, gm_n9068, gm_n81);
	nor (gm_n9070, gm_n45, gm_n62, gm_n47, gm_n9069, in_21);
	and (gm_n9071, gm_n49, in_12, in_11, gm_n3889, in_14);
	nand (gm_n9072, gm_n81, in_16, in_15, gm_n9071, gm_n47);
	nor (gm_n9073, in_21, gm_n45, gm_n62, gm_n9072);
	or (gm_n9074, in_13, in_12, in_11, gm_n7319, in_14);
	nor (gm_n9075, in_17, gm_n46, gm_n63, gm_n9074, in_18);
	nand (gm_n9076, gm_n71, in_20, in_19, gm_n9075);
	nand (gm_n9077, in_12, in_11, gm_n52, gm_n1688, gm_n49);
	nor (gm_n9078, gm_n46, in_15, gm_n50, gm_n9077, gm_n81);
	nand (gm_n9079, in_20, in_19, gm_n47, gm_n9078, in_21);
	nand (gm_n9080, in_12, in_11, gm_n52, gm_n1080, gm_n49);
	nor (gm_n9081, gm_n46, gm_n63, in_14, gm_n9080, in_17);
	nand (gm_n9082, in_20, gm_n62, gm_n47, gm_n9081, in_21);
	or (gm_n9083, gm_n48, gm_n53, in_10, gm_n6475, in_13);
	nor (gm_n9084, gm_n46, gm_n63, in_14, gm_n9083, gm_n81);
	nand (gm_n9085, gm_n45, gm_n62, gm_n47, gm_n9084, gm_n71);
	nand (gm_n9086, in_8, in_7, gm_n82, gm_n374, in_9);
	nor (gm_n9087, in_12, gm_n53, in_10, gm_n9086, in_13);
	nand (gm_n9088, gm_n46, in_15, in_14, gm_n9087, gm_n81);
	nor (gm_n9089, gm_n45, gm_n62, gm_n47, gm_n9088, in_21);
	nand (gm_n9090, in_11, gm_n52, in_9, gm_n3451, gm_n48);
	nor (gm_n9091, gm_n63, in_14, in_13, gm_n9090, in_16);
	nand (gm_n9092, in_19, in_18, gm_n81, gm_n9091, gm_n45);
	nor (gm_n9093, gm_n9092, in_21);
	nand (gm_n9094, in_16, gm_n63, gm_n50, gm_n8328, in_17);
	nor (gm_n9095, in_20, in_19, in_18, gm_n9094, in_21);
	nand (gm_n9096, gm_n81, in_16, in_15, gm_n4399, in_18);
	nor (gm_n9097, in_21, gm_n45, in_19, gm_n9096);
	nand (gm_n9098, in_13, gm_n48, in_11, gm_n8311, gm_n50);
	nor (gm_n9099, in_17, gm_n46, in_15, gm_n9098, gm_n47);
	nand (gm_n9100, gm_n71, gm_n45, in_19, gm_n9099);
	nand (gm_n9101, in_12, gm_n53, gm_n52, gm_n2001, in_13);
	nor (gm_n9102, gm_n46, gm_n63, in_14, gm_n9101, gm_n81);
	nand (gm_n9103, in_20, gm_n62, gm_n47, gm_n9102, gm_n71);
	or (gm_n9104, gm_n48, gm_n53, in_10, gm_n5620, gm_n49);
	nor (gm_n9105, in_16, in_15, in_14, gm_n9104, in_17);
	nand (gm_n9106, gm_n45, gm_n62, gm_n47, gm_n9105, in_21);
	nand (gm_n9107, in_14, gm_n49, in_12, gm_n5264, in_15);
	nor (gm_n9108, in_18, gm_n81, in_16, gm_n9107, in_19);
	nand (gm_n9109, gm_n9108, in_21, gm_n45);
	nand (gm_n9110, in_16, in_15, gm_n50, gm_n5038, gm_n81);
	nor (gm_n9111, gm_n45, gm_n62, in_18, gm_n9110, gm_n71);
	nand (gm_n9112, in_19, gm_n47, in_17, gm_n8904, gm_n45);
	nor (gm_n9113, gm_n9112, gm_n71);
	nor (gm_n9114, in_13, gm_n48, in_11, gm_n1908, in_14);
	nand (gm_n9115, gm_n81, gm_n46, in_15, gm_n9114, in_18);
	nor (gm_n9116, gm_n71, in_20, gm_n62, gm_n9115);
	nor (gm_n9117, gm_n48, gm_n53, in_10, gm_n1174, in_13);
	nand (gm_n9118, gm_n46, gm_n63, in_14, gm_n9117, in_17);
	nor (gm_n9119, gm_n45, gm_n62, gm_n47, gm_n9118, in_21);
	nand (gm_n9120, gm_n48, gm_n53, gm_n52, gm_n5375, gm_n49);
	nor (gm_n9121, gm_n46, in_15, gm_n50, gm_n9120, gm_n81);
	nand (gm_n9122, gm_n45, gm_n62, in_18, gm_n9121, gm_n71);
	nand (gm_n9123, gm_n50, in_13, gm_n48, gm_n298, in_15);
	nor (gm_n9124, in_18, gm_n81, in_16, gm_n9123, gm_n62);
	nand (gm_n9125, gm_n9124, gm_n71, gm_n45);
	and (gm_n9126, gm_n46, in_15, in_14, gm_n2974, in_17);
	nand (gm_n9127, gm_n45, gm_n62, in_18, gm_n9126, in_21);
	nand (gm_n9128, gm_n63, in_14, in_13, gm_n1710, gm_n46);
	nor (gm_n9129, gm_n62, in_18, gm_n81, gm_n9128, gm_n45);
	nand (gm_n9130, gm_n9129, gm_n71);
	nand (gm_n9131, in_16, in_15, in_14, gm_n1113, in_17);
	nor (gm_n9132, in_20, in_19, in_18, gm_n9131, in_21);
	nor (gm_n9133, in_15, gm_n50, in_13, gm_n6613, in_16);
	nand (gm_n9134, in_19, gm_n47, gm_n81, gm_n9133, gm_n45);
	nor (gm_n9135, gm_n9134, gm_n71);
	or (gm_n9136, in_16, gm_n63, in_14, gm_n3732, gm_n81);
	nor (gm_n9137, gm_n45, in_19, gm_n47, gm_n9136, in_21);
	nand (gm_n9138, in_16, in_15, gm_n50, gm_n7224, gm_n81);
	nor (gm_n9139, gm_n45, gm_n62, gm_n47, gm_n9138, gm_n71);
	nor (gm_n9140, in_9, in_8, in_7, gm_n463, in_10);
	nand (gm_n9141, in_13, in_12, gm_n53, gm_n9140, gm_n50);
	nor (gm_n9142, gm_n81, in_16, gm_n63, gm_n9141, in_18);
	nand (gm_n9143, gm_n71, gm_n45, in_19, gm_n9142);
	nand (gm_n9144, gm_n50, in_13, in_12, gm_n9008, in_15);
	nor (gm_n9145, in_18, in_17, in_16, gm_n9144, gm_n62);
	nand (gm_n9146, gm_n9145, in_21, in_20);
	and (gm_n9147, gm_n6996, in_13);
	and (gm_n9148, gm_n46, in_15, gm_n50, gm_n9147, in_17);
	nand (gm_n9149, in_20, in_19, in_18, gm_n9148, gm_n71);
	nand (gm_n9150, in_13, gm_n48, in_11, gm_n3920, in_14);
	nor (gm_n9151, gm_n81, in_16, gm_n63, gm_n9150, gm_n47);
	nand (gm_n9152, gm_n71, gm_n45, gm_n62, gm_n9151);
	nand (gm_n9153, gm_n691, in_9, gm_n64);
	nor (gm_n9154, gm_n48, gm_n53, gm_n52, gm_n9153, in_13);
	nand (gm_n9155, gm_n46, gm_n63, gm_n50, gm_n9154, in_17);
	nor (gm_n9156, gm_n45, gm_n62, in_18, gm_n9155, gm_n71);
	or (gm_n9157, in_10, gm_n51, in_8, gm_n2239, gm_n53);
	nor (gm_n9158, gm_n50, in_13, in_12, gm_n9157, in_15);
	nand (gm_n9159, gm_n47, gm_n81, gm_n46, gm_n9158, gm_n62);
	nor (gm_n9160, gm_n9159, gm_n71, gm_n45);
	or (gm_n9161, gm_n53, in_10, in_9, gm_n1957, in_12);
	nor (gm_n9162, in_15, in_14, in_13, gm_n9161, in_16);
	nand (gm_n9163, in_19, gm_n47, gm_n81, gm_n9162, gm_n45);
	nor (gm_n9164, gm_n9163, gm_n71);
	and (gm_n9165, gm_n49, gm_n48, in_11, gm_n6773, gm_n50);
	nand (gm_n9166, gm_n81, gm_n46, in_15, gm_n9165, gm_n47);
	nor (gm_n9167, gm_n71, in_20, gm_n62, gm_n9166);
	nor (gm_n9168, in_11, gm_n52, gm_n51, gm_n253, in_12);
	nand (gm_n9169, gm_n63, in_14, in_13, gm_n9168, in_16);
	nor (gm_n9170, in_19, gm_n47, gm_n81, gm_n9169, gm_n45);
	nand (gm_n9171, gm_n9170, in_21);
	nand (gm_n9172, gm_n49, gm_n48, gm_n53, gm_n5305, in_14);
	nor (gm_n9173, gm_n81, in_16, gm_n63, gm_n9172, gm_n47);
	nand (gm_n9174, in_21, gm_n45, in_19, gm_n9173);
	nand (gm_n9175, gm_n50, in_13, gm_n48, gm_n3760, in_15);
	nor (gm_n9176, gm_n47, gm_n81, gm_n46, gm_n9175, gm_n62);
	nand (gm_n9177, gm_n9176, in_21, in_20);
	nand (gm_n9178, in_12, gm_n53, in_10, gm_n8629, gm_n49);
	nor (gm_n9179, gm_n46, in_15, gm_n50, gm_n9178, in_17);
	nand (gm_n9180, gm_n45, in_19, in_18, gm_n9179, in_21);
	nor (gm_n9181, in_12, in_11, in_10, gm_n7235, in_13);
	nand (gm_n9182, gm_n46, in_15, in_14, gm_n9181, gm_n81);
	nor (gm_n9183, in_20, in_19, gm_n47, gm_n9182, gm_n71);
	nand (gm_n9184, gm_n46, gm_n63, gm_n50, gm_n4355, in_17);
	nor (gm_n9185, in_20, gm_n62, gm_n47, gm_n9184, gm_n71);
	nor (gm_n9186, in_13, in_12, in_11, gm_n6397, in_14);
	nand (gm_n9187, in_17, gm_n46, in_15, gm_n9186, in_18);
	nor (gm_n9188, in_21, gm_n45, gm_n62, gm_n9187);
	nor (gm_n9189, gm_n1052, gm_n52, in_9);
	and (gm_n9190, in_13, in_12, gm_n53, gm_n9189, in_14);
	nand (gm_n9191, gm_n81, gm_n46, in_15, gm_n9190, in_18);
	nor (gm_n9192, gm_n71, gm_n45, gm_n62, gm_n9191);
	nand (gm_n9193, gm_n50, gm_n49, gm_n48, gm_n8290, in_15);
	nor (gm_n9194, gm_n47, gm_n81, in_16, gm_n9193, gm_n62);
	nand (gm_n9195, gm_n9194, gm_n71, in_20);
	nand (gm_n9196, in_15, in_14, in_13, gm_n3272, in_16);
	nor (gm_n9197, in_19, gm_n47, in_17, gm_n9196, in_20);
	nand (gm_n9198, gm_n9197, gm_n71);
	or (gm_n9199, in_12, in_11, gm_n52, gm_n7154, gm_n49);
	nor (gm_n9200, gm_n46, gm_n63, gm_n50, gm_n9199, in_17);
	nand (gm_n9201, in_20, in_19, in_18, gm_n9200, in_21);
	nand (gm_n9202, in_13, in_12, in_11, gm_n7425, in_14);
	nor (gm_n9203, gm_n81, in_16, in_15, gm_n9202, in_18);
	nand (gm_n9204, gm_n71, in_20, in_19, gm_n9203);
	and (gm_n9205, gm_n50, gm_n49, in_12, gm_n1340, gm_n63);
	nand (gm_n9206, gm_n47, in_17, gm_n46, gm_n9205, gm_n62);
	nor (gm_n9207, gm_n9206, gm_n71, in_20);
	and (gm_n9208, gm_n48, in_11, in_10, gm_n3069, gm_n49);
	nand (gm_n9209, gm_n46, gm_n63, in_14, gm_n9208, gm_n81);
	nor (gm_n9210, gm_n45, gm_n62, gm_n47, gm_n9209, gm_n71);
	and (gm_n9211, in_14, in_13, in_12, gm_n2824, gm_n63);
	nand (gm_n9212, in_18, in_17, gm_n46, gm_n9211, in_19);
	nor (gm_n9213, gm_n9212, gm_n71, gm_n45);
	nor (gm_n9214, in_14, gm_n49, in_12, gm_n8113, in_15);
	nand (gm_n9215, gm_n47, in_17, in_16, gm_n9214, gm_n62);
	nor (gm_n9216, gm_n9215, gm_n71, in_20);
	nand (gm_n9217, gm_n48, gm_n53, in_10, gm_n5676, in_13);
	nor (gm_n9218, gm_n46, in_15, gm_n50, gm_n9217, gm_n81);
	nand (gm_n9219, gm_n45, in_19, in_18, gm_n9218, in_21);
	nand (gm_n9220, gm_n48, gm_n53, in_10, gm_n6668, in_13);
	nor (gm_n9221, in_16, in_15, gm_n50, gm_n9220, in_17);
	nand (gm_n9222, in_20, gm_n62, in_18, gm_n9221, gm_n71);
	nand (gm_n9223, gm_n48, gm_n53, in_10, gm_n3748, gm_n49);
	nor (gm_n9224, in_16, gm_n63, gm_n50, gm_n9223, in_17);
	nand (gm_n9225, gm_n45, gm_n62, in_18, gm_n9224, gm_n71);
	nor (gm_n9226, in_11, in_10, in_9, gm_n2266, in_12);
	nand (gm_n9227, in_15, in_14, gm_n49, gm_n9226, gm_n46);
	nor (gm_n9228, in_19, gm_n47, in_17, gm_n9227, in_20);
	nand (gm_n9229, gm_n9228, gm_n71);
	or (gm_n9230, gm_n46, in_15, gm_n50, gm_n5807, gm_n81);
	nor (gm_n9231, in_20, gm_n62, gm_n47, gm_n9230, gm_n71);
	and (gm_n9232, gm_n63, gm_n50, gm_n49, gm_n6804, in_16);
	nand (gm_n9233, gm_n62, gm_n47, in_17, gm_n9232, in_20);
	nor (gm_n9234, gm_n9233, in_21);
	and (gm_n9235, gm_n48, gm_n53, gm_n52, gm_n2555, in_13);
	nand (gm_n9236, in_16, in_15, in_14, gm_n9235, gm_n81);
	nor (gm_n9237, in_20, in_19, gm_n47, gm_n9236, in_21);
	nor (gm_n9238, in_14, gm_n49, in_12, gm_n2382, gm_n63);
	nand (gm_n9239, gm_n47, gm_n81, in_16, gm_n9238, gm_n62);
	nor (gm_n9240, gm_n9239, in_21, gm_n45);
	nand (gm_n9241, gm_n63, gm_n50, gm_n49, gm_n495, gm_n46);
	nor (gm_n9242, gm_n62, gm_n47, gm_n81, gm_n9241, gm_n45);
	nand (gm_n9243, gm_n9242, in_21);
	nand (gm_n9244, in_12, gm_n53, gm_n52, gm_n142, gm_n49);
	nor (gm_n9245, in_16, in_15, gm_n50, gm_n9244, gm_n81);
	nand (gm_n9246, gm_n45, gm_n62, gm_n47, gm_n9245, in_21);
	nand (gm_n9247, gm_n48, gm_n53, in_10, gm_n4570, in_13);
	nor (gm_n9248, gm_n46, in_15, in_14, gm_n9247, in_17);
	nand (gm_n9249, gm_n45, gm_n62, in_18, gm_n9248, gm_n71);
	nand (gm_n9250, gm_n48, in_11, gm_n52, gm_n654, gm_n49);
	nor (gm_n9251, in_16, gm_n63, in_14, gm_n9250, gm_n81);
	nand (gm_n9252, gm_n45, in_19, in_18, gm_n9251, in_21);
	and (gm_n9253, in_11, in_10, in_9, gm_n1279);
	and (gm_n9254, in_14, gm_n49, gm_n48, gm_n9253, gm_n63);
	nand (gm_n9255, in_18, gm_n81, in_16, gm_n9254, gm_n62);
	nor (gm_n9256, gm_n9255, gm_n71, gm_n45);
	nor (gm_n9257, gm_n50, gm_n49, gm_n48, gm_n3476, gm_n63);
	nand (gm_n9258, in_18, in_17, gm_n46, gm_n9257, in_19);
	nor (gm_n9259, gm_n9258, in_21, in_20);
	nand (gm_n9260, in_11, gm_n52, gm_n51, gm_n109, gm_n48);
	nor (gm_n9261, gm_n63, gm_n50, gm_n49, gm_n9260, in_16);
	nand (gm_n9262, gm_n62, in_18, in_17, gm_n9261, in_20);
	nor (gm_n9263, gm_n9262, in_21);
	nor (gm_n9264, gm_n50, in_13, in_12, gm_n613, in_15);
	nand (gm_n9265, in_18, gm_n81, gm_n46, gm_n9264, in_19);
	nor (gm_n9266, gm_n9265, in_21, gm_n45);
	and (gm_n9267, in_9, in_8, gm_n55, gm_n151, gm_n52);
	nand (gm_n9268, in_13, gm_n48, gm_n53, gm_n9267, gm_n50);
	nor (gm_n9269, gm_n81, gm_n46, gm_n63, gm_n9268, gm_n47);
	nand (gm_n9270, gm_n71, in_20, gm_n62, gm_n9269);
	nor (gm_n9271, in_11, in_10, in_9, gm_n1052, in_12);
	nand (gm_n9272, gm_n9271, gm_n50, gm_n49);
	nor (gm_n9273, gm_n81, in_16, in_15, gm_n9272, in_18);
	nand (gm_n9274, gm_n71, in_20, in_19, gm_n9273);
	nor (gm_n9275, in_16, gm_n63, gm_n50, gm_n4738, gm_n81);
	nand (gm_n9276, gm_n45, in_19, gm_n47, gm_n9275, in_21);
	nand (gm_n9277, gm_n63, in_14, in_13, gm_n4108, in_16);
	nor (gm_n9278, gm_n62, in_18, in_17, gm_n9277, gm_n45);
	nand (gm_n9279, gm_n9278, gm_n71);
	nand (gm_n9280, in_17, gm_n46, gm_n63, gm_n3263, gm_n47);
	nor (gm_n9281, in_21, gm_n45, gm_n62, gm_n9280);
	and (gm_n9282, gm_n63, in_14, gm_n49, gm_n6777, in_16);
	nand (gm_n9283, gm_n62, in_18, gm_n81, gm_n9282, in_20);
	nor (gm_n9284, gm_n9283, in_21);
	and (gm_n9285, in_14, in_13, gm_n48, gm_n3065, in_15);
	nand (gm_n9286, gm_n47, in_17, in_16, gm_n9285, gm_n62);
	nor (gm_n9287, gm_n9286, gm_n71, in_20);
	nand (gm_n9288, in_11, gm_n52, in_9, gm_n6549, in_12);
	nor (gm_n9289, in_15, gm_n50, in_13, gm_n9288, in_16);
	nand (gm_n9290, gm_n62, gm_n47, gm_n81, gm_n9289, gm_n45);
	nor (gm_n9291, gm_n9290, gm_n71);
	nor (gm_n9292, in_11, gm_n52, in_9, gm_n3146);
	nand (gm_n9293, in_14, in_13, in_12, gm_n9292, gm_n63);
	nor (gm_n9294, in_18, gm_n81, gm_n46, gm_n9293, gm_n62);
	nand (gm_n9295, gm_n9294, gm_n71, in_20);
	nand (gm_n9296, in_12, in_11, in_10, gm_n1365, in_13);
	nor (gm_n9297, in_16, gm_n63, gm_n50, gm_n9296, in_17);
	nand (gm_n9298, gm_n45, in_19, gm_n47, gm_n9297, in_21);
	and (gm_n9299, in_17, in_16, gm_n63, gm_n4508, in_18);
	nand (gm_n9300, in_21, in_20, in_19, gm_n9299);
	nor (gm_n9301, gm_n52, gm_n51, in_8, gm_n3077, in_11);
	nand (gm_n9302, in_14, gm_n49, gm_n48, gm_n9301, in_15);
	nor (gm_n9303, gm_n47, in_17, in_16, gm_n9302, gm_n62);
	nand (gm_n9304, gm_n9303, in_21, gm_n45);
	nor (gm_n9305, gm_n49, gm_n48, gm_n53, gm_n3833, gm_n50);
	nand (gm_n9306, in_17, in_16, gm_n63, gm_n9305, gm_n47);
	nor (gm_n9307, gm_n71, in_20, gm_n62, gm_n9306);
	nand (gm_n9308, gm_n81, in_16, gm_n63, gm_n9190, gm_n47);
	nor (gm_n9309, gm_n71, in_20, gm_n62, gm_n9308);
	nor (gm_n9310, in_15, gm_n50, gm_n49, gm_n2195, gm_n46);
	nand (gm_n9311, in_19, in_18, gm_n81, gm_n9310, gm_n45);
	nor (gm_n9312, gm_n9311, in_21);
	and (gm_n9313, in_13, gm_n48, gm_n53, gm_n7250, in_14);
	nand (gm_n9314, gm_n81, gm_n46, gm_n63, gm_n9313, in_18);
	nor (gm_n9315, in_21, in_20, gm_n62, gm_n9314);
	nand (gm_n9316, gm_n49, gm_n48, in_11, gm_n1865, in_14);
	nor (gm_n9317, in_17, gm_n46, gm_n63, gm_n9316, in_18);
	nand (gm_n9318, gm_n71, gm_n45, gm_n62, gm_n9317);
	nand (gm_n9319, gm_n48, gm_n53, in_10, gm_n4630, gm_n49);
	nor (gm_n9320, gm_n46, gm_n63, in_14, gm_n9319, gm_n81);
	nand (gm_n9321, gm_n45, in_19, gm_n47, gm_n9320, gm_n71);
	nor (gm_n9322, in_13, gm_n48, in_11, gm_n4972);
	and (gm_n9323, gm_n46, in_15, in_14, gm_n9322, in_17);
	nand (gm_n9324, gm_n45, gm_n62, gm_n47, gm_n9323, gm_n71);
	nand (gm_n9325, gm_n55, in_6, in_5, gm_n493, in_8);
	nor (gm_n9326, gm_n53, in_10, gm_n51, gm_n9325, in_12);
	nand (gm_n9327, gm_n63, in_14, gm_n49, gm_n9326, gm_n46);
	nor (gm_n9328, gm_n62, gm_n47, gm_n81, gm_n9327, gm_n45);
	nand (gm_n9329, gm_n9328, gm_n71);
	or (gm_n9330, gm_n53, in_10, in_9, gm_n8122, gm_n48);
	nor (gm_n9331, gm_n63, in_14, gm_n49, gm_n9330, in_16);
	nand (gm_n9332, gm_n62, gm_n47, gm_n81, gm_n9331, gm_n45);
	nor (gm_n9333, gm_n9332, gm_n71);
	nand (gm_n9334, in_12, in_11, in_10, gm_n4319, in_13);
	or (gm_n9335, in_16, in_15, in_14, gm_n9334, in_17);
	nor (gm_n9336, gm_n45, gm_n62, in_18, gm_n9335, gm_n71);
	or (gm_n9337, in_11, gm_n52, gm_n51, gm_n1879, in_12);
	nor (gm_n9338, in_15, in_14, gm_n49, gm_n9337, gm_n46);
	nand (gm_n9339, gm_n62, in_18, in_17, gm_n9338, in_20);
	nor (gm_n9340, gm_n9339, in_21);
	nor (gm_n9341, gm_n53, in_10, in_9, gm_n1750);
	and (gm_n9342, gm_n50, in_13, in_12, gm_n9341, in_15);
	nand (gm_n9343, in_18, gm_n81, in_16, gm_n9342, in_19);
	nor (gm_n9344, gm_n9343, gm_n71, gm_n45);
	nand (gm_n9345, in_14, gm_n49, in_12, gm_n7729, in_15);
	nor (gm_n9346, gm_n47, in_17, in_16, gm_n9345, in_19);
	nand (gm_n9347, gm_n9346, gm_n71, gm_n45);
	and (gm_n9348, gm_n46, in_15, in_14, gm_n8529, gm_n81);
	nand (gm_n9349, in_20, gm_n62, gm_n47, gm_n9348, gm_n71);
	nand (gm_n9350, in_12, in_11, in_10, gm_n1962, in_13);
	nor (gm_n9351, in_16, gm_n63, in_14, gm_n9350, gm_n81);
	nand (gm_n9352, in_20, in_19, gm_n47, gm_n9351, gm_n71);
	and (gm_n9353, gm_n53, gm_n52, gm_n51, gm_n2432, in_12);
	nand (gm_n9354, gm_n63, gm_n50, in_13, gm_n9353, in_16);
	nor (gm_n9355, gm_n62, gm_n47, gm_n81, gm_n9354, in_20);
	nand (gm_n9356, gm_n9355, gm_n71);
	nand (gm_n9357, gm_n1380, gm_n52, gm_n51);
	nor (gm_n9358, gm_n49, gm_n48, gm_n53, gm_n9357, gm_n50);
	nand (gm_n9359, in_17, gm_n46, in_15, gm_n9358, gm_n47);
	nor (gm_n9360, in_21, gm_n45, in_19, gm_n9359);
	nand (gm_n9361, in_11, in_10, gm_n51, gm_n4273, gm_n48);
	nor (gm_n9362, in_15, gm_n50, in_13, gm_n9361, gm_n46);
	nand (gm_n9363, in_19, in_18, in_17, gm_n9362, gm_n45);
	nor (gm_n9364, gm_n9363, gm_n71);
	nand (gm_n9365, in_11, in_10, in_9, gm_n2194, gm_n48);
	nor (gm_n9366, in_15, in_14, gm_n49, gm_n9365, in_16);
	nand (gm_n9367, in_19, in_18, in_17, gm_n9366, gm_n45);
	nor (gm_n9368, gm_n9367, gm_n71);
	nand (gm_n9369, gm_n46, in_15, gm_n50, gm_n5748, in_17);
	nor (gm_n9370, in_20, gm_n62, gm_n47, gm_n9369, gm_n71);
	nor (gm_n9371, in_11, gm_n52, in_9, gm_n410, in_12);
	nand (gm_n9372, gm_n63, gm_n50, gm_n49, gm_n9371, gm_n46);
	nor (gm_n9373, gm_n62, in_18, in_17, gm_n9372, in_20);
	nand (gm_n9374, gm_n9373, gm_n71);
	nor (gm_n9375, gm_n53, in_10, gm_n51, gm_n3542, in_12);
	nand (gm_n9376, in_15, gm_n50, gm_n49, gm_n9375, gm_n46);
	nor (gm_n9377, gm_n62, gm_n47, gm_n81, gm_n9376, in_20);
	nand (gm_n9378, gm_n9377, gm_n71);
	nand (gm_n9379, gm_n50, in_13, in_12, gm_n4154, gm_n63);
	nor (gm_n9380, gm_n47, gm_n81, in_16, gm_n9379, gm_n62);
	nand (gm_n9381, gm_n9380, in_21, gm_n45);
	nand (gm_n9382, gm_n48, in_11, gm_n52, gm_n4127, gm_n49);
	nor (gm_n9383, in_16, gm_n63, in_14, gm_n9382, in_17);
	nand (gm_n9384, in_20, in_19, gm_n47, gm_n9383, in_21);
	nand (gm_n9385, in_11, in_10, in_9, gm_n3214);
	nor (gm_n9386, in_14, gm_n49, gm_n48, gm_n9385);
	nand (gm_n9387, in_17, gm_n46, gm_n63, gm_n9386, in_18);
	nor (gm_n9388, in_21, in_20, gm_n62, gm_n9387);
	nand (gm_n9389, gm_n53, gm_n52, gm_n51, gm_n1788, gm_n48);
	nor (gm_n9390, in_15, gm_n50, in_13, gm_n9389, gm_n46);
	nand (gm_n9391, gm_n62, in_18, in_17, gm_n9390, in_20);
	nor (gm_n9392, gm_n9391, in_21);
	or (gm_n9393, in_11, gm_n52, gm_n51, gm_n1434, gm_n48);
	nor (gm_n9394, gm_n63, gm_n50, in_13, gm_n9393, in_16);
	nand (gm_n9395, in_19, in_18, gm_n81, gm_n9394, gm_n45);
	nor (gm_n9396, gm_n9395, gm_n71);
	nand (gm_n9397, in_11, gm_n52, gm_n51, gm_n1952, gm_n48);
	nor (gm_n9398, in_15, in_14, in_13, gm_n9397, in_16);
	nand (gm_n9399, in_19, in_18, in_17, gm_n9398, in_20);
	nor (gm_n9400, gm_n9399, in_21);
	nor (gm_n9401, in_10, in_9, gm_n64, gm_n3077, in_11);
	nand (gm_n9402, gm_n50, in_13, in_12, gm_n9401, gm_n63);
	nor (gm_n9403, in_18, in_17, gm_n46, gm_n9402, gm_n62);
	nand (gm_n9404, gm_n9403, in_21, in_20);
	nand (gm_n9405, in_14, in_13, gm_n48, gm_n4992, in_15);
	nor (gm_n9406, gm_n47, gm_n81, in_16, gm_n9405, in_19);
	nand (gm_n9407, gm_n9406, in_21, gm_n45);
	nand (gm_n9408, gm_n48, in_11, in_10, gm_n120, in_13);
	nor (gm_n9409, gm_n46, in_15, in_14, gm_n9408, in_17);
	nand (gm_n9410, gm_n45, gm_n62, in_18, gm_n9409, gm_n71);
	nor (gm_n9411, gm_n47, in_17, gm_n46, gm_n3136, in_19);
	nand (gm_n9412, gm_n9411, in_21, gm_n45);
	nor (gm_n9413, in_12, in_11, in_10, gm_n432, gm_n49);
	nand (gm_n9414, in_16, in_15, gm_n50, gm_n9413, gm_n81);
	nor (gm_n9415, gm_n45, gm_n62, in_18, gm_n9414, gm_n71);
	nand (gm_n9416, in_11, gm_n52, gm_n51, gm_n3856, gm_n48);
	nor (gm_n9417, in_15, gm_n50, in_13, gm_n9416, in_16);
	nand (gm_n9418, gm_n62, gm_n47, in_17, gm_n9417, in_20);
	nor (gm_n9419, gm_n9418, in_21);
	nor (gm_n9420, gm_n49, gm_n48, in_11, gm_n3655, in_14);
	nand (gm_n9421, gm_n81, in_16, in_15, gm_n9420, gm_n47);
	nor (gm_n9422, in_21, in_20, gm_n62, gm_n9421);
	nand (gm_n9423, gm_n46, gm_n63, gm_n50, gm_n5191, in_17);
	nor (gm_n9424, in_20, in_19, gm_n47, gm_n9423, in_21);
	or (gm_n9425, in_7, in_6, in_5, gm_n75, gm_n64);
	nor (gm_n9426, gm_n9425, gm_n51);
	nand (gm_n9427, gm_n48, in_11, in_10, gm_n9426, gm_n49);
	nor (gm_n9428, in_16, in_15, gm_n50, gm_n9427, in_17);
	nand (gm_n9429, gm_n45, in_19, gm_n47, gm_n9428, gm_n71);
	nand (gm_n9430, in_14, in_13, in_12, gm_n3276, gm_n63);
	nor (gm_n9431, gm_n47, in_17, in_16, gm_n9430, gm_n62);
	nand (gm_n9432, gm_n9431, in_21, gm_n45);
	or (gm_n9433, in_12, in_11, gm_n52, gm_n104, gm_n49);
	nor (gm_n9434, in_16, in_15, in_14, gm_n9433, in_17);
	nand (gm_n9435, in_20, in_19, in_18, gm_n9434, gm_n71);
	and (gm_n9436, in_10, gm_n51, gm_n64, gm_n338);
	nand (gm_n9437, gm_n49, in_12, gm_n53, gm_n9436, in_14);
	nor (gm_n9438, in_17, gm_n46, in_15, gm_n9437, gm_n47);
	nand (gm_n9439, gm_n71, gm_n45, gm_n62, gm_n9438);
	nand (gm_n9440, in_14, gm_n49, gm_n48, gm_n8064, gm_n63);
	nor (gm_n9441, in_18, gm_n81, in_16, gm_n9440, in_19);
	nand (gm_n9442, gm_n9441, in_21, in_20);
	nand (gm_n9443, gm_n9435, gm_n9432, gm_n9429, gm_n9442, gm_n9439);
	nor (gm_n9444, gm_n9422, gm_n9419, gm_n9415, gm_n9443, gm_n9424);
	nand (gm_n9445, gm_n9410, gm_n9407, gm_n9404, gm_n9444, gm_n9412);
	nor (gm_n9446, gm_n9396, gm_n9392, gm_n9388, gm_n9445, gm_n9400);
	nand (gm_n9447, gm_n9381, gm_n9378, gm_n9374, gm_n9446, gm_n9384);
	nor (gm_n9448, gm_n9368, gm_n9364, gm_n9360, gm_n9447, gm_n9370);
	nand (gm_n9449, gm_n9352, gm_n9349, gm_n9347, gm_n9448, gm_n9356);
	nor (gm_n9450, gm_n9340, gm_n9336, gm_n9333, gm_n9449, gm_n9344);
	nand (gm_n9451, gm_n9324, gm_n9321, gm_n9318, gm_n9450, gm_n9329);
	nor (gm_n9452, gm_n9312, gm_n9309, gm_n9307, gm_n9451, gm_n9315);
	nand (gm_n9453, gm_n9300, gm_n9298, gm_n9295, gm_n9452, gm_n9304);
	nor (gm_n9454, gm_n9287, gm_n9284, gm_n9281, gm_n9453, gm_n9291);
	nand (gm_n9455, gm_n9276, gm_n9274, gm_n9270, gm_n9454, gm_n9279);
	nor (gm_n9456, gm_n9263, gm_n9259, gm_n9256, gm_n9455, gm_n9266);
	nand (gm_n9457, gm_n9249, gm_n9246, gm_n9243, gm_n9456, gm_n9252);
	nor (gm_n9458, gm_n9237, gm_n9234, gm_n9231, gm_n9457, gm_n9240);
	nand (gm_n9459, gm_n9225, gm_n9222, gm_n9219, gm_n9458, gm_n9229);
	nor (gm_n9460, gm_n9213, gm_n9210, gm_n9207, gm_n9459, gm_n9216);
	nand (gm_n9461, gm_n9201, gm_n9198, gm_n9195, gm_n9460, gm_n9204);
	nor (gm_n9462, gm_n9188, gm_n9185, gm_n9183, gm_n9461, gm_n9192);
	nand (gm_n9463, gm_n9177, gm_n9174, gm_n9171, gm_n9462, gm_n9180);
	nor (gm_n9464, gm_n9164, gm_n9160, gm_n9156, gm_n9463, gm_n9167);
	nand (gm_n9465, gm_n9149, gm_n9146, gm_n9143, gm_n9464, gm_n9152);
	nor (gm_n9466, gm_n9137, gm_n9135, gm_n9132, gm_n9465, gm_n9139);
	nand (gm_n9467, gm_n9127, gm_n9125, gm_n9122, gm_n9466, gm_n9130);
	nor (gm_n9468, gm_n9116, gm_n9113, gm_n9111, gm_n9467, gm_n9119);
	nand (gm_n9469, gm_n9106, gm_n9103, gm_n9100, gm_n9468, gm_n9109);
	nor (gm_n9470, gm_n9095, gm_n9093, gm_n9089, gm_n9469, gm_n9097);
	nand (gm_n9471, gm_n9082, gm_n9079, gm_n9076, gm_n9470, gm_n9085);
	nor (gm_n9472, gm_n9070, gm_n9067, gm_n9064, gm_n9471, gm_n9073);
	nand (gm_n9473, gm_n9057, gm_n9054, gm_n9052, gm_n9472, gm_n9060);
	nor (gm_n9474, gm_n9046, gm_n9042, gm_n9039, gm_n9473, gm_n9049);
	nand (gm_n9475, gm_n9033, gm_n9029, gm_n9026, gm_n9474, gm_n9036);
	nor (gm_n9476, gm_n9019, gm_n9016, gm_n9013, gm_n9475, gm_n9023);
	nand (gm_n9477, gm_n9007, gm_n9004, gm_n9001, gm_n9476, gm_n9011);
	nor (gm_n9478, gm_n8993, gm_n8990, gm_n8988, gm_n9477, gm_n8997);
	nand (gm_n9479, gm_n8982, gm_n8979, gm_n8975, gm_n9478, gm_n8985);
	nor (out_15, gm_n9479, gm_n8972);
	nand (gm_n9481, gm_n53, in_10, gm_n51, gm_n1212, in_12);
	nor (gm_n9482, in_15, gm_n50, gm_n49, gm_n9481, gm_n46);
	nand (gm_n9483, gm_n62, in_18, in_17, gm_n9482, gm_n45);
	nor (gm_n9484, gm_n9483, gm_n71);
	nor (gm_n9485, gm_n53, gm_n52, gm_n51, gm_n1869);
	nand (gm_n9486, in_14, in_13, gm_n48, gm_n9485, in_15);
	nor (gm_n9487, gm_n47, in_17, gm_n46, gm_n9486, gm_n62);
	nand (gm_n9488, gm_n9487, gm_n71, in_20);
	nand (gm_n9489, gm_n48, in_11, gm_n52, gm_n7176, in_13);
	nor (gm_n9490, in_16, in_15, in_14, gm_n9489, gm_n81);
	nand (gm_n9491, in_20, in_19, gm_n47, gm_n9490, gm_n71);
	and (gm_n9492, gm_n1222, gm_n52, in_9);
	nand (gm_n9493, gm_n49, in_12, in_11, gm_n9492, in_14);
	nor (gm_n9494, gm_n81, gm_n46, in_15, gm_n9493, gm_n47);
	nand (gm_n9495, in_21, in_20, in_19, gm_n9494);
	nand (gm_n9496, in_13, gm_n48, in_11, gm_n9043, in_14);
	nor (gm_n9497, in_17, in_16, gm_n63, gm_n9496, in_18);
	nand (gm_n9498, gm_n71, gm_n45, in_19, gm_n9497);
	and (gm_n9499, in_12, gm_n53, gm_n52, gm_n2729, in_13);
	nand (gm_n9500, in_16, in_15, in_14, gm_n9499, gm_n81);
	nor (gm_n9501, gm_n45, gm_n62, in_18, gm_n9500, gm_n71);
	nand (gm_n9502, in_11, in_10, in_9, gm_n2254);
	nor (gm_n9503, in_14, gm_n49, in_12, gm_n9502, in_15);
	nand (gm_n9504, in_18, gm_n81, gm_n46, gm_n9503, in_19);
	nor (gm_n9505, gm_n9504, gm_n71, gm_n45);
	nor (gm_n9506, gm_n63, in_14, gm_n49, gm_n4191, gm_n46);
	nand (gm_n9507, gm_n62, gm_n47, gm_n81, gm_n9506, in_20);
	nor (gm_n9508, gm_n9507, gm_n71);
	and (gm_n9509, in_12, in_11, in_10, gm_n1688, in_13);
	nand (gm_n9510, gm_n46, gm_n63, gm_n50, gm_n9509, in_17);
	nor (gm_n9511, in_20, gm_n62, in_18, gm_n9510, gm_n71);
	nand (gm_n9512, in_12, in_11, in_10, gm_n6217, in_13);
	nor (gm_n9513, gm_n46, gm_n63, gm_n50, gm_n9512, in_17);
	nand (gm_n9514, in_20, in_19, gm_n47, gm_n9513, in_21);
	nand (gm_n9515, in_14, gm_n49, gm_n48, gm_n1772, in_15);
	nor (gm_n9516, gm_n47, in_17, in_16, gm_n9515, in_19);
	nand (gm_n9517, gm_n9516, in_21, gm_n45);
	and (gm_n9518, gm_n64, gm_n55, in_6, gm_n1075, gm_n51);
	nand (gm_n9519, gm_n48, in_11, in_10, gm_n9518, gm_n49);
	nor (gm_n9520, in_16, in_15, gm_n50, gm_n9519, gm_n81);
	nand (gm_n9521, gm_n45, gm_n62, in_18, gm_n9520, gm_n71);
	nor (gm_n9522, in_11, in_10, in_9, gm_n2077, gm_n48);
	nand (gm_n9523, gm_n63, gm_n50, gm_n49, gm_n9522, in_16);
	nor (gm_n9524, in_19, gm_n47, in_17, gm_n9523, gm_n45);
	nand (gm_n9525, gm_n9524, gm_n71);
	nor (gm_n9526, in_13, in_12, gm_n53, gm_n8276, in_14);
	nand (gm_n9527, in_17, gm_n46, in_15, gm_n9526, gm_n47);
	nor (gm_n9528, gm_n71, in_20, in_19, gm_n9527);
	or (gm_n9529, in_16, gm_n63, gm_n50, gm_n5673, gm_n81);
	nor (gm_n9530, gm_n45, gm_n62, gm_n47, gm_n9529, gm_n71);
	nor (gm_n9531, gm_n49, gm_n48, in_11, gm_n6305, gm_n50);
	nand (gm_n9532, gm_n81, in_16, gm_n63, gm_n9531, in_18);
	nor (gm_n9533, gm_n71, in_20, in_19, gm_n9532);
	nor (gm_n9534, in_12, in_11, gm_n52, gm_n104, in_13);
	nand (gm_n9535, gm_n46, gm_n63, gm_n50, gm_n9534, in_17);
	nor (gm_n9536, in_20, gm_n62, gm_n47, gm_n9535, in_21);
	nor (gm_n9537, gm_n64, gm_n55, in_6, gm_n96, in_9);
	nand (gm_n9538, in_12, in_11, in_10, gm_n9537, gm_n49);
	nor (gm_n9539, gm_n46, gm_n63, gm_n50, gm_n9538, in_17);
	nand (gm_n9540, in_20, gm_n62, gm_n47, gm_n9539, in_21);
	nor (gm_n9541, gm_n2300, gm_n52, in_9);
	nand (gm_n9542, gm_n49, gm_n48, gm_n53, gm_n9541, gm_n50);
	nor (gm_n9543, in_17, in_16, gm_n63, gm_n9542, in_18);
	nand (gm_n9544, in_21, gm_n45, in_19, gm_n9543);
	nand (gm_n9545, in_14, in_13, in_12, gm_n9253, in_15);
	nor (gm_n9546, gm_n47, in_17, in_16, gm_n9545, gm_n62);
	nand (gm_n9547, gm_n9546, gm_n71, in_20);
	and (gm_n9548, in_17, in_16, gm_n63, gm_n8736, in_18);
	nand (gm_n9549, in_21, gm_n45, gm_n62, gm_n9548);
	nor (gm_n9550, gm_n49, gm_n48, gm_n53, gm_n1844, in_14);
	nand (gm_n9551, in_17, gm_n46, in_15, gm_n9550, in_18);
	nor (gm_n9552, gm_n71, in_20, gm_n62, gm_n9551);
	nor (gm_n9553, in_13, in_12, gm_n53, gm_n5056, in_14);
	nand (gm_n9554, in_17, in_16, gm_n63, gm_n9553, in_18);
	nor (gm_n9555, gm_n71, in_20, in_19, gm_n9554);
	and (gm_n9556, gm_n49, in_12, gm_n53, gm_n7023, gm_n50);
	nand (gm_n9557, in_17, in_16, in_15, gm_n9556, in_18);
	nor (gm_n9558, gm_n71, in_20, gm_n62, gm_n9557);
	nor (gm_n9559, gm_n63, in_14, gm_n49, gm_n4406, gm_n46);
	nand (gm_n9560, gm_n62, gm_n47, gm_n81, gm_n9559, gm_n45);
	nor (gm_n9561, gm_n9560, gm_n71);
	nand (gm_n9562, in_12, in_11, in_10, gm_n2749, in_13);
	nor (gm_n9563, in_16, in_15, gm_n50, gm_n9562, gm_n81);
	nand (gm_n9564, in_20, gm_n62, gm_n47, gm_n9563, in_21);
	and (gm_n9565, gm_n49, gm_n48, gm_n53, gm_n3885, gm_n50);
	and (gm_n9566, gm_n81, in_16, gm_n63, gm_n9565, in_18);
	nand (gm_n9567, in_21, in_20, in_19, gm_n9566);
	nand (gm_n9568, in_15, gm_n50, gm_n49, gm_n5539, in_16);
	nor (gm_n9569, in_19, in_18, gm_n81, gm_n9568, gm_n45);
	nand (gm_n9570, gm_n9569, in_21);
	nor (gm_n9571, gm_n53, gm_n52, gm_n51, gm_n686, in_12);
	nand (gm_n9572, in_15, gm_n50, gm_n49, gm_n9571, in_16);
	nor (gm_n9573, gm_n62, in_18, in_17, gm_n9572, gm_n45);
	nand (gm_n9574, gm_n9573, gm_n71);
	nand (gm_n9575, gm_n46, gm_n63, gm_n50, gm_n7792, gm_n81);
	nor (gm_n9576, in_20, gm_n62, in_18, gm_n9575, in_21);
	nand (gm_n9577, in_16, in_15, gm_n50, gm_n8277, in_17);
	nor (gm_n9578, gm_n45, in_19, in_18, gm_n9577, gm_n71);
	nand (gm_n9579, in_11, gm_n52, in_9, gm_n5422, in_12);
	nor (gm_n9580, gm_n63, gm_n50, gm_n49, gm_n9579, gm_n46);
	nand (gm_n9581, gm_n62, gm_n47, in_17, gm_n9580, in_20);
	nor (gm_n9582, gm_n9581, gm_n71);
	nor (gm_n9583, gm_n50, in_13, in_12, gm_n2048, in_15);
	nand (gm_n9584, gm_n47, in_17, in_16, gm_n9583, gm_n62);
	nor (gm_n9585, gm_n9584, in_21, in_20);
	nand (gm_n9586, gm_n48, gm_n53, gm_n52, gm_n8629, in_13);
	nor (gm_n9587, in_16, gm_n63, gm_n50, gm_n9586, gm_n81);
	nand (gm_n9588, in_20, in_19, in_18, gm_n9587, gm_n71);
	nor (gm_n9589, in_10, gm_n51, gm_n64, gm_n3718);
	nand (gm_n9590, gm_n49, gm_n48, in_11, gm_n9589, in_14);
	nor (gm_n9591, gm_n81, gm_n46, gm_n63, gm_n9590, gm_n47);
	nand (gm_n9592, in_21, in_20, gm_n62, gm_n9591);
	nand (gm_n9593, in_12, gm_n53, in_10, gm_n654, gm_n49);
	nor (gm_n9594, in_16, gm_n63, in_14, gm_n9593, in_17);
	nand (gm_n9595, in_20, gm_n62, in_18, gm_n9594, in_21);
	nand (gm_n9596, gm_n48, gm_n53, gm_n52, gm_n3069, in_13);
	nor (gm_n9597, in_16, gm_n63, gm_n50, gm_n9596, gm_n81);
	nand (gm_n9598, gm_n45, in_19, gm_n47, gm_n9597, gm_n71);
	nor (gm_n9599, gm_n49, in_12, gm_n53, gm_n6609, gm_n50);
	nand (gm_n9600, gm_n81, gm_n46, in_15, gm_n9599, gm_n47);
	nor (gm_n9601, gm_n71, in_20, in_19, gm_n9600);
	nand (gm_n9602, gm_n53, gm_n52, in_9, gm_n3299);
	nor (gm_n9603, in_14, gm_n49, in_12, gm_n9602, in_15);
	nand (gm_n9604, in_18, in_17, in_16, gm_n9603, gm_n62);
	nor (gm_n9605, gm_n9604, gm_n71, gm_n45);
	and (gm_n9606, in_14, gm_n49, gm_n48, gm_n8138, gm_n63);
	nand (gm_n9607, gm_n47, gm_n81, in_16, gm_n9606, gm_n62);
	nor (gm_n9608, gm_n9607, gm_n71, in_20);
	or (gm_n9609, in_8, gm_n55, in_6, gm_n103, gm_n51);
	nor (gm_n9610, gm_n48, gm_n53, in_10, gm_n9609, gm_n49);
	nand (gm_n9611, gm_n46, in_15, in_14, gm_n9610, in_17);
	nor (gm_n9612, in_20, in_19, gm_n47, gm_n9611, gm_n71);
	and (gm_n9613, gm_n53, gm_n52, gm_n51, gm_n2601, in_12);
	nand (gm_n9614, in_15, in_14, gm_n49, gm_n9613, gm_n46);
	nor (gm_n9615, gm_n62, in_18, gm_n81, gm_n9614, gm_n45);
	nand (gm_n9616, gm_n9615, gm_n71);
	nor (gm_n9617, in_11, gm_n52, gm_n51, gm_n1098, gm_n48);
	nand (gm_n9618, gm_n63, in_14, in_13, gm_n9617, in_16);
	nor (gm_n9619, in_19, gm_n47, in_17, gm_n9618, gm_n45);
	nand (gm_n9620, gm_n9619, in_21);
	nor (gm_n9621, gm_n51, in_8, gm_n55, gm_n259, in_10);
	nand (gm_n9622, in_13, in_12, gm_n53, gm_n9621, gm_n50);
	nor (gm_n9623, gm_n81, in_16, in_15, gm_n9622, in_18);
	nand (gm_n9624, gm_n71, gm_n45, in_19, gm_n9623);
	nand (gm_n9625, in_15, gm_n50, gm_n49, gm_n6164, in_16);
	nor (gm_n9626, gm_n62, in_18, gm_n81, gm_n9625, in_20);
	nand (gm_n9627, gm_n9626, gm_n71);
	nor (gm_n9628, gm_n49, gm_n48, in_11, gm_n4410, in_14);
	nand (gm_n9629, in_17, gm_n46, in_15, gm_n9628, in_18);
	nor (gm_n9630, gm_n71, in_20, gm_n62, gm_n9629);
	nor (gm_n9631, in_12, in_11, gm_n52, gm_n1398, gm_n49);
	nand (gm_n9632, gm_n46, gm_n63, gm_n50, gm_n9631, gm_n81);
	nor (gm_n9633, gm_n45, in_19, gm_n47, gm_n9632, gm_n71);
	nor (gm_n9634, in_13, gm_n48, gm_n53, gm_n2677, in_14);
	nand (gm_n9635, gm_n81, in_16, gm_n63, gm_n9634, in_18);
	nor (gm_n9636, gm_n71, gm_n45, in_19, gm_n9635);
	nor (gm_n9637, gm_n48, in_11, gm_n52, gm_n2327, gm_n49);
	nand (gm_n9638, gm_n46, in_15, gm_n50, gm_n9637, gm_n81);
	nor (gm_n9639, gm_n45, gm_n62, gm_n47, gm_n9638, gm_n71);
	nor (gm_n9640, in_9, gm_n64, gm_n55, gm_n279, gm_n52);
	nand (gm_n9641, gm_n49, in_12, gm_n53, gm_n9640, gm_n50);
	nor (gm_n9642, in_17, in_16, gm_n63, gm_n9641, gm_n47);
	nand (gm_n9643, in_21, in_20, gm_n62, gm_n9642);
	nand (gm_n9644, in_13, in_12, gm_n53, gm_n1257, gm_n50);
	nor (gm_n9645, gm_n81, gm_n46, gm_n63, gm_n9644, gm_n47);
	nand (gm_n9646, in_21, in_20, gm_n62, gm_n9645);
	nand (gm_n9647, gm_n53, gm_n52, in_9, gm_n194, gm_n48);
	nor (gm_n9648, gm_n9647, gm_n49);
	and (gm_n9649, in_16, in_15, in_14, gm_n9648, gm_n81);
	nand (gm_n9650, gm_n45, in_19, gm_n47, gm_n9649, gm_n71);
	nand (gm_n9651, in_15, gm_n50, in_13, gm_n4860, in_16);
	nor (gm_n9652, gm_n62, gm_n47, gm_n81, gm_n9651, in_20);
	nand (gm_n9653, gm_n9652, gm_n71);
	and (gm_n9654, gm_n48, gm_n53, gm_n52, gm_n2877, in_13);
	nand (gm_n9655, in_16, gm_n63, in_14, gm_n9654, gm_n81);
	nor (gm_n9656, in_20, gm_n62, in_18, gm_n9655, gm_n71);
	nor (gm_n9657, gm_n48, in_11, gm_n52, gm_n7227, in_13);
	nand (gm_n9658, in_16, gm_n63, gm_n50, gm_n9657, in_17);
	nor (gm_n9659, in_20, gm_n62, gm_n47, gm_n9658, in_21);
	nand (gm_n9660, in_11, in_10, in_9, gm_n4388, in_12);
	nor (gm_n9661, gm_n63, gm_n50, gm_n49, gm_n9660, in_16);
	nand (gm_n9662, gm_n62, gm_n47, gm_n81, gm_n9661, gm_n45);
	nor (gm_n9663, gm_n9662, in_21);
	nand (gm_n9664, gm_n53, in_10, gm_n51, gm_n1469, in_12);
	nor (gm_n9665, in_15, gm_n50, gm_n49, gm_n9664, gm_n46);
	nand (gm_n9666, in_19, in_18, in_17, gm_n9665, in_20);
	nor (gm_n9667, gm_n9666, in_21);
	nand (gm_n9668, gm_n50, in_13, gm_n48, gm_n5034, gm_n63);
	nor (gm_n9669, gm_n47, in_17, in_16, gm_n9668, in_19);
	nand (gm_n9670, gm_n9669, in_21, gm_n45);
	and (gm_n9671, gm_n48, in_11, in_10, gm_n7115, gm_n49);
	and (gm_n9672, in_16, gm_n63, gm_n50, gm_n9671, in_17);
	nand (gm_n9673, gm_n45, gm_n62, gm_n47, gm_n9672, in_21);
	nor (gm_n9674, gm_n52, in_9, in_8, gm_n3077, in_11);
	nand (gm_n9675, gm_n50, gm_n49, gm_n48, gm_n9674, gm_n63);
	nor (gm_n9676, in_18, in_17, in_16, gm_n9675, in_19);
	nand (gm_n9677, gm_n9676, gm_n71, in_20);
	nor (gm_n9678, in_16, in_15, gm_n50, gm_n2556, in_17);
	nand (gm_n9679, gm_n45, in_19, in_18, gm_n9678, gm_n71);
	nand (gm_n9680, in_11, gm_n52, in_9, gm_n8063, gm_n48);
	nor (gm_n9681, in_15, gm_n50, gm_n49, gm_n9680, gm_n46);
	nand (gm_n9682, gm_n62, gm_n47, gm_n81, gm_n9681, gm_n45);
	nor (gm_n9683, gm_n9682, in_21);
	nor (gm_n9684, in_15, gm_n50, gm_n49, gm_n6508, in_16);
	nand (gm_n9685, in_19, gm_n47, gm_n81, gm_n9684, in_20);
	nor (gm_n9686, gm_n9685, in_21);
	and (gm_n9687, gm_n49, in_12, in_11, gm_n7695, in_14);
	nand (gm_n9688, gm_n81, in_16, in_15, gm_n9687, gm_n47);
	nor (gm_n9689, in_21, gm_n45, gm_n62, gm_n9688);
	nand (gm_n9690, in_10, gm_n51, gm_n64, gm_n1608, gm_n53);
	nor (gm_n9691, in_14, gm_n49, in_12, gm_n9690, in_15);
	nand (gm_n9692, in_18, in_17, gm_n46, gm_n9691, in_19);
	nor (gm_n9693, gm_n9692, in_21, in_20);
	nand (gm_n9694, in_12, gm_n53, in_10, gm_n2415, gm_n49);
	nor (gm_n9695, in_16, gm_n63, in_14, gm_n9694, gm_n81);
	nand (gm_n9696, in_20, gm_n62, gm_n47, gm_n9695, gm_n71);
	and (gm_n9697, gm_n46, gm_n63, in_14, gm_n8664, gm_n81);
	nand (gm_n9698, in_20, in_19, in_18, gm_n9697, in_21);
	nand (gm_n9699, in_14, gm_n49, in_12, gm_n5756, in_15);
	nor (gm_n9700, in_18, in_17, gm_n46, gm_n9699, in_19);
	nand (gm_n9701, gm_n9700, gm_n71, gm_n45);
	and (gm_n9702, in_17, gm_n46, gm_n63, gm_n8709, in_18);
	nand (gm_n9703, gm_n71, gm_n45, in_19, gm_n9702);
	nor (gm_n9704, in_14, gm_n49, in_12, gm_n7619, gm_n63);
	nand (gm_n9705, gm_n47, in_17, in_16, gm_n9704, in_19);
	nor (gm_n9706, gm_n9705, gm_n71, gm_n45);
	nor (gm_n9707, gm_n49, gm_n48, gm_n53, gm_n5272, in_14);
	nand (gm_n9708, gm_n81, in_16, gm_n63, gm_n9707, gm_n47);
	nor (gm_n9709, gm_n71, in_20, in_19, gm_n9708);
	nor (gm_n9710, in_12, in_11, in_10, gm_n3809, gm_n49);
	nand (gm_n9711, in_16, gm_n63, in_14, gm_n9710, gm_n81);
	nor (gm_n9712, in_20, in_19, gm_n47, gm_n9711, gm_n71);
	nor (gm_n9713, in_12, in_11, gm_n52, gm_n228, gm_n49);
	nand (gm_n9714, in_16, in_15, in_14, gm_n9713, in_17);
	nor (gm_n9715, gm_n45, gm_n62, in_18, gm_n9714, gm_n71);
	nand (gm_n9716, in_12, gm_n53, in_10, gm_n696, gm_n49);
	nor (gm_n9717, in_16, gm_n63, gm_n50, gm_n9716, in_17);
	nand (gm_n9718, gm_n45, in_19, gm_n47, gm_n9717, gm_n71);
	nand (gm_n9719, gm_n48, gm_n53, in_10, gm_n6139, in_13);
	nor (gm_n9720, in_16, in_15, gm_n50, gm_n9719, gm_n81);
	nand (gm_n9721, gm_n45, gm_n62, in_18, gm_n9720, gm_n71);
	nor (gm_n9722, gm_n2951, in_9);
	nand (gm_n9723, gm_n48, gm_n53, in_10, gm_n9722, gm_n49);
	nor (gm_n9724, gm_n46, gm_n63, in_14, gm_n9723, in_17);
	nand (gm_n9725, in_20, in_19, gm_n47, gm_n9724, gm_n71);
	and (gm_n9726, gm_n53, gm_n52, in_9, gm_n1293, in_12);
	nand (gm_n9727, gm_n63, gm_n50, gm_n49, gm_n9726, in_16);
	nor (gm_n9728, gm_n62, in_18, in_17, gm_n9727, in_20);
	nand (gm_n9729, gm_n9728, in_21);
	nand (gm_n9730, in_11, gm_n52, in_9, gm_n2047, gm_n48);
	nor (gm_n9731, in_15, in_14, gm_n49, gm_n9730, gm_n46);
	nand (gm_n9732, gm_n62, gm_n47, in_17, gm_n9731, in_20);
	nor (gm_n9733, gm_n9732, gm_n71);
	nor (gm_n9734, gm_n50, in_13, in_12, gm_n7122, in_15);
	nand (gm_n9735, gm_n47, gm_n81, gm_n46, gm_n9734, gm_n62);
	nor (gm_n9736, gm_n9735, gm_n71, gm_n45);
	nand (gm_n9737, gm_n53, gm_n52, gm_n51, gm_n1134, gm_n48);
	nor (gm_n9738, gm_n63, gm_n50, in_13, gm_n9737, gm_n46);
	nand (gm_n9739, in_19, gm_n47, gm_n81, gm_n9738, gm_n45);
	nor (gm_n9740, gm_n9739, gm_n71);
	nor (gm_n9741, gm_n50, gm_n49, gm_n48, gm_n9690, gm_n63);
	nand (gm_n9742, in_18, in_17, in_16, gm_n9741, gm_n62);
	nor (gm_n9743, gm_n9742, in_21, in_20);
	nor (gm_n9744, gm_n46, gm_n63, gm_n50, gm_n8215, gm_n81);
	nand (gm_n9745, gm_n45, gm_n62, gm_n47, gm_n9744, gm_n71);
	and (gm_n9746, gm_n658, gm_n51);
	nand (gm_n9747, gm_n48, gm_n53, gm_n52, gm_n9746, gm_n49);
	nor (gm_n9748, in_16, in_15, gm_n50, gm_n9747, gm_n81);
	nand (gm_n9749, gm_n45, gm_n62, in_18, gm_n9748, gm_n71);
	nand (gm_n9750, gm_n49, gm_n48, gm_n53, gm_n8854, gm_n50);
	nor (gm_n9751, in_17, gm_n46, in_15, gm_n9750, gm_n47);
	nand (gm_n9752, gm_n71, in_20, gm_n62, gm_n9751);
	nand (gm_n9753, gm_n50, gm_n49, gm_n48, gm_n3805, gm_n63);
	nor (gm_n9754, gm_n47, in_17, gm_n46, gm_n9753, gm_n62);
	nand (gm_n9755, gm_n9754, gm_n71, in_20);
	nor (gm_n9756, gm_n49, in_12, in_11, gm_n8152, in_14);
	nand (gm_n9757, gm_n81, gm_n46, in_15, gm_n9756, gm_n47);
	nor (gm_n9758, in_21, gm_n45, gm_n62, gm_n9757);
	nand (gm_n9759, in_16, gm_n63, gm_n50, gm_n1281, gm_n81);
	nor (gm_n9760, gm_n45, in_19, gm_n47, gm_n9759, gm_n71);
	nand (gm_n9761, in_11, in_10, gm_n51, gm_n114, in_12);
	nor (gm_n9762, gm_n63, in_14, gm_n49, gm_n9761, gm_n46);
	nand (gm_n9763, in_19, gm_n47, gm_n81, gm_n9762, gm_n45);
	nor (gm_n9764, gm_n9763, gm_n71);
	or (gm_n9765, in_11, gm_n52, in_9, gm_n3340, in_12);
	nor (gm_n9766, gm_n63, gm_n50, in_13, gm_n9765, in_16);
	nand (gm_n9767, in_19, gm_n47, in_17, gm_n9766, in_20);
	nor (gm_n9768, gm_n9767, gm_n71);
	nor (gm_n9769, in_9, in_8, gm_n55, gm_n525, in_10);
	nand (gm_n9770, in_13, gm_n48, gm_n53, gm_n9769, gm_n50);
	nor (gm_n9771, gm_n81, in_16, gm_n63, gm_n9770, in_18);
	nand (gm_n9772, gm_n71, in_20, in_19, gm_n9771);
	and (gm_n9773, in_16, gm_n63, gm_n50, gm_n6136, gm_n81);
	nand (gm_n9774, gm_n45, in_19, in_18, gm_n9773, gm_n71);
	nand (gm_n9775, gm_n50, in_13, gm_n48, gm_n2316, in_15);
	nor (gm_n9776, gm_n47, in_17, in_16, gm_n9775, gm_n62);
	nand (gm_n9777, gm_n9776, gm_n71, in_20);
	nor (gm_n9778, gm_n53, gm_n52, gm_n51, gm_n520);
	nand (gm_n9779, in_14, in_13, in_12, gm_n9778, gm_n63);
	nor (gm_n9780, in_18, in_17, gm_n46, gm_n9779, in_19);
	nand (gm_n9781, gm_n9780, in_21, in_20);
	nand (gm_n9782, gm_n53, gm_n52, in_9, gm_n5340, gm_n48);
	nor (gm_n9783, in_15, in_14, in_13, gm_n9782, gm_n46);
	nand (gm_n9784, in_19, in_18, in_17, gm_n9783, gm_n45);
	nor (gm_n9785, gm_n9784, gm_n71);
	and (gm_n9786, gm_n48, in_11, in_10, gm_n5375, in_13);
	nand (gm_n9787, gm_n46, gm_n63, in_14, gm_n9786, in_17);
	nor (gm_n9788, in_20, in_19, in_18, gm_n9787, in_21);
	nand (gm_n9789, gm_n46, gm_n63, gm_n50, gm_n4476, in_17);
	nor (gm_n9790, in_20, in_19, gm_n47, gm_n9789, in_21);
	or (gm_n9791, in_13, gm_n48, gm_n53, gm_n7096, gm_n50);
	or (gm_n9792, in_17, in_16, gm_n63, gm_n9791, gm_n47);
	nor (gm_n9793, gm_n71, in_20, in_19, gm_n9792);
	nand (gm_n9794, gm_n48, gm_n53, gm_n52, gm_n2482, gm_n49);
	nor (gm_n9795, gm_n46, gm_n63, gm_n50, gm_n9794, gm_n81);
	nand (gm_n9796, gm_n45, gm_n62, in_18, gm_n9795, in_21);
	and (gm_n9797, gm_n52, in_9, gm_n64, gm_n1608, in_11);
	nand (gm_n9798, gm_n50, gm_n49, in_12, gm_n9797, gm_n63);
	nor (gm_n9799, in_18, gm_n81, gm_n46, gm_n9798, gm_n62);
	nand (gm_n9800, gm_n9799, gm_n71, in_20);
	nor (gm_n9801, gm_n62, in_18, in_17, gm_n6379, in_20);
	nand (gm_n9802, gm_n9801, in_21);
	nand (gm_n9803, gm_n2446, gm_n49);
	nor (gm_n9804, gm_n46, in_15, in_14, gm_n9803, in_17);
	nand (gm_n9805, in_20, gm_n62, in_18, gm_n9804, in_21);
	or (gm_n9806, in_10, in_9, in_8, gm_n478, gm_n53);
	nor (gm_n9807, gm_n50, gm_n49, in_12, gm_n9806, gm_n63);
	nand (gm_n9808, gm_n47, in_17, gm_n46, gm_n9807, in_19);
	nor (gm_n9809, gm_n9808, in_21, in_20);
	nand (gm_n9810, gm_n53, gm_n52, in_9, gm_n1178, in_12);
	nor (gm_n9811, gm_n63, gm_n50, in_13, gm_n9810, gm_n46);
	nand (gm_n9812, in_19, gm_n47, gm_n81, gm_n9811, gm_n45);
	nor (gm_n9813, gm_n9812, in_21);
	nand (gm_n9814, gm_n46, gm_n63, gm_n50, gm_n360, in_17);
	nor (gm_n9815, gm_n45, gm_n62, in_18, gm_n9814, gm_n71);
	and (gm_n9816, gm_n49, in_12, gm_n53, gm_n1652, in_14);
	nand (gm_n9817, gm_n81, gm_n46, gm_n63, gm_n9816, gm_n47);
	nor (gm_n9818, in_21, in_20, gm_n62, gm_n9817);
	nand (gm_n9819, gm_n49, in_12, in_11, gm_n8854, gm_n50);
	nor (gm_n9820, in_17, gm_n46, in_15, gm_n9819, in_18);
	nand (gm_n9821, in_21, gm_n45, in_19, gm_n9820);
	nand (gm_n9822, gm_n48, in_11, gm_n52, gm_n3611, in_13);
	nor (gm_n9823, gm_n46, gm_n63, in_14, gm_n9822, gm_n81);
	nand (gm_n9824, gm_n45, gm_n62, in_18, gm_n9823, gm_n71);
	nor (gm_n9825, gm_n53, gm_n52, in_9, gm_n2902, gm_n48);
	nand (gm_n9826, in_15, gm_n50, in_13, gm_n9825, gm_n46);
	nor (gm_n9827, in_19, in_18, in_17, gm_n9826, gm_n45);
	nand (gm_n9828, gm_n9827, gm_n71);
	or (gm_n9829, in_14, gm_n49, in_12, gm_n7309, in_15);
	nor (gm_n9830, gm_n47, in_17, gm_n46, gm_n9829, in_19);
	nand (gm_n9831, gm_n9830, in_21, gm_n45);
	and (gm_n9832, gm_n49, gm_n48, in_11, gm_n9436, gm_n50);
	nand (gm_n9833, gm_n81, gm_n46, gm_n63, gm_n9832, in_18);
	nor (gm_n9834, gm_n71, gm_n45, in_19, gm_n9833);
	nor (gm_n9835, in_12, gm_n53, in_10, gm_n1621, gm_n49);
	nand (gm_n9836, gm_n46, in_15, gm_n50, gm_n9835, gm_n81);
	nor (gm_n9837, gm_n45, in_19, in_18, gm_n9836, in_21);
	nand (gm_n9838, gm_n53, gm_n52, gm_n51, gm_n717);
	nor (gm_n9839, gm_n50, in_13, in_12, gm_n9838, gm_n63);
	nand (gm_n9840, in_18, gm_n81, in_16, gm_n9839, in_19);
	nor (gm_n9841, gm_n9840, gm_n71, in_20);
	nand (gm_n9842, in_17, in_16, gm_n63, gm_n2802, in_18);
	nor (gm_n9843, in_21, gm_n45, in_19, gm_n9842);
	nand (gm_n9844, gm_n63, gm_n50, gm_n49, gm_n6992, gm_n46);
	nor (gm_n9845, in_19, gm_n47, gm_n81, gm_n9844, in_20);
	nand (gm_n9846, gm_n9845, in_21);
	and (gm_n9847, in_16, gm_n63, in_14, gm_n5550, gm_n81);
	nand (gm_n9848, gm_n45, gm_n62, gm_n47, gm_n9847, gm_n71);
	nor (gm_n9849, gm_n46, gm_n63, in_14, gm_n2928, gm_n81);
	nand (gm_n9850, in_20, in_19, in_18, gm_n9849, in_21);
	nand (gm_n9851, in_14, in_13, gm_n48, gm_n396, in_15);
	nor (gm_n9852, in_18, in_17, in_16, gm_n9851, gm_n62);
	nand (gm_n9853, gm_n9852, gm_n71, in_20);
	nand (gm_n9854, gm_n53, in_10, gm_n51, gm_n3091, gm_n48);
	nor (gm_n9855, gm_n63, gm_n50, gm_n49, gm_n9854, gm_n46);
	nand (gm_n9856, gm_n62, in_18, in_17, gm_n9855, gm_n45);
	nor (gm_n9857, gm_n9856, gm_n71);
	nand (gm_n9858, gm_n46, gm_n63, in_14, gm_n4644, in_17);
	nor (gm_n9859, in_20, gm_n62, in_18, gm_n9858, gm_n71);
	nand (gm_n9860, in_9, in_8, gm_n55, gm_n66, in_10);
	nor (gm_n9861, gm_n49, in_12, gm_n53, gm_n9860, gm_n50);
	nand (gm_n9862, gm_n81, in_16, gm_n63, gm_n9861, in_18);
	nor (gm_n9863, gm_n71, gm_n45, in_19, gm_n9862);
	and (gm_n9864, gm_n48, in_11, gm_n52, gm_n1201, gm_n49);
	nand (gm_n9865, gm_n46, gm_n63, gm_n50, gm_n9864, gm_n81);
	nor (gm_n9866, gm_n45, in_19, in_18, gm_n9865, gm_n71);
	nand (gm_n9867, in_8, gm_n55, in_6, gm_n2640, gm_n51);
	or (gm_n9868, gm_n48, in_11, gm_n52, gm_n9867, in_13);
	nor (gm_n9869, in_16, in_15, gm_n50, gm_n9868, in_17);
	nand (gm_n9870, gm_n45, in_19, in_18, gm_n9869, in_21);
	nand (gm_n9871, in_13, in_12, in_11, gm_n3082, gm_n50);
	nor (gm_n9872, in_17, in_16, in_15, gm_n9871, gm_n47);
	nand (gm_n9873, gm_n71, gm_n45, gm_n62, gm_n9872);
	or (gm_n9874, in_12, gm_n53, gm_n52, gm_n5605, in_13);
	nor (gm_n9875, in_16, gm_n63, gm_n50, gm_n9874, gm_n81);
	nand (gm_n9876, gm_n45, in_19, gm_n47, gm_n9875, gm_n71);
	and (gm_n9877, in_8, gm_n55, gm_n82, gm_n374, gm_n51);
	nand (gm_n9878, gm_n48, in_11, gm_n52, gm_n9877, gm_n49);
	nor (gm_n9879, gm_n46, in_15, gm_n50, gm_n9878, in_17);
	nand (gm_n9880, gm_n45, in_19, in_18, gm_n9879, gm_n71);
	nor (gm_n9881, in_15, gm_n50, in_13, gm_n7033, gm_n46);
	nand (gm_n9882, in_19, gm_n47, gm_n81, gm_n9881, in_20);
	nor (gm_n9883, gm_n9882, gm_n71);
	nand (gm_n9884, in_16, gm_n63, gm_n50, gm_n7792, gm_n81);
	nor (gm_n9885, in_20, in_19, in_18, gm_n9884, in_21);
	nand (gm_n9886, gm_n53, in_10, in_9, gm_n4168, gm_n48);
	nor (gm_n9887, gm_n63, gm_n50, gm_n49, gm_n9886, in_16);
	nand (gm_n9888, gm_n62, in_18, gm_n81, gm_n9887, in_20);
	nor (gm_n9889, gm_n9888, gm_n71);
	nand (gm_n9890, in_16, gm_n63, in_14, gm_n3578, gm_n81);
	nor (gm_n9891, in_20, in_19, gm_n47, gm_n9890, gm_n71);
	nand (gm_n9892, in_13, gm_n48, gm_n53, gm_n5601, gm_n50);
	nor (gm_n9893, in_17, in_16, gm_n63, gm_n9892, in_18);
	nand (gm_n9894, gm_n71, in_20, in_19, gm_n9893);
	nand (gm_n9895, in_14, in_13, gm_n48, gm_n8732, in_15);
	nor (gm_n9896, in_18, in_17, in_16, gm_n9895, gm_n62);
	nand (gm_n9897, gm_n9896, gm_n71, in_20);
	and (gm_n9898, gm_n52, gm_n51, gm_n64, gm_n4213, in_11);
	nand (gm_n9899, gm_n50, gm_n49, gm_n48, gm_n9898, gm_n63);
	nor (gm_n9900, in_18, in_17, gm_n46, gm_n9899, in_19);
	nand (gm_n9901, gm_n9900, gm_n71, gm_n45);
	and (gm_n9902, in_9, in_8, in_7, gm_n136);
	nand (gm_n9903, in_12, in_11, in_10, gm_n9902, gm_n49);
	nor (gm_n9904, in_16, gm_n63, gm_n50, gm_n9903, gm_n81);
	nand (gm_n9905, in_20, gm_n62, gm_n47, gm_n9904, gm_n71);
	or (gm_n9906, in_16, in_15, gm_n50, gm_n5700, in_17);
	nor (gm_n9907, in_20, gm_n62, gm_n47, gm_n9906, gm_n71);
	and (gm_n9908, gm_n48, gm_n53, gm_n52, gm_n912, in_13);
	nand (gm_n9909, in_16, in_15, in_14, gm_n9908, in_17);
	nor (gm_n9910, in_20, gm_n62, gm_n47, gm_n9909, gm_n71);
	nand (gm_n9911, gm_n52, in_9, gm_n64, gm_n2708, gm_n53);
	nor (gm_n9912, gm_n50, in_13, gm_n48, gm_n9911, gm_n63);
	nand (gm_n9913, gm_n47, in_17, in_16, gm_n9912, gm_n62);
	nor (gm_n9914, gm_n9913, gm_n71, gm_n45);
	nor (gm_n9915, gm_n50, in_13, in_12, gm_n701, in_15);
	nand (gm_n9916, in_18, gm_n81, in_16, gm_n9915, in_19);
	nor (gm_n9917, gm_n9916, in_21, in_20);
	nor (gm_n9918, in_18, in_17, in_16, gm_n5694, in_19);
	nand (gm_n9919, gm_n9918, gm_n71, in_20);
	nor (gm_n9920, in_11, in_10, in_9, gm_n5263, gm_n48);
	nand (gm_n9921, gm_n63, in_14, gm_n49, gm_n9920, gm_n46);
	nor (gm_n9922, gm_n62, in_18, in_17, gm_n9921, in_20);
	nand (gm_n9923, gm_n9922, gm_n71);
	nand (gm_n9924, gm_n49, gm_n48, in_11, gm_n4120, gm_n50);
	nor (gm_n9925, gm_n81, gm_n46, in_15, gm_n9924, in_18);
	nand (gm_n9926, in_21, gm_n45, in_19, gm_n9925);
	nor (gm_n9927, gm_n52, in_9, in_8, gm_n3174, gm_n53);
	nand (gm_n9928, gm_n50, in_13, gm_n48, gm_n9927, gm_n63);
	nor (gm_n9929, gm_n47, in_17, gm_n46, gm_n9928, in_19);
	nand (gm_n9930, gm_n9929, in_21, gm_n45);
	nor (gm_n9931, in_12, in_11, gm_n52, gm_n4692, in_13);
	nand (gm_n9932, gm_n46, gm_n63, in_14, gm_n9931, gm_n81);
	nor (gm_n9933, gm_n45, in_19, in_18, gm_n9932, gm_n71);
	nand (gm_n9934, gm_n62, in_18, in_17, gm_n4162, in_20);
	nor (gm_n9935, gm_n9934, gm_n71);
	nand (gm_n9936, gm_n46, in_15, in_14, gm_n3641, in_17);
	nor (gm_n9937, in_20, gm_n62, in_18, gm_n9936, in_21);
	nor (gm_n9938, in_12, in_11, in_10, gm_n531, gm_n49);
	nand (gm_n9939, gm_n46, gm_n63, gm_n50, gm_n9938, in_17);
	nor (gm_n9940, in_20, in_19, gm_n47, gm_n9939, gm_n71);
	nand (gm_n9941, gm_n50, in_13, gm_n48, gm_n8651, gm_n63);
	nor (gm_n9942, gm_n47, in_17, in_16, gm_n9941, gm_n62);
	nand (gm_n9943, gm_n9942, gm_n71, gm_n45);
	nand (gm_n9944, in_7, in_6, gm_n72, gm_n89, gm_n64);
	nor (gm_n9945, in_11, gm_n52, in_9, gm_n9944);
	nand (gm_n9946, gm_n50, gm_n49, gm_n48, gm_n9945, in_15);
	nor (gm_n9947, in_18, gm_n81, in_16, gm_n9946, gm_n62);
	nand (gm_n9948, gm_n9947, gm_n71, gm_n45);
	nand (gm_n9949, gm_n63, gm_n50, in_13, gm_n2565, in_16);
	nor (gm_n9950, in_19, in_18, gm_n81, gm_n9949, in_20);
	nand (gm_n9951, gm_n9950, in_21);
	nand (gm_n9952, in_14, gm_n49, in_12, gm_n6080, in_15);
	nor (gm_n9953, in_18, gm_n81, in_16, gm_n9952, in_19);
	nand (gm_n9954, gm_n9953, in_21, gm_n45);
	nor (gm_n9955, gm_n81, gm_n46, in_15, gm_n9791, gm_n47);
	nand (gm_n9956, in_21, in_20, gm_n62, gm_n9955);
	nand (gm_n9957, gm_n9951, gm_n9948, gm_n9943, gm_n9956, gm_n9954);
	nor (gm_n9958, gm_n9937, gm_n9935, gm_n9933, gm_n9957, gm_n9940);
	nand (gm_n9959, gm_n9926, gm_n9923, gm_n9919, gm_n9958, gm_n9930);
	nor (gm_n9960, gm_n9914, gm_n9910, gm_n9907, gm_n9959, gm_n9917);
	nand (gm_n9961, gm_n9901, gm_n9897, gm_n9894, gm_n9960, gm_n9905);
	nor (gm_n9962, gm_n9889, gm_n9885, gm_n9883, gm_n9961, gm_n9891);
	nand (gm_n9963, gm_n9876, gm_n9873, gm_n9870, gm_n9962, gm_n9880);
	nor (gm_n9964, gm_n9863, gm_n9859, gm_n9857, gm_n9963, gm_n9866);
	nand (gm_n9965, gm_n9850, gm_n9848, gm_n9846, gm_n9964, gm_n9853);
	nor (gm_n9966, gm_n9841, gm_n9837, gm_n9834, gm_n9965, gm_n9843);
	nand (gm_n9967, gm_n9828, gm_n9824, gm_n9821, gm_n9966, gm_n9831);
	nor (gm_n9968, gm_n9815, gm_n9813, gm_n9809, gm_n9967, gm_n9818);
	nand (gm_n9969, gm_n9802, gm_n9800, gm_n9796, gm_n9968, gm_n9805);
	nor (gm_n9970, gm_n9790, gm_n9788, gm_n9785, gm_n9969, gm_n9793);
	nand (gm_n9971, gm_n9777, gm_n9774, gm_n9772, gm_n9970, gm_n9781);
	nor (gm_n9972, gm_n9764, gm_n9760, gm_n9758, gm_n9971, gm_n9768);
	nand (gm_n9973, gm_n9752, gm_n9749, gm_n9745, gm_n9972, gm_n9755);
	nor (gm_n9974, gm_n9740, gm_n9736, gm_n9733, gm_n9973, gm_n9743);
	nand (gm_n9975, gm_n9725, gm_n9721, gm_n9718, gm_n9974, gm_n9729);
	nor (gm_n9976, gm_n9712, gm_n9709, gm_n9706, gm_n9975, gm_n9715);
	nand (gm_n9977, gm_n9701, gm_n9698, gm_n9696, gm_n9976, gm_n9703);
	nor (gm_n9978, gm_n9689, gm_n9686, gm_n9683, gm_n9977, gm_n9693);
	nand (gm_n9979, gm_n9677, gm_n9673, gm_n9670, gm_n9978, gm_n9679);
	nor (gm_n9980, gm_n9663, gm_n9659, gm_n9656, gm_n9979, gm_n9667);
	nand (gm_n9981, gm_n9650, gm_n9646, gm_n9643, gm_n9980, gm_n9653);
	nor (gm_n9982, gm_n9636, gm_n9633, gm_n9630, gm_n9981, gm_n9639);
	nand (gm_n9983, gm_n9624, gm_n9620, gm_n9616, gm_n9982, gm_n9627);
	nor (gm_n9984, gm_n9608, gm_n9605, gm_n9601, gm_n9983, gm_n9612);
	nand (gm_n9985, gm_n9595, gm_n9592, gm_n9588, gm_n9984, gm_n9598);
	nor (gm_n9986, gm_n9582, gm_n9578, gm_n9576, gm_n9985, gm_n9585);
	nand (gm_n9987, gm_n9570, gm_n9567, gm_n9564, gm_n9986, gm_n9574);
	nor (gm_n9988, gm_n9558, gm_n9555, gm_n9552, gm_n9987, gm_n9561);
	nand (gm_n9989, gm_n9547, gm_n9544, gm_n9540, gm_n9988, gm_n9549);
	nor (gm_n9990, gm_n9533, gm_n9530, gm_n9528, gm_n9989, gm_n9536);
	nand (gm_n9991, gm_n9521, gm_n9517, gm_n9514, gm_n9990, gm_n9525);
	nor (gm_n9992, gm_n9508, gm_n9505, gm_n9501, gm_n9991, gm_n9511);
	nand (gm_n9993, gm_n9495, gm_n9491, gm_n9488, gm_n9992, gm_n9498);
	nor (out_16, gm_n9993, gm_n9484);
	nor (gm_n9995, gm_n48, in_11, in_10, gm_n1524, in_13);
	nand (gm_n9996, in_16, gm_n63, gm_n50, gm_n9995, in_17);
	nor (gm_n9997, in_20, gm_n62, gm_n47, gm_n9996, gm_n71);
	nor (gm_n9998, gm_n50, gm_n49, gm_n48, gm_n5689, gm_n63);
	nand (gm_n9999, in_18, in_17, gm_n46, gm_n9998, in_19);
	nor (gm_n10000, gm_n9999, in_21, in_20);
	nor (gm_n10001, gm_n48, gm_n53, in_10, gm_n4547, in_13);
	nand (gm_n10002, gm_n46, gm_n63, gm_n50, gm_n10001, gm_n81);
	nor (gm_n10003, in_20, in_19, gm_n47, gm_n10002, gm_n71);
	nand (gm_n10004, gm_n49, gm_n48, gm_n53, gm_n1889, in_14);
	nor (gm_n10005, in_17, gm_n46, gm_n63, gm_n10004, in_18);
	nand (gm_n10006, gm_n71, gm_n45, gm_n62, gm_n10005);
	nand (gm_n10007, in_13, gm_n48, in_11, gm_n5048, gm_n50);
	nor (gm_n10008, in_17, gm_n46, gm_n63, gm_n10007, in_18);
	nand (gm_n10009, in_21, in_20, in_19, gm_n10008);
	and (gm_n10010, gm_n49, in_12, in_11, gm_n224);
	and (gm_n10011, in_16, in_15, gm_n50, gm_n10010, in_17);
	nand (gm_n10012, gm_n45, in_19, in_18, gm_n10011, gm_n71);
	nand (gm_n10013, gm_n48, gm_n53, in_10, gm_n4984, in_13);
	nor (gm_n10014, gm_n46, gm_n63, gm_n50, gm_n10013, in_17);
	nand (gm_n10015, gm_n45, gm_n62, gm_n47, gm_n10014, in_21);
	nand (gm_n10016, in_16, in_15, gm_n50, gm_n1530, in_17);
	nor (gm_n10017, in_20, gm_n62, gm_n47, gm_n10016, gm_n71);
	nand (gm_n10018, in_17, in_16, in_15, gm_n5330, gm_n47);
	nor (gm_n10019, gm_n71, gm_n45, in_19, gm_n10018);
	and (gm_n10020, gm_n50, in_13, in_12, gm_n7246, gm_n63);
	nand (gm_n10021, gm_n47, gm_n81, in_16, gm_n10020, gm_n62);
	nor (gm_n10022, gm_n10021, in_21, gm_n45);
	nand (gm_n10023, in_16, gm_n63, in_14, gm_n4344, gm_n81);
	nor (gm_n10024, gm_n45, gm_n62, in_18, gm_n10023, gm_n71);
	nor (gm_n10025, gm_n53, in_10, gm_n51, gm_n751);
	nand (gm_n10026, in_14, in_13, gm_n48, gm_n10025, gm_n63);
	nor (gm_n10027, gm_n47, in_17, in_16, gm_n10026, gm_n62);
	nand (gm_n10028, gm_n10027, in_21, in_20);
	nor (gm_n10029, in_9, gm_n64, in_7, gm_n1256, gm_n52);
	nand (gm_n10030, gm_n49, in_12, in_11, gm_n10029, in_14);
	nor (gm_n10031, in_17, gm_n46, in_15, gm_n10030, gm_n47);
	nand (gm_n10032, in_21, gm_n45, gm_n62, gm_n10031);
	nand (gm_n10033, in_14, in_13, in_12, gm_n5351, in_15);
	nor (gm_n10034, gm_n47, in_17, gm_n46, gm_n10033, gm_n62);
	nand (gm_n10035, gm_n10034, gm_n71, gm_n45);
	nand (gm_n10036, in_13, gm_n48, in_11, gm_n3420, in_14);
	nor (gm_n10037, gm_n81, gm_n46, in_15, gm_n10036, gm_n47);
	nand (gm_n10038, in_21, gm_n45, in_19, gm_n10037);
	and (gm_n10039, in_14, gm_n49, in_12, gm_n2881, gm_n63);
	nand (gm_n10040, in_18, gm_n81, in_16, gm_n10039, in_19);
	nor (gm_n10041, gm_n10040, in_21, in_20);
	or (gm_n10042, gm_n131, gm_n51);
	nor (gm_n10043, in_12, in_11, gm_n52, gm_n10042, in_13);
	nand (gm_n10044, in_16, in_15, in_14, gm_n10043, gm_n81);
	nor (gm_n10045, gm_n45, in_19, in_18, gm_n10044, gm_n71);
	nor (gm_n10046, gm_n45, in_19, in_18, gm_n4672, in_21);
	nor (gm_n10047, gm_n48, gm_n53, gm_n52, gm_n2841, gm_n49);
	nand (gm_n10048, gm_n46, in_15, in_14, gm_n10047, gm_n81);
	nor (gm_n10049, in_20, gm_n62, in_18, gm_n10048, gm_n71);
	nand (gm_n10050, gm_n48, in_11, gm_n52, gm_n7115, gm_n49);
	nor (gm_n10051, in_16, in_15, in_14, gm_n10050, in_17);
	nand (gm_n10052, in_20, gm_n62, gm_n47, gm_n10051, gm_n71);
	nand (gm_n10053, gm_n48, in_11, gm_n52, gm_n1413, gm_n49);
	nor (gm_n10054, in_16, in_15, in_14, gm_n10053, in_17);
	nand (gm_n10055, in_20, in_19, in_18, gm_n10054, in_21);
	nand (gm_n10056, gm_n48, gm_n53, in_10, gm_n2729, gm_n49);
	nor (gm_n10057, in_16, in_15, in_14, gm_n10056, gm_n81);
	nand (gm_n10058, gm_n45, in_19, in_18, gm_n10057, in_21);
	nand (gm_n10059, in_15, in_14, in_13, gm_n6426, in_16);
	nor (gm_n10060, in_19, in_18, gm_n81, gm_n10059, gm_n45);
	nand (gm_n10061, gm_n10060, in_21);
	nand (gm_n10062, in_11, in_10, gm_n51, gm_n5668, in_12);
	nor (gm_n10063, gm_n63, in_14, in_13, gm_n10062, gm_n46);
	nand (gm_n10064, in_19, in_18, in_17, gm_n10063, gm_n45);
	nor (gm_n10065, gm_n10064, in_21);
	nor (gm_n10066, gm_n48, gm_n53, in_10, gm_n264, gm_n49);
	nand (gm_n10067, in_16, in_15, gm_n50, gm_n10066, gm_n81);
	nor (gm_n10068, gm_n45, gm_n62, in_18, gm_n10067, in_21);
	and (gm_n10069, gm_n48, gm_n53, gm_n52, gm_n696, gm_n49);
	nand (gm_n10070, in_16, in_15, gm_n50, gm_n10069, gm_n81);
	nor (gm_n10071, in_20, in_19, in_18, gm_n10070, gm_n71);
	nor (gm_n10072, gm_n48, in_11, gm_n52, gm_n639, gm_n49);
	nand (gm_n10073, gm_n46, in_15, gm_n50, gm_n10072, gm_n81);
	nor (gm_n10074, in_20, gm_n62, gm_n47, gm_n10073, in_21);
	or (gm_n10075, gm_n48, gm_n53, gm_n52, gm_n6760, gm_n49);
	nor (gm_n10076, gm_n46, in_15, in_14, gm_n10075, gm_n81);
	nand (gm_n10077, gm_n45, in_19, gm_n47, gm_n10076, gm_n71);
	nand (gm_n10078, gm_n49, gm_n48, gm_n53, gm_n4813, in_14);
	nor (gm_n10079, gm_n81, in_16, in_15, gm_n10078, in_18);
	nand (gm_n10080, in_21, in_20, in_19, gm_n10079);
	nor (gm_n10081, in_11, gm_n52, gm_n51, gm_n2266, gm_n48);
	nand (gm_n10082, in_15, gm_n50, gm_n49, gm_n10081, in_16);
	nor (gm_n10083, gm_n62, gm_n47, gm_n81, gm_n10082, in_20);
	nand (gm_n10084, gm_n10083, gm_n71);
	nor (gm_n10085, in_11, gm_n52, in_9, gm_n4314, in_12);
	and (gm_n10086, gm_n63, gm_n50, gm_n49, gm_n10085, in_16);
	and (gm_n10087, in_19, in_18, gm_n81, gm_n10086, in_20);
	nand (gm_n10088, gm_n10087, in_21);
	and (gm_n10089, in_12, in_11, in_10, gm_n1671, gm_n49);
	nand (gm_n10090, in_16, in_15, in_14, gm_n10089, gm_n81);
	nor (gm_n10091, gm_n45, gm_n62, in_18, gm_n10090, gm_n71);
	and (gm_n10092, gm_n53, in_10, gm_n51, gm_n1142, in_12);
	and (gm_n10093, in_15, gm_n50, in_13, gm_n10092, gm_n46);
	nand (gm_n10094, in_19, gm_n47, gm_n81, gm_n10093, in_20);
	nor (gm_n10095, gm_n10094, gm_n71);
	and (gm_n10096, gm_n48, gm_n53, in_10, gm_n1332, in_13);
	nand (gm_n10097, in_16, gm_n63, gm_n50, gm_n10096, in_17);
	nor (gm_n10098, in_20, in_19, in_18, gm_n10097, in_21);
	nor (gm_n10099, in_14, in_13, gm_n48, gm_n1320, in_15);
	nand (gm_n10100, in_18, gm_n81, in_16, gm_n10099, in_19);
	nor (gm_n10101, gm_n10100, gm_n71, gm_n45);
	nand (gm_n10102, in_13, gm_n48, gm_n53, gm_n7103, in_14);
	nor (gm_n10103, gm_n81, in_16, gm_n63, gm_n10102, in_18);
	nand (gm_n10104, in_21, gm_n45, gm_n62, gm_n10103);
	nor (gm_n10105, in_16, gm_n63, in_14, gm_n2406, gm_n81);
	nand (gm_n10106, in_20, gm_n62, gm_n47, gm_n10105, gm_n71);
	or (gm_n10107, gm_n50, gm_n49, in_12, gm_n9385, gm_n63);
	nor (gm_n10108, in_18, in_17, gm_n46, gm_n10107, gm_n62);
	nand (gm_n10109, gm_n10108, gm_n71, in_20);
	or (gm_n10110, gm_n2610, in_9);
	or (gm_n10111, gm_n48, gm_n53, gm_n52, gm_n10110, gm_n49);
	nor (gm_n10112, gm_n46, in_15, gm_n50, gm_n10111, gm_n81);
	nand (gm_n10113, gm_n45, gm_n62, in_18, gm_n10112, in_21);
	nor (gm_n10114, gm_n50, in_13, gm_n48, gm_n2739, gm_n63);
	nand (gm_n10115, in_18, in_17, in_16, gm_n10114, gm_n62);
	nor (gm_n10116, gm_n10115, gm_n71, in_20);
	and (gm_n10117, in_12, in_11, in_10, gm_n4876, gm_n49);
	nand (gm_n10118, gm_n46, in_15, in_14, gm_n10117, gm_n81);
	nor (gm_n10119, in_20, in_19, gm_n47, gm_n10118, in_21);
	and (gm_n10120, in_10, gm_n51, in_8, gm_n838);
	and (gm_n10121, gm_n49, in_12, in_11, gm_n10120, gm_n50);
	nand (gm_n10122, gm_n81, in_16, in_15, gm_n10121, gm_n47);
	nor (gm_n10123, in_21, in_20, gm_n62, gm_n10122);
	nor (gm_n10124, in_12, in_11, in_10, gm_n2931, in_13);
	nand (gm_n10125, in_16, in_15, gm_n50, gm_n10124, gm_n81);
	nor (gm_n10126, in_20, gm_n62, in_18, gm_n10125, in_21);
	nor (gm_n10127, in_16, in_15, gm_n50, gm_n1312, in_17);
	nand (gm_n10128, in_20, in_19, gm_n47, gm_n10127, gm_n71);
	nand (gm_n10129, gm_n50, gm_n49, gm_n48, gm_n8123, in_15);
	nor (gm_n10130, in_18, gm_n81, gm_n46, gm_n10129, in_19);
	nand (gm_n10131, gm_n10130, gm_n71, in_20);
	nor (gm_n10132, gm_n53, gm_n52, gm_n51, gm_n738, gm_n48);
	nand (gm_n10133, gm_n10132, gm_n49);
	nor (gm_n10134, in_16, gm_n63, gm_n50, gm_n10133, gm_n81);
	nand (gm_n10135, in_20, in_19, gm_n47, gm_n10134, gm_n71);
	nor (gm_n10136, gm_n53, in_10, gm_n51, gm_n5586, gm_n48);
	nand (gm_n10137, in_15, gm_n50, gm_n49, gm_n10136, gm_n46);
	nor (gm_n10138, in_19, in_18, gm_n81, gm_n10137, in_20);
	nand (gm_n10139, gm_n10138, gm_n71);
	and (gm_n10140, in_12, in_11, in_10, gm_n6430, in_13);
	nand (gm_n10141, in_16, in_15, in_14, gm_n10140, gm_n81);
	nor (gm_n10142, gm_n45, gm_n62, gm_n47, gm_n10141, in_21);
	nand (gm_n10143, in_16, gm_n63, in_14, gm_n9671, in_17);
	nor (gm_n10144, in_20, in_19, in_18, gm_n10143, in_21);
	nand (gm_n10145, in_17, in_16, gm_n63, gm_n6222, gm_n47);
	nor (gm_n10146, in_21, in_20, in_19, gm_n10145);
	nand (gm_n10147, gm_n81, in_16, in_15, gm_n9565, in_18);
	nor (gm_n10148, in_21, gm_n45, in_19, gm_n10147);
	or (gm_n10149, gm_n49, in_12, in_11, gm_n3332, in_14);
	nor (gm_n10150, in_17, in_16, in_15, gm_n10149, in_18);
	nand (gm_n10151, in_21, in_20, gm_n62, gm_n10150);
	nand (gm_n10152, in_12, in_11, in_10, gm_n2685, gm_n49);
	nor (gm_n10153, in_16, gm_n63, in_14, gm_n10152, gm_n81);
	nand (gm_n10154, in_20, in_19, gm_n47, gm_n10153, in_21);
	or (gm_n10155, in_12, in_11, gm_n52, gm_n2845, gm_n49);
	nor (gm_n10156, gm_n46, in_15, in_14, gm_n10155, gm_n81);
	nand (gm_n10157, gm_n45, gm_n62, in_18, gm_n10156, in_21);
	nand (gm_n10158, gm_n48, in_11, in_10, gm_n7172, gm_n49);
	nor (gm_n10159, in_16, in_15, gm_n50, gm_n10158, in_17);
	nand (gm_n10160, in_20, gm_n62, gm_n47, gm_n10159, gm_n71);
	and (gm_n10161, gm_n48, gm_n53, in_10, gm_n2334, gm_n49);
	nand (gm_n10162, in_16, gm_n63, gm_n50, gm_n10161, in_17);
	nor (gm_n10163, gm_n45, gm_n62, gm_n47, gm_n10162, in_21);
	nor (gm_n10164, in_12, in_11, in_10, gm_n5268, gm_n49);
	nand (gm_n10165, gm_n46, in_15, gm_n50, gm_n10164, gm_n81);
	nor (gm_n10166, in_20, gm_n62, in_18, gm_n10165, gm_n71);
	nor (gm_n10167, in_12, in_11, in_10, gm_n1152, gm_n49);
	nand (gm_n10168, in_16, in_15, gm_n50, gm_n10167, gm_n81);
	nor (gm_n10169, in_20, gm_n62, in_18, gm_n10168, in_21);
	nand (gm_n10170, in_16, in_15, gm_n50, gm_n8513, gm_n81);
	nor (gm_n10171, in_20, in_19, in_18, gm_n10170, gm_n71);
	nor (gm_n10172, in_16, gm_n63, gm_n50, gm_n7082, gm_n81);
	nand (gm_n10173, in_20, in_19, gm_n47, gm_n10172, gm_n71);
	nand (gm_n10174, gm_n50, in_13, in_12, gm_n7270, in_15);
	nor (gm_n10175, in_18, in_17, in_16, gm_n10174, gm_n62);
	nand (gm_n10176, gm_n10175, gm_n71, in_20);
	nand (gm_n10177, gm_n63, gm_n50, in_13, gm_n1556, gm_n46);
	nor (gm_n10178, gm_n62, in_18, gm_n81, gm_n10177, gm_n45);
	nand (gm_n10179, gm_n10178, in_21);
	nor (gm_n10180, gm_n8790, in_9);
	nand (gm_n10181, gm_n48, in_11, gm_n52, gm_n10180, gm_n49);
	nor (gm_n10182, gm_n46, in_15, in_14, gm_n10181, gm_n81);
	nand (gm_n10183, gm_n45, in_19, in_18, gm_n10182, in_21);
	or (gm_n10184, gm_n46, gm_n63, in_14, gm_n780, gm_n81);
	nor (gm_n10185, gm_n45, gm_n62, in_18, gm_n10184, gm_n71);
	nor (gm_n10186, in_14, in_13, gm_n48, gm_n6120, gm_n63);
	nand (gm_n10187, in_18, in_17, in_16, gm_n10186, in_19);
	nor (gm_n10188, gm_n10187, in_21, gm_n45);
	or (gm_n10189, in_8, gm_n55, gm_n82, gm_n141, in_9);
	nor (gm_n10190, in_12, gm_n53, gm_n52, gm_n10189, in_13);
	nand (gm_n10191, in_16, gm_n63, in_14, gm_n10190, gm_n81);
	nor (gm_n10192, in_20, gm_n62, gm_n47, gm_n10191, in_21);
	nand (gm_n10193, in_11, in_10, gm_n51, gm_n3489, gm_n48);
	nor (gm_n10194, gm_n63, in_14, in_13, gm_n10193, in_16);
	nand (gm_n10195, gm_n62, in_18, gm_n81, gm_n10194, in_20);
	nor (gm_n10196, gm_n10195, in_21);
	nand (gm_n10197, in_12, in_11, gm_n52, gm_n200, in_13);
	nor (gm_n10198, gm_n46, in_15, in_14, gm_n10197, gm_n81);
	nand (gm_n10199, gm_n45, in_19, gm_n47, gm_n10198, in_21);
	nor (gm_n10200, in_16, gm_n63, in_14, gm_n9334, in_17);
	nand (gm_n10201, in_20, in_19, in_18, gm_n10200, in_21);
	or (gm_n10202, gm_n48, gm_n53, in_10, gm_n9086, in_13);
	nor (gm_n10203, in_16, in_15, gm_n50, gm_n10202, in_17);
	nand (gm_n10204, gm_n45, gm_n62, in_18, gm_n10203, gm_n71);
	nand (gm_n10205, in_14, gm_n49, gm_n48, gm_n9341, in_15);
	nor (gm_n10206, gm_n47, in_17, in_16, gm_n10205, in_19);
	nand (gm_n10207, gm_n10206, gm_n71, in_20);
	and (gm_n10208, in_13, in_12, in_11, gm_n7939, in_14);
	nand (gm_n10209, in_17, in_16, in_15, gm_n10208, in_18);
	nor (gm_n10210, gm_n71, in_20, in_19, gm_n10209);
	nor (gm_n10211, in_8, in_7, gm_n82, gm_n530, gm_n51);
	and (gm_n10212, in_12, in_11, in_10, gm_n10211, in_13);
	nand (gm_n10213, in_16, in_15, in_14, gm_n10212, gm_n81);
	nor (gm_n10214, gm_n45, gm_n62, gm_n47, gm_n10213, gm_n71);
	nor (gm_n10215, in_15, gm_n50, in_13, gm_n2636, gm_n46);
	nand (gm_n10216, in_19, in_18, in_17, gm_n10215, gm_n45);
	nor (gm_n10217, gm_n10216, in_21);
	nand (gm_n10218, gm_n46, in_15, gm_n50, gm_n7647, in_17);
	nor (gm_n10219, gm_n45, in_19, gm_n47, gm_n10218, gm_n71);
	nand (gm_n10220, gm_n48, in_11, gm_n52, gm_n2522, in_13);
	nor (gm_n10221, gm_n46, gm_n63, gm_n50, gm_n10220, gm_n81);
	nand (gm_n10222, gm_n45, in_19, in_18, gm_n10221, in_21);
	nand (gm_n10223, gm_n48, gm_n53, gm_n52, gm_n3659, in_13);
	nor (gm_n10224, in_16, gm_n63, gm_n50, gm_n10223, gm_n81);
	nand (gm_n10225, in_20, in_19, in_18, gm_n10224, in_21);
	nor (gm_n10226, in_11, in_10, in_9, gm_n4489, in_12);
	nand (gm_n10227, in_15, in_14, in_13, gm_n10226, gm_n46);
	nor (gm_n10228, in_19, in_18, in_17, gm_n10227, in_20);
	nand (gm_n10229, gm_n10228, gm_n71);
	and (gm_n10230, in_11, in_10, gm_n51, gm_n2699, gm_n48);
	nand (gm_n10231, in_15, in_14, gm_n49, gm_n10230, in_16);
	nor (gm_n10232, in_19, gm_n47, in_17, gm_n10231, gm_n45);
	nand (gm_n10233, gm_n10232, in_21);
	and (gm_n10234, in_13, gm_n48, in_11, gm_n7611, in_14);
	nand (gm_n10235, gm_n81, gm_n46, in_15, gm_n10234, in_18);
	nor (gm_n10236, gm_n71, gm_n45, in_19, gm_n10235);
	and (gm_n10237, gm_n50, in_13, in_12, gm_n3194, gm_n63);
	nand (gm_n10238, in_18, in_17, gm_n46, gm_n10237, gm_n62);
	nor (gm_n10239, gm_n10238, in_21, gm_n45);
	and (gm_n10240, gm_n48, in_11, in_10, gm_n2749, in_13);
	nand (gm_n10241, in_16, in_15, in_14, gm_n10240, gm_n81);
	nor (gm_n10242, in_20, in_19, in_18, gm_n10241, in_21);
	nand (gm_n10243, gm_n46, gm_n63, in_14, gm_n3125, in_17);
	nor (gm_n10244, in_20, in_19, in_18, gm_n10243, gm_n71);
	nand (gm_n10245, in_12, in_11, gm_n52, gm_n3909, gm_n49);
	nor (gm_n10246, in_16, gm_n63, in_14, gm_n10245, in_17);
	nand (gm_n10247, in_20, in_19, in_18, gm_n10246, gm_n71);
	nand (gm_n10248, gm_n48, gm_n53, gm_n52, gm_n1675, gm_n49);
	nor (gm_n10249, in_16, in_15, in_14, gm_n10248, gm_n81);
	nand (gm_n10250, in_20, in_19, gm_n47, gm_n10249, gm_n71);
	nor (gm_n10251, in_17, in_16, gm_n63, gm_n9272, gm_n47);
	nand (gm_n10252, gm_n71, gm_n45, in_19, gm_n10251);
	nor (gm_n10253, gm_n51, gm_n64, gm_n55, gm_n843, in_10);
	nand (gm_n10254, in_13, in_12, in_11, gm_n10253, in_14);
	nor (gm_n10255, gm_n81, in_16, gm_n63, gm_n10254, gm_n47);
	nand (gm_n10256, in_21, gm_n45, gm_n62, gm_n10255);
	nand (gm_n10257, in_9, gm_n64, gm_n55, gm_n136, gm_n52);
	nor (gm_n10258, in_13, in_12, gm_n53, gm_n10257, gm_n50);
	nand (gm_n10259, gm_n81, in_16, gm_n63, gm_n10258, gm_n47);
	nor (gm_n10260, gm_n71, in_20, in_19, gm_n10259);
	nor (gm_n10261, gm_n49, gm_n48, in_11, gm_n9357, gm_n50);
	nand (gm_n10262, gm_n81, gm_n46, in_15, gm_n10261, gm_n47);
	nor (gm_n10263, gm_n71, in_20, in_19, gm_n10262);
	and (gm_n10264, in_12, in_11, in_10, gm_n9746, gm_n49);
	nand (gm_n10265, in_16, gm_n63, in_14, gm_n10264, in_17);
	nor (gm_n10266, gm_n45, gm_n62, gm_n47, gm_n10265, gm_n71);
	and (gm_n10267, in_13, gm_n48, gm_n53, gm_n5509, gm_n50);
	nand (gm_n10268, gm_n81, in_16, in_15, gm_n10267, in_18);
	nor (gm_n10269, in_21, gm_n45, in_19, gm_n10268);
	nand (gm_n10270, gm_n50, in_13, in_12, gm_n7060);
	nor (gm_n10271, in_17, gm_n46, in_15, gm_n10270, gm_n47);
	nand (gm_n10272, gm_n71, gm_n45, in_19, gm_n10271);
	nand (gm_n10273, gm_n63, in_14, gm_n49, gm_n4428, in_16);
	nor (gm_n10274, in_19, gm_n47, in_17, gm_n10273, in_20);
	nand (gm_n10275, gm_n10274, in_21);
	nand (gm_n10276, gm_n49, in_12, gm_n53, gm_n5116, in_14);
	nor (gm_n10277, gm_n81, in_16, gm_n63, gm_n10276, gm_n47);
	nand (gm_n10278, in_21, gm_n45, gm_n62, gm_n10277);
	nand (gm_n10279, in_13, in_12, gm_n53, gm_n5928, gm_n50);
	nor (gm_n10280, gm_n81, gm_n46, in_15, gm_n10279, in_18);
	nand (gm_n10281, in_21, gm_n45, in_19, gm_n10280);
	and (gm_n10282, gm_n48, in_11, in_10, gm_n9902, in_13);
	nand (gm_n10283, gm_n46, in_15, gm_n50, gm_n10282, in_17);
	nor (gm_n10284, gm_n45, in_19, gm_n47, gm_n10283, in_21);
	and (gm_n10285, in_14, gm_n49, in_12, gm_n8409, gm_n63);
	nand (gm_n10286, gm_n47, in_17, in_16, gm_n10285, in_19);
	nor (gm_n10287, gm_n10286, in_21, gm_n45);
	nor (gm_n10288, gm_n45, gm_n62, in_18, gm_n9136, gm_n71);
	nor (gm_n10289, in_12, gm_n53, gm_n52, gm_n4715, in_13);
	nand (gm_n10290, gm_n46, in_15, in_14, gm_n10289, gm_n81);
	nor (gm_n10291, in_20, in_19, in_18, gm_n10290, gm_n71);
	nand (gm_n10292, in_13, gm_n48, gm_n53, gm_n4310, gm_n50);
	nor (gm_n10293, gm_n81, gm_n46, in_15, gm_n10292, gm_n47);
	nand (gm_n10294, gm_n71, gm_n45, gm_n62, gm_n10293);
	nand (gm_n10295, gm_n49, gm_n48, gm_n53, gm_n6313, gm_n50);
	nor (gm_n10296, gm_n81, gm_n46, in_15, gm_n10295, in_18);
	nand (gm_n10297, in_21, in_20, gm_n62, gm_n10296);
	nand (gm_n10298, in_12, in_11, gm_n52, gm_n380, gm_n49);
	nor (gm_n10299, gm_n46, in_15, gm_n50, gm_n10298, gm_n81);
	nand (gm_n10300, gm_n45, gm_n62, gm_n47, gm_n10299, gm_n71);
	nand (gm_n10301, in_14, in_13, gm_n48, gm_n1789, in_15);
	nor (gm_n10302, in_18, gm_n81, gm_n46, gm_n10301, gm_n62);
	nand (gm_n10303, gm_n10302, in_21, in_20);
	nor (gm_n10304, in_15, in_14, gm_n49, gm_n5612, in_16);
	nand (gm_n10305, in_19, in_18, in_17, gm_n10304, in_20);
	nor (gm_n10306, gm_n10305, in_21);
	nand (gm_n10307, in_11, gm_n52, in_9, gm_n6643, gm_n48);
	nor (gm_n10308, in_15, gm_n50, in_13, gm_n10307, gm_n46);
	nand (gm_n10309, in_19, gm_n47, in_17, gm_n10308, gm_n45);
	nor (gm_n10310, gm_n10309, gm_n71);
	nor (gm_n10311, in_14, in_13, gm_n48, gm_n4402, in_15);
	nand (gm_n10312, in_18, in_17, gm_n46, gm_n10311, in_19);
	nor (gm_n10313, gm_n10312, in_21, gm_n45);
	nor (gm_n10314, gm_n63, gm_n50, in_13, gm_n275, in_16);
	nand (gm_n10315, in_19, in_18, in_17, gm_n10314, gm_n45);
	nor (gm_n10316, gm_n10315, gm_n71);
	nor (gm_n10317, gm_n53, in_10, in_9, gm_n1239, gm_n48);
	nand (gm_n10318, gm_n63, in_14, in_13, gm_n10317, gm_n46);
	nor (gm_n10319, gm_n62, gm_n47, gm_n81, gm_n10318, gm_n45);
	nand (gm_n10320, gm_n10319, gm_n71);
	or (gm_n10321, in_13, gm_n48, gm_n53, gm_n2518, in_14);
	nor (gm_n10322, gm_n81, in_16, in_15, gm_n10321, in_18);
	nand (gm_n10323, in_21, in_20, gm_n62, gm_n10322);
	nand (gm_n10324, gm_n48, gm_n53, gm_n52, gm_n6539, gm_n49);
	nor (gm_n10325, gm_n46, gm_n63, gm_n50, gm_n10324, gm_n81);
	nand (gm_n10326, gm_n45, gm_n62, in_18, gm_n10325, in_21);
	nor (gm_n10327, in_11, gm_n52, gm_n51, gm_n2823, gm_n48);
	nand (gm_n10328, gm_n63, in_14, gm_n49, gm_n10327, gm_n46);
	nor (gm_n10329, in_19, in_18, in_17, gm_n10328, in_20);
	nand (gm_n10330, gm_n10329, in_21);
	and (gm_n10331, gm_n5185, in_9);
	and (gm_n10332, in_12, in_11, in_10, gm_n10331, in_13);
	nand (gm_n10333, gm_n46, in_15, gm_n50, gm_n10332, gm_n81);
	nor (gm_n10334, in_20, gm_n62, gm_n47, gm_n10333, gm_n71);
	and (gm_n10335, gm_n50, in_13, gm_n48, gm_n8537, in_15);
	nand (gm_n10336, in_18, gm_n81, in_16, gm_n10335, in_19);
	nor (gm_n10337, gm_n10336, in_21, in_20);
	nor (gm_n10338, in_14, gm_n49, gm_n48, gm_n3175, in_15);
	nand (gm_n10339, gm_n47, in_17, in_16, gm_n10338, in_19);
	nor (gm_n10340, gm_n10339, in_21, in_20);
	and (gm_n10341, gm_n49, gm_n48, gm_n53, gm_n2186, in_14);
	nand (gm_n10342, gm_n81, in_16, in_15, gm_n10341, gm_n47);
	nor (gm_n10343, in_21, gm_n45, in_19, gm_n10342);
	nor (gm_n10344, gm_n3743, in_10, gm_n51);
	nand (gm_n10345, in_13, in_12, gm_n53, gm_n10344, in_14);
	nor (gm_n10346, in_17, in_16, in_15, gm_n10345, gm_n47);
	nand (gm_n10347, in_21, in_20, gm_n62, gm_n10346);
	nand (gm_n10348, in_13, in_12, in_11, gm_n5003, in_14);
	nor (gm_n10349, in_17, gm_n46, gm_n63, gm_n10348, in_18);
	nand (gm_n10350, gm_n71, in_20, gm_n62, gm_n10349);
	nor (gm_n10351, in_11, gm_n52, gm_n51, gm_n520);
	nand (gm_n10352, in_14, gm_n49, gm_n48, gm_n10351, in_15);
	nor (gm_n10353, gm_n47, in_17, in_16, gm_n10352, in_19);
	nand (gm_n10354, gm_n10353, gm_n71, gm_n45);
	and (gm_n10355, in_11, gm_n52, gm_n51, gm_n1192);
	nand (gm_n10356, gm_n10355, in_13, gm_n48);
	nor (gm_n10357, in_16, in_15, in_14, gm_n10356, gm_n81);
	nand (gm_n10358, in_20, in_19, in_18, gm_n10357, gm_n71);
	and (gm_n10359, gm_n49, in_12, in_11, gm_n6576, in_14);
	nand (gm_n10360, in_17, gm_n46, gm_n63, gm_n10359, gm_n47);
	nor (gm_n10361, in_21, gm_n45, gm_n62, gm_n10360);
	and (gm_n10362, gm_n49, in_12, in_11, gm_n1609, in_14);
	nand (gm_n10363, in_17, in_16, gm_n63, gm_n10362, gm_n47);
	nor (gm_n10364, in_21, in_20, gm_n62, gm_n10363);
	nor (gm_n10365, gm_n48, in_11, in_10, gm_n3249, gm_n49);
	nand (gm_n10366, in_16, gm_n63, in_14, gm_n10365, gm_n81);
	nor (gm_n10367, gm_n45, in_19, in_18, gm_n10366, gm_n71);
	and (gm_n10368, gm_n48, in_11, in_10, gm_n1755, in_13);
	nand (gm_n10369, gm_n46, in_15, gm_n50, gm_n10368, gm_n81);
	nor (gm_n10370, gm_n45, in_19, gm_n47, gm_n10369, gm_n71);
	and (gm_n10371, gm_n53, in_10, gm_n51, gm_n4293, in_12);
	nand (gm_n10372, in_15, in_14, in_13, gm_n10371, gm_n46);
	nor (gm_n10373, gm_n62, gm_n47, in_17, gm_n10372, gm_n45);
	nand (gm_n10374, gm_n10373, in_21);
	nand (gm_n10375, in_13, in_12, in_11, gm_n903, gm_n50);
	nor (gm_n10376, in_17, gm_n46, gm_n63, gm_n10375, in_18);
	nand (gm_n10377, gm_n71, gm_n45, in_19, gm_n10376);
	nand (gm_n10378, gm_n48, in_11, in_10, gm_n934, in_13);
	nor (gm_n10379, gm_n46, gm_n63, gm_n50, gm_n10378, in_17);
	nand (gm_n10380, in_20, gm_n62, in_18, gm_n10379, in_21);
	nor (gm_n10381, in_17, in_16, gm_n63, gm_n10270, in_18);
	nand (gm_n10382, gm_n71, in_20, in_19, gm_n10381);
	and (gm_n10383, gm_n63, gm_n50, gm_n49, gm_n9168, in_16);
	nand (gm_n10384, in_19, in_18, gm_n81, gm_n10383, gm_n45);
	nor (gm_n10385, gm_n10384, gm_n71);
	and (gm_n10386, in_10, gm_n51, in_8, gm_n691);
	and (gm_n10387, in_13, gm_n48, in_11, gm_n10386, gm_n50);
	nand (gm_n10388, in_17, in_16, gm_n63, gm_n10387, in_18);
	nor (gm_n10389, in_21, gm_n45, in_19, gm_n10388);
	nand (gm_n10390, in_16, in_15, gm_n50, gm_n1067, in_17);
	nor (gm_n10391, gm_n45, in_19, in_18, gm_n10390, gm_n71);
	or (gm_n10392, gm_n53, gm_n52, in_9, gm_n1763, in_12);
	nor (gm_n10393, in_15, gm_n50, gm_n49, gm_n10392, in_16);
	nand (gm_n10394, gm_n62, in_18, in_17, gm_n10393, in_20);
	nor (gm_n10395, gm_n10394, in_21);
	and (gm_n10396, in_11, gm_n52, gm_n51, gm_n4723, gm_n48);
	nand (gm_n10397, in_15, gm_n50, gm_n49, gm_n10396, in_16);
	nor (gm_n10398, in_19, in_18, gm_n81, gm_n10397, in_20);
	nand (gm_n10399, gm_n10398, gm_n71);
	nand (gm_n10400, in_13, in_12, in_11, gm_n2078, in_14);
	nor (gm_n10401, gm_n81, in_16, in_15, gm_n10400, gm_n47);
	nand (gm_n10402, gm_n71, in_20, gm_n62, gm_n10401);
	nand (gm_n10403, in_12, gm_n53, gm_n52, gm_n5893, in_13);
	nor (gm_n10404, gm_n46, gm_n63, gm_n50, gm_n10403, in_17);
	nand (gm_n10405, gm_n45, in_19, in_18, gm_n10404, gm_n71);
	nand (gm_n10406, gm_n48, gm_n53, gm_n52, gm_n200, gm_n49);
	nor (gm_n10407, in_16, gm_n63, gm_n50, gm_n10406, gm_n81);
	nand (gm_n10408, gm_n45, gm_n62, in_18, gm_n10407, gm_n71);
	nor (gm_n10409, in_12, gm_n53, gm_n52, gm_n893, in_13);
	nand (gm_n10410, in_16, in_15, in_14, gm_n10409, in_17);
	nor (gm_n10411, gm_n45, in_19, gm_n47, gm_n10410, gm_n71);
	nand (gm_n10412, gm_n46, in_15, in_14, gm_n7496, gm_n81);
	nor (gm_n10413, in_20, gm_n62, in_18, gm_n10412, in_21);
	nor (gm_n10414, gm_n50, in_13, in_12, gm_n317, in_15);
	nand (gm_n10415, in_18, in_17, in_16, gm_n10414, gm_n62);
	nor (gm_n10416, gm_n10415, in_21, gm_n45);
	nand (gm_n10417, in_17, gm_n46, gm_n63, gm_n623, gm_n47);
	nor (gm_n10418, gm_n71, in_20, gm_n62, gm_n10417);
	nand (gm_n10419, in_12, in_11, in_10, gm_n2877, gm_n49);
	nor (gm_n10420, gm_n46, gm_n63, gm_n50, gm_n10419, gm_n81);
	nand (gm_n10421, in_20, gm_n62, gm_n47, gm_n10420, in_21);
	nor (gm_n10422, in_19, in_18, gm_n81, gm_n6481, gm_n45);
	nand (gm_n10423, gm_n10422, gm_n71);
	nand (gm_n10424, gm_n50, gm_n49, gm_n48, gm_n4370, in_15);
	nor (gm_n10425, in_18, gm_n81, gm_n46, gm_n10424, in_19);
	nand (gm_n10426, gm_n10425, in_21, gm_n45);
	and (gm_n10427, gm_n53, in_10, in_9, gm_n1222, gm_n48);
	nand (gm_n10428, gm_n63, in_14, in_13, gm_n10427, in_16);
	nor (gm_n10429, in_19, gm_n47, gm_n81, gm_n10428, in_20);
	nand (gm_n10430, gm_n10429, gm_n71);
	nand (gm_n10431, in_9, gm_n64, in_7, gm_n504, in_10);
	nor (gm_n10432, in_13, gm_n48, gm_n53, gm_n10431, gm_n50);
	nand (gm_n10433, gm_n81, gm_n46, in_15, gm_n10432, in_18);
	nor (gm_n10434, in_21, gm_n45, in_19, gm_n10433);
	nor (gm_n10435, gm_n63, in_14, gm_n49, gm_n334, in_16);
	nand (gm_n10436, gm_n62, in_18, in_17, gm_n10435, in_20);
	nor (gm_n10437, gm_n10436, gm_n71);
	or (gm_n10438, in_11, in_10, gm_n51, gm_n3557, gm_n48);
	nor (gm_n10439, in_15, gm_n50, in_13, gm_n10438, in_16);
	nand (gm_n10440, gm_n10439, gm_n47, gm_n81);
	nor (gm_n10441, in_21, gm_n45, in_19, gm_n10440);
	nor (gm_n10442, gm_n50, gm_n49, in_12, gm_n4790, gm_n63);
	nand (gm_n10443, in_18, in_17, gm_n46, gm_n10442, in_19);
	nor (gm_n10444, gm_n10443, gm_n71, gm_n45);
	or (gm_n10445, gm_n50, gm_n49, gm_n48, gm_n6120, in_15);
	nor (gm_n10446, gm_n47, in_17, in_16, gm_n10445, in_19);
	nand (gm_n10447, gm_n10446, gm_n71, gm_n45);
	or (gm_n10448, in_12, in_11, in_10, gm_n7400, gm_n49);
	nor (gm_n10449, in_16, gm_n63, gm_n50, gm_n10448, in_17);
	nand (gm_n10450, gm_n45, in_19, in_18, gm_n10449, gm_n71);
	nand (gm_n10451, gm_n50, gm_n49, gm_n48, gm_n2039, gm_n63);
	nor (gm_n10452, gm_n47, in_17, gm_n46, gm_n10451, in_19);
	nand (gm_n10453, gm_n10452, in_21, gm_n45);
	nand (gm_n10454, gm_n10453, gm_n10450, gm_n10447);
	nor (gm_n10455, gm_n10441, gm_n10437, gm_n10434, gm_n10454, gm_n10444);
	nand (gm_n10456, gm_n10426, gm_n10423, gm_n10421, gm_n10455, gm_n10430);
	nor (gm_n10457, gm_n10416, gm_n10413, gm_n10411, gm_n10456, gm_n10418);
	nand (gm_n10458, gm_n10405, gm_n10402, gm_n10399, gm_n10457, gm_n10408);
	nor (gm_n10459, gm_n10391, gm_n10389, gm_n10385, gm_n10458, gm_n10395);
	nand (gm_n10460, gm_n10380, gm_n10377, gm_n10374, gm_n10459, gm_n10382);
	nor (gm_n10461, gm_n10367, gm_n10364, gm_n10361, gm_n10460, gm_n10370);
	nand (gm_n10462, gm_n10354, gm_n10350, gm_n10347, gm_n10461, gm_n10358);
	nor (gm_n10463, gm_n10340, gm_n10337, gm_n10334, gm_n10462, gm_n10343);
	nand (gm_n10464, gm_n10326, gm_n10323, gm_n10320, gm_n10463, gm_n10330);
	nor (gm_n10465, gm_n10313, gm_n10310, gm_n10306, gm_n10464, gm_n10316);
	nand (gm_n10466, gm_n10300, gm_n10297, gm_n10294, gm_n10465, gm_n10303);
	nor (gm_n10467, gm_n10288, gm_n10287, gm_n10284, gm_n10466, gm_n10291);
	nand (gm_n10468, gm_n10278, gm_n10275, gm_n10272, gm_n10467, gm_n10281);
	nor (gm_n10469, gm_n10266, gm_n10263, gm_n10260, gm_n10468, gm_n10269);
	nand (gm_n10470, gm_n10252, gm_n10250, gm_n10247, gm_n10469, gm_n10256);
	nor (gm_n10471, gm_n10242, gm_n10239, gm_n10236, gm_n10470, gm_n10244);
	nand (gm_n10472, gm_n10229, gm_n10225, gm_n10222, gm_n10471, gm_n10233);
	nor (gm_n10473, gm_n10217, gm_n10214, gm_n10210, gm_n10472, gm_n10219);
	nand (gm_n10474, gm_n10204, gm_n10201, gm_n10199, gm_n10473, gm_n10207);
	nor (gm_n10475, gm_n10192, gm_n10188, gm_n10185, gm_n10474, gm_n10196);
	nand (gm_n10476, gm_n10179, gm_n10176, gm_n10173, gm_n10475, gm_n10183);
	nor (gm_n10477, gm_n10169, gm_n10166, gm_n10163, gm_n10476, gm_n10171);
	nand (gm_n10478, gm_n10157, gm_n10154, gm_n10151, gm_n10477, gm_n10160);
	nor (gm_n10479, gm_n10146, gm_n10144, gm_n10142, gm_n10478, gm_n10148);
	nand (gm_n10480, gm_n10135, gm_n10131, gm_n10128, gm_n10479, gm_n10139);
	nor (gm_n10481, gm_n10123, gm_n10119, gm_n10116, gm_n10480, gm_n10126);
	nand (gm_n10482, gm_n10109, gm_n10106, gm_n10104, gm_n10481, gm_n10113);
	nor (gm_n10483, gm_n10098, gm_n10095, gm_n10091, gm_n10482, gm_n10101);
	nand (gm_n10484, gm_n10084, gm_n10080, gm_n10077, gm_n10483, gm_n10088);
	nor (gm_n10485, gm_n10071, gm_n10068, gm_n10065, gm_n10484, gm_n10074);
	nand (gm_n10486, gm_n10058, gm_n10055, gm_n10052, gm_n10485, gm_n10061);
	nor (gm_n10487, gm_n10046, gm_n10045, gm_n10041, gm_n10486, gm_n10049);
	nand (gm_n10488, gm_n10035, gm_n10032, gm_n10028, gm_n10487, gm_n10038);
	nor (gm_n10489, gm_n10022, gm_n10019, gm_n10017, gm_n10488, gm_n10024);
	nand (gm_n10490, gm_n10012, gm_n10009, gm_n10006, gm_n10489, gm_n10015);
	nor (out_17, gm_n10003, gm_n10000, gm_n9997, gm_n10490);
	and (gm_n10492, in_14, in_13, gm_n48, gm_n7514, in_15);
	nand (gm_n10493, in_18, gm_n81, in_16, gm_n10492, gm_n62);
	nor (gm_n10494, gm_n10493, gm_n71, gm_n45);
	nand (gm_n10495, in_15, gm_n50, in_13, gm_n8232, gm_n46);
	nor (gm_n10496, in_19, in_18, gm_n81, gm_n10495, gm_n45);
	nand (gm_n10497, gm_n10496, in_21);
	nand (gm_n10498, gm_n49, in_12, in_11, gm_n5858, gm_n50);
	nor (gm_n10499, gm_n81, gm_n46, in_15, gm_n10498, gm_n47);
	nand (gm_n10500, in_21, gm_n45, gm_n62, gm_n10499);
	nand (gm_n10501, gm_n49, in_12, gm_n53, gm_n9589, gm_n50);
	nor (gm_n10502, gm_n81, gm_n46, gm_n63, gm_n10501, gm_n47);
	nand (gm_n10503, in_21, in_20, gm_n62, gm_n10502);
	or (gm_n10504, gm_n49, gm_n48, gm_n53, gm_n4432, in_14);
	nor (gm_n10505, in_17, in_16, gm_n63, gm_n10504, gm_n47);
	nand (gm_n10506, gm_n71, in_20, gm_n62, gm_n10505);
	and (gm_n10507, in_13, in_12, gm_n53, gm_n2276, gm_n50);
	nand (gm_n10508, in_17, gm_n46, gm_n63, gm_n10507, gm_n47);
	nor (gm_n10509, gm_n71, gm_n45, in_19, gm_n10508);
	nand (gm_n10510, gm_n53, in_10, in_9, gm_n1421, gm_n48);
	nor (gm_n10511, gm_n63, gm_n50, in_13, gm_n10510, gm_n46);
	nand (gm_n10512, in_19, in_18, gm_n81, gm_n10511, in_20);
	nor (gm_n10513, gm_n10512, in_21);
	nand (gm_n10514, in_11, gm_n52, in_9, gm_n1936, gm_n48);
	nor (gm_n10515, in_15, in_14, in_13, gm_n10514, gm_n46);
	nand (gm_n10516, in_19, in_18, in_17, gm_n10515, in_20);
	nor (gm_n10517, gm_n10516, gm_n71);
	nor (gm_n10518, in_12, in_11, in_10, gm_n9867, in_13);
	nand (gm_n10519, in_16, gm_n63, in_14, gm_n10518, in_17);
	nor (gm_n10520, gm_n45, in_19, in_18, gm_n10519, gm_n71);
	nor (gm_n10521, gm_n53, in_10, gm_n51, gm_n218, gm_n48);
	nand (gm_n10522, gm_n63, gm_n50, gm_n49, gm_n10521, gm_n46);
	nor (gm_n10523, gm_n62, gm_n47, in_17, gm_n10522, gm_n45);
	nand (gm_n10524, gm_n10523, gm_n71);
	and (gm_n10525, in_11, in_10, gm_n51, gm_n4388);
	nand (gm_n10526, gm_n50, in_13, gm_n48, gm_n10525, in_15);
	nor (gm_n10527, gm_n47, in_17, in_16, gm_n10526, gm_n62);
	nand (gm_n10528, gm_n10527, in_21, in_20);
	nor (gm_n10529, in_16, gm_n63, gm_n50, gm_n4210, in_17);
	nand (gm_n10530, gm_n45, in_19, gm_n47, gm_n10529, gm_n71);
	nand (gm_n10531, gm_n48, in_11, gm_n52, gm_n912, in_13);
	nor (gm_n10532, gm_n46, in_15, in_14, gm_n10531, gm_n81);
	nand (gm_n10533, gm_n45, in_19, gm_n47, gm_n10532, gm_n71);
	nand (gm_n10534, gm_n46, gm_n63, gm_n50, gm_n6985, gm_n81);
	nor (gm_n10535, in_20, in_19, gm_n47, gm_n10534, in_21);
	nor (gm_n10536, in_12, in_11, in_10, gm_n6309, gm_n49);
	nand (gm_n10537, in_16, in_15, in_14, gm_n10536, in_17);
	nor (gm_n10538, in_20, gm_n62, gm_n47, gm_n10537, gm_n71);
	nand (gm_n10539, gm_n81, gm_n46, in_15, gm_n2505, gm_n47);
	nor (gm_n10540, gm_n71, in_20, gm_n62, gm_n10539);
	nor (gm_n10541, in_13, gm_n48, in_11, gm_n5423, in_14);
	nand (gm_n10542, gm_n81, gm_n46, gm_n63, gm_n10541, in_18);
	nor (gm_n10543, gm_n71, in_20, in_19, gm_n10542);
	nand (gm_n10544, gm_n48, gm_n53, in_10, gm_n6217, in_13);
	nor (gm_n10545, gm_n46, in_15, in_14, gm_n10544, in_17);
	nand (gm_n10546, in_20, gm_n62, in_18, gm_n10545, in_21);
	nor (gm_n10547, in_11, in_10, gm_n51, gm_n1709, gm_n48);
	nand (gm_n10548, gm_n63, gm_n50, gm_n49, gm_n10547, in_16);
	nor (gm_n10549, gm_n62, gm_n47, gm_n81, gm_n10548, in_20);
	nand (gm_n10550, gm_n10549, in_21);
	nand (gm_n10551, in_14, gm_n49, in_12, gm_n2433, in_15);
	nor (gm_n10552, in_18, in_17, gm_n46, gm_n10551, gm_n62);
	nand (gm_n10553, gm_n10552, in_21, gm_n45);
	nand (gm_n10554, gm_n49, gm_n48, in_11, gm_n2218, gm_n50);
	nor (gm_n10555, gm_n81, gm_n46, in_15, gm_n10554, gm_n47);
	nand (gm_n10556, in_21, in_20, in_19, gm_n10555);
	nand (gm_n10557, gm_n53, gm_n52, gm_n51, gm_n3043, in_12);
	nor (gm_n10558, in_15, in_14, in_13, gm_n10557, in_16);
	nand (gm_n10559, in_19, gm_n47, gm_n81, gm_n10558, in_20);
	nor (gm_n10560, gm_n10559, gm_n71);
	and (gm_n10561, gm_n48, gm_n53, in_10, gm_n9518, gm_n49);
	nand (gm_n10562, in_16, gm_n63, gm_n50, gm_n10561, in_17);
	nor (gm_n10563, gm_n45, gm_n62, gm_n47, gm_n10562, gm_n71);
	and (gm_n10564, in_12, in_11, in_10, gm_n4266, gm_n49);
	nand (gm_n10565, gm_n46, gm_n63, gm_n50, gm_n10564, in_17);
	nor (gm_n10566, in_20, in_19, gm_n47, gm_n10565, gm_n71);
	nor (gm_n10567, gm_n48, in_11, in_10, gm_n1076, gm_n49);
	nand (gm_n10568, in_16, in_15, gm_n50, gm_n10567, in_17);
	nor (gm_n10569, gm_n45, in_19, in_18, gm_n10568, in_21);
	nand (gm_n10570, gm_n49, gm_n48, in_11, gm_n2305, in_14);
	nor (gm_n10571, in_17, in_16, in_15, gm_n10570, gm_n47);
	nand (gm_n10572, gm_n71, gm_n45, in_19, gm_n10571);
	nand (gm_n10573, gm_n49, in_12, gm_n53, gm_n8676, in_14);
	nor (gm_n10574, gm_n81, gm_n46, gm_n63, gm_n10573, in_18);
	nand (gm_n10575, in_21, gm_n45, gm_n62, gm_n10574);
	nand (gm_n10576, in_15, gm_n50, gm_n49, gm_n10092, in_16);
	nor (gm_n10577, gm_n62, gm_n47, gm_n81, gm_n10576, in_20);
	nand (gm_n10578, gm_n10577, gm_n71);
	nor (gm_n10579, in_11, in_10, in_9, gm_n2345);
	nand (gm_n10580, in_14, in_13, gm_n48, gm_n10579, gm_n63);
	nor (gm_n10581, gm_n47, in_17, in_16, gm_n10580, gm_n62);
	nand (gm_n10582, gm_n10581, in_21, in_20);
	nand (gm_n10583, gm_n47, in_17, gm_n46, gm_n8977, in_19);
	nor (gm_n10584, gm_n10583, gm_n71, in_20);
	nor (gm_n10585, in_13, in_12, gm_n53, gm_n6135, in_14);
	nand (gm_n10586, gm_n81, gm_n46, gm_n63, gm_n10585, gm_n47);
	nor (gm_n10587, gm_n71, in_20, in_19, gm_n10586);
	and (gm_n10588, in_13, gm_n48, in_11, gm_n5289, gm_n50);
	nand (gm_n10589, gm_n81, in_16, in_15, gm_n10588, gm_n47);
	nor (gm_n10590, in_21, gm_n45, in_19, gm_n10589);
	nand (gm_n10591, gm_n53, in_10, gm_n51, gm_n6549, in_12);
	nor (gm_n10592, gm_n63, gm_n50, in_13, gm_n10591, gm_n46);
	nand (gm_n10593, in_19, gm_n47, gm_n81, gm_n10592, gm_n45);
	nor (gm_n10594, gm_n10593, gm_n71);
	nor (gm_n10595, in_9, gm_n64, gm_n55, gm_n525, gm_n52);
	nand (gm_n10596, gm_n49, gm_n48, gm_n53, gm_n10595, gm_n50);
	nor (gm_n10597, gm_n81, in_16, gm_n63, gm_n10596, in_18);
	nand (gm_n10598, gm_n71, gm_n45, gm_n62, gm_n10597);
	or (gm_n10599, in_12, gm_n53, gm_n52, gm_n5268, gm_n49);
	nor (gm_n10600, in_16, in_15, gm_n50, gm_n10599, gm_n81);
	nand (gm_n10601, gm_n45, in_19, in_18, gm_n10600, in_21);
	and (gm_n10602, gm_n53, gm_n52, gm_n51, gm_n1156, in_12);
	nand (gm_n10603, in_15, gm_n50, gm_n49, gm_n10602, in_16);
	nor (gm_n10604, gm_n62, gm_n47, in_17, gm_n10603, in_20);
	nand (gm_n10605, gm_n10604, in_21);
	nor (gm_n10606, in_16, gm_n63, gm_n50, gm_n6887, in_17);
	nand (gm_n10607, gm_n45, in_19, gm_n47, gm_n10606, in_21);
	and (gm_n10608, in_12, gm_n53, gm_n52, gm_n5676, gm_n49);
	nand (gm_n10609, in_16, gm_n63, gm_n50, gm_n10608, in_17);
	nor (gm_n10610, gm_n45, gm_n62, gm_n47, gm_n10609, in_21);
	nor (gm_n10611, in_12, in_11, in_10, gm_n3515, gm_n49);
	nand (gm_n10612, in_16, gm_n63, in_14, gm_n10611, gm_n81);
	nor (gm_n10613, gm_n45, in_19, in_18, gm_n10612, gm_n71);
	nand (gm_n10614, gm_n46, gm_n63, in_14, gm_n10089, gm_n81);
	nor (gm_n10615, gm_n45, in_19, in_18, gm_n10614, in_21);
	nor (gm_n10616, in_12, gm_n53, gm_n52, gm_n639, gm_n49);
	nand (gm_n10617, in_16, gm_n63, in_14, gm_n10616, in_17);
	nor (gm_n10618, in_20, gm_n62, in_18, gm_n10617, in_21);
	and (gm_n10619, gm_n53, gm_n52, gm_n51, gm_n3064, gm_n48);
	nand (gm_n10620, gm_n63, in_14, gm_n49, gm_n10619, gm_n46);
	nor (gm_n10621, in_19, in_18, in_17, gm_n10620, gm_n45);
	nand (gm_n10622, gm_n10621, in_21);
	nand (gm_n10623, gm_n48, in_11, in_10, gm_n2641, in_13);
	nor (gm_n10624, gm_n46, gm_n63, in_14, gm_n10623, in_17);
	nand (gm_n10625, gm_n45, in_19, gm_n47, gm_n10624, in_21);
	nand (gm_n10626, in_12, in_11, gm_n52, gm_n311, in_13);
	nor (gm_n10627, in_16, in_15, in_14, gm_n10626, in_17);
	nand (gm_n10628, gm_n45, in_19, in_18, gm_n10627, gm_n71);
	nand (gm_n10629, in_13, in_12, gm_n53, gm_n2127, in_14);
	nor (gm_n10630, gm_n81, in_16, in_15, gm_n10629, in_18);
	nand (gm_n10631, in_21, gm_n45, gm_n62, gm_n10630);
	nor (gm_n10632, in_12, in_11, gm_n52, gm_n2043, gm_n49);
	nand (gm_n10633, gm_n46, gm_n63, in_14, gm_n10632, in_17);
	nor (gm_n10634, in_20, in_19, gm_n47, gm_n10633, in_21);
	nor (gm_n10635, in_12, gm_n53, in_10, gm_n2845, in_13);
	nand (gm_n10636, in_16, in_15, in_14, gm_n10635, in_17);
	nor (gm_n10637, gm_n45, gm_n62, gm_n47, gm_n10636, gm_n71);
	and (gm_n10638, gm_n49, gm_n48, gm_n53, gm_n3460, gm_n50);
	nand (gm_n10639, gm_n81, in_16, gm_n63, gm_n10638, in_18);
	nor (gm_n10640, in_21, gm_n45, in_19, gm_n10639);
	nor (gm_n10641, gm_n63, gm_n50, gm_n49, gm_n8002, in_16);
	nand (gm_n10642, in_19, gm_n47, gm_n81, gm_n10641, gm_n45);
	nor (gm_n10643, gm_n10642, gm_n71);
	nand (gm_n10644, gm_n50, gm_n49, in_12, gm_n5225, in_15);
	nor (gm_n10645, in_18, in_17, in_16, gm_n10644, gm_n62);
	nand (gm_n10646, gm_n10645, gm_n71, gm_n45);
	nand (gm_n10647, in_13, gm_n48, in_11, gm_n9769, gm_n50);
	nor (gm_n10648, gm_n81, in_16, gm_n63, gm_n10647, in_18);
	nand (gm_n10649, in_21, in_20, in_19, gm_n10648);
	nand (gm_n10650, in_13, in_12, gm_n53, gm_n8870, gm_n50);
	nor (gm_n10651, in_17, gm_n46, in_15, gm_n10650, in_18);
	nand (gm_n10652, in_21, gm_n45, gm_n62, gm_n10651);
	or (gm_n10653, gm_n49, gm_n48, in_11, gm_n5041, gm_n50);
	nor (gm_n10654, gm_n81, gm_n46, in_15, gm_n10653, in_18);
	nand (gm_n10655, in_21, gm_n45, gm_n62, gm_n10654);
	and (gm_n10656, in_12, gm_n53, in_10, gm_n8038, gm_n49);
	nand (gm_n10657, in_16, in_15, gm_n50, gm_n10656, in_17);
	nor (gm_n10658, gm_n45, in_19, in_18, gm_n10657, gm_n71);
	and (gm_n10659, in_12, gm_n53, gm_n52, gm_n449, in_13);
	nand (gm_n10660, in_16, gm_n63, in_14, gm_n10659, gm_n81);
	nor (gm_n10661, gm_n45, in_19, in_18, gm_n10660, gm_n71);
	nor (gm_n10662, gm_n48, gm_n53, gm_n52, gm_n7400, gm_n49);
	nand (gm_n10663, gm_n46, gm_n63, in_14, gm_n10662, in_17);
	nor (gm_n10664, in_20, in_19, in_18, gm_n10663, gm_n71);
	nand (gm_n10665, gm_n46, in_15, gm_n50, gm_n9648, gm_n81);
	nor (gm_n10666, in_20, gm_n62, gm_n47, gm_n10665, in_21);
	or (gm_n10667, gm_n48, gm_n53, in_10, gm_n1398, in_13);
	nor (gm_n10668, in_16, in_15, gm_n50, gm_n10667, in_17);
	nand (gm_n10669, in_20, in_19, gm_n47, gm_n10668, in_21);
	or (gm_n10670, in_12, gm_n53, gm_n52, gm_n2931, gm_n49);
	nor (gm_n10671, in_16, in_15, gm_n50, gm_n10670, gm_n81);
	nand (gm_n10672, in_20, in_19, in_18, gm_n10671, in_21);
	nand (gm_n10673, in_12, gm_n53, in_10, gm_n4752, gm_n49);
	nor (gm_n10674, in_16, gm_n63, in_14, gm_n10673, gm_n81);
	nand (gm_n10675, gm_n45, in_19, in_18, gm_n10674, gm_n71);
	nand (gm_n10676, in_12, in_11, in_10, gm_n1227, in_13);
	nor (gm_n10677, gm_n46, in_15, gm_n50, gm_n10676, gm_n81);
	nand (gm_n10678, gm_n45, in_19, gm_n47, gm_n10677, in_21);
	nand (gm_n10679, in_11, gm_n52, in_9, gm_n3804, in_12);
	nor (gm_n10680, in_15, in_14, in_13, gm_n10679, gm_n46);
	nand (gm_n10681, gm_n62, in_18, gm_n81, gm_n10680, in_20);
	nor (gm_n10682, gm_n10681, in_21);
	and (gm_n10683, in_14, gm_n49, gm_n48, gm_n5099, in_15);
	nand (gm_n10684, gm_n47, gm_n81, gm_n46, gm_n10683, gm_n62);
	nor (gm_n10685, gm_n10684, gm_n71, in_20);
	nor (gm_n10686, in_12, in_11, gm_n52, gm_n4366, gm_n49);
	nand (gm_n10687, gm_n46, in_15, gm_n50, gm_n10686, in_17);
	nor (gm_n10688, gm_n45, in_19, in_18, gm_n10687, in_21);
	nor (gm_n10689, gm_n63, in_14, gm_n49, gm_n7492, gm_n46);
	nand (gm_n10690, in_19, in_18, in_17, gm_n10689, gm_n45);
	nor (gm_n10691, gm_n10690, in_21);
	and (gm_n10692, gm_n46, gm_n63, gm_n50, gm_n10089, gm_n81);
	nand (gm_n10693, gm_n45, in_19, in_18, gm_n10692, gm_n71);
	nor (gm_n10694, in_16, gm_n63, gm_n50, gm_n10356, in_17);
	nand (gm_n10695, gm_n45, gm_n62, gm_n47, gm_n10694, in_21);
	nand (gm_n10696, in_13, in_12, gm_n53, gm_n1328, gm_n50);
	nor (gm_n10697, in_17, in_16, gm_n63, gm_n10696, in_18);
	nand (gm_n10698, gm_n71, gm_n45, in_19, gm_n10697);
	or (gm_n10699, gm_n1735, in_10, in_9);
	or (gm_n10700, in_13, gm_n48, in_11, gm_n10699, in_14);
	nor (gm_n10701, in_17, gm_n46, in_15, gm_n10700, in_18);
	nand (gm_n10702, in_21, in_20, gm_n62, gm_n10701);
	nor (gm_n10703, in_13, in_12, in_11, gm_n3184, in_14);
	nand (gm_n10704, gm_n81, in_16, in_15, gm_n10703, gm_n47);
	nor (gm_n10705, in_21, in_20, in_19, gm_n10704);
	and (gm_n10706, in_15, in_14, gm_n49, gm_n3978, gm_n46);
	nand (gm_n10707, gm_n62, gm_n47, in_17, gm_n10706, in_20);
	nor (gm_n10708, gm_n10707, gm_n71);
	nor (gm_n10709, gm_n48, in_11, in_10, gm_n6475, in_13);
	nand (gm_n10710, in_16, gm_n63, in_14, gm_n10709, in_17);
	nor (gm_n10711, in_20, gm_n62, gm_n47, gm_n10710, gm_n71);
	nor (gm_n10712, gm_n63, in_14, in_13, gm_n7126, gm_n46);
	nand (gm_n10713, in_19, gm_n47, in_17, gm_n10712, in_20);
	nor (gm_n10714, gm_n10713, gm_n71);
	nand (gm_n10715, in_13, in_12, gm_n53, gm_n1298, gm_n50);
	nor (gm_n10716, gm_n81, in_16, gm_n63, gm_n10715, in_18);
	nand (gm_n10717, in_21, gm_n45, in_19, gm_n10716);
	or (gm_n10718, gm_n49, in_12, gm_n53, gm_n4351, in_14);
	nor (gm_n10719, gm_n81, in_16, in_15, gm_n10718, gm_n47);
	nand (gm_n10720, in_21, gm_n45, in_19, gm_n10719);
	nor (gm_n10721, in_9, in_8, in_7, gm_n843, in_10);
	nand (gm_n10722, gm_n49, in_12, in_11, gm_n10721, in_14);
	nor (gm_n10723, in_17, in_16, in_15, gm_n10722, in_18);
	nand (gm_n10724, gm_n71, in_20, gm_n62, gm_n10723);
	nor (gm_n10725, gm_n363, gm_n51);
	nand (gm_n10726, in_12, in_11, in_10, gm_n10725, in_13);
	nor (gm_n10727, gm_n46, in_15, in_14, gm_n10726, gm_n81);
	nand (gm_n10728, in_20, gm_n62, gm_n47, gm_n10727, gm_n71);
	nor (gm_n10729, gm_n48, gm_n53, in_10, gm_n7154, gm_n49);
	nand (gm_n10730, in_16, in_15, gm_n50, gm_n10729, gm_n81);
	nor (gm_n10731, gm_n45, in_19, gm_n47, gm_n10730, in_21);
	nor (gm_n10732, gm_n53, gm_n52, in_9, gm_n395);
	and (gm_n10733, in_14, gm_n49, gm_n48, gm_n10732, in_15);
	nand (gm_n10734, in_18, gm_n81, gm_n46, gm_n10733, gm_n62);
	nor (gm_n10735, gm_n10734, gm_n71, in_20);
	nor (gm_n10736, in_12, in_11, gm_n52, gm_n898, in_13);
	nand (gm_n10737, in_16, in_15, in_14, gm_n10736, in_17);
	nor (gm_n10738, gm_n45, gm_n62, in_18, gm_n10737, in_21);
	nor (gm_n10739, in_14, gm_n49, in_12, gm_n922, gm_n63);
	nand (gm_n10740, in_18, gm_n81, in_16, gm_n10739, in_19);
	nor (gm_n10741, gm_n10740, gm_n71, in_20);
	nand (gm_n10742, gm_n49, in_12, gm_n53, gm_n1696, in_14);
	nor (gm_n10743, gm_n81, in_16, gm_n63, gm_n10742, gm_n47);
	nand (gm_n10744, in_21, gm_n45, gm_n62, gm_n10743);
	and (gm_n10745, gm_n53, in_10, in_9, gm_n194, gm_n48);
	nand (gm_n10746, gm_n63, in_14, gm_n49, gm_n10745, in_16);
	nor (gm_n10747, gm_n62, in_18, gm_n81, gm_n10746, gm_n45);
	nand (gm_n10748, gm_n10747, in_21);
	nand (gm_n10749, gm_n48, in_11, gm_n52, gm_n1840, gm_n49);
	nor (gm_n10750, gm_n46, gm_n63, gm_n50, gm_n10749, in_17);
	nand (gm_n10751, gm_n45, in_19, in_18, gm_n10750, gm_n71);
	nand (gm_n10752, gm_n63, gm_n50, in_13, gm_n2960, gm_n46);
	nor (gm_n10753, gm_n62, gm_n47, in_17, gm_n10752, in_20);
	nand (gm_n10754, gm_n10753, in_21);
	and (gm_n10755, gm_n63, in_14, gm_n49, gm_n5253, gm_n46);
	nand (gm_n10756, in_19, gm_n47, gm_n81, gm_n10755, in_20);
	nor (gm_n10757, gm_n10756, gm_n71);
	or (gm_n10758, gm_n51, in_8, in_7, gm_n897, in_10);
	nor (gm_n10759, gm_n10758, in_11);
	and (gm_n10760, gm_n50, gm_n49, gm_n48, gm_n10759, gm_n63);
	nand (gm_n10761, in_18, in_17, gm_n46, gm_n10760, gm_n62);
	nor (gm_n10762, gm_n10761, gm_n71, in_20);
	nand (gm_n10763, gm_n51, in_8, in_7, gm_n151, gm_n52);
	nor (gm_n10764, in_13, in_12, in_11, gm_n10763, gm_n50);
	nand (gm_n10765, gm_n81, gm_n46, gm_n63, gm_n10764, gm_n47);
	nor (gm_n10766, in_21, in_20, gm_n62, gm_n10765);
	and (gm_n10767, in_14, gm_n49, in_12, gm_n2023, gm_n63);
	nand (gm_n10768, in_18, gm_n81, gm_n46, gm_n10767, in_19);
	nor (gm_n10769, gm_n10768, in_21, in_20);
	nor (gm_n10770, gm_n51, gm_n64, in_7, gm_n463, gm_n52);
	nand (gm_n10771, in_13, gm_n48, gm_n53, gm_n10770, gm_n50);
	nor (gm_n10772, in_17, gm_n46, gm_n63, gm_n10771, gm_n47);
	nand (gm_n10773, in_21, in_20, gm_n62, gm_n10772);
	and (gm_n10774, in_8, in_7, in_6, gm_n2640, in_9);
	nand (gm_n10775, gm_n48, in_11, gm_n52, gm_n10774, gm_n49);
	nor (gm_n10776, in_16, gm_n63, in_14, gm_n10775, in_17);
	nand (gm_n10777, gm_n45, gm_n62, in_18, gm_n10776, gm_n71);
	nor (gm_n10778, in_11, gm_n52, in_9, gm_n1098);
	nand (gm_n10779, in_14, gm_n49, gm_n48, gm_n10778, gm_n63);
	nor (gm_n10780, gm_n47, gm_n81, in_16, gm_n10779, in_19);
	nand (gm_n10781, gm_n10780, in_21, gm_n45);
	nand (gm_n10782, in_15, in_14, gm_n49, gm_n4243, gm_n46);
	nor (gm_n10783, in_19, in_18, in_17, gm_n10782, gm_n45);
	nand (gm_n10784, gm_n10783, in_21);
	nand (gm_n10785, in_8, in_7, gm_n82, gm_n1075, in_9);
	nor (gm_n10786, in_12, in_11, gm_n52, gm_n10785, in_13);
	nand (gm_n10787, gm_n46, in_15, in_14, gm_n10786, gm_n81);
	nor (gm_n10788, gm_n45, gm_n62, gm_n47, gm_n10787, in_21);
	and (gm_n10789, gm_n48, gm_n53, gm_n52, gm_n8163, in_13);
	nand (gm_n10790, gm_n46, gm_n63, gm_n50, gm_n10789, in_17);
	nor (gm_n10791, gm_n45, in_19, gm_n47, gm_n10790, gm_n71);
	and (gm_n10792, in_15, in_14, in_13, gm_n718, gm_n46);
	nand (gm_n10793, gm_n62, gm_n47, in_17, gm_n10792, gm_n45);
	nor (gm_n10794, gm_n10793, in_21);
	and (gm_n10795, gm_n49, gm_n48, in_11, gm_n1135, gm_n50);
	nand (gm_n10796, gm_n81, in_16, gm_n63, gm_n10795, gm_n47);
	nor (gm_n10797, gm_n71, gm_n45, in_19, gm_n10796);
	nor (gm_n10798, gm_n51, in_8, gm_n55, gm_n223, in_10);
	nand (gm_n10799, gm_n49, in_12, gm_n53, gm_n10798, in_14);
	nor (gm_n10800, gm_n81, gm_n46, in_15, gm_n10799, gm_n47);
	nand (gm_n10801, gm_n71, gm_n45, in_19, gm_n10800);
	and (gm_n10802, gm_n81, gm_n46, in_15, gm_n4433, in_18);
	nand (gm_n10803, in_21, in_20, in_19, gm_n10802);
	nand (gm_n10804, in_13, in_12, gm_n53, gm_n2725, in_14);
	nor (gm_n10805, gm_n81, in_16, gm_n63, gm_n10804, gm_n47);
	nand (gm_n10806, in_21, gm_n45, in_19, gm_n10805);
	nand (gm_n10807, in_13, gm_n48, gm_n53, gm_n5181, in_14);
	nor (gm_n10808, gm_n81, gm_n46, gm_n63, gm_n10807, gm_n47);
	nand (gm_n10809, gm_n71, in_20, in_19, gm_n10808);
	or (gm_n10810, gm_n53, gm_n52, gm_n51, gm_n955);
	nor (gm_n10811, gm_n50, gm_n49, in_12, gm_n10810, gm_n63);
	nand (gm_n10812, in_18, in_17, gm_n46, gm_n10811, in_19);
	nor (gm_n10813, gm_n10812, in_21, gm_n45);
	nor (gm_n10814, in_14, gm_n49, gm_n48, gm_n5084, in_15);
	nand (gm_n10815, in_18, in_17, in_16, gm_n10814, gm_n62);
	nor (gm_n10816, gm_n10815, gm_n71, gm_n45);
	nand (gm_n10817, in_11, in_10, in_9, gm_n1147, in_12);
	nor (gm_n10818, gm_n63, in_14, gm_n49, gm_n10817, gm_n46);
	nand (gm_n10819, gm_n62, in_18, in_17, gm_n10818, in_20);
	nor (gm_n10820, gm_n10819, in_21);
	and (gm_n10821, gm_n48, in_11, in_10, gm_n1307, gm_n49);
	nand (gm_n10822, gm_n46, gm_n63, gm_n50, gm_n10821, gm_n81);
	nor (gm_n10823, in_20, in_19, gm_n47, gm_n10822, in_21);
	nand (gm_n10824, in_12, in_11, gm_n52, gm_n5375, in_13);
	nor (gm_n10825, in_16, gm_n63, in_14, gm_n10824, in_17);
	nand (gm_n10826, in_20, in_19, gm_n47, gm_n10825, gm_n71);
	nand (gm_n10827, gm_n49, gm_n48, in_11, gm_n8105, in_14);
	nor (gm_n10828, gm_n81, gm_n46, in_15, gm_n10827, gm_n47);
	nand (gm_n10829, gm_n71, gm_n45, in_19, gm_n10828);
	nand (gm_n10830, gm_n63, gm_n50, in_13, gm_n3945, in_16);
	nor (gm_n10831, in_19, in_18, in_17, gm_n10830, gm_n45);
	nand (gm_n10832, gm_n10831, gm_n71);
	nand (gm_n10833, gm_n49, gm_n48, gm_n53, gm_n4209, in_14);
	nor (gm_n10834, in_17, gm_n46, gm_n63, gm_n10833, in_18);
	nand (gm_n10835, in_21, gm_n45, gm_n62, gm_n10834);
	nand (gm_n10836, gm_n53, in_10, gm_n51, gm_n2653, gm_n48);
	nor (gm_n10837, gm_n63, gm_n50, in_13, gm_n10836, gm_n46);
	nand (gm_n10838, gm_n62, in_18, in_17, gm_n10837, gm_n45);
	nor (gm_n10839, gm_n10838, in_21);
	and (gm_n10840, gm_n48, gm_n53, gm_n52, gm_n2067, gm_n49);
	nand (gm_n10841, in_16, in_15, in_14, gm_n10840, gm_n81);
	nor (gm_n10842, in_20, in_19, gm_n47, gm_n10841, in_21);
	and (gm_n10843, gm_n63, gm_n50, in_13, gm_n849, in_16);
	nand (gm_n10844, in_19, in_18, in_17, gm_n10843, gm_n45);
	nor (gm_n10845, gm_n10844, gm_n71);
	nand (gm_n10846, in_11, in_10, gm_n51, gm_n3519, gm_n48);
	nor (gm_n10847, gm_n63, gm_n50, in_13, gm_n10846, in_16);
	nand (gm_n10848, in_19, in_18, in_17, gm_n10847, in_20);
	nor (gm_n10849, gm_n10848, in_21);
	nand (gm_n10850, gm_n63, in_14, in_13, gm_n2190, in_16);
	nor (gm_n10851, in_19, in_18, in_17, gm_n10850, gm_n45);
	nand (gm_n10852, gm_n10851, gm_n71);
	and (gm_n10853, in_11, gm_n52, in_9, gm_n3193, in_12);
	nand (gm_n10854, gm_n63, in_14, gm_n49, gm_n10853, in_16);
	nor (gm_n10855, in_19, in_18, in_17, gm_n10854, gm_n45);
	nand (gm_n10856, gm_n10855, gm_n71);
	nand (gm_n10857, gm_n49, in_12, in_11, gm_n4677, gm_n50);
	nor (gm_n10858, gm_n81, gm_n46, in_15, gm_n10857, in_18);
	nand (gm_n10859, gm_n71, gm_n45, gm_n62, gm_n10858);
	nand (gm_n10860, in_15, in_14, gm_n49, gm_n5764, gm_n46);
	nor (gm_n10861, gm_n62, in_18, in_17, gm_n10860, in_20);
	nand (gm_n10862, gm_n10861, gm_n71);
	nand (gm_n10863, gm_n51, in_8, in_7, gm_n66, gm_n52);
	nor (gm_n10864, in_13, gm_n48, in_11, gm_n10863, in_14);
	nand (gm_n10865, gm_n81, in_16, gm_n63, gm_n10864, gm_n47);
	nor (gm_n10866, in_21, in_20, gm_n62, gm_n10865);
	or (gm_n10867, gm_n53, gm_n52, in_9, gm_n5263, gm_n48);
	nor (gm_n10868, gm_n63, gm_n50, gm_n49, gm_n10867, in_16);
	nand (gm_n10869, gm_n62, gm_n47, in_17, gm_n10868, in_20);
	nor (gm_n10870, gm_n10869, in_21);
	nor (gm_n10871, gm_n48, gm_n53, gm_n52, gm_n1152, in_13);
	nand (gm_n10872, gm_n46, gm_n63, gm_n50, gm_n10871, in_17);
	nor (gm_n10873, in_20, in_19, in_18, gm_n10872, gm_n71);
	and (gm_n10874, gm_n50, gm_n49, gm_n48, gm_n9778, in_15);
	nand (gm_n10875, gm_n47, gm_n81, gm_n46, gm_n10874, gm_n62);
	nor (gm_n10876, gm_n10875, in_21, gm_n45);
	nand (gm_n10877, in_13, in_12, in_11, gm_n219, in_14);
	nor (gm_n10878, gm_n81, gm_n46, in_15, gm_n10877, in_18);
	nand (gm_n10879, in_21, gm_n45, in_19, gm_n10878);
	nand (gm_n10880, gm_n49, in_12, in_11, gm_n6853, gm_n50);
	nor (gm_n10881, in_17, gm_n46, gm_n63, gm_n10880, in_18);
	nand (gm_n10882, gm_n71, in_20, in_19, gm_n10881);
	nor (gm_n10883, gm_n53, in_10, in_9, gm_n599, gm_n48);
	nand (gm_n10884, gm_n63, in_14, gm_n49, gm_n10883, gm_n46);
	nor (gm_n10885, gm_n62, in_18, in_17, gm_n10884, gm_n45);
	nand (gm_n10886, gm_n10885, in_21);
	or (gm_n10887, gm_n50, gm_n49, in_12, gm_n1460, in_15);
	nor (gm_n10888, gm_n47, gm_n81, gm_n46, gm_n10887, gm_n62);
	nand (gm_n10889, gm_n10888, gm_n71, gm_n45);
	nand (gm_n10890, in_11, in_10, in_9, gm_n1469, gm_n48);
	nor (gm_n10891, gm_n10890, in_14, in_13);
	nand (gm_n10892, in_17, in_16, gm_n63, gm_n10891, in_18);
	nor (gm_n10893, in_21, gm_n45, in_19, gm_n10892);
	nand (gm_n10894, in_17, gm_n46, gm_n63, gm_n4814, in_18);
	nor (gm_n10895, gm_n71, gm_n45, in_19, gm_n10894);
	nor (gm_n10896, gm_n63, gm_n50, gm_n49, gm_n1143, in_16);
	nand (gm_n10897, in_19, gm_n47, in_17, gm_n10896, gm_n45);
	nor (gm_n10898, gm_n10897, gm_n71);
	nor (gm_n10899, gm_n48, gm_n53, gm_n52, gm_n2052, in_13);
	nand (gm_n10900, gm_n46, in_15, in_14, gm_n10899, gm_n81);
	nor (gm_n10901, gm_n45, in_19, in_18, gm_n10900, in_21);
	nand (gm_n10902, in_12, gm_n53, in_10, gm_n1262, in_13);
	nor (gm_n10903, in_16, in_15, in_14, gm_n10902, in_17);
	nand (gm_n10904, in_20, gm_n62, gm_n47, gm_n10903, in_21);
	nand (gm_n10905, in_15, gm_n50, in_13, gm_n9375, gm_n46);
	nor (gm_n10906, gm_n62, in_18, in_17, gm_n10905, gm_n45);
	nand (gm_n10907, gm_n10906, in_21);
	nor (gm_n10908, gm_n81, in_16, gm_n63, gm_n455, gm_n47);
	nand (gm_n10909, gm_n71, gm_n45, in_19, gm_n10908);
	nand (gm_n10910, in_15, gm_n50, gm_n49, gm_n7044, in_16);
	nor (gm_n10911, gm_n62, gm_n47, gm_n81, gm_n10910, in_20);
	nand (gm_n10912, gm_n10911, gm_n71);
	nor (gm_n10913, in_14, gm_n49, gm_n48, gm_n4864, in_15);
	nand (gm_n10914, gm_n47, in_17, in_16, gm_n10913, gm_n62);
	nor (gm_n10915, gm_n10914, in_21, in_20);
	nor (gm_n10916, in_13, gm_n48, in_11, gm_n3360, gm_n50);
	nand (gm_n10917, gm_n81, gm_n46, in_15, gm_n10916, gm_n47);
	nor (gm_n10918, in_21, gm_n45, gm_n62, gm_n10917);
	nor (gm_n10919, gm_n50, gm_n49, gm_n48, gm_n7953, gm_n63);
	nand (gm_n10920, gm_n47, in_17, in_16, gm_n10919, in_19);
	nor (gm_n10921, gm_n10920, gm_n71, in_20);
	nor (gm_n10922, gm_n63, in_14, gm_n49, gm_n4134, in_16);
	nand (gm_n10923, in_19, gm_n47, gm_n81, gm_n10922, gm_n45);
	nor (gm_n10924, gm_n10923, gm_n71);
	nand (gm_n10925, in_15, in_14, in_13, gm_n4055, gm_n46);
	nor (gm_n10926, in_19, gm_n47, in_17, gm_n10925, in_20);
	nand (gm_n10927, gm_n10926, in_21);
	and (gm_n10928, gm_n53, in_10, in_9, gm_n189, in_12);
	nand (gm_n10929, in_15, gm_n50, gm_n49, gm_n10928, in_16);
	nor (gm_n10930, in_19, in_18, in_17, gm_n10929, in_20);
	nand (gm_n10931, gm_n10930, in_21);
	nand (gm_n10932, in_14, gm_n49, gm_n48, gm_n1857, in_15);
	nor (gm_n10933, in_18, gm_n81, gm_n46, gm_n10932, gm_n62);
	nand (gm_n10934, gm_n10933, gm_n71, in_20);
	nor (gm_n10935, in_16, in_15, in_14, gm_n6144, gm_n81);
	nand (gm_n10936, in_20, in_19, gm_n47, gm_n10935, in_21);
	nor (gm_n10937, in_13, gm_n48, in_11, gm_n5966, gm_n50);
	nand (gm_n10938, in_17, in_16, gm_n63, gm_n10937, gm_n47);
	nor (gm_n10939, in_21, in_20, in_19, gm_n10938);
	nor (gm_n10940, in_15, in_14, in_13, gm_n8896, gm_n46);
	nand (gm_n10941, in_19, in_18, in_17, gm_n10940, gm_n45);
	nor (gm_n10942, gm_n10941, gm_n71);
	nand (gm_n10943, gm_n53, in_10, gm_n51, gm_n3519, gm_n48);
	nor (gm_n10944, in_15, gm_n50, in_13, gm_n10943, in_16);
	nand (gm_n10945, gm_n62, in_18, in_17, gm_n10944, gm_n45);
	nor (gm_n10946, gm_n10945, in_21);
	nor (gm_n10947, gm_n49, gm_n48, gm_n53, gm_n6605, gm_n50);
	nand (gm_n10948, gm_n81, gm_n46, gm_n63, gm_n10947, in_18);
	nor (gm_n10949, in_21, gm_n45, in_19, gm_n10948);
	nand (gm_n10950, gm_n48, in_11, gm_n52, gm_n6714, gm_n49);
	nor (gm_n10951, gm_n46, gm_n63, gm_n50, gm_n10950, in_17);
	nand (gm_n10952, gm_n45, in_19, in_18, gm_n10951, in_21);
	nor (gm_n10953, in_11, gm_n52, gm_n51, gm_n1957, gm_n48);
	nand (gm_n10954, in_15, gm_n50, gm_n49, gm_n10953, in_16);
	nor (gm_n10955, gm_n62, gm_n47, in_17, gm_n10954, gm_n45);
	nand (gm_n10956, gm_n10955, gm_n71);
	nor (gm_n10957, gm_n62, gm_n47, in_17, gm_n3115, gm_n45);
	nand (gm_n10958, gm_n10957, in_21);
	nor (gm_n10959, in_11, gm_n52, in_9, gm_n8224, gm_n48);
	nand (gm_n10960, gm_n63, in_14, in_13, gm_n10959, in_16);
	nor (gm_n10961, in_19, gm_n47, in_17, gm_n10960, in_20);
	nand (gm_n10962, gm_n10961, in_21);
	nand (gm_n10963, in_14, in_13, in_12, gm_n10759, gm_n63);
	nor (gm_n10964, in_18, gm_n81, in_16, gm_n10963, in_19);
	nand (gm_n10965, gm_n10964, in_21, gm_n45);
	nand (gm_n10966, gm_n10958, gm_n10956, gm_n10952, gm_n10965, gm_n10962);
	nor (gm_n10967, gm_n10946, gm_n10942, gm_n10939, gm_n10966, gm_n10949);
	nand (gm_n10968, gm_n10934, gm_n10931, gm_n10927, gm_n10967, gm_n10936);
	nor (gm_n10969, gm_n10921, gm_n10918, gm_n10915, gm_n10968, gm_n10924);
	nand (gm_n10970, gm_n10909, gm_n10907, gm_n10904, gm_n10969, gm_n10912);
	nor (gm_n10971, gm_n10898, gm_n10895, gm_n10893, gm_n10970, gm_n10901);
	nand (gm_n10972, gm_n10886, gm_n10882, gm_n10879, gm_n10971, gm_n10889);
	nor (gm_n10973, gm_n10873, gm_n10870, gm_n10866, gm_n10972, gm_n10876);
	nand (gm_n10974, gm_n10859, gm_n10856, gm_n10852, gm_n10973, gm_n10862);
	nor (gm_n10975, gm_n10845, gm_n10842, gm_n10839, gm_n10974, gm_n10849);
	nand (gm_n10976, gm_n10832, gm_n10829, gm_n10826, gm_n10975, gm_n10835);
	nor (gm_n10977, gm_n10820, gm_n10816, gm_n10813, gm_n10976, gm_n10823);
	nand (gm_n10978, gm_n10806, gm_n10803, gm_n10801, gm_n10977, gm_n10809);
	nor (gm_n10979, gm_n10794, gm_n10791, gm_n10788, gm_n10978, gm_n10797);
	nand (gm_n10980, gm_n10781, gm_n10777, gm_n10773, gm_n10979, gm_n10784);
	nor (gm_n10981, gm_n10766, gm_n10762, gm_n10757, gm_n10980, gm_n10769);
	nand (gm_n10982, gm_n10751, gm_n10748, gm_n10744, gm_n10981, gm_n10754);
	nor (gm_n10983, gm_n10738, gm_n10735, gm_n10731, gm_n10982, gm_n10741);
	nand (gm_n10984, gm_n10724, gm_n10720, gm_n10717, gm_n10983, gm_n10728);
	nor (gm_n10985, gm_n10711, gm_n10708, gm_n10705, gm_n10984, gm_n10714);
	nand (gm_n10986, gm_n10698, gm_n10695, gm_n10693, gm_n10985, gm_n10702);
	nor (gm_n10987, gm_n10688, gm_n10685, gm_n10682, gm_n10986, gm_n10691);
	nand (gm_n10988, gm_n10675, gm_n10672, gm_n10669, gm_n10987, gm_n10678);
	nor (gm_n10989, gm_n10664, gm_n10661, gm_n10658, gm_n10988, gm_n10666);
	nand (gm_n10990, gm_n10652, gm_n10649, gm_n10646, gm_n10989, gm_n10655);
	nor (gm_n10991, gm_n10640, gm_n10637, gm_n10634, gm_n10990, gm_n10643);
	nand (gm_n10992, gm_n10628, gm_n10625, gm_n10622, gm_n10991, gm_n10631);
	nor (gm_n10993, gm_n10615, gm_n10613, gm_n10610, gm_n10992, gm_n10618);
	nand (gm_n10994, gm_n10605, gm_n10601, gm_n10598, gm_n10993, gm_n10607);
	nor (gm_n10995, gm_n10590, gm_n10587, gm_n10584, gm_n10994, gm_n10594);
	nand (gm_n10996, gm_n10578, gm_n10575, gm_n10572, gm_n10995, gm_n10582);
	nor (gm_n10997, gm_n10566, gm_n10563, gm_n10560, gm_n10996, gm_n10569);
	nand (gm_n10998, gm_n10553, gm_n10550, gm_n10546, gm_n10997, gm_n10556);
	nor (gm_n10999, gm_n10540, gm_n10538, gm_n10535, gm_n10998, gm_n10543);
	nand (gm_n11000, gm_n10530, gm_n10528, gm_n10524, gm_n10999, gm_n10533);
	nor (gm_n11001, gm_n10517, gm_n10513, gm_n10509, gm_n11000, gm_n10520);
	nand (gm_n11002, gm_n10503, gm_n10500, gm_n10497, gm_n11001, gm_n10506);
	nor (out_18, gm_n11002, gm_n10494);
	nor (gm_n11004, in_12, gm_n53, in_10, gm_n531, in_13);
	nand (gm_n11005, in_16, in_15, gm_n50, gm_n11004, in_17);
	nor (gm_n11006, in_20, in_19, gm_n47, gm_n11005, in_21);
	nand (gm_n11007, in_12, in_11, in_10, gm_n7134, in_13);
	nor (gm_n11008, in_16, gm_n63, in_14, gm_n11007, gm_n81);
	nand (gm_n11009, in_20, in_19, in_18, gm_n11008, in_21);
	nand (gm_n11010, in_12, gm_n53, gm_n52, gm_n6857, in_13);
	nor (gm_n11011, in_16, in_15, in_14, gm_n11010, gm_n81);
	nand (gm_n11012, gm_n45, gm_n62, gm_n47, gm_n11011, in_21);
	and (gm_n11013, gm_n81, in_16, gm_n63, gm_n8658, in_18);
	nand (gm_n11014, in_21, gm_n45, gm_n62, gm_n11013);
	nand (gm_n11015, in_13, gm_n48, gm_n53, gm_n1551, in_14);
	nor (gm_n11016, gm_n81, in_16, in_15, gm_n11015, in_18);
	nand (gm_n11017, in_21, gm_n45, gm_n62, gm_n11016);
	nor (gm_n11018, in_12, gm_n53, in_10, gm_n7154, in_13);
	nand (gm_n11019, gm_n46, gm_n63, in_14, gm_n11018, gm_n81);
	nor (gm_n11020, in_20, gm_n62, in_18, gm_n11019, in_21);
	nor (gm_n11021, in_12, in_11, gm_n52, gm_n2327, gm_n49);
	nand (gm_n11022, in_16, gm_n63, in_14, gm_n11021, in_17);
	nor (gm_n11023, in_20, gm_n62, in_18, gm_n11022, gm_n71);
	nand (gm_n11024, gm_n46, in_15, in_14, gm_n5424, gm_n81);
	nor (gm_n11025, in_20, gm_n62, in_18, gm_n11024, gm_n71);
	and (gm_n11026, in_13, in_12, in_11, gm_n6975, in_14);
	nand (gm_n11027, in_17, gm_n46, gm_n63, gm_n11026, gm_n47);
	nor (gm_n11028, gm_n71, gm_n45, gm_n62, gm_n11027);
	nand (gm_n11029, in_13, gm_n48, gm_n53, gm_n10120, in_14);
	nor (gm_n11030, gm_n81, in_16, in_15, gm_n11029, in_18);
	nand (gm_n11031, in_21, in_20, gm_n62, gm_n11030);
	and (gm_n11032, gm_n53, gm_n52, in_9, gm_n1874, gm_n48);
	nand (gm_n11033, in_15, in_14, gm_n49, gm_n11032, gm_n46);
	nor (gm_n11034, gm_n62, in_18, in_17, gm_n11033, gm_n45);
	nand (gm_n11035, gm_n11034, gm_n71);
	and (gm_n11036, in_10, gm_n51, gm_n64, gm_n302, in_11);
	nand (gm_n11037, in_14, gm_n49, gm_n48, gm_n11036, in_15);
	nor (gm_n11038, gm_n47, in_17, gm_n46, gm_n11037, in_19);
	nand (gm_n11039, gm_n11038, gm_n71, gm_n45);
	nor (gm_n11040, gm_n53, gm_n52, gm_n51, gm_n395);
	nand (gm_n11041, in_14, gm_n49, gm_n48, gm_n11040, in_15);
	nor (gm_n11042, in_18, gm_n81, gm_n46, gm_n11041, gm_n62);
	nand (gm_n11043, gm_n11042, gm_n71, gm_n45);
	and (gm_n11044, gm_n48, gm_n53, in_10, gm_n2555, gm_n49);
	nand (gm_n11045, gm_n46, gm_n63, in_14, gm_n11044, in_17);
	nor (gm_n11046, gm_n45, gm_n62, in_18, gm_n11045, gm_n71);
	and (gm_n11047, gm_n49, in_12, gm_n53, gm_n3291, in_14);
	nand (gm_n11048, in_17, gm_n46, gm_n63, gm_n11047, gm_n47);
	nor (gm_n11049, gm_n71, gm_n45, gm_n62, gm_n11048);
	and (gm_n11050, in_7, gm_n82, in_5, gm_n296, gm_n64);
	nand (gm_n11051, gm_n53, in_10, in_9, gm_n11050, in_12);
	nor (gm_n11052, in_15, gm_n50, in_13, gm_n11051, in_16);
	nand (gm_n11053, in_19, gm_n47, in_17, gm_n11052, in_20);
	nor (gm_n11054, gm_n11053, gm_n71);
	nand (gm_n11055, in_17, in_16, gm_n63, gm_n9114, in_18);
	nor (gm_n11056, in_21, in_20, in_19, gm_n11055);
	nand (gm_n11057, in_15, in_14, in_13, gm_n9371, in_16);
	nor (gm_n11058, in_19, in_18, gm_n81, gm_n11057, gm_n45);
	nand (gm_n11059, gm_n11058, in_21);
	nand (gm_n11060, gm_n49, in_12, in_11, gm_n579, in_14);
	nor (gm_n11061, in_17, gm_n46, gm_n63, gm_n11060, gm_n47);
	nand (gm_n11062, gm_n71, in_20, in_19, gm_n11061);
	nand (gm_n11063, in_12, gm_n53, gm_n52, gm_n7186, gm_n49);
	nor (gm_n11064, in_16, in_15, gm_n50, gm_n11063, gm_n81);
	nand (gm_n11065, gm_n45, in_19, gm_n47, gm_n11064, in_21);
	nand (gm_n11066, gm_n50, in_13, gm_n48, gm_n2035, gm_n63);
	nor (gm_n11067, in_18, in_17, in_16, gm_n11066, in_19);
	nand (gm_n11068, gm_n11067, in_21, in_20);
	and (gm_n11069, gm_n50, in_13, in_12, gm_n4090, gm_n63);
	nand (gm_n11070, in_18, gm_n81, gm_n46, gm_n11069, in_19);
	nor (gm_n11071, gm_n11070, in_21, in_20);
	and (gm_n11072, in_13, in_12, in_11, gm_n4447, gm_n50);
	nand (gm_n11073, gm_n81, in_16, gm_n63, gm_n11072, gm_n47);
	nor (gm_n11074, in_21, gm_n45, gm_n62, gm_n11073);
	and (gm_n11075, in_15, gm_n50, in_13, gm_n10521, in_16);
	nand (gm_n11076, gm_n62, in_18, gm_n81, gm_n11075, gm_n45);
	nor (gm_n11077, gm_n11076, gm_n71);
	nor (gm_n11078, gm_n50, gm_n49, gm_n48, gm_n10810, gm_n63);
	nand (gm_n11079, in_18, gm_n81, gm_n46, gm_n11078, gm_n62);
	nor (gm_n11080, gm_n11079, in_21, gm_n45);
	nand (gm_n11081, gm_n48, gm_n53, gm_n52, gm_n3566, in_13);
	nor (gm_n11082, in_16, in_15, gm_n50, gm_n11081, gm_n81);
	nand (gm_n11083, in_20, gm_n62, gm_n47, gm_n11082, in_21);
	nand (gm_n11084, gm_n48, in_11, in_10, gm_n3941, gm_n49);
	nor (gm_n11085, in_16, gm_n63, in_14, gm_n11084, in_17);
	nand (gm_n11086, gm_n45, in_19, gm_n47, gm_n11085, gm_n71);
	and (gm_n11087, gm_n47, in_17, in_16, gm_n2447, in_19);
	nand (gm_n11088, gm_n11087, gm_n71, gm_n45);
	nand (gm_n11089, in_13, gm_n48, in_11, gm_n3350, gm_n50);
	nor (gm_n11090, in_17, in_16, gm_n63, gm_n11089, gm_n47);
	nand (gm_n11091, in_21, gm_n45, gm_n62, gm_n11090);
	and (gm_n11092, gm_n50, gm_n49, gm_n48, gm_n7459, gm_n63);
	nand (gm_n11093, in_18, gm_n81, in_16, gm_n11092, in_19);
	nor (gm_n11094, gm_n11093, gm_n71, gm_n45);
	and (gm_n11095, gm_n50, gm_n49, in_12, gm_n4961, gm_n63);
	nand (gm_n11096, in_18, in_17, in_16, gm_n11095, in_19);
	nor (gm_n11097, gm_n11096, in_21, in_20);
	and (gm_n11098, gm_n49, gm_n48, in_11, gm_n6124, gm_n50);
	nand (gm_n11099, in_17, in_16, in_15, gm_n11098, gm_n47);
	nor (gm_n11100, gm_n71, in_20, gm_n62, gm_n11099);
	nand (gm_n11101, gm_n62, in_18, in_17, gm_n10086, in_20);
	nor (gm_n11102, gm_n11101, gm_n71);
	nand (gm_n11103, gm_n63, in_14, gm_n49, gm_n608, in_16);
	nor (gm_n11104, in_19, in_18, gm_n81, gm_n11103, gm_n45);
	nand (gm_n11105, gm_n11104, gm_n71);
	nor (gm_n11106, gm_n53, in_10, in_9, gm_n453, gm_n48);
	nand (gm_n11107, gm_n63, gm_n50, gm_n49, gm_n11106, gm_n46);
	nor (gm_n11108, in_19, gm_n47, gm_n81, gm_n11107, in_20);
	nand (gm_n11109, gm_n11108, in_21);
	nor (gm_n11110, gm_n81, in_16, in_15, gm_n776, gm_n47);
	nand (gm_n11111, gm_n71, in_20, gm_n62, gm_n11110);
	nand (gm_n11112, gm_n48, in_11, gm_n52, gm_n10331, in_13);
	nor (gm_n11113, in_16, in_15, in_14, gm_n11112, gm_n81);
	nand (gm_n11114, gm_n45, in_19, in_18, gm_n11113, gm_n71);
	and (gm_n11115, gm_n50, gm_n49, in_12, gm_n2627, gm_n63);
	nand (gm_n11116, in_18, gm_n81, gm_n46, gm_n11115, gm_n62);
	nor (gm_n11117, gm_n11116, gm_n71, in_20);
	nand (gm_n11118, in_18, in_17, in_16, gm_n5239, in_19);
	nor (gm_n11119, gm_n11118, gm_n71, gm_n45);
	nor (gm_n11120, in_14, in_13, in_12, gm_n2898, in_15);
	nand (gm_n11121, gm_n47, in_17, in_16, gm_n11120, in_19);
	nor (gm_n11122, gm_n11121, gm_n71, in_20);
	and (gm_n11123, in_14, gm_n49, gm_n48, gm_n5993, gm_n63);
	nand (gm_n11124, gm_n47, gm_n81, in_16, gm_n11123, in_19);
	nor (gm_n11125, gm_n11124, gm_n71, in_20);
	nand (gm_n11126, in_14, in_13, in_12, gm_n11040, in_15);
	nor (gm_n11127, in_18, in_17, gm_n46, gm_n11126, in_19);
	nand (gm_n11128, gm_n11127, in_21, in_20);
	nand (gm_n11129, gm_n50, in_13, in_12, gm_n10351, gm_n63);
	nor (gm_n11130, in_18, gm_n81, gm_n46, gm_n11129, in_19);
	nand (gm_n11131, gm_n11130, in_21, gm_n45);
	nand (gm_n11132, in_14, gm_n49, gm_n48, gm_n8516, gm_n63);
	nor (gm_n11133, gm_n47, in_17, in_16, gm_n11132, in_19);
	nand (gm_n11134, gm_n11133, in_21, in_20);
	nand (gm_n11135, in_12, in_11, in_10, gm_n8786, in_13);
	nor (gm_n11136, gm_n46, in_15, in_14, gm_n11135, gm_n81);
	nand (gm_n11137, in_20, in_19, gm_n47, gm_n11136, in_21);
	nor (gm_n11138, in_13, in_12, gm_n53, gm_n4398, gm_n50);
	nand (gm_n11139, gm_n81, in_16, gm_n63, gm_n11138, gm_n47);
	nor (gm_n11140, in_21, gm_n45, in_19, gm_n11139);
	and (gm_n11141, gm_n48, gm_n53, in_10, gm_n1700, gm_n49);
	nand (gm_n11142, gm_n46, in_15, in_14, gm_n11141, in_17);
	nor (gm_n11143, gm_n45, in_19, gm_n47, gm_n11142, gm_n71);
	and (gm_n11144, gm_n50, in_13, gm_n48, gm_n1016, gm_n63);
	nand (gm_n11145, gm_n47, in_17, in_16, gm_n11144, gm_n62);
	nor (gm_n11146, gm_n11145, gm_n71, in_20);
	and (gm_n11147, gm_n49, in_12, in_11, gm_n1298, in_14);
	nand (gm_n11148, gm_n81, gm_n46, gm_n63, gm_n11147, in_18);
	nor (gm_n11149, gm_n71, in_20, in_19, gm_n11148);
	nand (gm_n11150, in_13, in_12, gm_n53, gm_n998, in_14);
	nor (gm_n11151, in_17, gm_n46, gm_n63, gm_n11150, gm_n47);
	nand (gm_n11152, gm_n71, gm_n45, in_19, gm_n11151);
	and (gm_n11153, gm_n46, in_15, in_14, gm_n5117, gm_n81);
	nand (gm_n11154, in_20, gm_n62, in_18, gm_n11153, gm_n71);
	and (gm_n11155, in_16, in_15, in_14, gm_n3152, in_17);
	nand (gm_n11156, in_20, in_19, in_18, gm_n11155, gm_n71);
	nand (gm_n11157, in_15, in_14, in_13, gm_n976, gm_n46);
	nor (gm_n11158, gm_n62, in_18, gm_n81, gm_n11157, in_20);
	nand (gm_n11159, gm_n11158, gm_n71);
	nand (gm_n11160, gm_n81, gm_n46, in_15, gm_n771, gm_n47);
	nor (gm_n11161, in_21, in_20, in_19, gm_n11160);
	or (gm_n11162, in_11, in_10, in_9, gm_n4314, gm_n48);
	nor (gm_n11163, gm_n63, in_14, gm_n49, gm_n11162, in_16);
	nand (gm_n11164, in_19, gm_n47, in_17, gm_n11163, in_20);
	nor (gm_n11165, gm_n11164, gm_n71);
	and (gm_n11166, in_14, gm_n49, in_12, gm_n9485, in_15);
	nand (gm_n11167, gm_n47, in_17, in_16, gm_n11166, gm_n62);
	nor (gm_n11168, gm_n11167, in_21, in_20);
	and (gm_n11169, in_13, gm_n48, in_11, gm_n10344, in_14);
	nand (gm_n11170, in_17, in_16, in_15, gm_n11169, in_18);
	nor (gm_n11171, in_21, gm_n45, in_19, gm_n11170);
	and (gm_n11172, gm_n46, in_15, in_14, gm_n1837, in_17);
	nand (gm_n11173, gm_n45, gm_n62, gm_n47, gm_n11172, gm_n71);
	nand (gm_n11174, gm_n49, gm_n48, in_11, gm_n6950, in_14);
	nor (gm_n11175, gm_n81, in_16, in_15, gm_n11174, gm_n47);
	nand (gm_n11176, gm_n71, gm_n45, in_19, gm_n11175);
	nand (gm_n11177, in_13, gm_n48, in_11, gm_n3937, gm_n50);
	nor (gm_n11178, in_17, gm_n46, in_15, gm_n11177, gm_n47);
	nand (gm_n11179, in_21, in_20, gm_n62, gm_n11178);
	nand (gm_n11180, gm_n55, in_6, in_5, gm_n284, in_8);
	nor (gm_n11181, gm_n11180, in_9);
	nand (gm_n11182, in_12, in_11, in_10, gm_n11181, gm_n49);
	nor (gm_n11183, gm_n46, gm_n63, in_14, gm_n11182, in_17);
	nand (gm_n11184, in_20, gm_n62, in_18, gm_n11183, in_21);
	nand (gm_n11185, in_11, in_10, gm_n51, gm_n792, in_12);
	nor (gm_n11186, in_15, gm_n50, gm_n49, gm_n11185, in_16);
	nand (gm_n11187, gm_n62, gm_n47, in_17, gm_n11186, in_20);
	nor (gm_n11188, gm_n11187, in_21);
	nor (gm_n11189, in_12, gm_n53, in_10, gm_n1617, gm_n49);
	nand (gm_n11190, gm_n46, gm_n63, in_14, gm_n11189, gm_n81);
	nor (gm_n11191, in_20, gm_n62, in_18, gm_n11190, in_21);
	nor (gm_n11192, in_8, gm_n55, in_6, gm_n119, in_9);
	and (gm_n11193, gm_n48, in_11, gm_n52, gm_n11192, in_13);
	nand (gm_n11194, gm_n46, in_15, in_14, gm_n11193, gm_n81);
	nor (gm_n11195, gm_n45, gm_n62, in_18, gm_n11194, in_21);
	nor (gm_n11196, in_15, in_14, gm_n49, gm_n7418, gm_n46);
	nand (gm_n11197, in_19, in_18, in_17, gm_n11196, gm_n45);
	nor (gm_n11198, gm_n11197, gm_n71);
	or (gm_n11199, gm_n64, gm_n55, in_6, gm_n141, gm_n51);
	nor (gm_n11200, gm_n11199, in_11, gm_n52);
	nand (gm_n11201, in_14, in_13, in_12, gm_n11200, gm_n63);
	nor (gm_n11202, gm_n47, in_17, in_16, gm_n11201, in_19);
	nand (gm_n11203, gm_n11202, in_21, in_20);
	nand (gm_n11204, gm_n48, gm_n53, in_10, gm_n4319, in_13);
	nor (gm_n11205, in_16, in_15, in_14, gm_n11204, in_17);
	nand (gm_n11206, gm_n45, in_19, gm_n47, gm_n11205, in_21);
	nand (gm_n11207, gm_n49, in_12, gm_n53, gm_n3480, in_14);
	nor (gm_n11208, in_17, gm_n46, gm_n63, gm_n11207, gm_n47);
	nand (gm_n11209, in_21, gm_n45, in_19, gm_n11208);
	nand (gm_n11210, in_12, in_11, gm_n52, gm_n11181, gm_n49);
	nor (gm_n11211, gm_n46, gm_n63, gm_n50, gm_n11210, in_17);
	nand (gm_n11212, in_20, gm_n62, in_18, gm_n11211, in_21);
	nor (gm_n11213, in_13, in_12, in_11, gm_n2602, in_14);
	nand (gm_n11214, gm_n81, gm_n46, gm_n63, gm_n11213, gm_n47);
	nor (gm_n11215, in_21, in_20, in_19, gm_n11214);
	nor (gm_n11216, gm_n48, gm_n53, in_10, gm_n4362, in_13);
	nand (gm_n11217, in_16, gm_n63, gm_n50, gm_n11216, in_17);
	nor (gm_n11218, in_20, in_19, gm_n47, gm_n11217, gm_n71);
	nor (gm_n11219, in_13, in_12, in_11, gm_n5877, in_14);
	nand (gm_n11220, gm_n81, gm_n46, in_15, gm_n11219, gm_n47);
	nor (gm_n11221, in_21, gm_n45, in_19, gm_n11220);
	nand (gm_n11222, in_11, in_10, gm_n51, gm_n4050, gm_n48);
	nor (gm_n11223, in_15, in_14, in_13, gm_n11222, gm_n46);
	nand (gm_n11224, in_19, gm_n47, gm_n81, gm_n11223, in_20);
	nor (gm_n11225, gm_n11224, in_21);
	nand (gm_n11226, in_13, gm_n48, gm_n53, gm_n7788, gm_n50);
	nor (gm_n11227, in_17, in_16, gm_n63, gm_n11226, in_18);
	nand (gm_n11228, in_21, gm_n45, gm_n62, gm_n11227);
	or (gm_n11229, gm_n50, in_13, gm_n48, gm_n2832, in_15);
	nor (gm_n11230, gm_n47, gm_n81, in_16, gm_n11229, gm_n62);
	nand (gm_n11231, gm_n11230, gm_n71, in_20);
	nand (gm_n11232, gm_n48, in_11, gm_n52, gm_n2619, in_13);
	nor (gm_n11233, gm_n46, gm_n63, in_14, gm_n11232, gm_n81);
	nand (gm_n11234, in_20, gm_n62, gm_n47, gm_n11233, in_21);
	and (gm_n11235, in_16, in_15, in_14, gm_n2079, in_17);
	nand (gm_n11236, gm_n45, gm_n62, in_18, gm_n11235, gm_n71);
	nor (gm_n11237, in_14, gm_n49, gm_n48, gm_n1103, in_15);
	nand (gm_n11238, in_18, in_17, gm_n46, gm_n11237, in_19);
	nor (gm_n11239, gm_n11238, gm_n71, in_20);
	nand (gm_n11240, in_17, gm_n46, in_15, gm_n2231, gm_n47);
	nor (gm_n11241, in_21, in_20, gm_n62, gm_n11240);
	nor (gm_n11242, gm_n48, gm_n53, in_10, gm_n2837, gm_n49);
	nand (gm_n11243, in_16, gm_n63, gm_n50, gm_n11242, in_17);
	nor (gm_n11244, in_20, gm_n62, gm_n47, gm_n11243, gm_n71);
	nor (gm_n11245, gm_n48, in_11, in_10, gm_n6518, gm_n49);
	nand (gm_n11246, in_16, gm_n63, in_14, gm_n11245, in_17);
	nor (gm_n11247, in_20, in_19, in_18, gm_n11246, in_21);
	nand (gm_n11248, in_12, gm_n53, in_10, gm_n3785, gm_n49);
	nor (gm_n11249, gm_n46, gm_n63, in_14, gm_n11248, gm_n81);
	nand (gm_n11250, in_20, in_19, in_18, gm_n11249, in_21);
	nand (gm_n11251, gm_n48, gm_n53, gm_n52, gm_n2661, in_13);
	nor (gm_n11252, in_16, gm_n63, in_14, gm_n11251, in_17);
	nand (gm_n11253, in_20, gm_n62, gm_n47, gm_n11252, gm_n71);
	nand (gm_n11254, in_12, gm_n53, gm_n52, gm_n343, gm_n49);
	nor (gm_n11255, gm_n46, gm_n63, gm_n50, gm_n11254, in_17);
	nand (gm_n11256, in_20, in_19, gm_n47, gm_n11255, gm_n71);
	or (gm_n11257, gm_n48, in_11, gm_n52, gm_n1524, in_13);
	nor (gm_n11258, gm_n46, in_15, in_14, gm_n11257, in_17);
	nand (gm_n11259, gm_n45, gm_n62, in_18, gm_n11258, gm_n71);
	nand (gm_n11260, in_11, in_10, gm_n51, gm_n8063, in_12);
	nor (gm_n11261, gm_n63, gm_n50, in_13, gm_n11260, in_16);
	nand (gm_n11262, in_19, in_18, in_17, gm_n11261, in_20);
	nor (gm_n11263, gm_n11262, gm_n71);
	and (gm_n11264, gm_n49, gm_n48, in_11, gm_n7991, gm_n50);
	nand (gm_n11265, gm_n81, in_16, gm_n63, gm_n11264, in_18);
	nor (gm_n11266, in_21, gm_n45, in_19, gm_n11265);
	nand (gm_n11267, in_11, in_10, in_9, gm_n2631, in_12);
	nor (gm_n11268, gm_n63, in_14, in_13, gm_n11267, gm_n46);
	nand (gm_n11269, gm_n62, gm_n47, in_17, gm_n11268, gm_n45);
	nor (gm_n11270, gm_n11269, gm_n71);
	nor (gm_n11271, gm_n49, in_12, gm_n53, gm_n6702, in_14);
	nand (gm_n11272, gm_n81, gm_n46, gm_n63, gm_n11271, in_18);
	nor (gm_n11273, gm_n71, gm_n45, in_19, gm_n11272);
	nand (gm_n11274, gm_n49, in_12, gm_n53, gm_n687, in_14);
	nor (gm_n11275, gm_n81, gm_n46, gm_n63, gm_n11274, in_18);
	nand (gm_n11276, gm_n71, in_20, gm_n62, gm_n11275);
	nand (gm_n11277, in_15, gm_n50, in_13, gm_n2346, in_16);
	nor (gm_n11278, gm_n62, gm_n47, in_17, gm_n11277, in_20);
	nand (gm_n11279, gm_n11278, in_21);
	nor (gm_n11280, in_11, in_10, in_9, gm_n6155, in_12);
	nand (gm_n11281, in_15, in_14, gm_n49, gm_n11280, gm_n46);
	nor (gm_n11282, gm_n62, in_18, in_17, gm_n11281, gm_n45);
	nand (gm_n11283, gm_n11282, in_21);
	nand (gm_n11284, in_12, gm_n53, gm_n52, gm_n1365, gm_n49);
	nor (gm_n11285, in_16, gm_n63, gm_n50, gm_n11284, gm_n81);
	nand (gm_n11286, gm_n45, gm_n62, in_18, gm_n11285, in_21);
	or (gm_n11287, gm_n53, gm_n52, in_9, gm_n3198, in_12);
	nor (gm_n11288, gm_n63, gm_n50, gm_n49, gm_n11287, gm_n46);
	nand (gm_n11289, gm_n62, gm_n47, in_17, gm_n11288, in_20);
	nor (gm_n11290, gm_n11289, in_21);
	nand (gm_n11291, in_16, in_15, gm_n50, gm_n5592, gm_n81);
	nor (gm_n11292, gm_n45, in_19, in_18, gm_n11291, in_21);
	and (gm_n11293, in_14, gm_n49, in_12, gm_n10778, gm_n63);
	nand (gm_n11294, gm_n47, in_17, gm_n46, gm_n11293, in_19);
	nor (gm_n11295, gm_n11294, gm_n71, in_20);
	nor (gm_n11296, gm_n48, in_11, gm_n52, gm_n264, gm_n49);
	nand (gm_n11297, gm_n46, in_15, in_14, gm_n11296, in_17);
	nor (gm_n11298, in_20, gm_n62, in_18, gm_n11297, gm_n71);
	and (gm_n11299, in_11, gm_n52, in_9, gm_n1279, gm_n48);
	nand (gm_n11300, gm_n63, in_14, gm_n49, gm_n11299, gm_n46);
	nor (gm_n11301, in_19, in_18, in_17, gm_n11300, gm_n45);
	nand (gm_n11302, gm_n11301, gm_n71);
	nand (gm_n11303, gm_n50, gm_n49, in_12, gm_n5064, gm_n63);
	nor (gm_n11304, in_18, in_17, in_16, gm_n11303, in_19);
	nand (gm_n11305, gm_n11304, in_21, gm_n45);
	and (gm_n11306, in_16, gm_n63, gm_n50, gm_n437, gm_n81);
	nand (gm_n11307, gm_n45, in_19, gm_n47, gm_n11306, gm_n71);
	nor (gm_n11308, in_11, in_10, gm_n51, gm_n3428, gm_n48);
	nand (gm_n11309, gm_n63, gm_n50, gm_n49, gm_n11308, gm_n46);
	nor (gm_n11310, in_19, gm_n47, in_17, gm_n11309, in_20);
	nand (gm_n11311, gm_n11310, in_21);
	nand (gm_n11312, gm_n53, in_10, in_9, gm_n2229, in_12);
	nor (gm_n11313, in_15, in_14, in_13, gm_n11312, in_16);
	nand (gm_n11314, gm_n62, gm_n47, gm_n81, gm_n11313, gm_n45);
	nor (gm_n11315, gm_n11314, gm_n71);
	or (gm_n11316, gm_n46, in_15, in_14, gm_n5700, in_17);
	nor (gm_n11317, gm_n45, in_19, in_18, gm_n11316, in_21);
	nand (gm_n11318, gm_n52, in_9, gm_n64, gm_n338, in_11);
	nor (gm_n11319, in_14, in_13, in_12, gm_n11318, gm_n63);
	nand (gm_n11320, in_18, in_17, in_16, gm_n11319, in_19);
	nor (gm_n11321, gm_n11320, in_21, gm_n45);
	and (gm_n11322, gm_n48, in_11, gm_n52, gm_n2685, in_13);
	nand (gm_n11323, gm_n46, in_15, gm_n50, gm_n11322, gm_n81);
	nor (gm_n11324, in_20, gm_n62, in_18, gm_n11323, gm_n71);
	and (gm_n11325, gm_n53, in_10, gm_n51, gm_n2234, in_12);
	nand (gm_n11326, in_15, gm_n50, gm_n49, gm_n11325, in_16);
	nor (gm_n11327, in_19, gm_n47, gm_n81, gm_n11326, in_20);
	nand (gm_n11328, gm_n11327, gm_n71);
	nand (gm_n11329, in_12, gm_n53, in_10, gm_n6905, in_13);
	nor (gm_n11330, in_16, in_15, gm_n50, gm_n11329, gm_n81);
	nand (gm_n11331, in_20, in_19, in_18, gm_n11330, in_21);
	nor (gm_n11332, gm_n46, in_15, gm_n50, gm_n7116, gm_n81);
	nand (gm_n11333, in_20, in_19, gm_n47, gm_n11332, in_21);
	or (gm_n11334, in_12, gm_n53, gm_n52, gm_n97, gm_n49);
	nor (gm_n11335, gm_n46, in_15, in_14, gm_n11334, gm_n81);
	nand (gm_n11336, in_20, in_19, in_18, gm_n11335, in_21);
	or (gm_n11337, in_10, in_9, gm_n64, gm_n907, gm_n53);
	nor (gm_n11338, in_14, in_13, in_12, gm_n11337, in_15);
	nand (gm_n11339, in_18, gm_n81, gm_n46, gm_n11338, in_19);
	nor (gm_n11340, gm_n11339, in_21, in_20);
	nand (gm_n11341, in_11, gm_n52, in_9, gm_n4119, gm_n48);
	nor (gm_n11342, in_15, gm_n50, gm_n49, gm_n11341, in_16);
	nand (gm_n11343, in_19, gm_n47, in_17, gm_n11342, gm_n45);
	nor (gm_n11344, gm_n11343, gm_n71);
	or (gm_n11345, gm_n3844, gm_n52, gm_n51);
	nor (gm_n11346, in_13, in_12, gm_n53, gm_n11345, gm_n50);
	nand (gm_n11347, in_17, in_16, gm_n63, gm_n11346, in_18);
	nor (gm_n11348, gm_n71, gm_n45, in_19, gm_n11347);
	nor (gm_n11349, in_12, gm_n53, in_10, gm_n5519, gm_n49);
	nand (gm_n11350, gm_n46, gm_n63, gm_n50, gm_n11349, in_17);
	nor (gm_n11351, gm_n45, gm_n62, gm_n47, gm_n11350, in_21);
	or (gm_n11352, gm_n49, gm_n48, in_11, gm_n1588, gm_n50);
	nor (gm_n11353, in_17, gm_n46, in_15, gm_n11352, gm_n47);
	nand (gm_n11354, gm_n71, gm_n45, in_19, gm_n11353);
	nand (gm_n11355, gm_n48, in_11, in_10, gm_n8256, gm_n49);
	nor (gm_n11356, in_16, in_15, gm_n50, gm_n11355, gm_n81);
	nand (gm_n11357, gm_n45, gm_n62, in_18, gm_n11356, gm_n71);
	nand (gm_n11358, gm_n49, in_12, gm_n53, gm_n7579, in_14);
	nor (gm_n11359, gm_n81, gm_n46, gm_n63, gm_n11358, gm_n47);
	nand (gm_n11360, in_21, gm_n45, gm_n62, gm_n11359);
	nand (gm_n11361, in_12, in_11, gm_n52, gm_n6668, gm_n49);
	nor (gm_n11362, in_16, gm_n63, gm_n50, gm_n11361, gm_n81);
	nand (gm_n11363, gm_n45, gm_n62, gm_n47, gm_n11362, gm_n71);
	and (gm_n11364, gm_n48, in_11, in_10, gm_n2056, in_13);
	nand (gm_n11365, in_16, gm_n63, in_14, gm_n11364, gm_n81);
	nor (gm_n11366, in_20, gm_n62, in_18, gm_n11365, gm_n71);
	nor (gm_n11367, in_12, in_11, in_10, gm_n1076, gm_n49);
	nand (gm_n11368, gm_n46, gm_n63, in_14, gm_n11367, in_17);
	nor (gm_n11369, in_20, gm_n62, in_18, gm_n11368, in_21);
	nand (gm_n11370, gm_n53, gm_n52, in_9, gm_n868, gm_n48);
	nor (gm_n11371, gm_n63, gm_n50, gm_n49, gm_n11370, in_16);
	nand (gm_n11372, in_19, gm_n47, gm_n81, gm_n11371, gm_n45);
	nor (gm_n11373, gm_n11372, in_21);
	nor (gm_n11374, gm_n63, in_14, in_13, gm_n3336, in_16);
	nand (gm_n11375, in_19, in_18, gm_n81, gm_n11374, in_20);
	nor (gm_n11376, gm_n11375, gm_n71);
	and (gm_n11377, gm_n53, in_10, in_9, gm_n1986);
	nand (gm_n11378, gm_n50, gm_n49, gm_n48, gm_n11377, gm_n63);
	nor (gm_n11379, gm_n47, in_17, gm_n46, gm_n11378, gm_n62);
	nand (gm_n11380, gm_n11379, in_21, in_20);
	and (gm_n11381, in_16, in_15, in_14, gm_n5903, gm_n81);
	nand (gm_n11382, gm_n45, gm_n62, gm_n47, gm_n11381, in_21);
	or (gm_n11383, in_12, in_11, gm_n52, gm_n6056, gm_n49);
	nor (gm_n11384, gm_n46, in_15, in_14, gm_n11383, in_17);
	nand (gm_n11385, in_20, gm_n62, gm_n47, gm_n11384, gm_n71);
	nand (gm_n11386, in_13, gm_n48, gm_n53, gm_n2464, gm_n50);
	nor (gm_n11387, in_17, gm_n46, gm_n63, gm_n11386, gm_n47);
	nand (gm_n11388, gm_n71, in_20, in_19, gm_n11387);
	nor (gm_n11389, gm_n49, gm_n48, in_11, gm_n11345, gm_n50);
	nand (gm_n11390, in_17, gm_n46, in_15, gm_n11389, gm_n47);
	nor (gm_n11391, in_21, gm_n45, gm_n62, gm_n11390);
	nand (gm_n11392, gm_n46, gm_n63, gm_n50, gm_n7817, gm_n81);
	nor (gm_n11393, gm_n45, gm_n62, gm_n47, gm_n11392, gm_n71);
	and (gm_n11394, gm_n50, in_13, gm_n48, gm_n7358, gm_n63);
	nand (gm_n11395, gm_n47, in_17, gm_n46, gm_n11394, gm_n62);
	nor (gm_n11396, gm_n11395, in_21, in_20);
	nor (gm_n11397, in_13, in_12, gm_n53, gm_n2015, in_14);
	nand (gm_n11398, gm_n81, gm_n46, gm_n63, gm_n11397, gm_n47);
	nor (gm_n11399, in_21, gm_n45, in_19, gm_n11398);
	nor (gm_n11400, in_11, gm_n52, in_9, gm_n2564, gm_n48);
	nand (gm_n11401, in_15, gm_n50, in_13, gm_n11400, gm_n46);
	nor (gm_n11402, gm_n62, in_18, in_17, gm_n11401, gm_n45);
	nand (gm_n11403, gm_n11402, in_21);
	nand (gm_n11404, in_12, gm_n53, in_10, gm_n200, gm_n49);
	nor (gm_n11405, gm_n46, in_15, in_14, gm_n11404, gm_n81);
	nand (gm_n11406, in_20, in_19, gm_n47, gm_n11405, gm_n71);
	or (gm_n11407, gm_n50, gm_n49, in_12, gm_n11337, gm_n63);
	nor (gm_n11408, in_18, gm_n81, in_16, gm_n11407, in_19);
	nand (gm_n11409, gm_n11408, gm_n71, gm_n45);
	nand (gm_n11410, gm_n48, in_11, in_10, gm_n3287, gm_n49);
	nor (gm_n11411, gm_n46, gm_n63, gm_n50, gm_n11410, in_17);
	nand (gm_n11412, in_20, in_19, gm_n47, gm_n11411, gm_n71);
	or (gm_n11413, in_16, in_15, in_14, gm_n7644, gm_n81);
	nor (gm_n11414, in_20, in_19, gm_n47, gm_n11413, in_21);
	nor (gm_n11415, in_14, in_13, gm_n48, gm_n9602, gm_n63);
	nand (gm_n11416, in_18, gm_n81, gm_n46, gm_n11415, in_19);
	nor (gm_n11417, gm_n11416, in_21, gm_n45);
	nand (gm_n11418, gm_n53, gm_n52, gm_n51, gm_n2034, in_12);
	nor (gm_n11419, in_15, in_14, gm_n49, gm_n11418, in_16);
	nand (gm_n11420, gm_n62, in_18, gm_n81, gm_n11419, gm_n45);
	nor (gm_n11421, gm_n11420, gm_n71);
	nor (gm_n11422, gm_n50, in_13, gm_n48, gm_n6917, in_15);
	nand (gm_n11423, gm_n47, in_17, in_16, gm_n11422, in_19);
	nor (gm_n11424, gm_n11423, gm_n71, gm_n45);
	nand (gm_n11425, gm_n49, in_12, gm_n53, gm_n5881, in_14);
	nor (gm_n11426, gm_n81, gm_n46, gm_n63, gm_n11425, gm_n47);
	nand (gm_n11427, gm_n71, in_20, in_19, gm_n11426);
	nor (gm_n11428, gm_n81, gm_n46, gm_n63, gm_n5566, in_18);
	nand (gm_n11429, gm_n71, gm_n45, in_19, gm_n11428);
	nor (gm_n11430, gm_n46, gm_n63, in_14, gm_n1983, gm_n81);
	nand (gm_n11431, in_20, in_19, gm_n47, gm_n11430, gm_n71);
	nor (gm_n11432, in_18, gm_n81, gm_n46, gm_n7085, in_19);
	nand (gm_n11433, gm_n11432, in_21, in_20);
	nand (gm_n11434, in_11, in_10, gm_n51, gm_n355, in_12);
	nor (gm_n11435, in_15, gm_n50, in_13, gm_n11434, in_16);
	nand (gm_n11436, gm_n62, gm_n47, gm_n81, gm_n11435, gm_n45);
	nor (gm_n11437, gm_n11436, in_21);
	nor (gm_n11438, in_12, gm_n53, in_10, gm_n10110, gm_n49);
	nand (gm_n11439, gm_n46, gm_n63, in_14, gm_n11438, gm_n81);
	nor (gm_n11440, in_20, in_19, gm_n47, gm_n11439, gm_n71);
	and (gm_n11441, gm_n48, gm_n53, gm_n52, gm_n2097, in_13);
	nand (gm_n11442, gm_n46, gm_n63, gm_n50, gm_n11441, in_17);
	nor (gm_n11443, gm_n45, in_19, gm_n47, gm_n11442, gm_n71);
	nor (gm_n11444, gm_n49, in_12, gm_n53, gm_n2428, in_14);
	nand (gm_n11445, in_17, in_16, in_15, gm_n11444, in_18);
	nor (gm_n11446, in_21, gm_n45, gm_n62, gm_n11445);
	nand (gm_n11447, in_13, gm_n48, in_11, gm_n8012, gm_n50);
	nor (gm_n11448, gm_n81, in_16, in_15, gm_n11447, gm_n47);
	nand (gm_n11449, in_21, in_20, in_19, gm_n11448);
	and (gm_n11450, gm_n548, gm_n51);
	nand (gm_n11451, gm_n48, in_11, in_10, gm_n11450, in_13);
	nor (gm_n11452, gm_n46, gm_n63, in_14, gm_n11451, gm_n81);
	nand (gm_n11453, gm_n45, gm_n62, in_18, gm_n11452, gm_n71);
	nand (gm_n11454, gm_n49, in_12, gm_n53, gm_n8881, gm_n50);
	nor (gm_n11455, in_17, gm_n46, gm_n63, gm_n11454, in_18);
	nand (gm_n11456, in_21, gm_n45, in_19, gm_n11455);
	nor (gm_n11457, gm_n53, gm_n52, gm_n51, gm_n1803, in_12);
	nand (gm_n11458, in_15, in_14, gm_n49, gm_n11457, gm_n46);
	nor (gm_n11459, in_19, in_18, in_17, gm_n11458, gm_n45);
	nand (gm_n11460, gm_n11459, gm_n71);
	nand (gm_n11461, gm_n50, gm_n49, in_12, gm_n10732, in_15);
	nor (gm_n11462, in_18, gm_n81, in_16, gm_n11461, in_19);
	nand (gm_n11463, gm_n11462, gm_n71, gm_n45);
	nand (gm_n11464, gm_n11456, gm_n11453, gm_n11449, gm_n11463, gm_n11460);
	nor (gm_n11465, gm_n11443, gm_n11440, gm_n11437, gm_n11464, gm_n11446);
	nand (gm_n11466, gm_n11431, gm_n11429, gm_n11427, gm_n11465, gm_n11433);
	nor (gm_n11467, gm_n11421, gm_n11417, gm_n11414, gm_n11466, gm_n11424);
	nand (gm_n11468, gm_n11409, gm_n11406, gm_n11403, gm_n11467, gm_n11412);
	nor (gm_n11469, gm_n11396, gm_n11393, gm_n11391, gm_n11468, gm_n11399);
	nand (gm_n11470, gm_n11385, gm_n11382, gm_n11380, gm_n11469, gm_n11388);
	nor (gm_n11471, gm_n11373, gm_n11369, gm_n11366, gm_n11470, gm_n11376);
	nand (gm_n11472, gm_n11360, gm_n11357, gm_n11354, gm_n11471, gm_n11363);
	nor (gm_n11473, gm_n11348, gm_n11344, gm_n11340, gm_n11472, gm_n11351);
	nand (gm_n11474, gm_n11333, gm_n11331, gm_n11328, gm_n11473, gm_n11336);
	nor (gm_n11475, gm_n11321, gm_n11317, gm_n11315, gm_n11474, gm_n11324);
	nand (gm_n11476, gm_n11307, gm_n11305, gm_n11302, gm_n11475, gm_n11311);
	nor (gm_n11477, gm_n11295, gm_n11292, gm_n11290, gm_n11476, gm_n11298);
	nand (gm_n11478, gm_n11283, gm_n11279, gm_n11276, gm_n11477, gm_n11286);
	nor (gm_n11479, gm_n11270, gm_n11266, gm_n11263, gm_n11478, gm_n11273);
	nand (gm_n11480, gm_n11256, gm_n11253, gm_n11250, gm_n11479, gm_n11259);
	nor (gm_n11481, gm_n11244, gm_n11241, gm_n11239, gm_n11480, gm_n11247);
	nand (gm_n11482, gm_n11234, gm_n11231, gm_n11228, gm_n11481, gm_n11236);
	nor (gm_n11483, gm_n11221, gm_n11218, gm_n11215, gm_n11482, gm_n11225);
	nand (gm_n11484, gm_n11209, gm_n11206, gm_n11203, gm_n11483, gm_n11212);
	nor (gm_n11485, gm_n11195, gm_n11191, gm_n11188, gm_n11484, gm_n11198);
	nand (gm_n11486, gm_n11179, gm_n11176, gm_n11173, gm_n11485, gm_n11184);
	nor (gm_n11487, gm_n11168, gm_n11165, gm_n11161, gm_n11486, gm_n11171);
	nand (gm_n11488, gm_n11156, gm_n11154, gm_n11152, gm_n11487, gm_n11159);
	nor (gm_n11489, gm_n11146, gm_n11143, gm_n11140, gm_n11488, gm_n11149);
	nand (gm_n11490, gm_n11134, gm_n11131, gm_n11128, gm_n11489, gm_n11137);
	nor (gm_n11491, gm_n11122, gm_n11119, gm_n11117, gm_n11490, gm_n11125);
	nand (gm_n11492, gm_n11111, gm_n11109, gm_n11105, gm_n11491, gm_n11114);
	nor (gm_n11493, gm_n11100, gm_n11097, gm_n11094, gm_n11492, gm_n11102);
	nand (gm_n11494, gm_n11088, gm_n11086, gm_n11083, gm_n11493, gm_n11091);
	nor (gm_n11495, gm_n11077, gm_n11074, gm_n11071, gm_n11494, gm_n11080);
	nand (gm_n11496, gm_n11065, gm_n11062, gm_n11059, gm_n11495, gm_n11068);
	nor (gm_n11497, gm_n11054, gm_n11049, gm_n11046, gm_n11496, gm_n11056);
	nand (gm_n11498, gm_n11039, gm_n11035, gm_n11031, gm_n11497, gm_n11043);
	nor (gm_n11499, gm_n11025, gm_n11023, gm_n11020, gm_n11498, gm_n11028);
	nand (gm_n11500, gm_n11014, gm_n11012, gm_n11009, gm_n11499, gm_n11017);
	nor (out_19, gm_n11500, gm_n11006);
	and (gm_n11502, gm_n49, in_12, gm_n53, gm_n2305, gm_n50);
	nand (gm_n11503, in_17, in_16, gm_n63, gm_n11502, in_18);
	nor (gm_n11504, gm_n71, in_20, gm_n62, gm_n11503);
	nand (gm_n11505, in_20, gm_n62, in_18, gm_n7050, gm_n71);
	nand (gm_n11506, gm_n49, in_12, gm_n53, gm_n2262, in_14);
	nor (gm_n11507, gm_n81, in_16, in_15, gm_n11506, gm_n47);
	nand (gm_n11508, gm_n71, gm_n45, gm_n62, gm_n11507);
	and (gm_n11509, in_17, gm_n46, in_15, gm_n10891, in_18);
	nand (gm_n11510, gm_n71, in_20, in_19, gm_n11509);
	nand (gm_n11511, in_12, in_11, gm_n52, gm_n9426, gm_n49);
	nor (gm_n11512, gm_n46, in_15, in_14, gm_n11511, gm_n81);
	nand (gm_n11513, in_20, gm_n62, in_18, gm_n11512, in_21);
	and (gm_n11514, in_12, in_11, gm_n52, gm_n1759, in_13);
	nand (gm_n11515, in_16, gm_n63, gm_n50, gm_n11514, in_17);
	nor (gm_n11516, in_20, gm_n62, in_18, gm_n11515, gm_n71);
	nor (gm_n11517, gm_n3844, gm_n52, in_9);
	and (gm_n11518, gm_n49, gm_n48, gm_n53, gm_n11517, in_14);
	nand (gm_n11519, gm_n81, gm_n46, gm_n63, gm_n11518, in_18);
	nor (gm_n11520, in_21, in_20, in_19, gm_n11519);
	nand (gm_n11521, gm_n46, in_15, gm_n50, gm_n9322, gm_n81);
	nor (gm_n11522, in_20, gm_n62, gm_n47, gm_n11521, in_21);
	and (gm_n11523, gm_n48, in_11, gm_n52, gm_n10725, in_13);
	nand (gm_n11524, in_16, in_15, in_14, gm_n11523, in_17);
	nor (gm_n11525, gm_n45, in_19, in_18, gm_n11524, in_21);
	nand (gm_n11526, gm_n48, gm_n53, gm_n52, gm_n5206, gm_n49);
	nor (gm_n11527, gm_n46, gm_n63, in_14, gm_n11526, gm_n81);
	nand (gm_n11528, in_20, in_19, in_18, gm_n11527, gm_n71);
	nand (gm_n11529, gm_n48, in_11, in_10, gm_n4876, gm_n49);
	nor (gm_n11530, gm_n46, in_15, gm_n50, gm_n11529, in_17);
	nand (gm_n11531, gm_n45, in_19, in_18, gm_n11530, in_21);
	nor (gm_n11532, in_18, in_17, gm_n46, gm_n3946, in_19);
	nand (gm_n11533, gm_n11532, gm_n71, gm_n45);
	nand (gm_n11534, in_15, gm_n50, gm_n49, gm_n3558, in_16);
	nor (gm_n11535, gm_n62, gm_n47, in_17, gm_n11534, in_20);
	nand (gm_n11536, gm_n11535, in_21);
	and (gm_n11537, gm_n50, in_13, in_12, gm_n10525, in_15);
	nand (gm_n11538, in_18, in_17, in_16, gm_n11537, gm_n62);
	nor (gm_n11539, gm_n11538, gm_n71, in_20);
	or (gm_n11540, in_16, in_15, gm_n50, gm_n6736, gm_n81);
	nor (gm_n11541, in_20, in_19, gm_n47, gm_n11540, gm_n71);
	nand (gm_n11542, gm_n53, gm_n52, in_9, gm_n1212, in_12);
	nor (gm_n11543, in_15, in_14, gm_n49, gm_n11542, in_16);
	nand (gm_n11544, gm_n62, in_18, gm_n81, gm_n11543, in_20);
	nor (gm_n11545, gm_n11544, gm_n71);
	nor (gm_n11546, in_12, gm_n53, gm_n52, gm_n6672, in_13);
	nand (gm_n11547, gm_n46, in_15, gm_n50, gm_n11546, gm_n81);
	nor (gm_n11548, in_20, gm_n62, gm_n47, gm_n11547, gm_n71);
	and (gm_n11549, gm_n53, in_10, gm_n51, gm_n114, gm_n48);
	nand (gm_n11550, in_15, gm_n50, in_13, gm_n11549, gm_n46);
	nor (gm_n11551, gm_n62, in_18, gm_n81, gm_n11550, gm_n45);
	nand (gm_n11552, gm_n11551, in_21);
	nand (gm_n11553, in_14, gm_n49, gm_n48, gm_n6069, in_15);
	nor (gm_n11554, in_18, in_17, gm_n46, gm_n11553, in_19);
	nand (gm_n11555, gm_n11554, in_21, gm_n45);
	nand (gm_n11556, gm_n50, gm_n49, in_12, gm_n10025, in_15);
	nor (gm_n11557, gm_n47, in_17, in_16, gm_n11556, in_19);
	nand (gm_n11558, gm_n11557, gm_n71, in_20);
	nand (gm_n11559, in_12, gm_n53, in_10, gm_n1394, in_13);
	nor (gm_n11560, in_16, gm_n63, gm_n50, gm_n11559, gm_n81);
	nand (gm_n11561, gm_n45, in_19, in_18, gm_n11560, in_21);
	nand (gm_n11562, in_16, in_15, gm_n50, gm_n3765, in_17);
	nor (gm_n11563, in_20, gm_n62, in_18, gm_n11562, gm_n71);
	nor (gm_n11564, in_13, gm_n48, gm_n53, gm_n5414, gm_n50);
	nand (gm_n11565, gm_n81, gm_n46, in_15, gm_n11564, in_18);
	nor (gm_n11566, gm_n71, gm_n45, gm_n62, gm_n11565);
	and (gm_n11567, in_11, in_10, gm_n51, gm_n2508, gm_n48);
	nand (gm_n11568, gm_n11567, in_14, gm_n49);
	or (gm_n11569, in_17, gm_n46, in_15, gm_n11568, in_18);
	nor (gm_n11570, gm_n71, in_20, gm_n62, gm_n11569);
	nor (gm_n11571, in_12, gm_n53, in_10, gm_n1744, in_13);
	nand (gm_n11572, in_16, in_15, gm_n50, gm_n11571, gm_n81);
	nor (gm_n11573, in_20, gm_n62, in_18, gm_n11572, in_21);
	nand (gm_n11574, gm_n48, gm_n53, gm_n52, gm_n7765, in_13);
	nor (gm_n11575, in_16, in_15, gm_n50, gm_n11574, gm_n81);
	nand (gm_n11576, in_20, gm_n62, in_18, gm_n11575, gm_n71);
	nand (gm_n11577, gm_n48, gm_n53, gm_n52, gm_n10211, in_13);
	nor (gm_n11578, gm_n46, in_15, in_14, gm_n11577, in_17);
	nand (gm_n11579, in_20, in_19, in_18, gm_n11578, gm_n71);
	or (gm_n11580, in_12, in_11, gm_n52, gm_n4262, gm_n49);
	nor (gm_n11581, gm_n46, in_15, gm_n50, gm_n11580, in_17);
	nand (gm_n11582, gm_n45, gm_n62, in_18, gm_n11581, in_21);
	and (gm_n11583, in_11, gm_n52, in_9, gm_n538, in_12);
	nand (gm_n11584, gm_n63, gm_n50, in_13, gm_n11583, in_16);
	nor (gm_n11585, gm_n62, gm_n47, gm_n81, gm_n11584, gm_n45);
	nand (gm_n11586, gm_n11585, gm_n71);
	nor (gm_n11587, in_13, gm_n48, gm_n53, gm_n7319, gm_n50);
	nand (gm_n11588, gm_n81, in_16, in_15, gm_n11587, gm_n47);
	nor (gm_n11589, in_21, gm_n45, in_19, gm_n11588);
	and (gm_n11590, gm_n49, in_12, gm_n53, gm_n9492, gm_n50);
	nand (gm_n11591, gm_n81, in_16, gm_n63, gm_n11590, gm_n47);
	nor (gm_n11592, in_21, in_20, gm_n62, gm_n11591);
	nand (gm_n11593, gm_n46, gm_n63, gm_n50, gm_n8160, in_17);
	nor (gm_n11594, in_20, in_19, in_18, gm_n11593, gm_n71);
	nor (gm_n11595, gm_n50, in_13, gm_n48, gm_n9502, in_15);
	nand (gm_n11596, in_18, in_17, gm_n46, gm_n11595, in_19);
	nor (gm_n11597, gm_n11596, in_21, in_20);
	and (gm_n11598, in_11, gm_n52, gm_n51, gm_n1070, in_12);
	nand (gm_n11599, in_15, in_14, in_13, gm_n11598, in_16);
	nor (gm_n11600, gm_n62, gm_n47, in_17, gm_n11599, gm_n45);
	nand (gm_n11601, gm_n11600, gm_n71);
	nand (gm_n11602, in_12, gm_n53, in_10, gm_n6294, in_13);
	nor (gm_n11603, gm_n46, in_15, in_14, gm_n11602, gm_n81);
	nand (gm_n11604, gm_n45, gm_n62, in_18, gm_n11603, gm_n71);
	nand (gm_n11605, gm_n50, in_13, in_12, gm_n10579, in_15);
	nor (gm_n11606, gm_n47, gm_n81, gm_n46, gm_n11605, in_19);
	nand (gm_n11607, gm_n11606, gm_n71, gm_n45);
	nand (gm_n11608, in_13, gm_n48, in_11, gm_n5315, in_14);
	nor (gm_n11609, in_17, gm_n46, in_15, gm_n11608, in_18);
	nand (gm_n11610, in_21, in_20, in_19, gm_n11609);
	nor (gm_n11611, in_12, in_11, in_10, gm_n6056, in_13);
	nand (gm_n11612, in_16, in_15, in_14, gm_n11611, gm_n81);
	nor (gm_n11613, gm_n45, gm_n62, in_18, gm_n11612, in_21);
	and (gm_n11614, in_12, in_11, in_10, gm_n380, gm_n49);
	nand (gm_n11615, in_16, in_15, in_14, gm_n11614, in_17);
	nor (gm_n11616, gm_n45, in_19, gm_n47, gm_n11615, gm_n71);
	and (gm_n11617, in_14, gm_n49, gm_n48, gm_n5595, in_15);
	nand (gm_n11618, in_18, in_17, gm_n46, gm_n11617, gm_n62);
	nor (gm_n11619, gm_n11618, in_21, gm_n45);
	and (gm_n11620, in_12, in_11, in_10, gm_n3553, gm_n49);
	nand (gm_n11621, in_16, gm_n63, in_14, gm_n11620, in_17);
	nor (gm_n11622, in_20, gm_n62, gm_n47, gm_n11621, in_21);
	and (gm_n11623, in_18, in_17, gm_n46, gm_n2302, gm_n62);
	nand (gm_n11624, gm_n11623, in_21, gm_n45);
	nand (gm_n11625, gm_n49, in_12, in_11, gm_n6401, in_14);
	nor (gm_n11626, gm_n81, in_16, gm_n63, gm_n11625, in_18);
	nand (gm_n11627, in_21, in_20, in_19, gm_n11626);
	nand (gm_n11628, gm_n48, in_11, gm_n52, gm_n3562, in_13);
	nor (gm_n11629, gm_n46, gm_n63, in_14, gm_n11628, gm_n81);
	nand (gm_n11630, gm_n45, gm_n62, gm_n47, gm_n11629, gm_n71);
	nand (gm_n11631, gm_n48, gm_n53, gm_n52, gm_n7984, gm_n49);
	nor (gm_n11632, gm_n46, gm_n63, gm_n50, gm_n11631, gm_n81);
	nand (gm_n11633, in_20, in_19, in_18, gm_n11632, gm_n71);
	or (gm_n11634, in_17, gm_n46, in_15, gm_n8918, in_18);
	nor (gm_n11635, in_21, gm_n45, gm_n62, gm_n11634);
	nor (gm_n11636, in_9, gm_n64, in_7, gm_n588, in_10);
	and (gm_n11637, gm_n49, in_12, in_11, gm_n11636, in_14);
	nand (gm_n11638, gm_n81, in_16, in_15, gm_n11637, in_18);
	nor (gm_n11639, gm_n71, in_20, gm_n62, gm_n11638);
	and (gm_n11640, gm_n48, gm_n53, in_10, gm_n6539, gm_n49);
	nand (gm_n11641, gm_n46, in_15, gm_n50, gm_n11640, gm_n81);
	nor (gm_n11642, in_20, in_19, gm_n47, gm_n11641, in_21);
	and (gm_n11643, in_13, in_12, in_11, gm_n1799, gm_n50);
	nand (gm_n11644, gm_n81, in_16, gm_n63, gm_n11643, in_18);
	nor (gm_n11645, gm_n71, in_20, gm_n62, gm_n11644);
	and (gm_n11646, in_11, in_10, gm_n51, gm_n7055, in_12);
	nand (gm_n11647, in_15, in_14, in_13, gm_n11646, gm_n46);
	nor (gm_n11648, in_19, in_18, in_17, gm_n11647, gm_n45);
	nand (gm_n11649, gm_n11648, gm_n71);
	nand (gm_n11650, gm_n50, gm_n49, gm_n48, gm_n9292, in_15);
	nor (gm_n11651, gm_n47, in_17, in_16, gm_n11650, in_19);
	nand (gm_n11652, gm_n11651, in_21, in_20);
	and (gm_n11653, in_10, gm_n51, gm_n64, gm_n5788, gm_n53);
	nand (gm_n11654, gm_n50, gm_n49, gm_n48, gm_n11653, in_15);
	nor (gm_n11655, in_18, in_17, in_16, gm_n11654, in_19);
	nand (gm_n11656, gm_n11655, in_21, in_20);
	nand (gm_n11657, in_13, gm_n48, gm_n53, gm_n3480, gm_n50);
	nor (gm_n11658, in_17, in_16, in_15, gm_n11657, gm_n47);
	nand (gm_n11659, gm_n71, in_20, in_19, gm_n11658);
	and (gm_n11660, gm_n71, in_20, in_19, gm_n1641);
	nand (gm_n11661, in_18, in_17, gm_n46, gm_n7565, gm_n62);
	nor (gm_n11662, gm_n11661, in_21, gm_n45);
	nor (gm_n11663, gm_n48, in_11, in_10, gm_n10042, gm_n49);
	nand (gm_n11664, gm_n46, in_15, in_14, gm_n11663, in_17);
	nor (gm_n11665, gm_n45, gm_n62, in_18, gm_n11664, in_21);
	nand (gm_n11666, in_11, in_10, gm_n51, gm_n1156, gm_n48);
	nor (gm_n11667, gm_n63, in_14, gm_n49, gm_n11666, gm_n46);
	nand (gm_n11668, in_19, in_18, in_17, gm_n11667, gm_n45);
	nor (gm_n11669, gm_n11668, in_21);
	nand (gm_n11670, in_15, in_14, in_13, gm_n6514, in_16);
	nor (gm_n11671, in_19, gm_n47, gm_n81, gm_n11670, in_20);
	nand (gm_n11672, gm_n11671, gm_n71);
	nand (gm_n11673, gm_n50, in_13, in_12, gm_n9945, in_15);
	nor (gm_n11674, in_18, gm_n81, in_16, gm_n11673, in_19);
	nand (gm_n11675, gm_n11674, gm_n71, gm_n45);
	and (gm_n11676, in_18, in_17, in_16, gm_n11338, in_19);
	nand (gm_n11677, gm_n11676, in_21, in_20);
	nor (gm_n11678, in_9, gm_n64, in_7, gm_n897, gm_n52);
	nand (gm_n11679, gm_n49, in_12, in_11, gm_n11678, in_14);
	nor (gm_n11680, in_17, gm_n46, in_15, gm_n11679, gm_n47);
	nand (gm_n11681, in_21, gm_n45, in_19, gm_n11680);
	nand (gm_n11682, in_17, gm_n46, in_15, gm_n9386, gm_n47);
	nor (gm_n11683, in_21, gm_n45, in_19, gm_n11682);
	and (gm_n11684, in_12, gm_n53, gm_n52, gm_n9722, in_13);
	nand (gm_n11685, in_16, gm_n63, gm_n50, gm_n11684, in_17);
	nor (gm_n11686, in_20, gm_n62, in_18, gm_n11685, in_21);
	nor (gm_n11687, gm_n50, in_13, in_12, gm_n8994, in_15);
	nand (gm_n11688, gm_n47, gm_n81, in_16, gm_n11687, in_19);
	nor (gm_n11689, gm_n11688, in_21, in_20);
	nor (gm_n11690, in_13, in_12, gm_n53, gm_n5816, in_14);
	nand (gm_n11691, in_17, in_16, in_15, gm_n11690, gm_n47);
	nor (gm_n11692, in_21, in_20, gm_n62, gm_n11691);
	nor (gm_n11693, in_8, gm_n55, gm_n82, gm_n530, in_9);
	nand (gm_n11694, gm_n48, in_11, in_10, gm_n11693, in_13);
	nor (gm_n11695, in_16, in_15, in_14, gm_n11694, gm_n81);
	nand (gm_n11696, gm_n45, in_19, in_18, gm_n11695, gm_n71);
	nor (gm_n11697, in_11, gm_n52, in_9, gm_n2503, in_12);
	nand (gm_n11698, gm_n63, in_14, gm_n49, gm_n11697, in_16);
	nor (gm_n11699, gm_n62, gm_n47, in_17, gm_n11698, gm_n45);
	nand (gm_n11700, gm_n11699, in_21);
	and (gm_n11701, gm_n47, in_17, gm_n46, gm_n3148, in_19);
	nand (gm_n11702, gm_n11701, gm_n71, gm_n45);
	or (gm_n11703, in_12, in_11, in_10, gm_n3809, in_13);
	nor (gm_n11704, in_16, in_15, gm_n50, gm_n11703, gm_n81);
	nand (gm_n11705, gm_n45, gm_n62, in_18, gm_n11704, gm_n71);
	and (gm_n11706, in_12, gm_n53, in_10, gm_n10180, gm_n49);
	nand (gm_n11707, in_16, gm_n63, in_14, gm_n11706, in_17);
	nor (gm_n11708, gm_n45, gm_n62, in_18, gm_n11707, gm_n71);
	nor (gm_n11709, in_13, in_12, gm_n53, gm_n7823, in_14);
	nand (gm_n11710, in_17, gm_n46, in_15, gm_n11709, in_18);
	nor (gm_n11711, gm_n71, gm_n45, in_19, gm_n11710);
	nor (gm_n11712, gm_n49, gm_n48, in_11, gm_n5760, gm_n50);
	nand (gm_n11713, in_17, gm_n46, in_15, gm_n11712, gm_n47);
	nor (gm_n11714, gm_n71, gm_n45, in_19, gm_n11713);
	nor (gm_n11715, gm_n49, in_12, gm_n53, gm_n7206, gm_n50);
	nand (gm_n11716, in_17, in_16, gm_n63, gm_n11715, gm_n47);
	nor (gm_n11717, in_21, in_20, gm_n62, gm_n11716);
	nand (gm_n11718, in_12, gm_n53, gm_n52, gm_n2555, in_13);
	nor (gm_n11719, in_16, in_15, gm_n50, gm_n11718, in_17);
	nand (gm_n11720, in_20, gm_n62, gm_n47, gm_n11719, in_21);
	nand (gm_n11721, gm_n49, gm_n48, in_11, gm_n7661, in_14);
	nor (gm_n11722, gm_n81, in_16, in_15, gm_n11721, in_18);
	nand (gm_n11723, gm_n71, in_20, gm_n62, gm_n11722);
	nand (gm_n11724, in_12, gm_n53, gm_n52, gm_n380, in_13);
	nor (gm_n11725, in_16, gm_n63, in_14, gm_n11724, in_17);
	nand (gm_n11726, in_20, gm_n62, in_18, gm_n11725, in_21);
	nand (gm_n11727, in_13, in_12, in_11, gm_n9189, in_14);
	nor (gm_n11728, in_17, in_16, gm_n63, gm_n11727, gm_n47);
	nand (gm_n11729, gm_n71, gm_n45, gm_n62, gm_n11728);
	nor (gm_n11730, in_13, in_12, in_11, gm_n1003, in_14);
	nand (gm_n11731, in_17, in_16, gm_n63, gm_n11730, in_18);
	nor (gm_n11732, gm_n71, gm_n45, in_19, gm_n11731);
	nand (gm_n11733, in_11, gm_n52, gm_n51, gm_n3183, gm_n48);
	nor (gm_n11734, in_15, gm_n50, in_13, gm_n11733, gm_n46);
	nand (gm_n11735, in_19, gm_n47, in_17, gm_n11734, in_20);
	nor (gm_n11736, gm_n11735, in_21);
	nor (gm_n11737, gm_n48, gm_n53, gm_n52, gm_n3781, in_13);
	nand (gm_n11738, in_16, gm_n63, gm_n50, gm_n11737, gm_n81);
	nor (gm_n11739, gm_n45, gm_n62, gm_n47, gm_n11738, gm_n71);
	nand (gm_n11740, gm_n46, gm_n63, in_14, gm_n9147, gm_n81);
	nor (gm_n11741, in_20, in_19, gm_n47, gm_n11740, in_21);
	nand (gm_n11742, in_15, in_14, gm_n49, gm_n2320, in_16);
	nor (gm_n11743, in_19, gm_n47, in_17, gm_n11742, gm_n45);
	nand (gm_n11744, gm_n11743, gm_n71);
	nand (gm_n11745, gm_n49, gm_n48, gm_n53, gm_n713, gm_n50);
	nor (gm_n11746, in_17, gm_n46, gm_n63, gm_n11745, in_18);
	nand (gm_n11747, gm_n71, gm_n45, gm_n62, gm_n11746);
	nand (gm_n11748, in_13, in_12, in_11, gm_n8071, gm_n50);
	nor (gm_n11749, in_17, gm_n46, in_15, gm_n11748, gm_n47);
	nand (gm_n11750, in_21, gm_n45, gm_n62, gm_n11749);
	nor (gm_n11751, gm_n53, gm_n52, in_9, gm_n4177);
	nand (gm_n11752, in_14, gm_n49, gm_n48, gm_n11751, gm_n63);
	nor (gm_n11753, gm_n47, in_17, gm_n46, gm_n11752, gm_n62);
	nand (gm_n11754, gm_n11753, gm_n71, gm_n45);
	nand (gm_n11755, in_18, gm_n81, gm_n46, gm_n8114, in_19);
	nor (gm_n11756, gm_n11755, in_21, in_20);
	nand (gm_n11757, in_11, in_10, gm_n51, gm_n1274, gm_n48);
	nor (gm_n11758, in_15, gm_n50, in_13, gm_n11757, in_16);
	nand (gm_n11759, gm_n62, in_18, in_17, gm_n11758, in_20);
	nor (gm_n11760, gm_n11759, in_21);
	nand (gm_n11761, gm_n53, gm_n52, in_9, gm_n1856, gm_n48);
	nor (gm_n11762, gm_n63, gm_n50, gm_n49, gm_n11761, in_16);
	nand (gm_n11763, in_19, in_18, gm_n81, gm_n11762, in_20);
	nor (gm_n11764, gm_n11763, in_21);
	nor (gm_n11765, in_13, gm_n48, in_11, gm_n10431, gm_n50);
	nand (gm_n11766, gm_n81, gm_n46, in_15, gm_n11765, gm_n47);
	nor (gm_n11767, gm_n71, in_20, in_19, gm_n11766);
	nor (gm_n11768, gm_n47, in_17, gm_n46, gm_n6687, gm_n62);
	nand (gm_n11769, gm_n11768, in_21, in_20);
	nand (gm_n11770, gm_n48, gm_n53, gm_n52, gm_n311, in_13);
	nor (gm_n11771, gm_n46, in_15, in_14, gm_n11770, in_17);
	nand (gm_n11772, in_20, gm_n62, gm_n47, gm_n11771, in_21);
	and (gm_n11773, in_17, gm_n46, gm_n63, gm_n8878, in_18);
	nand (gm_n11774, gm_n71, gm_n45, in_19, gm_n11773);
	nand (gm_n11775, in_12, in_11, gm_n52, gm_n3239, gm_n49);
	nor (gm_n11776, in_16, in_15, in_14, gm_n11775, in_17);
	nand (gm_n11777, in_20, in_19, gm_n47, gm_n11776, gm_n71);
	nor (gm_n11778, gm_n63, gm_n50, in_13, gm_n9330, in_16);
	nand (gm_n11779, in_19, in_18, gm_n81, gm_n11778, in_20);
	nor (gm_n11780, gm_n11779, in_21);
	and (gm_n11781, gm_n50, gm_n49, in_12, gm_n11377, gm_n63);
	nand (gm_n11782, gm_n47, gm_n81, gm_n46, gm_n11781, in_19);
	nor (gm_n11783, gm_n11782, in_21, in_20);
	nand (gm_n11784, gm_n46, gm_n63, in_14, gm_n3097, gm_n81);
	nor (gm_n11785, in_20, gm_n62, in_18, gm_n11784, in_21);
	nor (gm_n11786, gm_n48, in_11, in_10, gm_n7154, in_13);
	nand (gm_n11787, gm_n46, in_15, gm_n50, gm_n11786, gm_n81);
	nor (gm_n11788, in_20, gm_n62, in_18, gm_n11787, gm_n71);
	nand (gm_n11789, in_12, in_11, gm_n52, gm_n1719, in_13);
	nor (gm_n11790, in_16, in_15, in_14, gm_n11789, gm_n81);
	nand (gm_n11791, in_20, gm_n62, gm_n47, gm_n11790, gm_n71);
	nor (gm_n11792, in_11, gm_n52, gm_n51, gm_n368, in_12);
	nand (gm_n11793, in_15, in_14, gm_n49, gm_n11792, gm_n46);
	nor (gm_n11794, gm_n62, in_18, in_17, gm_n11793, gm_n45);
	nand (gm_n11795, gm_n11794, in_21);
	nand (gm_n11796, gm_n49, in_12, gm_n53, gm_n2947, in_14);
	nor (gm_n11797, gm_n81, gm_n46, gm_n63, gm_n11796, in_18);
	nand (gm_n11798, gm_n71, gm_n45, gm_n62, gm_n11797);
	nor (gm_n11799, gm_n4393, in_9);
	nand (gm_n11800, in_12, gm_n53, gm_n52, gm_n11799, gm_n49);
	nor (gm_n11801, gm_n46, gm_n63, in_14, gm_n11800, in_17);
	nand (gm_n11802, gm_n45, gm_n62, in_18, gm_n11801, in_21);
	and (gm_n11803, in_13, gm_n48, in_11, gm_n6076, in_14);
	and (gm_n11804, in_17, gm_n46, gm_n63, gm_n11803, in_18);
	and (gm_n11805, gm_n71, gm_n45, gm_n62, gm_n11804);
	and (gm_n11806, gm_n48, in_11, in_10, gm_n10774, gm_n49);
	nand (gm_n11807, in_16, in_15, gm_n50, gm_n11806, in_17);
	nor (gm_n11808, gm_n45, in_19, gm_n47, gm_n11807, gm_n71);
	nand (gm_n11809, in_17, gm_n46, gm_n63, gm_n8362, in_18);
	nor (gm_n11810, in_21, gm_n45, gm_n62, gm_n11809);
	nor (gm_n11811, in_12, in_11, in_10, gm_n2052, gm_n49);
	nand (gm_n11812, in_16, gm_n63, gm_n50, gm_n11811, in_17);
	nor (gm_n11813, gm_n45, gm_n62, gm_n47, gm_n11812, gm_n71);
	nand (gm_n11814, in_15, in_14, in_13, gm_n8924, in_16);
	nor (gm_n11815, gm_n62, in_18, gm_n81, gm_n11814, gm_n45);
	nand (gm_n11816, gm_n11815, gm_n71);
	nand (gm_n11817, gm_n49, in_12, in_11, gm_n1053, in_14);
	nor (gm_n11818, gm_n81, in_16, gm_n63, gm_n11817, in_18);
	nand (gm_n11819, gm_n71, gm_n45, in_19, gm_n11818);
	nand (gm_n11820, gm_n50, gm_n49, in_12, gm_n6913, in_15);
	nor (gm_n11821, gm_n47, in_17, gm_n46, gm_n11820, in_19);
	nand (gm_n11822, gm_n11821, in_21, gm_n45);
	nand (gm_n11823, gm_n49, gm_n48, in_11, gm_n11636, in_14);
	nor (gm_n11824, in_17, gm_n46, gm_n63, gm_n11823, gm_n47);
	nand (gm_n11825, in_21, in_20, gm_n62, gm_n11824);
	nand (gm_n11826, gm_n53, in_10, in_9, gm_n548, gm_n48);
	nor (gm_n11827, gm_n63, in_14, gm_n49, gm_n11826, gm_n46);
	nand (gm_n11828, in_19, in_18, in_17, gm_n11827, in_20);
	nor (gm_n11829, gm_n11828, in_21);
	nand (gm_n11830, in_11, in_10, gm_n51, gm_n1192, gm_n48);
	nor (gm_n11831, gm_n11830, in_13);
	nand (gm_n11832, gm_n46, in_15, gm_n50, gm_n11831, gm_n81);
	nor (gm_n11833, gm_n45, gm_n62, in_18, gm_n11832, in_21);
	nor (gm_n11834, in_12, gm_n53, in_10, gm_n9153, gm_n49);
	nand (gm_n11835, in_16, gm_n63, gm_n50, gm_n11834, in_17);
	nor (gm_n11836, gm_n45, in_19, gm_n47, gm_n11835, gm_n71);
	nand (gm_n11837, in_11, in_10, gm_n51, gm_n1116, in_12);
	nor (gm_n11838, gm_n63, gm_n50, in_13, gm_n11837, gm_n46);
	nand (gm_n11839, gm_n62, gm_n47, gm_n81, gm_n11838, gm_n45);
	nor (gm_n11840, gm_n11839, gm_n71);
	or (gm_n11841, gm_n48, in_11, in_10, gm_n1372, gm_n49);
	nor (gm_n11842, gm_n46, in_15, in_14, gm_n11841, in_17);
	nand (gm_n11843, in_20, in_19, in_18, gm_n11842, in_21);
	nand (gm_n11844, gm_n48, in_11, gm_n52, gm_n2681, in_13);
	nor (gm_n11845, in_16, in_15, gm_n50, gm_n11844, gm_n81);
	nand (gm_n11846, in_20, gm_n62, gm_n47, gm_n11845, gm_n71);
	nand (gm_n11847, in_14, gm_n49, in_12, gm_n9945, gm_n63);
	nor (gm_n11848, gm_n47, in_17, gm_n46, gm_n11847, gm_n62);
	nand (gm_n11849, gm_n11848, in_21, gm_n45);
	and (gm_n11850, in_14, in_13, gm_n48, gm_n1924);
	and (gm_n11851, in_17, in_16, in_15, gm_n11850, in_18);
	nand (gm_n11852, in_21, gm_n45, in_19, gm_n11851);
	or (gm_n11853, in_16, gm_n63, gm_n50, gm_n2128, gm_n81);
	nor (gm_n11854, in_20, in_19, in_18, gm_n11853, gm_n71);
	nor (gm_n11855, gm_n48, gm_n53, gm_n52, gm_n4366, gm_n49);
	nand (gm_n11856, in_16, gm_n63, in_14, gm_n11855, in_17);
	nor (gm_n11857, gm_n45, gm_n62, gm_n47, gm_n11856, in_21);
	or (gm_n11858, in_11, gm_n52, in_9, gm_n1709, in_12);
	nor (gm_n11859, gm_n63, gm_n50, gm_n49, gm_n11858, gm_n46);
	nand (gm_n11860, in_19, gm_n47, in_17, gm_n11859, in_20);
	nor (gm_n11861, gm_n11860, in_21);
	nor (gm_n11862, in_12, gm_n53, in_10, gm_n4097, in_13);
	nand (gm_n11863, in_16, in_15, gm_n50, gm_n11862, gm_n81);
	nor (gm_n11864, gm_n45, in_19, in_18, gm_n11863, in_21);
	nand (gm_n11865, in_13, in_12, in_11, gm_n4703, gm_n50);
	nor (gm_n11866, gm_n81, in_16, gm_n63, gm_n11865, in_18);
	nand (gm_n11867, in_21, in_20, in_19, gm_n11866);
	nand (gm_n11868, gm_n49, in_12, in_11, gm_n329, in_14);
	nor (gm_n11869, in_17, gm_n46, in_15, gm_n11868, in_18);
	nand (gm_n11870, gm_n71, gm_n45, gm_n62, gm_n11869);
	nand (gm_n11871, in_12, gm_n53, in_10, gm_n3309, gm_n49);
	nor (gm_n11872, gm_n46, in_15, gm_n50, gm_n11871, gm_n81);
	nand (gm_n11873, gm_n45, in_19, in_18, gm_n11872, gm_n71);
	and (gm_n11874, gm_n64, gm_n55, in_6, gm_n638, in_9);
	nand (gm_n11875, gm_n48, gm_n53, gm_n52, gm_n11874, in_13);
	nor (gm_n11876, gm_n46, gm_n63, gm_n50, gm_n11875, in_17);
	nand (gm_n11877, gm_n45, in_19, in_18, gm_n11876, gm_n71);
	and (gm_n11878, in_15, in_14, gm_n49, gm_n6764, in_16);
	nand (gm_n11879, gm_n62, gm_n47, gm_n81, gm_n11878, in_20);
	nor (gm_n11880, gm_n11879, gm_n71);
	nor (gm_n11881, in_14, gm_n49, gm_n48, gm_n5362, in_15);
	nand (gm_n11882, in_18, in_17, gm_n46, gm_n11881, gm_n62);
	nor (gm_n11883, gm_n11882, in_21, gm_n45);
	or (gm_n11884, gm_n53, in_10, gm_n51, gm_n2419, in_12);
	nor (gm_n11885, in_15, gm_n50, in_13, gm_n11884, in_16);
	nand (gm_n11886, gm_n62, gm_n47, in_17, gm_n11885, in_20);
	nor (gm_n11887, gm_n11886, gm_n71);
	nor (gm_n11888, gm_n50, gm_n49, gm_n48, gm_n3962, in_15);
	nand (gm_n11889, in_18, in_17, gm_n46, gm_n11888, in_19);
	nor (gm_n11890, gm_n11889, in_21, in_20);
	nand (gm_n11891, gm_n48, in_11, gm_n52, gm_n3416, in_13);
	nor (gm_n11892, in_16, in_15, in_14, gm_n11891, in_17);
	nand (gm_n11893, in_20, gm_n62, gm_n47, gm_n11892, gm_n71);
	nand (gm_n11894, gm_n48, in_11, gm_n52, gm_n1671, gm_n49);
	nor (gm_n11895, gm_n46, gm_n63, gm_n50, gm_n11894, in_17);
	nand (gm_n11896, in_20, gm_n62, in_18, gm_n11895, gm_n71);
	nand (gm_n11897, in_13, gm_n48, gm_n53, gm_n1062, gm_n50);
	nor (gm_n11898, gm_n81, gm_n46, gm_n63, gm_n11897, in_18);
	nand (gm_n11899, gm_n71, in_20, in_19, gm_n11898);
	nor (gm_n11900, in_11, gm_n52, gm_n51, gm_n1217, in_12);
	nand (gm_n11901, in_15, gm_n50, gm_n49, gm_n11900, in_16);
	nor (gm_n11902, gm_n62, gm_n47, gm_n81, gm_n11901, in_20);
	nand (gm_n11903, gm_n11902, gm_n71);
	nand (gm_n11904, gm_n51, in_8, gm_n55, gm_n66, gm_n52);
	nor (gm_n11905, in_13, in_12, in_11, gm_n11904, gm_n50);
	nand (gm_n11906, gm_n81, gm_n46, in_15, gm_n11905, in_18);
	nor (gm_n11907, in_21, in_20, in_19, gm_n11906);
	nor (gm_n11908, in_14, in_13, in_12, gm_n7998, in_15);
	nand (gm_n11909, gm_n47, in_17, gm_n46, gm_n11908, gm_n62);
	nor (gm_n11910, gm_n11909, gm_n71, in_20);
	nor (gm_n11911, in_13, gm_n48, gm_n53, gm_n3433, in_14);
	nand (gm_n11912, in_17, gm_n46, in_15, gm_n11911, gm_n47);
	nor (gm_n11913, gm_n71, gm_n45, gm_n62, gm_n11912);
	nand (gm_n11914, in_11, in_10, gm_n51, gm_n1555, gm_n48);
	nor (gm_n11915, gm_n63, gm_n50, in_13, gm_n11914);
	nand (gm_n11916, gm_n47, in_17, gm_n46, gm_n11915, in_19);
	nor (gm_n11917, gm_n11916, in_21, in_20);
	nand (gm_n11918, gm_n63, gm_n50, gm_n49, gm_n7484, gm_n46);
	nor (gm_n11919, gm_n62, in_18, in_17, gm_n11918, gm_n45);
	nand (gm_n11920, gm_n11919, in_21);
	nand (gm_n11921, in_12, in_11, in_10, gm_n3677, in_13);
	nor (gm_n11922, gm_n46, gm_n63, in_14, gm_n11921, in_17);
	nand (gm_n11923, gm_n45, gm_n62, gm_n47, gm_n11922, in_21);
	nor (gm_n11924, in_17, in_16, gm_n63, gm_n11568, gm_n47);
	nand (gm_n11925, gm_n71, in_20, in_19, gm_n11924);
	nor (gm_n11926, gm_n46, in_15, in_14, gm_n10133, in_17);
	nand (gm_n11927, in_20, in_19, gm_n47, gm_n11926, gm_n71);
	nand (gm_n11928, in_11, in_10, gm_n51, gm_n3064, gm_n48);
	nor (gm_n11929, in_15, in_14, in_13, gm_n11928, gm_n46);
	nand (gm_n11930, gm_n62, gm_n47, gm_n81, gm_n11929, in_20);
	nor (gm_n11931, gm_n11930, gm_n71);
	nand (gm_n11932, in_11, gm_n52, in_9, gm_n1643, gm_n48);
	nor (gm_n11933, gm_n63, in_14, in_13, gm_n11932, gm_n46);
	nand (gm_n11934, in_19, in_18, in_17, gm_n11933, in_20);
	nor (gm_n11935, gm_n11934, in_21);
	nand (gm_n11936, gm_n53, in_10, in_9, gm_n2508, gm_n48);
	nor (gm_n11937, gm_n63, in_14, in_13, gm_n11936, in_16);
	nand (gm_n11938, gm_n62, gm_n47, in_17, gm_n11937, gm_n45);
	nor (gm_n11939, gm_n11938, gm_n71);
	nor (gm_n11940, in_13, gm_n48, gm_n53, gm_n10699, in_14);
	nand (gm_n11941, gm_n81, in_16, in_15, gm_n11940, in_18);
	nor (gm_n11942, gm_n71, gm_n45, in_19, gm_n11941);
	or (gm_n11943, in_13, gm_n48, in_11, gm_n1920, in_14);
	nor (gm_n11944, gm_n81, in_16, gm_n63, gm_n11943, gm_n47);
	nand (gm_n11945, gm_n71, in_20, in_19, gm_n11944);
	or (gm_n11946, gm_n48, in_11, in_10, gm_n7068, gm_n49);
	nor (gm_n11947, in_16, gm_n63, in_14, gm_n11946, gm_n81);
	nand (gm_n11948, in_20, gm_n62, in_18, gm_n11947, in_21);
	nand (gm_n11949, gm_n63, in_14, gm_n49, gm_n1639, in_16);
	nor (gm_n11950, in_19, in_18, gm_n81, gm_n11949, in_20);
	nand (gm_n11951, gm_n11950, gm_n71);
	nor (gm_n11952, gm_n53, in_10, in_9, gm_n8122, in_12);
	nand (gm_n11953, gm_n63, gm_n50, in_13, gm_n11952, in_16);
	nor (gm_n11954, gm_n62, in_18, gm_n81, gm_n11953, gm_n45);
	nand (gm_n11955, gm_n11954, gm_n71);
	nand (gm_n11956, gm_n48, in_11, in_10, gm_n8570, gm_n49);
	nor (gm_n11957, gm_n46, gm_n63, gm_n50, gm_n11956, in_17);
	nand (gm_n11958, gm_n45, gm_n62, in_18, gm_n11957, in_21);
	nand (gm_n11959, gm_n11951, gm_n11948, gm_n11945, gm_n11958, gm_n11955);
	nor (gm_n11960, gm_n11939, gm_n11935, gm_n11931, gm_n11959, gm_n11942);
	nand (gm_n11961, gm_n11925, gm_n11923, gm_n11920, gm_n11960, gm_n11927);
	nor (gm_n11962, gm_n11913, gm_n11910, gm_n11907, gm_n11961, gm_n11917);
	nand (gm_n11963, gm_n11899, gm_n11896, gm_n11893, gm_n11962, gm_n11903);
	nor (gm_n11964, gm_n11887, gm_n11883, gm_n11880, gm_n11963, gm_n11890);
	nand (gm_n11965, gm_n11873, gm_n11870, gm_n11867, gm_n11964, gm_n11877);
	nor (gm_n11966, gm_n11861, gm_n11857, gm_n11854, gm_n11965, gm_n11864);
	nand (gm_n11967, gm_n11849, gm_n11846, gm_n11843, gm_n11966, gm_n11852);
	nor (gm_n11968, gm_n11836, gm_n11833, gm_n11829, gm_n11967, gm_n11840);
	nand (gm_n11969, gm_n11822, gm_n11819, gm_n11816, gm_n11968, gm_n11825);
	nor (gm_n11970, gm_n11810, gm_n11808, gm_n11805, gm_n11969, gm_n11813);
	nand (gm_n11971, gm_n11798, gm_n11795, gm_n11791, gm_n11970, gm_n11802);
	nor (gm_n11972, gm_n11785, gm_n11783, gm_n11780, gm_n11971, gm_n11788);
	nand (gm_n11973, gm_n11774, gm_n11772, gm_n11769, gm_n11972, gm_n11777);
	nor (gm_n11974, gm_n11764, gm_n11760, gm_n11756, gm_n11973, gm_n11767);
	nand (gm_n11975, gm_n11750, gm_n11747, gm_n11744, gm_n11974, gm_n11754);
	nor (gm_n11976, gm_n11739, gm_n11736, gm_n11732, gm_n11975, gm_n11741);
	nand (gm_n11977, gm_n11726, gm_n11723, gm_n11720, gm_n11976, gm_n11729);
	nor (gm_n11978, gm_n11714, gm_n11711, gm_n11708, gm_n11977, gm_n11717);
	nand (gm_n11979, gm_n11702, gm_n11700, gm_n11696, gm_n11978, gm_n11705);
	nor (gm_n11980, gm_n11689, gm_n11686, gm_n11683, gm_n11979, gm_n11692);
	nand (gm_n11981, gm_n11677, gm_n11675, gm_n11672, gm_n11980, gm_n11681);
	nor (gm_n11982, gm_n11665, gm_n11662, gm_n11660, gm_n11981, gm_n11669);
	nand (gm_n11983, gm_n11656, gm_n11652, gm_n11649, gm_n11982, gm_n11659);
	nor (gm_n11984, gm_n11642, gm_n11639, gm_n11635, gm_n11983, gm_n11645);
	nand (gm_n11985, gm_n11630, gm_n11627, gm_n11624, gm_n11984, gm_n11633);
	nor (gm_n11986, gm_n11619, gm_n11616, gm_n11613, gm_n11985, gm_n11622);
	nand (gm_n11987, gm_n11607, gm_n11604, gm_n11601, gm_n11986, gm_n11610);
	nor (gm_n11988, gm_n11594, gm_n11592, gm_n11589, gm_n11987, gm_n11597);
	nand (gm_n11989, gm_n11582, gm_n11579, gm_n11576, gm_n11988, gm_n11586);
	nor (gm_n11990, gm_n11570, gm_n11566, gm_n11563, gm_n11989, gm_n11573);
	nand (gm_n11991, gm_n11558, gm_n11555, gm_n11552, gm_n11990, gm_n11561);
	nor (gm_n11992, gm_n11545, gm_n11541, gm_n11539, gm_n11991, gm_n11548);
	nand (gm_n11993, gm_n11533, gm_n11531, gm_n11528, gm_n11992, gm_n11536);
	nor (gm_n11994, gm_n11522, gm_n11520, gm_n11516, gm_n11993, gm_n11525);
	nand (gm_n11995, gm_n11510, gm_n11508, gm_n11505, gm_n11994, gm_n11513);
	nor (out_20, gm_n11995, gm_n11504);
	and (gm_n11997, gm_n48, in_11, in_10, gm_n8194, in_13);
	nand (gm_n11998, in_16, in_15, in_14, gm_n11997, in_17);
	nor (gm_n11999, gm_n45, in_19, gm_n47, gm_n11998, gm_n71);
	nand (gm_n12000, in_16, in_15, gm_n50, gm_n6339, gm_n81);
	nor (gm_n12001, gm_n45, in_19, in_18, gm_n12000, gm_n71);
	or (gm_n12002, in_8, gm_n55, gm_n82, gm_n156, in_9);
	nor (gm_n12003, in_12, in_11, in_10, gm_n12002, gm_n49);
	nand (gm_n12004, gm_n46, gm_n63, in_14, gm_n12003, gm_n81);
	nor (gm_n12005, gm_n45, gm_n62, gm_n47, gm_n12004, gm_n71);
	nand (gm_n12006, in_13, in_12, in_11, gm_n3226, in_14);
	nor (gm_n12007, in_17, gm_n46, in_15, gm_n12006, in_18);
	nand (gm_n12008, in_21, gm_n45, gm_n62, gm_n12007);
	or (gm_n12009, gm_n49, in_12, gm_n53, gm_n7319, gm_n50);
	nor (gm_n12010, gm_n81, gm_n46, in_15, gm_n12009, in_18);
	nand (gm_n12011, in_21, in_20, in_19, gm_n12010);
	nand (gm_n12012, gm_n50, in_13, gm_n48, gm_n3524, in_15);
	nor (gm_n12013, in_18, in_17, in_16, gm_n12012, in_19);
	nand (gm_n12014, gm_n12013, in_21, gm_n45);
	nand (gm_n12015, in_14, in_13, in_12, gm_n5392, in_15);
	nor (gm_n12016, gm_n47, in_17, gm_n46, gm_n12015, in_19);
	nand (gm_n12017, gm_n12016, gm_n71, gm_n45);
	nor (gm_n12018, in_15, gm_n50, in_13, gm_n11370, gm_n46);
	nand (gm_n12019, in_19, in_18, in_17, gm_n12018, gm_n45);
	nor (gm_n12020, gm_n12019, in_21);
	nor (gm_n12021, in_12, in_11, gm_n52, gm_n4809, gm_n49);
	nand (gm_n12022, gm_n46, gm_n63, gm_n50, gm_n12021, in_17);
	nor (gm_n12023, gm_n45, gm_n62, in_18, gm_n12022, in_21);
	and (gm_n12024, in_12, gm_n53, gm_n52, gm_n11450, gm_n49);
	nand (gm_n12025, gm_n46, in_15, in_14, gm_n12024, gm_n81);
	nor (gm_n12026, in_20, gm_n62, gm_n47, gm_n12025, gm_n71);
	and (gm_n12027, gm_n50, gm_n49, gm_n48, gm_n7746, gm_n63);
	nand (gm_n12028, gm_n47, in_17, in_16, gm_n12027, in_19);
	nor (gm_n12029, gm_n12028, gm_n71, in_20);
	nor (gm_n12030, in_11, gm_n52, gm_n51, gm_n3340, gm_n48);
	nand (gm_n12031, in_15, in_14, in_13, gm_n12030, in_16);
	nor (gm_n12032, in_19, gm_n47, gm_n81, gm_n12031, in_20);
	nand (gm_n12033, gm_n12032, in_21);
	or (gm_n12034, gm_n48, gm_n53, gm_n52, gm_n4554, gm_n49);
	nor (gm_n12035, gm_n46, in_15, gm_n50, gm_n12034, gm_n81);
	nand (gm_n12036, gm_n45, gm_n62, in_18, gm_n12035, in_21);
	and (gm_n12037, in_11, in_10, gm_n51, gm_n792, gm_n48);
	nand (gm_n12038, gm_n63, in_14, in_13, gm_n12037, gm_n46);
	nor (gm_n12039, in_19, in_18, gm_n81, gm_n12038, gm_n45);
	nand (gm_n12040, gm_n12039, gm_n71);
	nand (gm_n12041, in_13, gm_n48, in_11, gm_n7510, in_14);
	nor (gm_n12042, in_17, in_16, in_15, gm_n12041, in_18);
	nand (gm_n12043, gm_n71, in_20, in_19, gm_n12042);
	and (gm_n12044, gm_n63, gm_n50, gm_n49, gm_n12037, gm_n46);
	nand (gm_n12045, in_19, in_18, in_17, gm_n12044, gm_n45);
	nor (gm_n12046, gm_n12045, gm_n71);
	nand (gm_n12047, gm_n53, in_10, in_9, gm_n3043, gm_n48);
	nor (gm_n12048, in_15, in_14, in_13, gm_n12047, gm_n46);
	nand (gm_n12049, in_19, in_18, gm_n81, gm_n12048, gm_n45);
	nor (gm_n12050, gm_n12049, gm_n71);
	or (gm_n12051, gm_n53, in_10, in_9, gm_n2926, in_12);
	nor (gm_n12052, in_15, in_14, in_13, gm_n12051, gm_n46);
	nand (gm_n12053, in_19, gm_n47, gm_n81, gm_n12052, gm_n45);
	nor (gm_n12054, gm_n12053, in_21);
	nor (gm_n12055, gm_n48, gm_n53, gm_n52, gm_n9867, gm_n49);
	nand (gm_n12056, gm_n46, in_15, in_14, gm_n12055, gm_n81);
	nor (gm_n12057, in_20, in_19, in_18, gm_n12056, gm_n71);
	nor (gm_n12058, in_11, gm_n52, in_9, gm_n368, gm_n48);
	nand (gm_n12059, gm_n63, in_14, gm_n49, gm_n12058, gm_n46);
	nor (gm_n12060, in_19, in_18, in_17, gm_n12059, gm_n45);
	nand (gm_n12061, gm_n12060, gm_n71);
	nand (gm_n12062, in_13, in_12, gm_n53, gm_n4043, gm_n50);
	nor (gm_n12063, in_17, gm_n46, gm_n63, gm_n12062, gm_n47);
	nand (gm_n12064, gm_n71, in_20, in_19, gm_n12063);
	nor (gm_n12065, gm_n51, in_8, gm_n55, gm_n843, in_10);
	nand (gm_n12066, in_13, in_12, in_11, gm_n12065, gm_n50);
	nor (gm_n12067, in_17, in_16, in_15, gm_n12066, in_18);
	nand (gm_n12068, in_21, gm_n45, gm_n62, gm_n12067);
	nand (gm_n12069, in_14, gm_n49, in_12, gm_n1987, gm_n63);
	nor (gm_n12070, gm_n47, gm_n81, in_16, gm_n12069, gm_n62);
	nand (gm_n12071, gm_n12070, in_21, in_20);
	and (gm_n12072, gm_n63, gm_n50, in_13, gm_n9030, gm_n46);
	nand (gm_n12073, gm_n62, in_18, gm_n81, gm_n12072, gm_n45);
	nor (gm_n12074, gm_n12073, in_21);
	nor (gm_n12075, in_14, gm_n49, in_12, gm_n650, gm_n63);
	nand (gm_n12076, in_18, in_17, gm_n46, gm_n12075, gm_n62);
	nor (gm_n12077, gm_n12076, gm_n71, gm_n45);
	nor (gm_n12078, in_14, in_13, in_12, gm_n1071, gm_n63);
	nand (gm_n12079, gm_n47, in_17, gm_n46, gm_n12078, gm_n62);
	nor (gm_n12080, gm_n12079, gm_n71, gm_n45);
	nand (gm_n12081, in_11, in_10, gm_n51, gm_n673, in_12);
	nor (gm_n12082, gm_n63, gm_n50, gm_n49, gm_n12081, gm_n46);
	nand (gm_n12083, in_19, gm_n47, in_17, gm_n12082, gm_n45);
	nor (gm_n12084, gm_n12083, gm_n71);
	nand (gm_n12085, gm_n48, in_11, in_10, gm_n1406, gm_n49);
	nor (gm_n12086, gm_n46, gm_n63, gm_n50, gm_n12085, in_17);
	nand (gm_n12087, gm_n45, gm_n62, in_18, gm_n12086, in_21);
	and (gm_n12088, in_18, in_17, gm_n46, gm_n3342, in_19);
	nand (gm_n12089, gm_n12088, gm_n71, in_20);
	nand (gm_n12090, gm_n50, gm_n49, in_12, gm_n1740, in_15);
	nor (gm_n12091, gm_n47, gm_n81, in_16, gm_n12090, gm_n62);
	nand (gm_n12092, gm_n12091, in_21, in_20);
	nand (gm_n12093, gm_n49, gm_n48, gm_n53, gm_n11636, in_14);
	nor (gm_n12094, gm_n81, in_16, in_15, gm_n12093, gm_n47);
	nand (gm_n12095, gm_n71, in_20, in_19, gm_n12094);
	nand (gm_n12096, in_11, gm_n52, gm_n51, gm_n2181, gm_n48);
	nor (gm_n12097, gm_n63, gm_n50, gm_n49, gm_n12096, gm_n46);
	nand (gm_n12098, in_19, gm_n47, in_17, gm_n12097, in_20);
	nor (gm_n12099, gm_n12098, gm_n71);
	nand (gm_n12100, gm_n53, in_10, gm_n51, gm_n3606, in_12);
	nor (gm_n12101, gm_n63, gm_n50, gm_n49, gm_n12100, gm_n46);
	nand (gm_n12102, gm_n62, in_18, gm_n81, gm_n12101, gm_n45);
	nor (gm_n12103, gm_n12102, in_21);
	and (gm_n12104, in_15, gm_n50, gm_n49, gm_n211, gm_n46);
	nand (gm_n12105, gm_n62, gm_n47, in_17, gm_n12104, gm_n45);
	nor (gm_n12106, gm_n12105, gm_n71);
	and (gm_n12107, in_12, gm_n53, in_10, gm_n7305, gm_n49);
	nand (gm_n12108, in_16, gm_n63, in_14, gm_n12107, in_17);
	nor (gm_n12109, in_20, gm_n62, gm_n47, gm_n12108, in_21);
	nand (gm_n12110, in_13, in_12, in_11, gm_n5358, gm_n50);
	nor (gm_n12111, in_17, in_16, gm_n63, gm_n12110, in_18);
	nand (gm_n12112, in_21, in_20, gm_n62, gm_n12111);
	nand (gm_n12113, in_12, gm_n53, in_10, gm_n6342, in_13);
	nor (gm_n12114, in_16, in_15, in_14, gm_n12113, in_17);
	nand (gm_n12115, gm_n45, in_19, gm_n47, gm_n12114, in_21);
	nand (gm_n12116, gm_n48, in_11, in_10, gm_n11192, gm_n49);
	nor (gm_n12117, in_16, in_15, gm_n50, gm_n12116, gm_n81);
	nand (gm_n12118, in_20, in_19, gm_n47, gm_n12117, gm_n71);
	nor (gm_n12119, gm_n53, gm_n52, in_9, gm_n2005, gm_n48);
	nand (gm_n12120, gm_n63, in_14, in_13, gm_n12119, in_16);
	nor (gm_n12121, in_19, gm_n47, gm_n81, gm_n12120, gm_n45);
	nand (gm_n12122, gm_n12121, gm_n71);
	nor (gm_n12123, in_13, in_12, in_11, gm_n2389, gm_n50);
	nand (gm_n12124, gm_n81, gm_n46, gm_n63, gm_n12123, gm_n47);
	nor (gm_n12125, gm_n71, in_20, in_19, gm_n12124);
	nor (gm_n12126, in_12, gm_n53, in_10, gm_n1174, gm_n49);
	nand (gm_n12127, gm_n46, gm_n63, in_14, gm_n12126, in_17);
	nor (gm_n12128, gm_n45, in_19, in_18, gm_n12127, in_21);
	nand (gm_n12129, in_16, gm_n63, in_14, gm_n10010, in_17);
	nor (gm_n12130, gm_n45, gm_n62, gm_n47, gm_n12129, in_21);
	nor (gm_n12131, gm_n48, gm_n53, gm_n52, gm_n9086, in_13);
	nand (gm_n12132, gm_n46, in_15, gm_n50, gm_n12131, gm_n81);
	nor (gm_n12133, in_20, gm_n62, gm_n47, gm_n12132, gm_n71);
	nor (gm_n12134, in_11, gm_n52, in_9, gm_n3557, gm_n48);
	nand (gm_n12135, in_15, in_14, in_13, gm_n12134, gm_n46);
	nor (gm_n12136, in_19, in_18, in_17, gm_n12135, gm_n45);
	nand (gm_n12137, gm_n12136, gm_n71);
	nand (gm_n12138, in_21, gm_n45, in_19, gm_n11804);
	nand (gm_n12139, gm_n48, in_11, gm_n52, gm_n142, gm_n49);
	nor (gm_n12140, in_16, in_15, gm_n50, gm_n12139, gm_n81);
	nand (gm_n12141, gm_n45, gm_n62, in_18, gm_n12140, in_21);
	and (gm_n12142, gm_n46, gm_n63, in_14, gm_n11831, in_17);
	nand (gm_n12143, gm_n45, in_19, gm_n47, gm_n12142, in_21);
	nor (gm_n12144, in_14, in_13, gm_n48, gm_n9838, gm_n63);
	nand (gm_n12145, in_18, in_17, gm_n46, gm_n12144, gm_n62);
	nor (gm_n12146, gm_n12145, in_21, in_20);
	nor (gm_n12147, gm_n71, in_20, gm_n62, gm_n10440);
	and (gm_n12148, in_12, gm_n53, gm_n52, gm_n4418, in_13);
	nand (gm_n12149, in_16, gm_n63, gm_n50, gm_n12148, in_17);
	nor (gm_n12150, in_20, gm_n62, gm_n47, gm_n12149, gm_n71);
	and (gm_n12151, in_12, gm_n53, gm_n52, gm_n4266, in_13);
	nand (gm_n12152, gm_n46, gm_n63, gm_n50, gm_n12151, gm_n81);
	nor (gm_n12153, in_20, gm_n62, gm_n47, gm_n12152, gm_n71);
	nand (gm_n12154, gm_n48, in_11, in_10, gm_n1413, in_13);
	nor (gm_n12155, in_16, gm_n63, in_14, gm_n12154, in_17);
	nand (gm_n12156, in_20, in_19, gm_n47, gm_n12155, gm_n71);
	nand (gm_n12157, in_13, in_12, gm_n53, gm_n10386, gm_n50);
	nor (gm_n12158, in_17, in_16, gm_n63, gm_n12157, gm_n47);
	nand (gm_n12159, in_21, in_20, gm_n62, gm_n12158);
	nand (gm_n12160, in_15, in_14, in_13, gm_n5010, gm_n46);
	nor (gm_n12161, gm_n62, in_18, gm_n81, gm_n12160, gm_n45);
	nand (gm_n12162, gm_n12161, gm_n71);
	nor (gm_n12163, gm_n53, in_10, gm_n51, gm_n8122, gm_n48);
	nand (gm_n12164, in_15, gm_n50, in_13, gm_n12163, gm_n46);
	nor (gm_n12165, gm_n62, in_18, gm_n81, gm_n12164, in_20);
	nand (gm_n12166, gm_n12165, in_21);
	nor (gm_n12167, in_12, in_11, in_10, gm_n5322, gm_n49);
	nand (gm_n12168, in_16, gm_n63, in_14, gm_n12167, in_17);
	nor (gm_n12169, gm_n45, gm_n62, gm_n47, gm_n12168, gm_n71);
	nor (gm_n12170, in_12, gm_n53, in_10, gm_n3683, in_13);
	nand (gm_n12171, in_16, gm_n63, gm_n50, gm_n12170, gm_n81);
	nor (gm_n12172, in_20, in_19, in_18, gm_n12171, in_21);
	nand (gm_n12173, in_9, in_8, in_7, gm_n66, gm_n52);
	nor (gm_n12174, in_13, in_12, gm_n53, gm_n12173, gm_n50);
	nand (gm_n12175, gm_n81, gm_n46, in_15, gm_n12174, in_18);
	nor (gm_n12176, in_21, in_20, in_19, gm_n12175);
	nor (gm_n12177, gm_n49, in_12, gm_n53, gm_n2575, in_14);
	nand (gm_n12178, gm_n81, gm_n46, gm_n63, gm_n12177, gm_n47);
	nor (gm_n12179, gm_n71, gm_n45, in_19, gm_n12178);
	nor (gm_n12180, gm_n46, in_15, gm_n50, gm_n9803, gm_n81);
	nand (gm_n12181, in_20, gm_n62, in_18, gm_n12180, in_21);
	nand (gm_n12182, in_13, in_12, in_11, gm_n11517, in_14);
	nor (gm_n12183, gm_n81, gm_n46, gm_n63, gm_n12182, gm_n47);
	nand (gm_n12184, gm_n71, gm_n45, gm_n62, gm_n12183);
	nand (gm_n12185, gm_n48, in_11, gm_n52, gm_n6883, gm_n49);
	nor (gm_n12186, gm_n46, in_15, in_14, gm_n12185, gm_n81);
	nand (gm_n12187, in_20, gm_n62, in_18, gm_n12186, gm_n71);
	nand (gm_n12188, gm_n1215, gm_n71, gm_n45);
	and (gm_n12189, gm_n63, in_14, gm_n49, gm_n11646, in_16);
	nand (gm_n12190, gm_n62, gm_n47, gm_n81, gm_n12189, in_20);
	nor (gm_n12191, gm_n12190, gm_n71);
	and (gm_n12192, in_12, gm_n53, in_10, gm_n11799, gm_n49);
	nand (gm_n12193, gm_n46, gm_n63, gm_n50, gm_n12192, in_17);
	nor (gm_n12194, gm_n45, in_19, in_18, gm_n12193, gm_n71);
	nor (gm_n12195, in_12, gm_n53, gm_n52, gm_n7154, in_13);
	nand (gm_n12196, gm_n46, in_15, gm_n50, gm_n12195, gm_n81);
	nor (gm_n12197, gm_n45, gm_n62, in_18, gm_n12196, gm_n71);
	nor (gm_n12198, in_15, gm_n50, in_13, gm_n9647, in_16);
	nand (gm_n12199, gm_n62, gm_n47, gm_n81, gm_n12198, gm_n45);
	nor (gm_n12200, gm_n12199, gm_n71);
	nand (gm_n12201, in_13, gm_n48, in_11, gm_n7250, in_14);
	nor (gm_n12202, in_17, in_16, in_15, gm_n12201, in_18);
	nand (gm_n12203, in_21, gm_n45, in_19, gm_n12202);
	nand (gm_n12204, in_12, in_11, in_10, gm_n3069, gm_n49);
	nor (gm_n12205, in_16, gm_n63, gm_n50, gm_n12204, gm_n81);
	nand (gm_n12206, gm_n45, gm_n62, gm_n47, gm_n12205, in_21);
	and (gm_n12207, gm_n46, in_15, gm_n50, gm_n8991, in_17);
	nand (gm_n12208, in_20, in_19, gm_n47, gm_n12207, in_21);
	and (gm_n12209, gm_n46, in_15, gm_n50, gm_n1913, in_17);
	nand (gm_n12210, gm_n45, in_19, gm_n47, gm_n12209, in_21);
	and (gm_n12211, gm_n48, gm_n53, in_10, gm_n3723, in_13);
	nand (gm_n12212, in_16, in_15, in_14, gm_n12211, in_17);
	nor (gm_n12213, gm_n45, gm_n62, in_18, gm_n12212, in_21);
	and (gm_n12214, in_14, in_13, gm_n48, gm_n286, gm_n63);
	nand (gm_n12215, gm_n47, gm_n81, in_16, gm_n12214, gm_n62);
	nor (gm_n12216, gm_n12215, in_21, in_20);
	nand (gm_n12217, in_16, gm_n63, in_14, gm_n215, in_17);
	nor (gm_n12218, in_20, gm_n62, gm_n47, gm_n12217, gm_n71);
	and (gm_n12219, in_12, in_11, gm_n52, gm_n2641, in_13);
	nand (gm_n12220, gm_n46, gm_n63, gm_n50, gm_n12219, in_17);
	nor (gm_n12221, gm_n45, gm_n62, in_18, gm_n12220, in_21);
	or (gm_n12222, gm_n48, gm_n53, gm_n52, gm_n347, gm_n49);
	nor (gm_n12223, in_16, gm_n63, gm_n50, gm_n12222, gm_n81);
	nand (gm_n12224, gm_n45, gm_n62, in_18, gm_n12223, gm_n71);
	and (gm_n12225, in_11, gm_n52, gm_n51, gm_n2601, in_12);
	nand (gm_n12226, in_15, gm_n50, in_13, gm_n12225, in_16);
	nor (gm_n12227, in_19, gm_n47, gm_n81, gm_n12226, in_20);
	nand (gm_n12228, gm_n12227, in_21);
	nand (gm_n12229, gm_n48, gm_n53, in_10, gm_n200, in_13);
	nor (gm_n12230, gm_n46, in_15, gm_n50, gm_n12229, gm_n81);
	nand (gm_n12231, gm_n45, in_19, gm_n47, gm_n12230, gm_n71);
	and (gm_n12232, in_11, gm_n52, gm_n51, gm_n644, gm_n48);
	nand (gm_n12233, in_15, gm_n50, in_13, gm_n12232, gm_n46);
	nor (gm_n12234, gm_n62, gm_n47, gm_n81, gm_n12233, in_20);
	nand (gm_n12235, gm_n12234, gm_n71);
	nor (gm_n12236, in_12, in_11, gm_n52, gm_n730, in_13);
	nand (gm_n12237, in_16, in_15, in_14, gm_n12236, in_17);
	nor (gm_n12238, in_20, in_19, gm_n47, gm_n12237, in_21);
	and (gm_n12239, gm_n63, in_14, in_13, gm_n3813, in_16);
	nand (gm_n12240, in_19, gm_n47, in_17, gm_n12239, gm_n45);
	nor (gm_n12241, gm_n12240, gm_n71);
	nand (gm_n12242, in_11, gm_n52, gm_n51, gm_n1279, gm_n48);
	nor (gm_n12243, gm_n63, gm_n50, gm_n49, gm_n12242, in_16);
	nand (gm_n12244, in_19, in_18, gm_n81, gm_n12243, gm_n45);
	nor (gm_n12245, gm_n12244, in_21);
	nand (gm_n12246, in_17, gm_n46, gm_n63, gm_n1589, in_18);
	nor (gm_n12247, gm_n71, gm_n45, gm_n62, gm_n12246);
	and (gm_n12248, in_10, in_9, gm_n64, gm_n838, in_11);
	nand (gm_n12249, gm_n50, gm_n49, in_12, gm_n12248, in_15);
	nor (gm_n12250, gm_n47, in_17, gm_n46, gm_n12249, in_19);
	nand (gm_n12251, gm_n12250, gm_n71, gm_n45);
	and (gm_n12252, in_16, in_15, in_14, gm_n1118, in_17);
	nand (gm_n12253, in_20, in_19, gm_n47, gm_n12252, gm_n71);
	nand (gm_n12254, in_13, gm_n48, gm_n53, gm_n5591, gm_n50);
	nor (gm_n12255, gm_n81, in_16, in_15, gm_n12254, gm_n47);
	nand (gm_n12256, gm_n71, gm_n45, gm_n62, gm_n12255);
	nand (gm_n12257, gm_n49, in_12, gm_n53, gm_n416, in_14);
	nor (gm_n12258, in_17, in_16, in_15, gm_n12257, gm_n47);
	nand (gm_n12259, in_21, gm_n45, gm_n62, gm_n12258);
	and (gm_n12260, gm_n50, in_13, in_12, gm_n11751, in_15);
	nand (gm_n12261, in_18, in_17, in_16, gm_n12260, gm_n62);
	nor (gm_n12262, gm_n12261, in_21, in_20);
	nand (gm_n12263, gm_n53, gm_n52, in_9, gm_n1986, in_12);
	nor (gm_n12264, in_15, gm_n50, in_13, gm_n12263, gm_n46);
	nand (gm_n12265, gm_n62, in_18, in_17, gm_n12264, gm_n45);
	nor (gm_n12266, gm_n12265, gm_n71);
	nor (gm_n12267, in_12, gm_n53, gm_n52, gm_n6518, in_13);
	nand (gm_n12268, gm_n46, gm_n63, gm_n50, gm_n12267, in_17);
	nor (gm_n12269, gm_n45, in_19, in_18, gm_n12268, in_21);
	nor (gm_n12270, in_13, in_12, in_11, gm_n7520, gm_n50);
	nand (gm_n12271, in_17, in_16, in_15, gm_n12270, in_18);
	nor (gm_n12272, in_21, gm_n45, in_19, gm_n12271);
	or (gm_n12273, in_20, gm_n62, gm_n47, gm_n6959, gm_n71);
	or (gm_n12274, in_12, in_11, in_10, gm_n3924, in_13);
	nor (gm_n12275, gm_n46, gm_n63, in_14, gm_n12274, gm_n81);
	nand (gm_n12276, in_20, gm_n62, in_18, gm_n12275, gm_n71);
	nand (gm_n12277, in_13, gm_n48, in_11, gm_n8809, gm_n50);
	nor (gm_n12278, gm_n81, in_16, in_15, gm_n12277, in_18);
	nand (gm_n12279, in_21, in_20, gm_n62, gm_n12278);
	nand (gm_n12280, in_20, in_19, in_18, gm_n6248, in_21);
	and (gm_n12281, gm_n48, in_11, gm_n52, gm_n380, in_13);
	nand (gm_n12282, in_16, in_15, in_14, gm_n12281, gm_n81);
	nor (gm_n12283, in_20, gm_n62, in_18, gm_n12282, gm_n71);
	and (gm_n12284, gm_n50, gm_n49, gm_n48, gm_n6236, in_15);
	nand (gm_n12285, in_18, gm_n81, in_16, gm_n12284, gm_n62);
	nor (gm_n12286, gm_n12285, in_21, gm_n45);
	and (gm_n12287, in_13, in_12, in_11, gm_n4907, gm_n50);
	nand (gm_n12288, gm_n81, gm_n46, gm_n63, gm_n12287, gm_n47);
	nor (gm_n12289, gm_n71, in_20, in_19, gm_n12288);
	and (gm_n12290, in_14, in_13, gm_n48, gm_n6156, gm_n63);
	nand (gm_n12291, gm_n47, gm_n81, in_16, gm_n12290, gm_n62);
	nor (gm_n12292, gm_n12291, gm_n71, gm_n45);
	and (gm_n12293, gm_n52, in_9, in_8, gm_n1088, in_11);
	nand (gm_n12294, gm_n50, gm_n49, gm_n48, gm_n12293, in_15);
	nor (gm_n12295, in_18, gm_n81, gm_n46, gm_n12294, in_19);
	nand (gm_n12296, gm_n12295, gm_n71, gm_n45);
	nand (gm_n12297, in_12, in_11, gm_n52, gm_n1307, gm_n49);
	nor (gm_n12298, gm_n46, gm_n63, in_14, gm_n12297, gm_n81);
	nand (gm_n12299, gm_n45, in_19, gm_n47, gm_n12298, gm_n71);
	nand (gm_n12300, in_14, in_13, in_12, gm_n5772, in_15);
	nor (gm_n12301, in_18, gm_n81, in_16, gm_n12300, in_19);
	nand (gm_n12302, gm_n12301, in_21, gm_n45);
	nand (gm_n12303, in_12, gm_n53, gm_n52, gm_n400, in_13);
	nor (gm_n12304, gm_n46, gm_n63, in_14, gm_n12303, gm_n81);
	nand (gm_n12305, gm_n45, in_19, gm_n47, gm_n12304, in_21);
	nand (gm_n12306, gm_n46, in_15, gm_n50, gm_n4753, in_17);
	nor (gm_n12307, gm_n45, in_19, in_18, gm_n12306, in_21);
	or (gm_n12308, gm_n51, gm_n64, in_7, gm_n84, in_10);
	nor (gm_n12309, in_13, gm_n48, in_11, gm_n12308, gm_n50);
	nand (gm_n12310, gm_n81, gm_n46, in_15, gm_n12309, in_18);
	nor (gm_n12311, gm_n71, in_20, gm_n62, gm_n12310);
	and (gm_n12312, gm_n50, in_13, gm_n48, gm_n11200, in_15);
	nand (gm_n12313, gm_n47, gm_n81, in_16, gm_n12312, gm_n62);
	nor (gm_n12314, gm_n12313, in_21, gm_n45);
	and (gm_n12315, in_13, in_12, in_11, gm_n5644, in_14);
	nand (gm_n12316, in_17, in_16, gm_n63, gm_n12315, in_18);
	nor (gm_n12317, gm_n71, gm_n45, gm_n62, gm_n12316);
	nand (gm_n12318, gm_n48, gm_n53, in_10, gm_n2877, in_13);
	nor (gm_n12319, gm_n46, in_15, in_14, gm_n12318, gm_n81);
	nand (gm_n12320, in_20, gm_n62, gm_n47, gm_n12319, in_21);
	or (gm_n12321, in_12, gm_n53, in_10, gm_n6056, gm_n49);
	nor (gm_n12322, gm_n46, in_15, gm_n50, gm_n12321, in_17);
	nand (gm_n12323, gm_n45, gm_n62, gm_n47, gm_n12322, in_21);
	nand (gm_n12324, in_13, gm_n48, gm_n53, gm_n1036, in_14);
	nor (gm_n12325, in_17, gm_n46, gm_n63, gm_n12324, gm_n47);
	nand (gm_n12326, gm_n71, in_20, gm_n62, gm_n12325);
	and (gm_n12327, gm_n47, in_17, in_16, gm_n11915, gm_n62);
	nand (gm_n12328, gm_n12327, gm_n71, in_20);
	or (gm_n12329, gm_n46, gm_n63, in_14, gm_n9427, in_17);
	nor (gm_n12330, gm_n45, gm_n62, in_18, gm_n12329, gm_n71);
	nand (gm_n12331, gm_n81, in_16, in_15, gm_n2590, in_18);
	nor (gm_n12332, in_21, gm_n45, in_19, gm_n12331);
	and (gm_n12333, in_15, in_14, gm_n49, gm_n3817, gm_n46);
	nand (gm_n12334, gm_n62, gm_n47, in_17, gm_n12333, gm_n45);
	nor (gm_n12335, gm_n12334, in_21);
	nor (gm_n12336, in_12, gm_n53, in_10, gm_n9609, gm_n49);
	nand (gm_n12337, in_16, in_15, in_14, gm_n12336, in_17);
	nor (gm_n12338, in_20, gm_n62, in_18, gm_n12337, gm_n71);
	nand (gm_n12339, gm_n48, in_11, in_10, gm_n3909, in_13);
	nor (gm_n12340, gm_n46, gm_n63, gm_n50, gm_n12339, gm_n81);
	nand (gm_n12341, gm_n45, in_19, in_18, gm_n12340, gm_n71);
	or (gm_n12342, in_13, gm_n48, in_11, gm_n464, in_14);
	nor (gm_n12343, gm_n81, gm_n46, in_15, gm_n12342, gm_n47);
	nand (gm_n12344, gm_n71, in_20, in_19, gm_n12343);
	and (gm_n12345, in_16, gm_n63, in_14, gm_n7187, gm_n81);
	nand (gm_n12346, in_20, gm_n62, gm_n47, gm_n12345, in_21);
	or (gm_n12347, gm_n48, gm_n53, gm_n52, gm_n1452, in_13);
	nor (gm_n12348, gm_n46, gm_n63, gm_n50, gm_n12347, gm_n81);
	nand (gm_n12349, gm_n45, gm_n62, in_18, gm_n12348, gm_n71);
	nor (gm_n12350, in_12, gm_n53, gm_n52, gm_n3159, in_13);
	nand (gm_n12351, gm_n46, in_15, in_14, gm_n12350, gm_n81);
	nor (gm_n12352, gm_n45, gm_n62, gm_n47, gm_n12351, gm_n71);
	nor (gm_n12353, gm_n48, gm_n53, in_10, gm_n6760, gm_n49);
	nand (gm_n12354, gm_n46, in_15, in_14, gm_n12353, gm_n81);
	nor (gm_n12355, gm_n45, gm_n62, in_18, gm_n12354, in_21);
	nor (gm_n12356, gm_n48, gm_n53, in_10, gm_n2845, gm_n49);
	nand (gm_n12357, in_16, gm_n63, gm_n50, gm_n12356, gm_n81);
	nor (gm_n12358, gm_n45, in_19, in_18, gm_n12357, in_21);
	nand (gm_n12359, in_17, gm_n46, gm_n63, gm_n11850, gm_n47);
	nor (gm_n12360, in_21, gm_n45, gm_n62, gm_n12359);
	nor (gm_n12361, in_11, gm_n52, in_9, gm_n3475, in_12);
	nand (gm_n12362, in_15, gm_n50, gm_n49, gm_n12361, gm_n46);
	nor (gm_n12363, gm_n62, gm_n47, in_17, gm_n12362, in_20);
	nand (gm_n12364, gm_n12363, gm_n71);
	and (gm_n12365, in_16, gm_n63, gm_n50, gm_n10821, gm_n81);
	nand (gm_n12366, gm_n45, in_19, gm_n47, gm_n12365, gm_n71);
	nand (gm_n12367, gm_n50, gm_n49, gm_n48, gm_n956, in_15);
	nor (gm_n12368, in_18, in_17, gm_n46, gm_n12367, gm_n62);
	nand (gm_n12369, gm_n12368, gm_n71, gm_n45);
	nand (gm_n12370, in_12, gm_n53, in_10, gm_n2956, in_13);
	nor (gm_n12371, in_16, gm_n63, gm_n50, gm_n12370, in_17);
	nand (gm_n12372, in_20, gm_n62, in_18, gm_n12371, in_21);
	and (gm_n12373, in_15, gm_n50, in_13, gm_n2210, in_16);
	nand (gm_n12374, in_19, in_18, in_17, gm_n12373, gm_n45);
	nor (gm_n12375, gm_n12374, gm_n71);
	nor (gm_n12376, in_15, gm_n50, gm_n49, gm_n9393, gm_n46);
	nand (gm_n12377, in_19, gm_n47, in_17, gm_n12376, in_20);
	nor (gm_n12378, gm_n12377, in_21);
	or (gm_n12379, in_9, gm_n64, gm_n55, gm_n843, in_10);
	nor (gm_n12380, in_13, in_12, gm_n53, gm_n12379, gm_n50);
	nand (gm_n12381, in_17, gm_n46, gm_n63, gm_n12380, gm_n47);
	nor (gm_n12382, gm_n71, in_20, in_19, gm_n12381);
	nor (gm_n12383, gm_n48, gm_n53, in_10, gm_n6897, gm_n49);
	nand (gm_n12384, gm_n46, gm_n63, gm_n50, gm_n12383, in_17);
	nor (gm_n12385, gm_n45, in_19, gm_n47, gm_n12384, in_21);
	nor (gm_n12386, gm_n53, gm_n52, in_9, gm_n333, gm_n48);
	nand (gm_n12387, gm_n63, gm_n50, in_13, gm_n12386, gm_n46);
	nor (gm_n12388, gm_n62, in_18, in_17, gm_n12387, gm_n45);
	nand (gm_n12389, gm_n12388, gm_n71);
	nand (gm_n12390, in_14, in_13, gm_n48, gm_n6550, in_15);
	nor (gm_n12391, gm_n47, gm_n81, gm_n46, gm_n12390, gm_n62);
	nand (gm_n12392, gm_n12391, in_21, gm_n45);
	nand (gm_n12393, in_14, gm_n49, in_12, gm_n10355, in_15);
	nor (gm_n12394, gm_n47, gm_n81, in_16, gm_n12393, in_19);
	nand (gm_n12395, gm_n12394, in_21, in_20);
	nand (gm_n12396, gm_n48, gm_n53, in_10, gm_n3731, gm_n49);
	nor (gm_n12397, in_16, gm_n63, gm_n50, gm_n12396, in_17);
	nand (gm_n12398, gm_n45, gm_n62, gm_n47, gm_n12397, gm_n71);
	and (gm_n12399, in_12, gm_n53, in_10, gm_n1365, in_13);
	nand (gm_n12400, in_16, gm_n63, in_14, gm_n12399, in_17);
	nor (gm_n12401, gm_n45, gm_n62, in_18, gm_n12400, in_21);
	nand (gm_n12402, gm_n64, gm_n55, in_6, gm_n374, in_9);
	nor (gm_n12403, in_12, gm_n53, gm_n52, gm_n12402, gm_n49);
	nand (gm_n12404, gm_n46, gm_n63, gm_n50, gm_n12403, gm_n81);
	nor (gm_n12405, in_20, in_19, in_18, gm_n12404, gm_n71);
	nor (gm_n12406, gm_n48, in_11, gm_n52, gm_n3012, gm_n49);
	nand (gm_n12407, gm_n46, gm_n63, gm_n50, gm_n12406, gm_n81);
	nor (gm_n12408, in_20, gm_n62, in_18, gm_n12407, gm_n71);
	nor (gm_n12409, gm_n50, gm_n49, gm_n48, gm_n8095, gm_n63);
	nand (gm_n12410, gm_n47, gm_n81, in_16, gm_n12409, gm_n62);
	nor (gm_n12411, gm_n12410, gm_n71, gm_n45);
	or (gm_n12412, gm_n45, in_19, in_18, gm_n4754, gm_n71);
	nand (gm_n12413, gm_n48, in_11, gm_n52, gm_n2984, in_13);
	nor (gm_n12414, in_16, gm_n63, in_14, gm_n12413, in_17);
	nand (gm_n12415, in_20, gm_n62, gm_n47, gm_n12414, gm_n71);
	nand (gm_n12416, gm_n48, gm_n53, in_10, gm_n205, gm_n49);
	nor (gm_n12417, in_16, in_15, gm_n50, gm_n12416, gm_n81);
	nand (gm_n12418, gm_n45, gm_n62, in_18, gm_n12417, gm_n71);
	nand (gm_n12419, in_12, in_11, gm_n52, gm_n9518, gm_n49);
	nor (gm_n12420, gm_n46, in_15, gm_n50, gm_n12419, in_17);
	nand (gm_n12421, gm_n45, in_19, in_18, gm_n12420, in_21);
	nor (gm_n12422, gm_n63, gm_n50, gm_n49, gm_n4501, gm_n46);
	nand (gm_n12423, gm_n62, gm_n47, gm_n81, gm_n12422, gm_n45);
	nor (gm_n12424, gm_n12423, gm_n71);
	nor (gm_n12425, in_15, in_14, gm_n49, gm_n2027, in_16);
	nand (gm_n12426, in_19, in_18, gm_n81, gm_n12425, gm_n45);
	nor (gm_n12427, gm_n12426, gm_n71);
	nor (gm_n12428, in_13, in_12, in_11, gm_n989, gm_n50);
	nand (gm_n12429, gm_n81, gm_n46, gm_n63, gm_n12428, in_18);
	nor (gm_n12430, in_21, in_20, gm_n62, gm_n12429);
	nor (gm_n12431, gm_n63, gm_n50, gm_n49, gm_n3607, gm_n46);
	nand (gm_n12432, in_19, gm_n47, in_17, gm_n12431, in_20);
	nor (gm_n12433, gm_n12432, in_21);
	nor (gm_n12434, gm_n52, in_9, gm_n64, gm_n4079, gm_n53);
	nand (gm_n12435, in_14, gm_n49, in_12, gm_n12434, in_15);
	nor (gm_n12436, in_18, in_17, gm_n46, gm_n12435, in_19);
	nand (gm_n12437, gm_n12436, in_21, in_20);
	and (gm_n12438, in_8, gm_n55, gm_n82, gm_n379, gm_n51);
	nand (gm_n12439, in_12, gm_n53, in_10, gm_n12438, gm_n49);
	nor (gm_n12440, gm_n46, gm_n63, gm_n50, gm_n12439, in_17);
	nand (gm_n12441, in_20, in_19, in_18, gm_n12440, in_21);
	nand (gm_n12442, in_13, gm_n48, in_11, gm_n9541, in_14);
	nor (gm_n12443, gm_n81, in_16, gm_n63, gm_n12442, gm_n47);
	nand (gm_n12444, gm_n71, gm_n45, gm_n62, gm_n12443);
	nand (gm_n12445, gm_n12444, gm_n12441, gm_n12437);
	nor (gm_n12446, gm_n12430, gm_n12427, gm_n12424, gm_n12445, gm_n12433);
	nand (gm_n12447, gm_n12418, gm_n12415, gm_n12412, gm_n12446, gm_n12421);
	nor (gm_n12448, gm_n12408, gm_n12405, gm_n12401, gm_n12447, gm_n12411);
	nand (gm_n12449, gm_n12395, gm_n12392, gm_n12389, gm_n12448, gm_n12398);
	nor (gm_n12450, gm_n12382, gm_n12378, gm_n12375, gm_n12449, gm_n12385);
	nand (gm_n12451, gm_n12369, gm_n12366, gm_n12364, gm_n12450, gm_n12372);
	nor (gm_n12452, gm_n12358, gm_n12355, gm_n12352, gm_n12451, gm_n12360);
	nand (gm_n12453, gm_n12346, gm_n12344, gm_n12341, gm_n12452, gm_n12349);
	nor (gm_n12454, gm_n12335, gm_n12332, gm_n12330, gm_n12453, gm_n12338);
	nand (gm_n12455, gm_n12326, gm_n12323, gm_n12320, gm_n12454, gm_n12328);
	nor (gm_n12456, gm_n12314, gm_n12311, gm_n12307, gm_n12455, gm_n12317);
	nand (gm_n12457, gm_n12302, gm_n12299, gm_n12296, gm_n12456, gm_n12305);
	nor (gm_n12458, gm_n12289, gm_n12286, gm_n12283, gm_n12457, gm_n12292);
	nand (gm_n12459, gm_n12279, gm_n12276, gm_n12273, gm_n12458, gm_n12280);
	nor (gm_n12460, gm_n12269, gm_n12266, gm_n12262, gm_n12459, gm_n12272);
	nand (gm_n12461, gm_n12256, gm_n12253, gm_n12251, gm_n12460, gm_n12259);
	nor (gm_n12462, gm_n12245, gm_n12241, gm_n12238, gm_n12461, gm_n12247);
	nand (gm_n12463, gm_n12231, gm_n12228, gm_n12224, gm_n12462, gm_n12235);
	nor (gm_n12464, gm_n12218, gm_n12216, gm_n12213, gm_n12463, gm_n12221);
	nand (gm_n12465, gm_n12208, gm_n12206, gm_n12203, gm_n12464, gm_n12210);
	nor (gm_n12466, gm_n12197, gm_n12194, gm_n12191, gm_n12465, gm_n12200);
	nand (gm_n12467, gm_n12187, gm_n12184, gm_n12181, gm_n12466, gm_n12188);
	nor (gm_n12468, gm_n12176, gm_n12172, gm_n12169, gm_n12467, gm_n12179);
	nand (gm_n12469, gm_n12162, gm_n12159, gm_n12156, gm_n12468, gm_n12166);
	nor (gm_n12470, gm_n12150, gm_n12147, gm_n12146, gm_n12469, gm_n12153);
	nand (gm_n12471, gm_n12141, gm_n12138, gm_n12137, gm_n12470, gm_n12143);
	nor (gm_n12472, gm_n12130, gm_n12128, gm_n12125, gm_n12471, gm_n12133);
	nand (gm_n12473, gm_n12118, gm_n12115, gm_n12112, gm_n12472, gm_n12122);
	nor (gm_n12474, gm_n12106, gm_n12103, gm_n12099, gm_n12473, gm_n12109);
	nand (gm_n12475, gm_n12092, gm_n12089, gm_n12087, gm_n12474, gm_n12095);
	nor (gm_n12476, gm_n12080, gm_n12077, gm_n12074, gm_n12475, gm_n12084);
	nand (gm_n12477, gm_n12068, gm_n12064, gm_n12061, gm_n12476, gm_n12071);
	nor (gm_n12478, gm_n12054, gm_n12050, gm_n12046, gm_n12477, gm_n12057);
	nand (gm_n12479, gm_n12040, gm_n12036, gm_n12033, gm_n12478, gm_n12043);
	nor (gm_n12480, gm_n12026, gm_n12023, gm_n12020, gm_n12479, gm_n12029);
	nand (gm_n12481, gm_n12014, gm_n12011, gm_n12008, gm_n12480, gm_n12017);
	nor (out_21, gm_n12005, gm_n12001, gm_n11999, gm_n12481);
endmodule
