module top ( g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 , g98 , g99 , g100 , g101 , g102 , g103 , g104 , g105 , g106 , g107 , g108 , g109 , g110 , g111 , g112 , g113 , g114 , g115 , g116 , g117 , g118 , g119 , g120 , g121 , g122 , g123 , g124 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g136 , g137 , g138 , g139 , g140 , g141 , g142 , g143 , g144 , g145 , g146 , g147 , g148 , g149 , g150 , g151 , g152 , g153 , g154 , g155 , g156 , g157 , g158 , g159 , g160 , g161 , g162 , g163 , g164 , g165 , g166 , g167 , g168 , g169 , g170 , g171 , g172 , g173 , g174 , g175 , g176 , g177 , g178 , g179 , g180 , g181 , g182 , g183 , g184 , g185 , g186 , g187 , g188 , g189 , g190 , g191 , g192 , g193 , g194 , g195 , g196 , g197 , g198 , g199 , g200 , g201 , g202 , g203 , g204 , g205 , g206 , g207 , g208 , g209 , g210 , g211 , g212 , g213 , g214 , g215 , g216 , g217 , g218 , g219 , g220 , g221 , g222 , g223 , g224 , g225 , g226 );
input g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 , g98 ;
output g99 , g100 , g101 , g102 , g103 , g104 , g105 , g106 , g107 , g108 , g109 , g110 , g111 , g112 , g113 , g114 , g115 , g116 , g117 , g118 , g119 , g120 , g121 , g122 , g123 , g124 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g136 , g137 , g138 , g139 , g140 , g141 , g142 , g143 , g144 , g145 , g146 , g147 , g148 , g149 , g150 , g151 , g152 , g153 , g154 , g155 , g156 , g157 , g158 , g159 , g160 , g161 , g162 , g163 , g164 , g165 , g166 , g167 , g168 , g169 , g170 , g171 , g172 , g173 , g174 , g175 , g176 , g177 , g178 , g179 , g180 , g181 , g182 , g183 , g184 , g185 , g186 , g187 , g188 , g189 , g190 , g191 , g192 , g193 , g194 , g195 , g196 , g197 , g198 , g199 , g200 , g201 , g202 , g203 , g204 , g205 , g206 , g207 , g208 , g209 , g210 , g211 , g212 , g213 , g214 , g215 , g216 , g217 , g218 , g219 , g220 , g221 , g222 , g223 , g224 , g225 , g226 ;

wire n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , 
     n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , 
     n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , 
     n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , 
     n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , 
     n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , 
     n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , 
     n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , 
     n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , 
     n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , 
     n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , 
     n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , 
     n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , 
     n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , 
     n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , 
     n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , 
     n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , 
     n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , 
     n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , 
     n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , 
     n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , 
     n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , 
     n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , 
     n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , 
     n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , 
     n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , 
     n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , 
     n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , 
     n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , 
     n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , 
     n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , 
     n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , 
     n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , 
     n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , 
     n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , 
     n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , 
     n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , 
     n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , 
     n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , 
     n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , 
     n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , 
     n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , 
     n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , 
     n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , 
     n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , 
     n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , 
     n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , 
     n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , 
     n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , 
     n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , 
     n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , 
     n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , 
     n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , 
     n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , 
     n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , 
     n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , 
     n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , 
     n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , 
     n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , 
     n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , 
     n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , 
     n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , 
     n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , 
     n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , 
     n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , 
     n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , 
     n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , 
     n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , 
     n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , 
     n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , 
     n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , 
     n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , 
     n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , 
     n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , 
     n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , 
     n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , 
     n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , 
     n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , 
     n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , 
     n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , 
     n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , 
     n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , 
     n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , 
     n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , 
     n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , 
     n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , 
     n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , 
     n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , 
     n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , 
     n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , 
     n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , 
     n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , 
     n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , 
     n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , 
     n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , 
     n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , 
     n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , 
     n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , 
     n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , 
     n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , 
     n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , 
     n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , 
     n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , 
     n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , 
     n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , 
     n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , 
     n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , 
     n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , 
     n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , 
     n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , 
     n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , 
     n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , 
     n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , 
     n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , 
     n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , 
     n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , 
     n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , 
     n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , 
     n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , 
     n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , 
     n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , 
     n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , 
     n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , 
     n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , 
     n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , 
     n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , 
     n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , 
     n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , 
     n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , 
     n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , 
     n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , 
     n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , 
     n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , 
     n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , 
     n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , 
     n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , 
     n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , 
     n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , 
     n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , 
     n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , 
     n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , 
     n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , 
     n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , 
     n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , 
     n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , 
     n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , 
     n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , 
     n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , 
     n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , 
     n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , 
     n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , 
     n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , 
     n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , 
     n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , 
     n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , 
     n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , 
     n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , 
     n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , 
     n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , 
     n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , 
     n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , 
     n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , 
     n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , 
     n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , 
     n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , 
     n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , 
     n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , 
     n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , 
     n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , 
     n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , 
     n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , 
     n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , 
     n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , 
     n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , 
     n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , 
     n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , 
     n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , 
     n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , 
     n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , 
     n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , 
     n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , 
     n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , 
     n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , 
     n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , 
     n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , 
     n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , 
     n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , 
     n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , 
     n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , 
     n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , 
     n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , 
     n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , 
     n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , 
     n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , 
     n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , 
     n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , 
     n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , 
     n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , 
     n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , 
     n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , 
     n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , 
     n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , 
     n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , 
     n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , 
     n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , 
     n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , 
     n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , 
     n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , 
     n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , 
     n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , 
     n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , 
     n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , 
     n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , 
     n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , 
     n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , 
     n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , 
     n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , 
     n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , 
     n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , 
     n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , 
     n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , 
     n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , 
     n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , 
     n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , 
     n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , 
     n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , 
     n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , 
     n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , 
     n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , 
     n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , 
     n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , 
     n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , 
     n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , 
     n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , 
     n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , 
     n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , 
     n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , 
     n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , 
     n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , 
     n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , 
     n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , 
     n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , 
     n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , 
     n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , 
     n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , 
     n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , 
     n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , 
     n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , 
     n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , 
     n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , 
     n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , 
     n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , 
     n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , 
     n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , 
     n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , 
     n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , 
     n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , 
     n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , 
     n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , 
     n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , 
     n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , 
     n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , 
     n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , 
     n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , 
     n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , 
     n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , 
     n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , 
     n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , 
     n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , 
     n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , 
     n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , 
     n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , 
     n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , 
     n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , 
     n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , 
     n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , 
     n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , 
     n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , 
     n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , 
     n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , 
     n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , 
     n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , 
     n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , 
     n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , 
     n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , 
     n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , 
     n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , 
     n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , 
     n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , 
     n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , 
     n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , 
     n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , 
     n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , 
     n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , 
     n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , 
     n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , 
     n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , 
     n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , 
     n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , 
     n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , 
     n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , 
     n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , 
     n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , 
     n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , 
     n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , 
     n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , 
     n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , 
     n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , 
     n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , 
     n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , 
     n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , 
     n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , 
     n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , 
     n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , 
     n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , 
     n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , 
     n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , 
     n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , 
     n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , 
     n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , 
     n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , 
     n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , 
     n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , 
     n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , 
     n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , 
     n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , 
     n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , 
     n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , 
     n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , 
     n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , 
     n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , 
     n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , 
     n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , 
     n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , 
     n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , 
     n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , 
     n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , 
     n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , 
     n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , 
     n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , 
     n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , 
     n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , 
     n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , 
     n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , 
     n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , 
     n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , 
     n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , 
     n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , 
     n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , 
     n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , 
     n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , 
     n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , 
     n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , 
     n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , 
     n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , 
     n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , 
     n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , 
     n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , 
     n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , 
     n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , 
     n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , 
     n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , 
     n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , 
     n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , 
     n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , 
     n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , 
     n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , 
     n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , 
     n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , 
     n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , 
     n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , 
     n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , 
     n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , 
     n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , 
     n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , 
     n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , 
     n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , 
     n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , 
     n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , 
     n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , 
     n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , 
     n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , 
     n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , 
     n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , 
     n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , 
     n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , 
     n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , 
     n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , 
     n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , 
     n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , 
     n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , 
     n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , 
     n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , 
     n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , 
     n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , 
     n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , 
     n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , 
     n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , 
     n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , 
     n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , 
     n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , 
     n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , 
     n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , 
     n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , 
     n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , 
     n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , 
     n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , 
     n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , 
     n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , 
     n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , 
     n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , 
     n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , 
     n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , 
     n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , 
     n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , 
     n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , 
     n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , 
     n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , 
     n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , 
     n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , 
     n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , 
     n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , 
     n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , 
     n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , 
     n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , 
     n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , 
     n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , 
     n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , 
     n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , 
     n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , 
     n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , 
     n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , 
     n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , 
     n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , 
     n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , 
     n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , 
     n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , 
     n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , 
     n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , 
     n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , 
     n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , 
     n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , 
     n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , 
     n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , 
     n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , 
     n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , 
     n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , 
     n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , 
     n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , 
     n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , 
     n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , 
     n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , 
     n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , 
     n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , 
     n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , 
     n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , 
     n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , 
     n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , 
     n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , 
     n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , 
     n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , 
     n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , 
     n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , 
     n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , 
     n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , 
     n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , 
     n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , 
     n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , 
     n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , 
     n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , 
     n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , 
     n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , 
     n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , 
     n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , 
     n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , 
     n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , 
     n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , 
     n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , 
     n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , 
     n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , 
     n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , 
     n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , 
     n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , 
     n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , 
     n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , 
     n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , 
     n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , 
     n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , 
     n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , 
     n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , 
     n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , 
     n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , 
     n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , 
     n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , 
     n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , 
     n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , 
     n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , 
     n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , 
     n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , 
     n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , 
     n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , 
     n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , 
     n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , 
     n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , 
     n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , 
     n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , 
     n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , 
     n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , 
     n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , 
     n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , 
     n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , 
     n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , 
     n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , 
     n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , 
     n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , 
     n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , 
     n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , 
     n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , 
     n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , 
     n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , 
     n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , 
     n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , 
     n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , 
     n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , 
     n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , 
     n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , 
     n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , 
     n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , 
     n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , 
     n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , 
     n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , 
     n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , 
     n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , 
     n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , 
     n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , 
     n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , 
     n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , 
     n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , 
     n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , 
     n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , 
     n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , 
     n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , 
     n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , 
     n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , 
     n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , 
     n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , 
     n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , 
     n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , 
     n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , 
     n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , 
     n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , 
     n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , 
     n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , 
     n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , 
     n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , 
     n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , 
     n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , 
     n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , 
     n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , 
     n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , 
     n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , 
     n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , 
     n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , 
     n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , 
     n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , 
     n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , 
     n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , 
     n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , 
     n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , 
     n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , 
     n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , 
     n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , 
     n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , 
     n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , 
     n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , 
     n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , 
     n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , 
     n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , 
     n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , 
     n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , 
     n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , 
     n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , 
     n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , 
     n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , 
     n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , 
     n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , 
     n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , 
     n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , 
     n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , 
     n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , 
     n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , 
     n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , 
     n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , 
     n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , 
     n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , 
     n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , 
     n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , 
     n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , 
     n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , 
     n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , 
     n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , 
     n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , 
     n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , 
     n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , 
     n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , 
     n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , 
     n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , 
     n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , 
     n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , 
     n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , 
     n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , 
     n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , 
     n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , 
     n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , 
     n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , 
     n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , 
     n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , 
     n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , 
     n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , 
     n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , 
     n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , 
     n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , 
     n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , 
     n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , 
     n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , 
     n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , 
     n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , 
     n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , 
     n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , 
     n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , 
     n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , 
     n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , 
     n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , 
     n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , 
     n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , 
     n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , 
     n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , 
     n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , 
     n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , 
     n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , 
     n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , 
     n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , 
     n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , 
     n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , 
     n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , 
     n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , 
     n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , 
     n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , 
     n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , 
     n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , 
     n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , 
     n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , 
     n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , 
     n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , 
     n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , 
     n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , 
     n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , 
     n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , 
     n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , 
     n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , 
     n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , 
     n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , 
     n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , 
     n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , 
     n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , 
     n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , 
     n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , 
     n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , 
     n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , 
     n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , 
     n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , 
     n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , 
     n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , 
     n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , 
     n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , 
     n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , 
     n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , 
     n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , 
     n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , 
     n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , 
     n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , 
     n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , 
     n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , 
     n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , 
     n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , 
     n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , 
     n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , 
     n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , 
     n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , 
     n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , 
     n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , 
     n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , 
     n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , 
     n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , 
     n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , 
     n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , 
     n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , 
     n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , 
     n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , 
     n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , 
     n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , 
     n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , 
     n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , 
     n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , 
     n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , 
     n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , 
     n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , 
     n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , 
     n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , 
     n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , 
     n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , 
     n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , 
     n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , 
     n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , 
     n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , 
     n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , 
     n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , 
     n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , 
     n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , 
     n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , 
     n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , 
     n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , 
     n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , 
     n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , 
     n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , 
     n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , 
     n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , 
     n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , 
     n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , 
     n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , 
     n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , 
     n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , 
     n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , 
     n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , 
     n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , 
     n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , 
     n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , 
     n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , 
     n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , 
     n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , 
     n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , 
     n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , 
     n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , 
     n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , 
     n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , 
     n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , 
     n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , 
     n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , 
     n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , 
     n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , 
     n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , 
     n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , 
     n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , 
     n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , 
     n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , 
     n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , 
     n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , 
     n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , 
     n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , 
     n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , 
     n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , 
     n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , 
     n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , 
     n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , 
     n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , 
     n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , 
     n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , 
     n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , 
     n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , 
     n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , 
     n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , 
     n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , 
     n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , 
     n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , 
     n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , 
     n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , 
     n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , 
     n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , 
     n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , 
     n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , 
     n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , 
     n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , 
     n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , 
     n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , 
     n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , 
     n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , 
     n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , 
     n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , 
     n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , 
     n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , 
     n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , 
     n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , 
     n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , 
     n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , 
     n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , 
     n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , 
     n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , 
     n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , 
     n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , 
     n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , 
     n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , 
     n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , 
     n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , 
     n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , 
     n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , 
     n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , 
     n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , 
     n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , 
     n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , 
     n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , 
     n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , 
     n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , 
     n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , 
     n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , 
     n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , 
     n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , 
     n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , 
     n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , 
     n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , 
     n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , 
     n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , 
     n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , 
     n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , 
     n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , 
     n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , 
     n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , 
     n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , 
     n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , 
     n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , 
     n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , 
     n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , 
     n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , 
     n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , 
     n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , 
     n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , 
     n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , 
     n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , 
     n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , 
     n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , 
     n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , 
     n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , 
     n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , 
     n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , 
     n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , 
     n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , 
     n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , 
     n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , 
     n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , 
     n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , 
     n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , 
     n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , 
     n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , 
     n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , 
     n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , 
     n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , 
     n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , 
     n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , 
     n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , 
     n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , 
     n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , 
     n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , 
     n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , 
     n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , 
     n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , 
     n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , 
     n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , 
     n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , 
     n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , 
     n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , 
     n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , 
     n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , 
     n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , 
     n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , 
     n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , 
     n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , 
     n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , 
     n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , 
     n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , 
     n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , 
     n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , 
     n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , 
     n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , 
     n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , 
     n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , 
     n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , 
     n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , 
     n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , 
     n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , 
     n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , 
     n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , 
     n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , 
     n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , 
     n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , 
     n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , 
     n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , 
     n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , 
     n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , 
     n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , 
     n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , 
     n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , 
     n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , 
     n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , 
     n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , 
     n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , 
     n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , 
     n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , 
     n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , 
     n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , 
     n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , 
     n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , 
     n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , 
     n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , 
     n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , 
     n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , 
     n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , 
     n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , 
     n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , 
     n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , 
     n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , 
     n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , 
     n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , 
     n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , 
     n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , 
     n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , 
     n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , 
     n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , 
     n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , 
     n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , 
     n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , 
     n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , 
     n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , 
     n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , 
     n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , 
     n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , 
     n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , 
     n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , 
     n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , 
     n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , 
     n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , 
     n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , 
     n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , 
     n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , 
     n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , 
     n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , 
     n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , 
     n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , 
     n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , 
     n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , 
     n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , 
     n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , 
     n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , 
     n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , 
     n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , 
     n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , 
     n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , 
     n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , 
     n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , 
     n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , 
     n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , 
     n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , 
     n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , 
     n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , 
     n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , 
     n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , 
     n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , 
     n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , 
     n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , 
     n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , 
     n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , 
     n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , 
     n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , 
     n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , 
     n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , 
     n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , 
     n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , 
     n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , 
     n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , 
     n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , 
     n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , 
     n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , 
     n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , 
     n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , 
     n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , 
     n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , 
     n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , 
     n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , 
     n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , 
     n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , 
     n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , 
     n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , 
     n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , 
     n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , 
     n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , 
     n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , 
     n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , 
     n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , 
     n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , 
     n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , 
     n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , 
     n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , 
     n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , 
     n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , 
     n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , 
     n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , 
     n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , 
     n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , 
     n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , 
     n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , 
     n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , 
     n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , 
     n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , 
     n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , 
     n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , 
     n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , 
     n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , 
     n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , 
     n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , 
     n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , 
     n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , 
     n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , 
     n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , 
     n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , 
     n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , 
     n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , 
     n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , 
     n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , 
     n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , 
     n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , 
     n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , 
     n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , 
     n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , 
     n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , 
     n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , 
     n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , 
     n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , 
     n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , 
     n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , 
     n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , 
     n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , 
     n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , 
     n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , 
     n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , 
     n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , 
     n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , 
     n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , 
     n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , 
     n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , 
     n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , 
     n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , 
     n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , 
     n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , 
     n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , 
     n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , 
     n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , 
     n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , 
     n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , 
     n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , 
     n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , 
     n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , 
     n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , 
     n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , 
     n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , 
     n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , 
     n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , 
     n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , 
     n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , 
     n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , 
     n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , 
     n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , 
     n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , 
     n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , 
     n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , 
     n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , 
     n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , 
     n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , 
     n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , 
     n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , 
     n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , 
     n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , 
     n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , 
     n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , 
     n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , 
     n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , 
     n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , 
     n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , 
     n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , 
     n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , 
     n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , 
     n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , 
     n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , 
     n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , 
     n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , 
     n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , 
     n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , 
     n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , 
     n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , 
     n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , 
     n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , 
     n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , 
     n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , 
     n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , 
     n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , 
     n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , 
     n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , 
     n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , 
     n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , 
     n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , 
     n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , 
     n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , 
     n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , 
     n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , 
     n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , 
     n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , 
     n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , 
     n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , 
     n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , 
     n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , 
     n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , 
     n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , 
     n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , 
     n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , 
     n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , 
     n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , 
     n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , 
     n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , 
     n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , 
     n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , 
     n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , 
     n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , 
     n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , 
     n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , 
     n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , 
     n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , 
     n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , 
     n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , 
     n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , 
     n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , 
     n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , 
     n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , 
     n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , 
     n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , 
     n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , 
     n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , 
     n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , 
     n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , 
     n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , 
     n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , 
     n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , 
     n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , 
     n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , 
     n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , 
     n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , 
     n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , 
     n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , 
     n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , 
     n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , 
     n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , 
     n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , 
     n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , 
     n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , 
     n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , 
     n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , 
     n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , 
     n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , 
     n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , 
     n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , 
     n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , 
     n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , 
     n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , 
     n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , 
     n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , 
     n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , 
     n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , 
     n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , 
     n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , 
     n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , 
     n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , 
     n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , 
     n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , 
     n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , 
     n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , 
     n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , 
     n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , 
     n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , 
     n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , 
     n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , 
     n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , 
     n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , 
     n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , 
     n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , 
     n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , 
     n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , 
     n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , 
     n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , 
     n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , 
     n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , 
     n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , 
     n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , 
     n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , 
     n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , 
     n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , 
     n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , 
     n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , 
     n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , 
     n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , 
     n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , 
     n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , 
     n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , 
     n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , 
     n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , 
     n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , 
     n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , 
     n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , 
     n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , 
     n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , 
     n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , 
     n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , 
     n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , 
     n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , 
     n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , 
     n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , 
     n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , 
     n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , 
     n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , 
     n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , 
     n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , 
     n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , 
     n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , 
     n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , 
     n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , 
     n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , 
     n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , 
     n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , 
     n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , 
     n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , 
     n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , 
     n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , 
     n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , 
     n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , 
     n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , 
     n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , 
     n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , 
     n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , 
     n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , 
     n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , 
     n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , 
     n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , 
     n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , 
     n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , 
     n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , 
     n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , 
     n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , 
     n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , 
     n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , 
     n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , 
     n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , 
     n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , 
     n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , 
     n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , 
     n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , 
     n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , 
     n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , 
     n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , 
     n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , 
     n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , 
     n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , 
     n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , 
     n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , 
     n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , 
     n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , 
     n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , 
     n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , 
     n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , 
     n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , 
     n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , 
     n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , 
     n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , 
     n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , 
     n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , 
     n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , 
     n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , 
     n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , 
     n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , 
     n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , 
     n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , 
     n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , 
     n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , 
     n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , 
     n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , 
     n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , 
     n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , 
     n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , 
     n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , 
     n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , 
     n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , 
     n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , 
     n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , 
     n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , 
     n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , 
     n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , 
     n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , 
     n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , 
     n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , 
     n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , 
     n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , 
     n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , 
     n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , 
     n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , 
     n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , 
     n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , 
     n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , 
     n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , 
     n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , 
     n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , 
     n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , 
     n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , 
     n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , 
     n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , 
     n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , 
     n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , 
     n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , 
     n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , 
     n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , 
     n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , 
     n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , 
     n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , 
     n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , 
     n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , 
     n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , 
     n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , 
     n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , 
     n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , 
     n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , 
     n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , 
     n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , 
     n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , 
     n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , 
     n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , 
     n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , 
     n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , 
     n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , 
     n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , 
     n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , 
     n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , 
     n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , 
     n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , 
     n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , 
     n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , 
     n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , 
     n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , 
     n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , 
     n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , 
     n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , 
     n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , 
     n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , 
     n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , 
     n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , 
     n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , 
     n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , 
     n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , 
     n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , 
     n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , 
     n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , 
     n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , 
     n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , 
     n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , 
     n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , 
     n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , 
     n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , 
     n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , 
     n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 ;
wire t_0 , t_1 ;
buf ( n1 , g0 );
buf ( n2 , g1 );
buf ( n3 , g2 );
buf ( n4 , g3 );
buf ( n5 , g4 );
buf ( n6 , g5 );
buf ( n7 , g6 );
buf ( n8 , g7 );
buf ( n9 , g8 );
buf ( n10 , g9 );
buf ( n11 , g10 );
buf ( n12 , g11 );
buf ( n13 , g12 );
buf ( n14 , g13 );
buf ( n15 , g14 );
buf ( n16 , g15 );
buf ( n17 , g16 );
buf ( n18 , g17 );
buf ( n19 , g18 );
buf ( n20 , g19 );
buf ( n21 , g20 );
buf ( n22 , g21 );
buf ( n23 , g22 );
buf ( n24 , g23 );
buf ( n25 , g24 );
buf ( n26 , g25 );
buf ( n27 , g26 );
buf ( n28 , g27 );
buf ( n29 , g28 );
buf ( n30 , g29 );
buf ( n31 , g30 );
buf ( n32 , g31 );
buf ( n33 , g32 );
buf ( n34 , g33 );
buf ( n35 , g34 );
buf ( n36 , g35 );
buf ( n37 , g36 );
buf ( n38 , g37 );
buf ( n39 , g38 );
buf ( n40 , g39 );
buf ( n41 , g40 );
buf ( n42 , g41 );
buf ( n43 , g42 );
buf ( n44 , g43 );
buf ( n45 , g44 );
buf ( n46 , g45 );
buf ( n47 , g46 );
buf ( n48 , g47 );
buf ( n49 , g48 );
buf ( n50 , g49 );
buf ( n51 , g50 );
buf ( n52 , g51 );
buf ( n53 , g52 );
buf ( n54 , g53 );
buf ( n55 , g54 );
buf ( n56 , g55 );
buf ( n57 , g56 );
buf ( n58 , g57 );
buf ( n59 , g58 );
buf ( n60 , g59 );
buf ( n61 , g60 );
buf ( n62 , g61 );
buf ( n63 , g62 );
buf ( n64 , g63 );
buf ( n65 , g64 );
buf ( n66 , g65 );
buf ( n67 , g66 );
buf ( n68 , g67 );
buf ( n69 , g68 );
buf ( n70 , g69 );
buf ( n71 , g70 );
buf ( n72 , g71 );
buf ( n73 , g72 );
buf ( n74 , g73 );
buf ( n75 , g74 );
buf ( n76 , g75 );
buf ( n77 , g76 );
buf ( n78 , g77 );
buf ( n79 , g78 );
buf ( n80 , g79 );
buf ( n81 , g80 );
buf ( n82 , g81 );
buf ( n83 , g82 );
buf ( n84 , g83 );
buf ( n85 , g84 );
buf ( n86 , g85 );
buf ( n87 , g86 );
buf ( n88 , g87 );
buf ( n89 , g88 );
buf ( n90 , g89 );
buf ( n91 , g90 );
buf ( n92 , g91 );
buf ( n93 , g92 );
buf ( n94 , g93 );
buf ( n95 , g94 );
buf ( n96 , g95 );
buf ( n97 , g96 );
buf ( n98 , g97 );
buf ( n99 , g98 );
buf ( g99 , n100 );
buf ( g100 , n101 );
buf ( g101 , n102 );
buf ( g102 , n103 );
buf ( g103 , n104 );
buf ( g104 , n105 );
buf ( g105 , n106 );
buf ( g106 , n107 );
buf ( g107 , n108 );
buf ( g108 , n109 );
buf ( g109 , n110 );
buf ( g110 , n111 );
buf ( g111 , n112 );
buf ( g112 , n113 );
buf ( g113 , n114 );
buf ( g114 , n115 );
buf ( g115 , n116 );
buf ( g116 , n117 );
buf ( g117 , n118 );
buf ( g118 , n119 );
buf ( g119 , n120 );
buf ( g120 , n121 );
buf ( g121 , n122 );
buf ( g122 , n123 );
buf ( g123 , n124 );
buf ( g124 , n125 );
buf ( g125 , n126 );
buf ( g126 , n127 );
buf ( g127 , n128 );
buf ( g128 , n129 );
buf ( g129 , n130 );
buf ( g130 , n131 );
buf ( g131 , n132 );
buf ( g132 , n133 );
buf ( g133 , n134 );
buf ( g134 , n135 );
buf ( g135 , n136 );
buf ( g136 , n137 );
buf ( g137 , n138 );
buf ( g138 , n139 );
buf ( g139 , n140 );
buf ( g140 , n141 );
buf ( g141 , n142 );
buf ( g142 , n143 );
buf ( g143 , n144 );
buf ( g144 , n145 );
buf ( g145 , n146 );
buf ( g146 , n147 );
buf ( g147 , n148 );
buf ( g148 , n149 );
buf ( g149 , n150 );
buf ( g150 , n151 );
buf ( g151 , n152 );
buf ( g152 , n153 );
buf ( g153 , n154 );
buf ( g154 , n155 );
buf ( g155 , n156 );
buf ( g156 , n157 );
buf ( g157 , n158 );
buf ( g158 , n159 );
buf ( g159 , n160 );
buf ( g160 , n161 );
buf ( g161 , n162 );
buf ( g162 , n163 );
buf ( g163 , n164 );
buf ( g164 , n165 );
buf ( g165 , n166 );
buf ( g166 , n167 );
buf ( g167 , n168 );
buf ( g168 , n169 );
buf ( g169 , n170 );
buf ( g170 , n171 );
buf ( g171 , n172 );
buf ( g172 , n173 );
buf ( g173 , n174 );
buf ( g174 , n175 );
buf ( g175 , n176 );
buf ( g176 , n177 );
buf ( g177 , n178 );
buf ( g178 , n179 );
buf ( g179 , n180 );
buf ( g180 , n181 );
buf ( g181 , n182 );
buf ( g182 , n183 );
buf ( g183 , n184 );
buf ( g184 , n185 );
buf ( g185 , n186 );
buf ( g186 , n187 );
buf ( g187 , n188 );
buf ( g188 , n189 );
buf ( g189 , n190 );
buf ( g190 , n191 );
buf ( g191 , n192 );
buf ( g192 , n193 );
buf ( g193 , n194 );
buf ( g194 , n195 );
buf ( g195 , n196 );
buf ( g196 , n197 );
buf ( g197 , n198 );
buf ( g198 , n199 );
buf ( g199 , n200 );
buf ( g200 , n201 );
buf ( g201 , n202 );
buf ( g202 , n203 );
buf ( g203 , n204 );
buf ( g204 , n205 );
buf ( g205 , n206 );
buf ( g206 , n207 );
buf ( g207 , n208 );
buf ( g208 , n209 );
buf ( g209 , n210 );
buf ( g210 , n211 );
buf ( g211 , n212 );
buf ( g212 , n213 );
buf ( g213 , n214 );
buf ( g214 , n215 );
buf ( g215 , n216 );
buf ( g216 , n217 );
buf ( g217 , n218 );
buf ( g218 , n219 );
buf ( g219 , n220 );
buf ( g220 , n221 );
buf ( g221 , n222 );
buf ( g222 , n223 );
buf ( g223 , n224 );
buf ( g224 , n225 );
buf ( g225 , n226 );
buf ( g226 , n227 );
buf ( n100 , n13705 );
buf ( n101 , n13705 );
buf ( n102 , n13704 );
buf ( n103 , n13704 );
buf ( n104 , n13704 );
buf ( n105 , n13705 );
buf ( n106 , n13705 );
buf ( n107 , n13705 );
buf ( n108 , n13704 );
buf ( n109 , n13704 );
buf ( n110 , n13704 );
buf ( n111 , n13705 );
buf ( n112 , n13705 );
buf ( n113 , n13704 );
buf ( n114 , n13704 );
buf ( n115 , n13704 );
buf ( n116 , n13705 );
buf ( n117 , n13705 );
buf ( n118 , n13705 );
buf ( n119 , n13705 );
buf ( n120 , n13704 );
buf ( n121 , n13704 );
buf ( n122 , n13705 );
buf ( n123 , n13704 );
buf ( n124 , n13705 );
buf ( n125 , n13705 );
buf ( n126 , n13704 );
buf ( n127 , n13704 );
buf ( n128 , n13704 );
buf ( n129 , n13705 );
buf ( n130 , n13704 );
buf ( n131 , n13705 );
buf ( n132 , n11070 );
buf ( n133 , n10406 );
buf ( n134 , n13080 );
buf ( n135 , n13124 );
buf ( n136 , n13120 );
buf ( n137 , n13155 );
buf ( n138 , n13157 );
buf ( n139 , n13706 );
buf ( n140 , n13351 );
buf ( n141 , n13359 );
buf ( n142 , n13406 );
buf ( n143 , n13375 );
buf ( n144 , n13376 );
buf ( n145 , n10796 );
buf ( n146 , n13379 );
buf ( n147 , n10620 );
buf ( n148 , n10696 );
buf ( n149 , n13504 );
buf ( n150 , n10643 );
buf ( n151 , n10448 );
buf ( n152 , n13541 );
buf ( n153 , n10576 );
buf ( n154 , n10551 );
buf ( n155 , n10463 );
buf ( n156 , n10486 );
buf ( n157 , n13607 );
buf ( n158 , n10503 );
buf ( n159 , n13665 );
buf ( n160 , n13677 );
buf ( n161 , n13685 );
buf ( n162 , n13690 );
buf ( n163 , n13699 );
buf ( n164 , 1'b0 );
buf ( n165 , 1'b0 );
buf ( n166 , 1'b0 );
buf ( n167 , 1'b0 );
buf ( n168 , 1'b0 );
buf ( n169 , 1'b0 );
buf ( n170 , 1'b0 );
buf ( n171 , n13390 );
buf ( n172 , n13374 );
buf ( n173 , n13374 );
buf ( n174 , n13374 );
buf ( n175 , n13374 );
buf ( n176 , n13374 );
buf ( n177 , n13374 );
buf ( n178 , n13374 );
buf ( n179 , n13374 );
buf ( n180 , n13374 );
buf ( n181 , n13374 );
buf ( n182 , n13374 );
buf ( n183 , n13374 );
buf ( n184 , n13374 );
buf ( n185 , n13374 );
buf ( n186 , n13374 );
buf ( n187 , n13374 );
buf ( n188 , n13374 );
buf ( n189 , n13374 );
buf ( n190 , n13374 );
buf ( n191 , n13374 );
buf ( n192 , n13374 );
buf ( n193 , n13374 );
buf ( n194 , n13374 );
buf ( n195 , n13374 );
buf ( n196 , n13374 );
buf ( n197 , n13374 );
buf ( n198 , n13307 );
buf ( n199 , n13328 );
buf ( n200 , n13213 );
buf ( n201 , n13068 );
buf ( n202 , n13153 );
buf ( n203 , n13090 );
buf ( n204 , n13128 );
buf ( n205 , n13338 );
buf ( n206 , n13178 );
buf ( n207 , n13237 );
buf ( n208 , n13403 );
buf ( n209 , n13373 );
buf ( n210 , n13417 );
buf ( n211 , n13703 );
buf ( n212 , n13444 );
buf ( n213 , n13461 );
buf ( n214 , n13470 );
buf ( n215 , n13480 );
buf ( n216 , n13495 );
buf ( n217 , n13502 );
buf ( n218 , n13513 );
buf ( n219 , n13528 );
buf ( n220 , n13540 );
buf ( n221 , n13553 );
buf ( n222 , n13566 );
buf ( n223 , n13584 );
buf ( n224 , n13602 );
buf ( n225 , n13650 );
buf ( n226 , n13621 );
buf ( n227 , n13654 );
not ( n237 , n1 );
not ( n238 , n237 );
nand ( n239 , n70 , n84 );
nand ( n240 , n69 , n85 );
nand ( n241 , n68 , n86 );
xnor ( n242 , n240 , n241 );
or ( n243 , n239 , n242 );
or ( n244 , n240 , n241 );
nand ( n245 , n243 , n244 );
and ( n246 , n68 , n85 );
not ( n247 , n69 );
not ( n248 , n84 );
nor ( n249 , n247 , n248 );
xor ( n250 , n246 , n249 );
xor ( n251 , n245 , n250 );
xor ( n252 , n242 , n239 );
nand ( n253 , n71 , n84 );
nand ( n254 , n69 , n86 );
nand ( n255 , n68 , n87 );
xnor ( n256 , n254 , n255 );
or ( n257 , n253 , n256 );
or ( n258 , n254 , n255 );
nand ( n259 , n257 , n258 );
xor ( n260 , n252 , n259 );
xor ( n261 , n256 , n253 );
nand ( n262 , n71 , n85 );
nand ( n263 , n69 , n87 );
nand ( n264 , n68 , n88 );
xnor ( n265 , n263 , n264 );
or ( n266 , n262 , n265 );
or ( n267 , n263 , n264 );
nand ( n268 , n266 , n267 );
not ( n269 , n70 );
not ( n270 , n85 );
nor ( n271 , n269 , n270 );
xor ( n272 , n268 , n271 );
and ( n273 , n261 , n272 );
and ( n274 , n271 , n268 );
nor ( n275 , n273 , n274 );
not ( n276 , n275 );
and ( n277 , n260 , n276 );
and ( n278 , n259 , n252 );
nor ( n279 , n277 , n278 );
not ( n280 , n279 );
nor ( n281 , n251 , n280 );
and ( n282 , n260 , n276 );
not ( n283 , n260 );
and ( n284 , n283 , n275 );
nor ( n285 , n282 , n284 );
nand ( n286 , n73 , n84 );
nand ( n287 , n72 , n85 );
nand ( n288 , n70 , n87 );
xnor ( n289 , n287 , n288 );
or ( n290 , n286 , n289 );
or ( n291 , n287 , n288 );
nand ( n292 , n290 , n291 );
not ( n293 , n72 );
nor ( n294 , n293 , n248 );
not ( n295 , n86 );
nor ( n296 , n269 , n295 );
xor ( n297 , n294 , n296 );
xor ( n298 , n292 , n297 );
xor ( n299 , n265 , n262 );
nand ( n300 , n71 , n86 );
nand ( n301 , n69 , n88 );
nand ( n302 , n68 , n89 );
xnor ( n303 , n301 , n302 );
or ( n304 , n300 , n303 );
or ( n305 , n301 , n302 );
nand ( n306 , n304 , n305 );
xor ( n307 , n299 , n306 );
and ( n308 , n298 , n307 );
and ( n309 , n306 , n299 );
nor ( n310 , n308 , n309 );
and ( n311 , n297 , n292 );
and ( n312 , n294 , n296 );
nor ( n313 , n311 , n312 );
xnor ( n314 , n261 , n272 );
xnor ( n315 , n313 , n314 );
or ( n316 , n310 , n315 );
or ( n317 , n313 , n314 );
nand ( n318 , n316 , n317 );
nor ( n319 , n285 , n318 );
nor ( n320 , n281 , n319 );
nand ( n321 , n72 , n89 );
nand ( n322 , n76 , n85 );
nand ( n323 , n75 , n86 );
xnor ( n324 , n322 , n323 );
xnor ( n325 , n321 , n324 );
nand ( n326 , n68 , n93 );
nand ( n327 , n69 , n92 );
not ( n328 , n327 );
and ( n329 , n326 , n328 );
not ( n330 , n326 );
and ( n331 , n330 , n327 );
nor ( n332 , n329 , n331 );
nand ( n333 , n71 , n90 );
and ( n334 , n332 , n333 );
not ( n335 , n332 );
not ( n336 , n333 );
and ( n337 , n335 , n336 );
nor ( n338 , n334 , n337 );
nand ( n339 , n70 , n92 );
nand ( n340 , n78 , n84 );
nand ( n341 , n77 , n85 );
xnor ( n342 , n340 , n341 );
or ( n343 , n339 , n342 );
or ( n344 , n340 , n341 );
nand ( n345 , n343 , n344 );
xnor ( n346 , n338 , n345 );
xnor ( n347 , n325 , n346 );
nand ( n348 , n74 , n87 );
not ( n349 , n348 );
and ( n350 , n71 , n91 );
not ( n351 , n350 );
nand ( n352 , n68 , n94 );
not ( n353 , n352 );
nand ( n354 , n69 , n93 );
not ( n355 , n354 );
not ( n356 , n355 );
or ( n357 , n353 , n356 );
or ( n358 , n355 , n352 );
nand ( n359 , n357 , n358 );
not ( n360 , n359 );
or ( n361 , n351 , n360 );
not ( n362 , n352 );
nand ( n363 , n362 , n355 );
nand ( n364 , n361 , n363 );
not ( n365 , n364 );
and ( n366 , n349 , n365 );
and ( n367 , n348 , n364 );
nor ( n368 , n366 , n367 );
and ( n369 , n72 , n90 );
not ( n370 , n369 );
nand ( n371 , n76 , n86 );
and ( n372 , n75 , n87 );
xnor ( n373 , n371 , n372 );
not ( n374 , n373 );
or ( n375 , n370 , n374 );
not ( n376 , n372 );
or ( n377 , n371 , n376 );
nand ( n378 , n375 , n377 );
xor ( n379 , n368 , n378 );
not ( n380 , n379 );
xor ( n381 , n359 , n350 );
not ( n382 , n381 );
and ( n383 , n342 , n339 );
not ( n384 , n342 );
not ( n385 , n339 );
and ( n386 , n384 , n385 );
nor ( n387 , n383 , n386 );
not ( n388 , n387 );
and ( n389 , n373 , n369 );
not ( n390 , n373 );
not ( n391 , n369 );
and ( n392 , n390 , n391 );
nor ( n393 , n389 , n392 );
not ( n394 , n393 );
not ( n395 , n394 );
or ( n396 , n388 , n395 );
not ( n397 , n387 );
nand ( n398 , n393 , n397 );
nand ( n399 , n396 , n398 );
not ( n400 , n399 );
or ( n401 , n382 , n400 );
not ( n402 , n394 );
nand ( n403 , n402 , n387 );
nand ( n404 , n401 , n403 );
not ( n405 , n404 );
and ( n406 , n380 , n405 );
and ( n407 , n379 , n404 );
nor ( n408 , n406 , n407 );
or ( n409 , n347 , n408 );
not ( n410 , n404 );
or ( n411 , n379 , n410 );
nand ( n412 , n409 , n411 );
and ( n413 , n73 , n89 );
and ( n414 , n74 , n88 );
xor ( n415 , n413 , n414 );
nand ( n416 , n74 , n89 );
not ( n417 , n416 );
not ( n418 , n417 );
nand ( n419 , n73 , n90 );
nand ( n420 , n79 , n84 );
xor ( n421 , n419 , n420 );
not ( n422 , n421 );
or ( n423 , n418 , n422 );
or ( n424 , n420 , n419 );
nand ( n425 , n423 , n424 );
and ( n426 , n415 , n425 );
and ( n427 , n414 , n413 );
nor ( n428 , n426 , n427 );
not ( n429 , n428 );
not ( n430 , n429 );
nand ( n431 , n70 , n93 );
nand ( n432 , n77 , n86 );
nand ( n433 , n78 , n85 );
xor ( n434 , n432 , n433 );
not ( n435 , n434 );
or ( n436 , n431 , n435 );
or ( n437 , n433 , n432 );
nand ( n438 , n436 , n437 );
not ( n439 , n438 );
nand ( n440 , n71 , n92 );
nand ( n441 , n68 , n95 );
nand ( n442 , n69 , n94 );
not ( n443 , n442 );
and ( n444 , n441 , n443 );
not ( n445 , n441 );
and ( n446 , n445 , n442 );
nor ( n447 , n444 , n446 );
or ( n448 , n440 , n447 );
not ( n449 , n443 );
or ( n450 , n449 , n441 );
nand ( n451 , n448 , n450 );
nand ( n452 , n72 , n91 );
not ( n453 , n452 );
not ( n454 , n453 );
nand ( n455 , n75 , n88 );
nand ( n456 , n76 , n87 );
and ( n457 , n455 , n456 );
not ( n458 , n455 );
nand ( n459 , n76 , n87 );
not ( n460 , n459 );
and ( n461 , n458 , n460 );
nor ( n462 , n457 , n461 );
not ( n463 , n462 );
or ( n464 , n454 , n463 );
not ( n465 , n455 );
nand ( n466 , n465 , n460 );
nand ( n467 , n464 , n466 );
xor ( n468 , n451 , n467 );
not ( n469 , n468 );
or ( n470 , n439 , n469 );
nand ( n471 , n467 , n451 );
nand ( n472 , n470 , n471 );
not ( n473 , n472 );
nand ( n474 , n73 , n88 );
nand ( n475 , n77 , n84 );
nand ( n476 , n70 , n91 );
xnor ( n477 , n475 , n476 );
xnor ( n478 , n474 , n477 );
and ( n479 , n473 , n478 );
not ( n480 , n473 );
not ( n481 , n478 );
and ( n482 , n480 , n481 );
nor ( n483 , n479 , n482 );
not ( n484 , n483 );
or ( n485 , n430 , n484 );
nand ( n486 , n481 , n472 );
nand ( n487 , n485 , n486 );
nand ( n488 , n69 , n91 );
nand ( n489 , n68 , n92 );
xnor ( n490 , n488 , n489 );
nand ( n491 , n71 , n89 );
xnor ( n492 , n490 , n491 );
nand ( n493 , n74 , n86 );
nand ( n494 , n70 , n90 );
not ( n495 , n494 );
nand ( n496 , n73 , n87 );
not ( n497 , n496 );
not ( n498 , n497 );
or ( n499 , n495 , n498 );
or ( n500 , n497 , n494 );
nand ( n501 , n499 , n500 );
xor ( n502 , n493 , n501 );
xor ( n503 , n492 , n502 );
nand ( n504 , n76 , n84 );
nand ( n505 , n75 , n85 );
xnor ( n506 , n504 , n505 );
nand ( n507 , n72 , n88 );
xor ( n508 , n506 , n507 );
xor ( n509 , n503 , n508 );
xnor ( n510 , n487 , n509 );
not ( n511 , n510 );
and ( n512 , n412 , n511 );
and ( n513 , n509 , n487 );
nor ( n514 , n512 , n513 );
not ( n515 , n501 );
or ( n516 , n493 , n515 );
or ( n517 , n496 , n494 );
nand ( n518 , n516 , n517 );
and ( n519 , n73 , n86 );
and ( n520 , n74 , n85 );
xor ( n521 , n519 , n520 );
xnor ( n522 , n518 , n521 );
nand ( n523 , n70 , n89 );
nand ( n524 , n75 , n84 );
nand ( n525 , n72 , n87 );
xnor ( n526 , n524 , n525 );
xnor ( n527 , n523 , n526 );
xnor ( n528 , n522 , n527 );
or ( n529 , n474 , n477 );
or ( n530 , n475 , n476 );
nand ( n531 , n529 , n530 );
or ( n532 , n321 , n324 );
or ( n533 , n322 , n323 );
nand ( n534 , n532 , n533 );
or ( n535 , n333 , n332 );
or ( n536 , n327 , n326 );
nand ( n537 , n535 , n536 );
xor ( n538 , n534 , n537 );
and ( n539 , n531 , n538 );
and ( n540 , n534 , n537 );
nor ( n541 , n539 , n540 );
xnor ( n542 , n528 , n541 );
not ( n543 , n502 );
not ( n544 , n492 );
and ( n545 , n543 , n544 );
and ( n546 , n508 , n503 );
nor ( n547 , n545 , n546 );
nand ( n548 , n69 , n90 );
nand ( n549 , n68 , n91 );
xnor ( n550 , n548 , n549 );
nand ( n551 , n71 , n88 );
xor ( n552 , n550 , n551 );
or ( n553 , n507 , n506 );
or ( n554 , n504 , n505 );
nand ( n555 , n553 , n554 );
or ( n556 , n491 , n490 );
or ( n557 , n488 , n489 );
nand ( n558 , n556 , n557 );
xor ( n559 , n555 , n558 );
xnor ( n560 , n552 , n559 );
xnor ( n561 , n547 , n560 );
xor ( n562 , n538 , n531 );
not ( n563 , n348 );
not ( n564 , n563 );
not ( n565 , n364 );
or ( n566 , n564 , n565 );
not ( n567 , n368 );
nand ( n568 , n378 , n567 );
nand ( n569 , n566 , n568 );
not ( n570 , n345 );
not ( n571 , n338 );
or ( n572 , n570 , n571 );
or ( n573 , n325 , n346 );
nand ( n574 , n572 , n573 );
xor ( n575 , n569 , n574 );
and ( n576 , n562 , n575 );
and ( n577 , n569 , n574 );
nor ( n578 , n576 , n577 );
xnor ( n579 , n561 , n578 );
xnor ( n580 , n542 , n579 );
xnor ( n581 , n514 , n580 );
xnor ( n582 , n347 , n408 );
not ( n583 , n428 );
not ( n584 , n483 );
and ( n585 , n583 , n584 );
and ( n586 , n428 , n483 );
nor ( n587 , n585 , n586 );
not ( n588 , n587 );
xor ( n589 , n468 , n438 );
not ( n590 , n589 );
nand ( n591 , n72 , n92 );
nand ( n592 , n76 , n88 );
nand ( n593 , n75 , n89 );
and ( n594 , n592 , n593 );
not ( n595 , n592 );
not ( n596 , n593 );
and ( n597 , n595 , n596 );
or ( n598 , n594 , n597 );
or ( n599 , n591 , n598 );
or ( n600 , n592 , n593 );
nand ( n601 , n599 , n600 );
not ( n602 , n601 );
and ( n603 , n71 , n93 );
not ( n604 , n603 );
nand ( n605 , n68 , n96 );
not ( n606 , n605 );
nand ( n607 , n69 , n95 );
not ( n608 , n607 );
not ( n609 , n608 );
or ( n610 , n606 , n609 );
or ( n611 , n608 , n605 );
nand ( n612 , n610 , n611 );
not ( n613 , n612 );
or ( n614 , n604 , n613 );
not ( n615 , n605 );
nand ( n616 , n615 , n608 );
nand ( n617 , n614 , n616 );
not ( n618 , n617 );
and ( n619 , n80 , n84 );
not ( n620 , n619 );
nand ( n621 , n73 , n91 );
not ( n622 , n621 );
nand ( n623 , n79 , n85 );
not ( n624 , n623 );
not ( n625 , n624 );
or ( n626 , n622 , n625 );
or ( n627 , n624 , n621 );
nand ( n628 , n626 , n627 );
not ( n629 , n628 );
or ( n630 , n620 , n629 );
not ( n631 , n621 );
nand ( n632 , n631 , n624 );
nand ( n633 , n630 , n632 );
not ( n634 , n633 );
not ( n635 , n634 );
or ( n636 , n618 , n635 );
or ( n637 , n634 , n617 );
nand ( n638 , n636 , n637 );
not ( n639 , n638 );
or ( n640 , n602 , n639 );
nand ( n641 , n633 , n617 );
nand ( n642 , n640 , n641 );
xor ( n643 , n425 , n415 );
xor ( n644 , n642 , n643 );
not ( n645 , n644 );
or ( n646 , n590 , n645 );
nand ( n647 , n643 , n642 );
nand ( n648 , n646 , n647 );
not ( n649 , n648 );
or ( n650 , n588 , n649 );
or ( n651 , n587 , n648 );
nand ( n652 , n650 , n651 );
not ( n653 , n652 );
or ( n654 , n582 , n653 );
not ( n655 , n648 );
or ( n656 , n587 , n655 );
nand ( n657 , n654 , n656 );
and ( n658 , n412 , n510 );
not ( n659 , n412 );
and ( n660 , n659 , n511 );
or ( n661 , n658 , n660 );
xor ( n662 , n562 , n575 );
xor ( n663 , n661 , n662 );
and ( n664 , n657 , n663 );
and ( n665 , n662 , n661 );
nor ( n666 , n664 , n665 );
nand ( n667 , n581 , n666 );
xnor ( n668 , n663 , n657 );
not ( n669 , n381 );
and ( n670 , n399 , n669 );
not ( n671 , n399 );
and ( n672 , n671 , n381 );
nor ( n673 , n670 , n672 );
xor ( n674 , n431 , n434 );
not ( n675 , n674 );
nand ( n676 , n70 , n94 );
not ( n677 , n676 );
not ( n678 , n677 );
nand ( n679 , n77 , n87 );
not ( n680 , n679 );
nand ( n681 , n78 , n86 );
not ( n682 , n681 );
not ( n683 , n682 );
or ( n684 , n680 , n683 );
or ( n685 , n682 , n679 );
nand ( n686 , n684 , n685 );
not ( n687 , n686 );
or ( n688 , n678 , n687 );
not ( n689 , n679 );
nand ( n690 , n689 , n682 );
nand ( n691 , n688 , n690 );
nand ( n692 , n675 , n691 );
and ( n693 , n421 , n416 );
not ( n694 , n421 );
and ( n695 , n694 , n417 );
nor ( n696 , n693 , n695 );
not ( n697 , n696 );
xnor ( n698 , n691 , n674 );
nand ( n699 , n697 , n698 );
and ( n700 , n692 , n699 );
xor ( n701 , n673 , n700 );
nand ( n702 , n80 , n85 );
nand ( n703 , n79 , n86 );
nand ( n704 , n73 , n92 );
xnor ( n705 , n703 , n704 );
or ( n706 , n702 , n705 );
or ( n707 , n703 , n704 );
nand ( n708 , n706 , n707 );
not ( n709 , n708 );
nand ( n710 , n74 , n90 );
and ( n711 , n70 , n95 );
not ( n712 , n711 );
nand ( n713 , n77 , n88 );
not ( n714 , n713 );
nand ( n715 , n78 , n87 );
not ( n716 , n715 );
not ( n717 , n716 );
or ( n718 , n714 , n717 );
or ( n719 , n716 , n713 );
nand ( n720 , n718 , n719 );
not ( n721 , n720 );
or ( n722 , n712 , n721 );
not ( n723 , n713 );
nand ( n724 , n723 , n716 );
nand ( n725 , n722 , n724 );
xnor ( n726 , n710 , n725 );
not ( n727 , n726 );
or ( n728 , n709 , n727 );
not ( n729 , n710 );
nand ( n730 , n729 , n725 );
nand ( n731 , n728 , n730 );
not ( n732 , n731 );
not ( n733 , n440 );
and ( n734 , n447 , n733 );
not ( n735 , n447 );
and ( n736 , n735 , n440 );
nor ( n737 , n734 , n736 );
and ( n738 , n462 , n452 );
not ( n739 , n462 );
and ( n740 , n739 , n453 );
nor ( n741 , n738 , n740 );
xnor ( n742 , n737 , n741 );
or ( n743 , n732 , n742 );
or ( n744 , n741 , n737 );
nand ( n745 , n743 , n744 );
xor ( n746 , n701 , n745 );
xor ( n747 , n598 , n591 );
not ( n748 , n747 );
and ( n749 , n686 , n676 );
not ( n750 , n686 );
and ( n751 , n750 , n677 );
nor ( n752 , n749 , n751 );
not ( n753 , n752 );
not ( n754 , n753 );
and ( n755 , n612 , n603 );
not ( n756 , n612 );
not ( n757 , n603 );
and ( n758 , n756 , n757 );
nor ( n759 , n755 , n758 );
not ( n760 , n759 );
not ( n761 , n760 );
or ( n762 , n754 , n761 );
nand ( n763 , n759 , n752 );
nand ( n764 , n762 , n763 );
not ( n765 , n764 );
or ( n766 , n748 , n765 );
nand ( n767 , n753 , n759 );
nand ( n768 , n766 , n767 );
not ( n769 , n768 );
xor ( n770 , n638 , n601 );
not ( n771 , n770 );
or ( n772 , n769 , n771 );
xor ( n773 , n628 , n619 );
and ( n774 , n72 , n93 );
not ( n775 , n774 );
nand ( n776 , n75 , n90 );
not ( n777 , n776 );
nand ( n778 , n76 , n89 );
not ( n779 , n778 );
not ( n780 , n779 );
or ( n781 , n777 , n780 );
or ( n782 , n779 , n776 );
nand ( n783 , n781 , n782 );
not ( n784 , n783 );
or ( n785 , n775 , n784 );
not ( n786 , n776 );
nand ( n787 , n786 , n779 );
nand ( n788 , n785 , n787 );
nand ( n789 , n71 , n94 );
not ( n790 , n789 );
not ( n791 , n790 );
nand ( n792 , n68 , n97 );
nand ( n793 , n69 , n96 );
not ( n794 , n793 );
xnor ( n795 , n792 , n794 );
not ( n796 , n795 );
or ( n797 , n791 , n796 );
not ( n798 , n792 );
nand ( n799 , n798 , n794 );
nand ( n800 , n797 , n799 );
xor ( n801 , n788 , n800 );
and ( n802 , n773 , n801 );
and ( n803 , n788 , n800 );
nor ( n804 , n802 , n803 );
not ( n805 , n804 );
not ( n806 , n768 );
not ( n807 , n806 );
not ( n808 , n770 );
or ( n809 , n807 , n808 );
not ( n810 , n770 );
nand ( n811 , n768 , n810 );
nand ( n812 , n809 , n811 );
nand ( n813 , n805 , n812 );
nand ( n814 , n772 , n813 );
and ( n815 , n644 , n589 );
not ( n816 , n644 );
not ( n817 , n589 );
and ( n818 , n816 , n817 );
nor ( n819 , n815 , n818 );
xor ( n820 , n814 , n819 );
and ( n821 , n746 , n820 );
and ( n822 , n819 , n814 );
nor ( n823 , n821 , n822 );
not ( n824 , n582 );
not ( n825 , n652 );
and ( n826 , n824 , n825 );
and ( n827 , n582 , n652 );
nor ( n828 , n826 , n827 );
not ( n829 , n745 );
not ( n830 , n701 );
or ( n831 , n829 , n830 );
or ( n832 , n700 , n673 );
nand ( n833 , n831 , n832 );
and ( n834 , n828 , n833 );
not ( n835 , n828 );
not ( n836 , n833 );
and ( n837 , n835 , n836 );
nor ( n838 , n834 , n837 );
or ( n839 , n823 , n838 );
or ( n840 , n836 , n828 );
nand ( n841 , n839 , n840 );
not ( n842 , n841 );
nand ( n843 , n668 , n842 );
nand ( n844 , n71 , n96 );
nand ( n845 , n83 , n84 );
nand ( n846 , n75 , n92 );
xnor ( n847 , n845 , n846 );
or ( n848 , n844 , n847 );
or ( n849 , n845 , n846 );
nand ( n850 , n848 , n849 );
nand ( n851 , n68 , n99 );
not ( n852 , n851 );
and ( n853 , n4 , n852 );
nand ( n854 , n82 , n85 );
not ( n855 , n854 );
not ( n856 , n855 );
nand ( n857 , n70 , n97 );
nand ( n858 , n74 , n93 );
and ( n859 , n857 , n858 );
not ( n860 , n857 );
nand ( n861 , n74 , n93 );
not ( n862 , n861 );
and ( n863 , n860 , n862 );
nor ( n864 , n859 , n863 );
not ( n865 , n864 );
or ( n866 , n856 , n865 );
not ( n867 , n862 );
or ( n868 , n867 , n857 );
nand ( n869 , n866 , n868 );
xor ( n870 , n853 , n869 );
xnor ( n871 , n850 , n870 );
nand ( n872 , n69 , n99 );
not ( n873 , n872 );
nand ( n874 , n873 , n5 );
not ( n875 , n874 );
xor ( n876 , n4 , n852 );
not ( n877 , n876 );
not ( n878 , n877 );
and ( n879 , n875 , n878 );
and ( n880 , n83 , n85 );
not ( n881 , n880 );
nand ( n882 , n75 , n93 );
nand ( n883 , n71 , n97 );
and ( n884 , n882 , n883 );
not ( n885 , n882 );
not ( n886 , n883 );
and ( n887 , n885 , n886 );
nor ( n888 , n884 , n887 );
not ( n889 , n888 );
or ( n890 , n881 , n889 );
not ( n891 , n882 );
nand ( n892 , n891 , n886 );
nand ( n893 , n890 , n892 );
and ( n894 , n874 , n876 );
not ( n895 , n874 );
and ( n896 , n895 , n877 );
or ( n897 , n894 , n896 );
and ( n898 , n893 , n897 );
nor ( n899 , n879 , n898 );
and ( n900 , n79 , n88 );
not ( n901 , n900 );
nand ( n902 , n72 , n95 );
not ( n903 , n902 );
nand ( n904 , n78 , n89 );
not ( n905 , n904 );
not ( n906 , n905 );
or ( n907 , n903 , n906 );
or ( n908 , n905 , n902 );
nand ( n909 , n907 , n908 );
not ( n910 , n909 );
or ( n911 , n901 , n910 );
not ( n912 , n902 );
nand ( n913 , n912 , n905 );
nand ( n914 , n911 , n913 );
nand ( n915 , n69 , n98 );
not ( n916 , n915 );
not ( n917 , n916 );
nand ( n918 , n76 , n91 );
not ( n919 , n918 );
nand ( n920 , n77 , n90 );
not ( n921 , n920 );
not ( n922 , n921 );
or ( n923 , n919 , n922 );
or ( n924 , n921 , n918 );
nand ( n925 , n923 , n924 );
not ( n926 , n925 );
or ( n927 , n917 , n926 );
not ( n928 , n918 );
nand ( n929 , n928 , n921 );
nand ( n930 , n927 , n929 );
xor ( n931 , n914 , n930 );
nand ( n932 , n81 , n86 );
nand ( n933 , n73 , n94 );
nand ( n934 , n80 , n87 );
xor ( n935 , n933 , n934 );
not ( n936 , n935 );
or ( n937 , n932 , n936 );
or ( n938 , n934 , n933 );
nand ( n939 , n937 , n938 );
and ( n940 , n931 , n939 );
not ( n941 , n931 );
not ( n942 , n939 );
and ( n943 , n941 , n942 );
nor ( n944 , n940 , n943 );
and ( n945 , n899 , n944 );
not ( n946 , n899 );
not ( n947 , n944 );
and ( n948 , n946 , n947 );
nor ( n949 , n945 , n948 );
or ( n950 , n871 , n949 );
or ( n951 , n899 , n947 );
nand ( n952 , n950 , n951 );
not ( n953 , n952 );
nand ( n954 , n79 , n87 );
nand ( n955 , n73 , n93 );
xor ( n956 , n954 , n955 );
nand ( n957 , n80 , n86 );
and ( n958 , n956 , n957 );
not ( n959 , n956 );
not ( n960 , n957 );
and ( n961 , n959 , n960 );
nor ( n962 , n958 , n961 );
nand ( n963 , n77 , n89 );
not ( n964 , n963 );
nand ( n965 , n78 , n88 );
not ( n966 , n965 );
not ( n967 , n966 );
or ( n968 , n964 , n967 );
or ( n969 , n966 , n963 );
nand ( n970 , n968 , n969 );
and ( n971 , n70 , n96 );
not ( n972 , n971 );
and ( n973 , n970 , n972 );
not ( n974 , n970 );
and ( n975 , n974 , n971 );
nor ( n976 , n973 , n975 );
not ( n977 , n976 );
and ( n978 , n962 , n977 );
not ( n979 , n962 );
and ( n980 , n979 , n976 );
nor ( n981 , n978 , n980 );
nand ( n982 , n74 , n94 );
not ( n983 , n982 );
not ( n984 , n983 );
nand ( n985 , n79 , n89 );
not ( n986 , n985 );
nand ( n987 , n80 , n88 );
not ( n988 , n987 );
not ( n989 , n988 );
or ( n990 , n986 , n989 );
not ( n991 , n987 );
or ( n992 , n991 , n985 );
nand ( n993 , n990 , n992 );
not ( n994 , n993 );
or ( n995 , n984 , n994 );
not ( n996 , n991 );
or ( n997 , n996 , n985 );
nand ( n998 , n995 , n997 );
not ( n999 , n998 );
nand ( n1000 , n77 , n91 );
not ( n1001 , n1000 );
not ( n1002 , n1001 );
nand ( n1003 , n72 , n96 );
not ( n1004 , n1003 );
nand ( n1005 , n76 , n92 );
not ( n1006 , n1005 );
not ( n1007 , n1006 );
or ( n1008 , n1004 , n1007 );
or ( n1009 , n1006 , n1003 );
nand ( n1010 , n1008 , n1009 );
not ( n1011 , n1010 );
or ( n1012 , n1002 , n1011 );
not ( n1013 , n1003 );
nand ( n1014 , n1013 , n1006 );
nand ( n1015 , n1012 , n1014 );
and ( n1016 , n73 , n95 );
not ( n1017 , n1016 );
nand ( n1018 , n78 , n90 );
not ( n1019 , n1018 );
nand ( n1020 , n70 , n98 );
not ( n1021 , n1020 );
not ( n1022 , n1021 );
or ( n1023 , n1019 , n1022 );
or ( n1024 , n1021 , n1018 );
nand ( n1025 , n1023 , n1024 );
not ( n1026 , n1025 );
or ( n1027 , n1017 , n1026 );
not ( n1028 , n1018 );
nand ( n1029 , n1028 , n1021 );
nand ( n1030 , n1027 , n1029 );
xor ( n1031 , n1015 , n1030 );
not ( n1032 , n1031 );
or ( n1033 , n999 , n1032 );
nand ( n1034 , n1015 , n1030 );
nand ( n1035 , n1033 , n1034 );
not ( n1036 , n1035 );
or ( n1037 , n981 , n1036 );
or ( n1038 , n976 , n962 );
nand ( n1039 , n1037 , n1038 );
nand ( n1040 , n72 , n94 );
not ( n1041 , n1040 );
not ( n1042 , n1041 );
nand ( n1043 , n76 , n90 );
not ( n1044 , n1043 );
nand ( n1045 , n75 , n91 );
not ( n1046 , n1045 );
not ( n1047 , n1046 );
or ( n1048 , n1044 , n1047 );
not ( n1049 , n1043 );
nand ( n1050 , n1045 , n1049 );
nand ( n1051 , n1048 , n1050 );
not ( n1052 , n1051 );
or ( n1053 , n1042 , n1052 );
not ( n1054 , n1043 );
nand ( n1055 , n1054 , n1046 );
nand ( n1056 , n1053 , n1055 );
not ( n1057 , n1056 );
not ( n1058 , n971 );
not ( n1059 , n970 );
or ( n1060 , n1058 , n1059 );
not ( n1061 , n963 );
nand ( n1062 , n1061 , n966 );
nand ( n1063 , n1060 , n1062 );
not ( n1064 , n1063 );
not ( n1065 , n1064 );
or ( n1066 , n1057 , n1065 );
or ( n1067 , n1064 , n1056 );
nand ( n1068 , n1066 , n1067 );
not ( n1069 , n960 );
not ( n1070 , n956 );
or ( n1071 , n1069 , n1070 );
or ( n1072 , n954 , n955 );
nand ( n1073 , n1071 , n1072 );
xnor ( n1074 , n1068 , n1073 );
and ( n1075 , n850 , n870 );
and ( n1076 , n853 , n869 );
nor ( n1077 , n1075 , n1076 );
not ( n1078 , n1077 );
not ( n1079 , n939 );
not ( n1080 , n931 );
or ( n1081 , n1079 , n1080 );
nand ( n1082 , n930 , n914 );
nand ( n1083 , n1081 , n1082 );
not ( n1084 , n1083 );
or ( n1085 , n1078 , n1084 );
or ( n1086 , n1077 , n1083 );
nand ( n1087 , n1085 , n1086 );
xor ( n1088 , n1074 , n1087 );
xnor ( n1089 , n1039 , n1088 );
not ( n1090 , n1089 );
or ( n1091 , n953 , n1090 );
not ( n1092 , n1088 );
nand ( n1093 , n1092 , n1039 );
nand ( n1094 , n1091 , n1093 );
not ( n1095 , n1094 );
xor ( n1096 , n702 , n705 );
xor ( n1097 , n711 , n720 );
xnor ( n1098 , n1096 , n1097 );
nand ( n1099 , n82 , n84 );
not ( n1100 , n1099 );
not ( n1101 , n1100 );
nand ( n1102 , n81 , n85 );
nand ( n1103 , n74 , n92 );
and ( n1104 , n1102 , n1103 );
not ( n1105 , n1102 );
not ( n1106 , n1103 );
and ( n1107 , n1105 , n1106 );
nor ( n1108 , n1104 , n1107 );
not ( n1109 , n1108 );
or ( n1110 , n1101 , n1109 );
not ( n1111 , n1102 );
nand ( n1112 , n1111 , n1106 );
nand ( n1113 , n1110 , n1112 );
and ( n1114 , n81 , n84 );
nand ( n1115 , n74 , n91 );
and ( n1116 , n1114 , n1115 );
not ( n1117 , n1114 );
not ( n1118 , n1115 );
and ( n1119 , n1117 , n1118 );
nor ( n1120 , n1116 , n1119 );
and ( n1121 , n1113 , n1120 );
not ( n1122 , n1113 );
not ( n1123 , n1120 );
and ( n1124 , n1122 , n1123 );
nor ( n1125 , n1121 , n1124 );
xor ( n1126 , n1098 , n1125 );
and ( n1127 , n1108 , n1100 );
not ( n1128 , n1108 );
and ( n1129 , n1128 , n1099 );
nor ( n1130 , n1127 , n1129 );
not ( n1131 , n1130 );
and ( n1132 , n1051 , n1040 );
not ( n1133 , n1051 );
and ( n1134 , n1133 , n1041 );
nor ( n1135 , n1132 , n1134 );
not ( n1136 , n1135 );
not ( n1137 , n1136 );
nand ( n1138 , n71 , n95 );
not ( n1139 , n1138 );
nand ( n1140 , n69 , n97 );
not ( n1141 , n1140 );
and ( n1142 , n68 , n98 );
not ( n1143 , n1142 );
or ( n1144 , n1141 , n1143 );
or ( n1145 , n1142 , n1140 );
nand ( n1146 , n1144 , n1145 );
not ( n1147 , n1146 );
or ( n1148 , n1139 , n1147 );
or ( n1149 , n1138 , n1146 );
nand ( n1150 , n1148 , n1149 );
not ( n1151 , n1150 );
not ( n1152 , n1151 );
or ( n1153 , n1137 , n1152 );
nand ( n1154 , n1150 , n1135 );
nand ( n1155 , n1153 , n1154 );
not ( n1156 , n1155 );
or ( n1157 , n1131 , n1156 );
nand ( n1158 , n1136 , n1150 );
nand ( n1159 , n1157 , n1158 );
not ( n1160 , n1138 );
not ( n1161 , n1160 );
not ( n1162 , n1146 );
or ( n1163 , n1161 , n1162 );
not ( n1164 , n1140 );
nand ( n1165 , n1164 , n1142 );
nand ( n1166 , n1163 , n1165 );
not ( n1167 , n1166 );
xnor ( n1168 , n774 , n783 );
not ( n1169 , n1168 );
or ( n1170 , n1167 , n1169 );
or ( n1171 , n1166 , n1168 );
nand ( n1172 , n1170 , n1171 );
and ( n1173 , n795 , n790 );
not ( n1174 , n795 );
and ( n1175 , n1174 , n789 );
nor ( n1176 , n1173 , n1175 );
and ( n1177 , n1172 , n1176 );
not ( n1178 , n1172 );
not ( n1179 , n1176 );
and ( n1180 , n1178 , n1179 );
nor ( n1181 , n1177 , n1180 );
xor ( n1182 , n1159 , n1181 );
and ( n1183 , n1126 , n1182 );
and ( n1184 , n1159 , n1181 );
nor ( n1185 , n1183 , n1184 );
xor ( n1186 , n764 , n747 );
not ( n1187 , n1176 );
not ( n1188 , n1172 );
or ( n1189 , n1187 , n1188 );
not ( n1190 , n1168 );
nand ( n1191 , n1166 , n1190 );
nand ( n1192 , n1189 , n1191 );
not ( n1193 , n1192 );
not ( n1194 , n1193 );
not ( n1195 , n773 );
not ( n1196 , n801 );
not ( n1197 , n1196 );
or ( n1198 , n1195 , n1197 );
not ( n1199 , n773 );
nand ( n1200 , n1199 , n801 );
nand ( n1201 , n1198 , n1200 );
not ( n1202 , n1201 );
or ( n1203 , n1194 , n1202 );
not ( n1204 , n1192 );
or ( n1205 , n1204 , n1201 );
nand ( n1206 , n1203 , n1205 );
xor ( n1207 , n1186 , n1206 );
xor ( n1208 , n1185 , n1207 );
or ( n1209 , n1095 , n1208 );
not ( n1210 , n1207 );
or ( n1211 , n1185 , n1210 );
nand ( n1212 , n1209 , n1211 );
not ( n1213 , n1212 );
not ( n1214 , n731 );
not ( n1215 , n742 );
or ( n1216 , n1214 , n1215 );
or ( n1217 , n731 , n742 );
nand ( n1218 , n1216 , n1217 );
not ( n1219 , n696 );
not ( n1220 , n698 );
or ( n1221 , n1219 , n1220 );
or ( n1222 , n696 , n698 );
nand ( n1223 , n1221 , n1222 );
xor ( n1224 , n1218 , n1223 );
xnor ( n1225 , n708 , n726 );
nand ( n1226 , n1063 , n1056 );
nand ( n1227 , n1073 , n1068 );
and ( n1228 , n1226 , n1227 );
and ( n1229 , n1123 , n1113 );
and ( n1230 , n1114 , n1118 );
nor ( n1231 , n1229 , n1230 );
not ( n1232 , n1231 );
and ( n1233 , n1228 , n1232 );
not ( n1234 , n1228 );
and ( n1235 , n1234 , n1231 );
nor ( n1236 , n1233 , n1235 );
or ( n1237 , n1225 , n1236 );
or ( n1238 , n1231 , n1228 );
nand ( n1239 , n1237 , n1238 );
xor ( n1240 , n1224 , n1239 );
not ( n1241 , n1125 );
not ( n1242 , n1098 );
and ( n1243 , n1241 , n1242 );
and ( n1244 , n1097 , n1096 );
nor ( n1245 , n1243 , n1244 );
not ( n1246 , n1245 );
not ( n1247 , n1246 );
not ( n1248 , n1074 );
not ( n1249 , n1248 );
not ( n1250 , n1087 );
or ( n1251 , n1249 , n1250 );
not ( n1252 , n1077 );
nand ( n1253 , n1252 , n1083 );
nand ( n1254 , n1251 , n1253 );
not ( n1255 , n1254 );
or ( n1256 , n1247 , n1255 );
and ( n1257 , n1236 , n1225 );
not ( n1258 , n1236 );
not ( n1259 , n1225 );
and ( n1260 , n1258 , n1259 );
nor ( n1261 , n1257 , n1260 );
xnor ( n1262 , n1245 , n1254 );
nand ( n1263 , n1261 , n1262 );
nand ( n1264 , n1256 , n1263 );
and ( n1265 , n812 , n805 );
not ( n1266 , n812 );
and ( n1267 , n1266 , n804 );
nor ( n1268 , n1265 , n1267 );
not ( n1269 , n1186 );
not ( n1270 , n1206 );
or ( n1271 , n1269 , n1270 );
not ( n1272 , n1201 );
or ( n1273 , n1204 , n1272 );
nand ( n1274 , n1271 , n1273 );
and ( n1275 , n1268 , n1274 );
not ( n1276 , n1268 );
not ( n1277 , n1274 );
and ( n1278 , n1276 , n1277 );
nor ( n1279 , n1275 , n1278 );
xor ( n1280 , n1264 , n1279 );
xor ( n1281 , n1240 , n1280 );
not ( n1282 , n1281 );
or ( n1283 , n1213 , n1282 );
nand ( n1284 , n1240 , n1280 );
nand ( n1285 , n1283 , n1284 );
not ( n1286 , n1285 );
xnor ( n1287 , n820 , n746 );
and ( n1288 , n1239 , n1224 );
and ( n1289 , n1223 , n1218 );
nor ( n1290 , n1288 , n1289 );
xnor ( n1291 , n1287 , n1290 );
and ( n1292 , n1264 , n1279 );
and ( n1293 , n1274 , n1268 );
nor ( n1294 , n1292 , n1293 );
xor ( n1295 , n1291 , n1294 );
not ( n1296 , n1295 );
nand ( n1297 , n1286 , n1296 );
not ( n1298 , n1297 );
xor ( n1299 , n838 , n823 );
or ( n1300 , n1294 , n1291 );
or ( n1301 , n1290 , n1287 );
nand ( n1302 , n1300 , n1301 );
nor ( n1303 , n1299 , n1302 );
nor ( n1304 , n1298 , n1303 );
xnor ( n1305 , n1155 , n1130 );
not ( n1306 , n1305 );
not ( n1307 , n1306 );
xor ( n1308 , n847 , n844 );
not ( n1309 , n1308 );
not ( n1310 , n932 );
not ( n1311 , n935 );
or ( n1312 , n1310 , n1311 );
or ( n1313 , n932 , n935 );
nand ( n1314 , n1312 , n1313 );
not ( n1315 , n1314 );
and ( n1316 , n864 , n854 );
not ( n1317 , n864 );
and ( n1318 , n1317 , n855 );
nor ( n1319 , n1316 , n1318 );
not ( n1320 , n1319 );
or ( n1321 , n1315 , n1320 );
not ( n1322 , n1319 );
not ( n1323 , n1314 );
nand ( n1324 , n1322 , n1323 );
nand ( n1325 , n1321 , n1324 );
not ( n1326 , n1325 );
or ( n1327 , n1309 , n1326 );
not ( n1328 , n1319 );
nand ( n1329 , n1328 , n1314 );
nand ( n1330 , n1327 , n1329 );
not ( n1331 , n1330 );
nand ( n1332 , n70 , n99 );
not ( n1333 , n1332 );
nand ( n1334 , n1333 , n6 );
nand ( n1335 , n81 , n87 );
nand ( n1336 , n82 , n86 );
not ( n1337 , n1336 );
and ( n1338 , n1335 , n1337 );
not ( n1339 , n1335 );
and ( n1340 , n1339 , n1336 );
nor ( n1341 , n1338 , n1340 );
or ( n1342 , n1334 , n1341 );
or ( n1343 , n1336 , n1335 );
nand ( n1344 , n1342 , n1343 );
and ( n1345 , n925 , n916 );
not ( n1346 , n925 );
and ( n1347 , n1346 , n915 );
nor ( n1348 , n1345 , n1347 );
and ( n1349 , n909 , n900 );
not ( n1350 , n909 );
not ( n1351 , n900 );
and ( n1352 , n1350 , n1351 );
nor ( n1353 , n1349 , n1352 );
xor ( n1354 , n1348 , n1353 );
and ( n1355 , n1344 , n1354 );
and ( n1356 , n1348 , n1353 );
nor ( n1357 , n1355 , n1356 );
and ( n1358 , n1331 , n1357 );
not ( n1359 , n1331 );
not ( n1360 , n1357 );
and ( n1361 , n1359 , n1360 );
nor ( n1362 , n1358 , n1361 );
not ( n1363 , n1362 );
or ( n1364 , n1307 , n1363 );
or ( n1365 , n1357 , n1331 );
nand ( n1366 , n1364 , n1365 );
and ( n1367 , n1182 , n1126 );
not ( n1368 , n1182 );
not ( n1369 , n1126 );
and ( n1370 , n1368 , n1369 );
nor ( n1371 , n1367 , n1370 );
not ( n1372 , n1371 );
and ( n1373 , n1366 , n1372 );
not ( n1374 , n1366 );
and ( n1375 , n1374 , n1371 );
nor ( n1376 , n1373 , n1375 );
not ( n1377 , n1376 );
not ( n1378 , n952 );
and ( n1379 , n1089 , n1378 );
not ( n1380 , n1089 );
and ( n1381 , n1380 , n952 );
nor ( n1382 , n1379 , n1381 );
not ( n1383 , n1382 );
and ( n1384 , n1377 , n1383 );
and ( n1385 , n1366 , n1371 );
nor ( n1386 , n1384 , n1385 );
not ( n1387 , n1261 );
not ( n1388 , n1262 );
not ( n1389 , n1388 );
and ( n1390 , n1387 , n1389 );
and ( n1391 , n1261 , n1388 );
nor ( n1392 , n1390 , n1391 );
not ( n1393 , n1094 );
not ( n1394 , n1208 );
and ( n1395 , n1393 , n1394 );
and ( n1396 , n1094 , n1208 );
nor ( n1397 , n1395 , n1396 );
xor ( n1398 , n1392 , n1397 );
not ( n1399 , n1398 );
or ( n1400 , n1386 , n1399 );
or ( n1401 , n1392 , n1397 );
nand ( n1402 , n1400 , n1401 );
not ( n1403 , n1402 );
xnor ( n1404 , n1212 , n1281 );
nand ( n1405 , n1403 , n1404 );
not ( n1406 , n1398 );
not ( n1407 , n1386 );
and ( n1408 , n1406 , n1407 );
and ( n1409 , n1386 , n1398 );
nor ( n1410 , n1408 , n1409 );
not ( n1411 , n949 );
and ( n1412 , n871 , n1411 );
not ( n1413 , n871 );
and ( n1414 , n1413 , n949 );
nor ( n1415 , n1412 , n1414 );
not ( n1416 , n1415 );
not ( n1417 , n1416 );
xnor ( n1418 , n1305 , n1362 );
not ( n1419 , n1418 );
or ( n1420 , n1417 , n1419 );
nand ( n1421 , n82 , n87 );
not ( n1422 , n1421 );
not ( n1423 , n1422 );
nand ( n1424 , n75 , n94 );
nand ( n1425 , n81 , n88 );
and ( n1426 , n1424 , n1425 );
not ( n1427 , n1424 );
nand ( n1428 , n81 , n88 );
not ( n1429 , n1428 );
and ( n1430 , n1427 , n1429 );
nor ( n1431 , n1426 , n1430 );
not ( n1432 , n1431 );
or ( n1433 , n1423 , n1432 );
not ( n1434 , n1424 );
nand ( n1435 , n1434 , n1429 );
nand ( n1436 , n1433 , n1435 );
nand ( n1437 , n80 , n89 );
not ( n1438 , n1437 );
not ( n1439 , n1438 );
nand ( n1440 , n71 , n98 );
nand ( n1441 , n74 , n95 );
and ( n1442 , n1440 , n1441 );
not ( n1443 , n1440 );
nand ( n1444 , n74 , n95 );
not ( n1445 , n1444 );
and ( n1446 , n1443 , n1445 );
nor ( n1447 , n1442 , n1446 );
not ( n1448 , n1447 );
or ( n1449 , n1439 , n1448 );
not ( n1450 , n1445 );
or ( n1451 , n1450 , n1440 );
nand ( n1452 , n1449 , n1451 );
xor ( n1453 , n1436 , n1452 );
xor ( n1454 , n888 , n880 );
xor ( n1455 , n1453 , n1454 );
not ( n1456 , n1455 );
nand ( n1457 , n77 , n92 );
nand ( n1458 , n76 , n93 );
nand ( n1459 , n72 , n97 );
xnor ( n1460 , n1458 , n1459 );
or ( n1461 , n1457 , n1460 );
or ( n1462 , n1458 , n1459 );
nand ( n1463 , n1461 , n1462 );
not ( n1464 , n5 );
not ( n1465 , n872 );
and ( n1466 , n1464 , n1465 );
and ( n1467 , n5 , n872 );
nor ( n1468 , n1466 , n1467 );
not ( n1469 , n1468 );
nand ( n1470 , n79 , n90 );
not ( n1471 , n1470 );
not ( n1472 , n1471 );
nand ( n1473 , n73 , n96 );
not ( n1474 , n1473 );
nand ( n1475 , n78 , n91 );
not ( n1476 , n1475 );
not ( n1477 , n1476 );
or ( n1478 , n1474 , n1477 );
or ( n1479 , n1476 , n1473 );
nand ( n1480 , n1478 , n1479 );
not ( n1481 , n1480 );
or ( n1482 , n1472 , n1481 );
not ( n1483 , n1473 );
nand ( n1484 , n1483 , n1476 );
nand ( n1485 , n1482 , n1484 );
not ( n1486 , n1485 );
or ( n1487 , n1469 , n1486 );
or ( n1488 , n1468 , n1485 );
nand ( n1489 , n1487 , n1488 );
not ( n1490 , n1489 );
and ( n1491 , n1463 , n1490 );
not ( n1492 , n1463 );
and ( n1493 , n1492 , n1489 );
nor ( n1494 , n1491 , n1493 );
not ( n1495 , n1494 );
not ( n1496 , n1495 );
xor ( n1497 , n1460 , n1457 );
not ( n1498 , n1497 );
nand ( n1499 , n81 , n89 );
not ( n1500 , n1499 );
not ( n1501 , n1500 );
nand ( n1502 , n75 , n95 );
not ( n1503 , n1502 );
nand ( n1504 , n72 , n98 );
not ( n1505 , n1504 );
not ( n1506 , n1505 );
or ( n1507 , n1503 , n1506 );
or ( n1508 , n1505 , n1502 );
nand ( n1509 , n1507 , n1508 );
not ( n1510 , n1509 );
or ( n1511 , n1501 , n1510 );
not ( n1512 , n1502 );
nand ( n1513 , n1512 , n1505 );
nand ( n1514 , n1511 , n1513 );
not ( n1515 , n1514 );
and ( n1516 , n1431 , n1421 );
not ( n1517 , n1431 );
and ( n1518 , n1517 , n1422 );
nor ( n1519 , n1516 , n1518 );
not ( n1520 , n1519 );
or ( n1521 , n1515 , n1520 );
not ( n1522 , n1514 );
not ( n1523 , n1519 );
nand ( n1524 , n1522 , n1523 );
nand ( n1525 , n1521 , n1524 );
not ( n1526 , n1525 );
or ( n1527 , n1498 , n1526 );
not ( n1528 , n1519 );
nand ( n1529 , n1528 , n1514 );
nand ( n1530 , n1527 , n1529 );
not ( n1531 , n1530 );
not ( n1532 , n1531 );
or ( n1533 , n1496 , n1532 );
nand ( n1534 , n1494 , n1530 );
nand ( n1535 , n1533 , n1534 );
not ( n1536 , n1535 );
or ( n1537 , n1456 , n1536 );
nand ( n1538 , n1495 , n1530 );
nand ( n1539 , n1537 , n1538 );
not ( n1540 , n1539 );
xnor ( n1541 , n1325 , n1308 );
not ( n1542 , n1541 );
nand ( n1543 , n83 , n87 );
nand ( n1544 , n76 , n94 );
nand ( n1545 , n82 , n88 );
not ( n1546 , n1545 );
and ( n1547 , n1544 , n1546 );
not ( n1548 , n1544 );
and ( n1549 , n1548 , n1545 );
nor ( n1550 , n1547 , n1549 );
or ( n1551 , n1543 , n1550 );
or ( n1552 , n1545 , n1544 );
nand ( n1553 , n1551 , n1552 );
not ( n1554 , n1553 );
nand ( n1555 , n78 , n92 );
not ( n1556 , n1555 );
not ( n1557 , n1556 );
nand ( n1558 , n73 , n97 );
nand ( n1559 , n77 , n93 );
and ( n1560 , n1558 , n1559 );
not ( n1561 , n1558 );
not ( n1562 , n1559 );
and ( n1563 , n1561 , n1562 );
nor ( n1564 , n1560 , n1563 );
not ( n1565 , n1564 );
or ( n1566 , n1557 , n1565 );
not ( n1567 , n1558 );
nand ( n1568 , n1567 , n1562 );
nand ( n1569 , n1566 , n1568 );
nand ( n1570 , n80 , n90 );
not ( n1571 , n1570 );
not ( n1572 , n1571 );
nand ( n1573 , n74 , n96 );
nand ( n1574 , n79 , n91 );
and ( n1575 , n1573 , n1574 );
not ( n1576 , n1573 );
not ( n1577 , n1574 );
and ( n1578 , n1576 , n1577 );
nor ( n1579 , n1575 , n1578 );
not ( n1580 , n1579 );
or ( n1581 , n1572 , n1580 );
not ( n1582 , n1573 );
nand ( n1583 , n1582 , n1577 );
nand ( n1584 , n1581 , n1583 );
xor ( n1585 , n1569 , n1584 );
not ( n1586 , n1585 );
or ( n1587 , n1554 , n1586 );
nand ( n1588 , n1584 , n1569 );
nand ( n1589 , n1587 , n1588 );
not ( n1590 , n1589 );
not ( n1591 , n7 );
nand ( n1592 , n71 , n99 );
nor ( n1593 , n1591 , n1592 );
not ( n1594 , n1593 );
nand ( n1595 , n83 , n86 );
not ( n1596 , n6 );
not ( n1597 , n1332 );
or ( n1598 , n1596 , n1597 );
or ( n1599 , n6 , n1332 );
nand ( n1600 , n1598 , n1599 );
xnor ( n1601 , n1595 , n1600 );
not ( n1602 , n1601 );
or ( n1603 , n1594 , n1602 );
not ( n1604 , n1595 );
nand ( n1605 , n1604 , n1600 );
nand ( n1606 , n1603 , n1605 );
xor ( n1607 , n1341 , n1334 );
xor ( n1608 , n1606 , n1607 );
not ( n1609 , n1608 );
or ( n1610 , n1590 , n1609 );
nand ( n1611 , n1607 , n1606 );
nand ( n1612 , n1610 , n1611 );
not ( n1613 , n1612 );
or ( n1614 , n1542 , n1613 );
or ( n1615 , n1541 , n1612 );
nand ( n1616 , n1614 , n1615 );
not ( n1617 , n1616 );
or ( n1618 , n1540 , n1617 );
not ( n1619 , n1541 );
nand ( n1620 , n1619 , n1612 );
nand ( n1621 , n1618 , n1620 );
not ( n1622 , n1621 );
not ( n1623 , n1622 );
not ( n1624 , n1416 );
not ( n1625 , n1418 );
not ( n1626 , n1625 );
or ( n1627 , n1624 , n1626 );
nand ( n1628 , n1415 , n1418 );
nand ( n1629 , n1627 , n1628 );
nand ( n1630 , n1623 , n1629 );
nand ( n1631 , n1420 , n1630 );
and ( n1632 , n1454 , n1453 );
and ( n1633 , n1436 , n1452 );
nor ( n1634 , n1632 , n1633 );
not ( n1635 , n1634 );
not ( n1636 , n998 );
not ( n1637 , n1636 );
not ( n1638 , n1031 );
and ( n1639 , n1637 , n1638 );
and ( n1640 , n1636 , n1031 );
nor ( n1641 , n1639 , n1640 );
not ( n1642 , n1641 );
and ( n1643 , n1635 , n1642 );
xor ( n1644 , n1354 , n1344 );
xnor ( n1645 , n1634 , n1641 );
not ( n1646 , n1645 );
and ( n1647 , n1644 , n1646 );
nor ( n1648 , n1643 , n1647 );
not ( n1649 , n1648 );
and ( n1650 , n993 , n982 );
not ( n1651 , n993 );
and ( n1652 , n1651 , n983 );
nor ( n1653 , n1650 , n1652 );
not ( n1654 , n1653 );
not ( n1655 , n1654 );
and ( n1656 , n1010 , n1001 );
not ( n1657 , n1010 );
not ( n1658 , n1001 );
and ( n1659 , n1657 , n1658 );
nor ( n1660 , n1656 , n1659 );
not ( n1661 , n1660 );
or ( n1662 , n1655 , n1661 );
xnor ( n1663 , n1025 , n1016 );
not ( n1664 , n1663 );
not ( n1665 , n1654 );
not ( n1666 , n1660 );
not ( n1667 , n1666 );
or ( n1668 , n1665 , n1667 );
nand ( n1669 , n1660 , n1653 );
nand ( n1670 , n1668 , n1669 );
nand ( n1671 , n1664 , n1670 );
nand ( n1672 , n1662 , n1671 );
not ( n1673 , n1672 );
xor ( n1674 , n893 , n897 );
not ( n1675 , n1674 );
not ( n1676 , n1463 );
not ( n1677 , n1489 );
or ( n1678 , n1676 , n1677 );
not ( n1679 , n1468 );
nand ( n1680 , n1679 , n1485 );
nand ( n1681 , n1678 , n1680 );
not ( n1682 , n1681 );
not ( n1683 , n1682 );
or ( n1684 , n1675 , n1683 );
not ( n1685 , n1674 );
nand ( n1686 , n1685 , n1681 );
nand ( n1687 , n1684 , n1686 );
not ( n1688 , n1687 );
or ( n1689 , n1673 , n1688 );
nand ( n1690 , n1674 , n1681 );
nand ( n1691 , n1689 , n1690 );
xor ( n1692 , n1036 , n981 );
not ( n1693 , n1692 );
and ( n1694 , n1691 , n1693 );
not ( n1695 , n1691 );
and ( n1696 , n1695 , n1692 );
nor ( n1697 , n1694 , n1696 );
not ( n1698 , n1697 );
and ( n1699 , n1649 , n1698 );
buf ( n1700 , n1692 );
and ( n1701 , n1700 , n1691 );
nor ( n1702 , n1699 , n1701 );
not ( n1703 , n1702 );
and ( n1704 , n1631 , n1703 );
not ( n1705 , n1631 );
and ( n1706 , n1705 , n1702 );
nor ( n1707 , n1704 , n1706 );
xor ( n1708 , n1382 , n1376 );
and ( n1709 , n1707 , n1708 );
and ( n1710 , n1703 , n1631 );
nor ( n1711 , n1709 , n1710 );
nand ( n1712 , n1410 , n1711 );
and ( n1713 , n79 , n92 );
not ( n1714 , n1713 );
nand ( n1715 , n74 , n97 );
and ( n1716 , n78 , n93 );
xnor ( n1717 , n1715 , n1716 );
not ( n1718 , n1717 );
or ( n1719 , n1714 , n1718 );
not ( n1720 , n1715 );
nand ( n1721 , n1720 , n1716 );
nand ( n1722 , n1719 , n1721 );
not ( n1723 , n1722 );
not ( n1724 , n8 );
nand ( n1725 , n72 , n99 );
nor ( n1726 , n1724 , n1725 );
xor ( n1727 , n1592 , n7 );
xor ( n1728 , n1726 , n1727 );
not ( n1729 , n1728 );
or ( n1730 , n1723 , n1729 );
or ( n1731 , n1722 , n1728 );
nand ( n1732 , n1730 , n1731 );
not ( n1733 , n1732 );
not ( n1734 , n8 );
not ( n1735 , n1725 );
and ( n1736 , n1734 , n1735 );
and ( n1737 , n8 , n1725 );
nor ( n1738 , n1736 , n1737 );
nand ( n1739 , n77 , n94 );
nand ( n1740 , n83 , n88 );
xnor ( n1741 , n1739 , n1740 );
or ( n1742 , n1738 , n1741 );
or ( n1743 , n1740 , n1739 );
nand ( n1744 , n1742 , n1743 );
nand ( n1745 , n83 , n89 );
not ( n1746 , n1745 );
not ( n1747 , n1746 );
nand ( n1748 , n74 , n98 );
not ( n1749 , n1748 );
nand ( n1750 , n77 , n95 );
not ( n1751 , n1750 );
not ( n1752 , n1751 );
or ( n1753 , n1749 , n1752 );
or ( n1754 , n1751 , n1748 );
nand ( n1755 , n1753 , n1754 );
not ( n1756 , n1755 );
or ( n1757 , n1747 , n1756 );
or ( n1758 , n1750 , n1748 );
nand ( n1759 , n1757 , n1758 );
not ( n1760 , n1759 );
nand ( n1761 , n73 , n99 );
not ( n1762 , n1761 );
nand ( n1763 , n1762 , n9 );
nand ( n1764 , n82 , n90 );
not ( n1765 , n1764 );
not ( n1766 , n1765 );
nand ( n1767 , n76 , n96 );
not ( n1768 , n1767 );
nand ( n1769 , n81 , n91 );
not ( n1770 , n1769 );
not ( n1771 , n1770 );
or ( n1772 , n1768 , n1771 );
or ( n1773 , n1770 , n1767 );
nand ( n1774 , n1772 , n1773 );
not ( n1775 , n1774 );
or ( n1776 , n1766 , n1775 );
not ( n1777 , n1767 );
nand ( n1778 , n1777 , n1770 );
nand ( n1779 , n1776 , n1778 );
xnor ( n1780 , n1763 , n1779 );
not ( n1781 , n1780 );
or ( n1782 , n1760 , n1781 );
not ( n1783 , n1763 );
nand ( n1784 , n1783 , n1779 );
nand ( n1785 , n1782 , n1784 );
xor ( n1786 , n1744 , n1785 );
not ( n1787 , n1786 );
or ( n1788 , n1733 , n1787 );
nand ( n1789 , n1744 , n1785 );
nand ( n1790 , n1788 , n1789 );
xor ( n1791 , n1585 , n1553 );
not ( n1792 , n1791 );
xnor ( n1793 , n1525 , n1497 );
not ( n1794 , n1793 );
or ( n1795 , n1792 , n1794 );
or ( n1796 , n1791 , n1793 );
nand ( n1797 , n1795 , n1796 );
xor ( n1798 , n1790 , n1797 );
not ( n1799 , n1798 );
and ( n1800 , n1717 , n1713 );
not ( n1801 , n1717 );
not ( n1802 , n1713 );
and ( n1803 , n1801 , n1802 );
nor ( n1804 , n1800 , n1803 );
not ( n1805 , n1804 );
and ( n1806 , n74 , n99 );
and ( n1807 , n10 , n1806 );
not ( n1808 , n1807 );
nand ( n1809 , n78 , n94 );
not ( n1810 , n9 );
not ( n1811 , n1761 );
or ( n1812 , n1810 , n1811 );
or ( n1813 , n9 , n1761 );
nand ( n1814 , n1812 , n1813 );
xnor ( n1815 , n1809 , n1814 );
not ( n1816 , n1815 );
or ( n1817 , n1808 , n1816 );
not ( n1818 , n1809 );
nand ( n1819 , n1818 , n1814 );
nand ( n1820 , n1817 , n1819 );
not ( n1821 , n1820 );
or ( n1822 , n1805 , n1821 );
xnor ( n1823 , n1741 , n1738 );
not ( n1824 , n1823 );
xor ( n1825 , n1804 , n1820 );
nand ( n1826 , n1824 , n1825 );
nand ( n1827 , n1822 , n1826 );
not ( n1828 , n1827 );
xor ( n1829 , n1780 , n1759 );
not ( n1830 , n1829 );
nand ( n1831 , n83 , n90 );
nand ( n1832 , n82 , n91 );
nand ( n1833 , n77 , n96 );
xnor ( n1834 , n1832 , n1833 );
or ( n1835 , n1831 , n1834 );
or ( n1836 , n1832 , n1833 );
nand ( n1837 , n1835 , n1836 );
not ( n1838 , n1837 );
nand ( n1839 , n81 , n92 );
not ( n1840 , n1839 );
not ( n1841 , n1840 );
nand ( n1842 , n76 , n97 );
not ( n1843 , n1842 );
nand ( n1844 , n80 , n93 );
not ( n1845 , n1844 );
not ( n1846 , n1845 );
or ( n1847 , n1843 , n1846 );
or ( n1848 , n1845 , n1842 );
nand ( n1849 , n1847 , n1848 );
not ( n1850 , n1849 );
or ( n1851 , n1841 , n1850 );
not ( n1852 , n1842 );
nand ( n1853 , n1852 , n1845 );
nand ( n1854 , n1851 , n1853 );
nand ( n1855 , n79 , n94 );
not ( n1856 , n1855 );
not ( n1857 , n1856 );
nand ( n1858 , n78 , n95 );
nand ( n1859 , n75 , n98 );
not ( n1860 , n1859 );
xnor ( n1861 , n1858 , n1860 );
not ( n1862 , n1861 );
or ( n1863 , n1857 , n1862 );
not ( n1864 , n1858 );
nand ( n1865 , n1864 , n1860 );
nand ( n1866 , n1863 , n1865 );
xor ( n1867 , n1854 , n1866 );
not ( n1868 , n1867 );
or ( n1869 , n1838 , n1868 );
nand ( n1870 , n1854 , n1866 );
nand ( n1871 , n1869 , n1870 );
not ( n1872 , n1871 );
not ( n1873 , n1872 );
nand ( n1874 , n75 , n97 );
not ( n1875 , n1874 );
nand ( n1876 , n79 , n93 );
not ( n1877 , n1876 );
not ( n1878 , n1877 );
or ( n1879 , n1875 , n1878 );
or ( n1880 , n1877 , n1874 );
nand ( n1881 , n1879 , n1880 );
and ( n1882 , n80 , n92 );
and ( n1883 , n1881 , n1882 );
not ( n1884 , n1881 );
not ( n1885 , n1882 );
and ( n1886 , n1884 , n1885 );
nor ( n1887 , n1883 , n1886 );
not ( n1888 , n1887 );
not ( n1889 , n1764 );
not ( n1890 , n1774 );
and ( n1891 , n1889 , n1890 );
and ( n1892 , n1764 , n1774 );
nor ( n1893 , n1891 , n1892 );
not ( n1894 , n1893 );
not ( n1895 , n1894 );
not ( n1896 , n1745 );
not ( n1897 , n1755 );
or ( n1898 , n1896 , n1897 );
or ( n1899 , n1745 , n1755 );
nand ( n1900 , n1898 , n1899 );
not ( n1901 , n1900 );
not ( n1902 , n1901 );
or ( n1903 , n1895 , n1902 );
nand ( n1904 , n1900 , n1893 );
nand ( n1905 , n1903 , n1904 );
not ( n1906 , n1905 );
or ( n1907 , n1888 , n1906 );
nand ( n1908 , n1894 , n1900 );
nand ( n1909 , n1907 , n1908 );
not ( n1910 , n1909 );
or ( n1911 , n1873 , n1910 );
or ( n1912 , n1872 , n1909 );
nand ( n1913 , n1911 , n1912 );
not ( n1914 , n1913 );
or ( n1915 , n1830 , n1914 );
nand ( n1916 , n1871 , n1909 );
nand ( n1917 , n1915 , n1916 );
not ( n1918 , n1917 );
or ( n1919 , n1828 , n1918 );
xor ( n1920 , n1732 , n1786 );
and ( n1921 , n1917 , n1827 );
not ( n1922 , n1917 );
not ( n1923 , n1827 );
and ( n1924 , n1922 , n1923 );
nor ( n1925 , n1921 , n1924 );
nand ( n1926 , n1920 , n1925 );
nand ( n1927 , n1919 , n1926 );
not ( n1928 , n1927 );
or ( n1929 , n1799 , n1928 );
and ( n1930 , n1509 , n1500 );
not ( n1931 , n1509 );
and ( n1932 , n1931 , n1499 );
nor ( n1933 , n1930 , n1932 );
not ( n1934 , n1933 );
and ( n1935 , n1564 , n1556 );
not ( n1936 , n1564 );
and ( n1937 , n1936 , n1555 );
nor ( n1938 , n1935 , n1937 );
not ( n1939 , n1938 );
and ( n1940 , n1579 , n1570 );
not ( n1941 , n1579 );
and ( n1942 , n1941 , n1571 );
nor ( n1943 , n1940 , n1942 );
not ( n1944 , n1943 );
or ( n1945 , n1939 , n1944 );
or ( n1946 , n1943 , n1938 );
nand ( n1947 , n1945 , n1946 );
not ( n1948 , n1947 );
or ( n1949 , n1934 , n1948 );
not ( n1950 , n1943 );
nand ( n1951 , n1950 , n1938 );
nand ( n1952 , n1949 , n1951 );
not ( n1953 , n1726 );
not ( n1954 , n1727 );
not ( n1955 , n1954 );
or ( n1956 , n1953 , n1955 );
not ( n1957 , n1728 );
nand ( n1958 , n1722 , n1957 );
nand ( n1959 , n1956 , n1958 );
xnor ( n1960 , n1952 , n1959 );
not ( n1961 , n1543 );
and ( n1962 , n1550 , n1961 );
not ( n1963 , n1550 );
and ( n1964 , n1963 , n1543 );
nor ( n1965 , n1962 , n1964 );
not ( n1966 , n1965 );
and ( n1967 , n82 , n89 );
not ( n1968 , n1967 );
nand ( n1969 , n76 , n95 );
not ( n1970 , n1969 );
nand ( n1971 , n73 , n98 );
not ( n1972 , n1971 );
not ( n1973 , n1972 );
or ( n1974 , n1970 , n1973 );
or ( n1975 , n1972 , n1969 );
nand ( n1976 , n1974 , n1975 );
not ( n1977 , n1976 );
or ( n1978 , n1968 , n1977 );
not ( n1979 , n1969 );
nand ( n1980 , n1979 , n1972 );
nand ( n1981 , n1978 , n1980 );
not ( n1982 , n1981 );
and ( n1983 , n81 , n90 );
not ( n1984 , n1983 );
nand ( n1985 , n75 , n96 );
not ( n1986 , n1985 );
nand ( n1987 , n80 , n91 );
not ( n1988 , n1987 );
not ( n1989 , n1988 );
or ( n1990 , n1986 , n1989 );
or ( n1991 , n1988 , n1985 );
nand ( n1992 , n1990 , n1991 );
not ( n1993 , n1992 );
or ( n1994 , n1984 , n1993 );
not ( n1995 , n1985 );
nand ( n1996 , n1995 , n1988 );
nand ( n1997 , n1994 , n1996 );
not ( n1998 , n1997 );
not ( n1999 , n1998 );
or ( n2000 , n1982 , n1999 );
or ( n2001 , n1998 , n1981 );
nand ( n2002 , n2000 , n2001 );
and ( n2003 , n1966 , n2002 );
and ( n2004 , n1997 , n1981 );
nor ( n2005 , n2003 , n2004 );
xor ( n2006 , n1960 , n2005 );
not ( n2007 , n2006 );
xor ( n2008 , n1947 , n1933 );
not ( n2009 , n2008 );
xor ( n2010 , n1992 , n1983 );
not ( n2011 , n2010 );
not ( n2012 , n1882 );
not ( n2013 , n1881 );
or ( n2014 , n2012 , n2013 );
not ( n2015 , n1874 );
nand ( n2016 , n2015 , n1877 );
nand ( n2017 , n2014 , n2016 );
not ( n2018 , n2017 );
xnor ( n2019 , n1967 , n1976 );
not ( n2020 , n2019 );
or ( n2021 , n2018 , n2020 );
or ( n2022 , n2017 , n2019 );
nand ( n2023 , n2021 , n2022 );
not ( n2024 , n2023 );
or ( n2025 , n2011 , n2024 );
not ( n2026 , n2019 );
nand ( n2027 , n2017 , n2026 );
nand ( n2028 , n2025 , n2027 );
not ( n2029 , n1965 );
not ( n2030 , n2002 );
or ( n2031 , n2029 , n2030 );
or ( n2032 , n1965 , n2002 );
nand ( n2033 , n2031 , n2032 );
xor ( n2034 , n2028 , n2033 );
not ( n2035 , n2034 );
or ( n2036 , n2009 , n2035 );
nand ( n2037 , n2028 , n2033 );
nand ( n2038 , n2036 , n2037 );
and ( n2039 , n1447 , n1437 );
not ( n2040 , n1447 );
and ( n2041 , n2040 , n1438 );
nor ( n2042 , n2039 , n2041 );
and ( n2043 , n1480 , n1471 );
not ( n2044 , n1480 );
and ( n2045 , n2044 , n1470 );
nor ( n2046 , n2043 , n2045 );
not ( n2047 , n2046 );
and ( n2048 , n2042 , n2047 );
not ( n2049 , n2042 );
and ( n2050 , n2049 , n2046 );
nor ( n2051 , n2048 , n2050 );
xor ( n2052 , n1601 , n1593 );
xor ( n2053 , n2051 , n2052 );
and ( n2054 , n2038 , n2053 );
not ( n2055 , n2038 );
not ( n2056 , n2053 );
and ( n2057 , n2055 , n2056 );
nor ( n2058 , n2054 , n2057 );
not ( n2059 , n2058 );
not ( n2060 , n2059 );
or ( n2061 , n2007 , n2060 );
or ( n2062 , n2006 , n2059 );
nand ( n2063 , n2061 , n2062 );
and ( n2064 , n1927 , n1798 );
not ( n2065 , n1927 );
and ( n2066 , n2065 , n1799 );
nor ( n2067 , n2064 , n2066 );
nand ( n2068 , n2063 , n2067 );
nand ( n2069 , n1929 , n2068 );
nand ( n2070 , n2053 , n2038 );
nand ( n2071 , n2006 , n2058 );
and ( n2072 , n2070 , n2071 );
xor ( n2073 , n1608 , n1589 );
not ( n2074 , n2047 );
not ( n2075 , n2042 );
and ( n2076 , n2074 , n2075 );
and ( n2077 , n2052 , n2051 );
nor ( n2078 , n2076 , n2077 );
not ( n2079 , n2078 );
not ( n2080 , n2079 );
not ( n2081 , n1670 );
and ( n2082 , n1663 , n2081 );
not ( n2083 , n1663 );
and ( n2084 , n2083 , n1670 );
nor ( n2085 , n2082 , n2084 );
not ( n2086 , n2085 );
not ( n2087 , n2086 );
or ( n2088 , n2080 , n2087 );
nand ( n2089 , n2078 , n2085 );
nand ( n2090 , n2088 , n2089 );
xnor ( n2091 , n2073 , n2090 );
not ( n2092 , n2091 );
and ( n2093 , n2072 , n2092 );
not ( n2094 , n2072 );
and ( n2095 , n2094 , n2091 );
nor ( n2096 , n2093 , n2095 );
xor ( n2097 , n1535 , n1455 );
or ( n2098 , n2005 , n1960 );
not ( n2099 , n1959 );
not ( n2100 , n1952 );
or ( n2101 , n2099 , n2100 );
nand ( n2102 , n2098 , n2101 );
xnor ( n2103 , n2097 , n2102 );
not ( n2104 , n1790 );
not ( n2105 , n1797 );
or ( n2106 , n2104 , n2105 );
not ( n2107 , n1793 );
nand ( n2108 , n1791 , n2107 );
nand ( n2109 , n2106 , n2108 );
not ( n2110 , n2109 );
xnor ( n2111 , n2103 , n2110 );
xor ( n2112 , n2096 , n2111 );
nand ( n2113 , n2069 , n2112 );
not ( n2114 , n2110 );
not ( n2115 , n2103 );
and ( n2116 , n2114 , n2115 );
and ( n2117 , n2102 , n2097 );
nor ( n2118 , n2116 , n2117 );
not ( n2119 , n2118 );
xor ( n2120 , n1539 , n1616 );
not ( n2121 , n2073 );
not ( n2122 , n2090 );
or ( n2123 , n2121 , n2122 );
or ( n2124 , n2078 , n2086 );
nand ( n2125 , n2123 , n2124 );
not ( n2126 , n2125 );
and ( n2127 , n1687 , n1672 );
not ( n2128 , n1687 );
not ( n2129 , n1672 );
and ( n2130 , n2128 , n2129 );
or ( n2131 , n2127 , n2130 );
not ( n2132 , n2131 );
not ( n2133 , n1644 );
not ( n2134 , n1645 );
or ( n2135 , n2133 , n2134 );
or ( n2136 , n1644 , n1645 );
nand ( n2137 , n2135 , n2136 );
not ( n2138 , n2137 );
and ( n2139 , n2132 , n2138 );
and ( n2140 , n2131 , n2137 );
nor ( n2141 , n2139 , n2140 );
not ( n2142 , n2141 );
and ( n2143 , n2126 , n2142 );
and ( n2144 , n2125 , n2141 );
nor ( n2145 , n2143 , n2144 );
xnor ( n2146 , n2120 , n2145 );
not ( n2147 , n2146 );
or ( n2148 , n2119 , n2147 );
or ( n2149 , n2118 , n2146 );
nand ( n2150 , n2148 , n2149 );
or ( n2151 , n2111 , n2096 );
or ( n2152 , n2091 , n2072 );
nand ( n2153 , n2151 , n2152 );
nor ( n2154 , n2150 , n2153 );
or ( n2155 , n2113 , n2154 );
nand ( n2156 , n2150 , n2153 );
nand ( n2157 , n2155 , n2156 );
not ( n2158 , n1622 );
not ( n2159 , n1629 );
and ( n2160 , n2158 , n2159 );
and ( n2161 , n1622 , n1629 );
nor ( n2162 , n2160 , n2161 );
not ( n2163 , n2162 );
xor ( n2164 , n1648 , n1697 );
not ( n2165 , n2164 );
not ( n2166 , n2125 );
or ( n2167 , n2166 , n2141 );
buf ( n2168 , n2131 );
not ( n2169 , n2137 );
or ( n2170 , n2168 , n2169 );
nand ( n2171 , n2167 , n2170 );
not ( n2172 , n2171 );
not ( n2173 , n2172 );
or ( n2174 , n2165 , n2173 );
not ( n2175 , n2164 );
nand ( n2176 , n2175 , n2171 );
nand ( n2177 , n2174 , n2176 );
not ( n2178 , n2177 );
or ( n2179 , n2163 , n2178 );
or ( n2180 , n2162 , n2177 );
nand ( n2181 , n2179 , n2180 );
not ( n2182 , n2118 );
not ( n2183 , n2182 );
not ( n2184 , n2146 );
or ( n2185 , n2183 , n2184 );
not ( n2186 , n2145 );
nand ( n2187 , n2186 , n2120 );
nand ( n2188 , n2185 , n2187 );
nor ( n2189 , n2181 , n2188 );
xor ( n2190 , n1707 , n1708 );
not ( n2191 , n2162 );
not ( n2192 , n2191 );
not ( n2193 , n2177 );
or ( n2194 , n2192 , n2193 );
not ( n2195 , n2172 );
nand ( n2196 , n2195 , n2164 );
nand ( n2197 , n2194 , n2196 );
nor ( n2198 , n2190 , n2197 );
nor ( n2199 , n2189 , n2198 );
nand ( n2200 , n1405 , n1712 , n2157 , n2199 );
nand ( n2201 , n2181 , n2188 );
or ( n2202 , n2198 , n2201 );
nand ( n2203 , n2190 , n2197 );
nand ( n2204 , n2202 , n2203 );
nand ( n2205 , n2204 , n1712 );
not ( n2206 , n1410 );
not ( n2207 , n1711 );
nand ( n2208 , n2206 , n2207 );
nand ( n2209 , n2205 , n2208 );
nand ( n2210 , n2209 , n1405 );
not ( n2211 , n1404 );
nand ( n2212 , n1402 , n2211 );
and ( n2213 , n2200 , n2210 , n2212 );
and ( n2214 , n2199 , n1712 );
not ( n2215 , n2069 );
not ( n2216 , n2112 );
nand ( n2217 , n2215 , n2216 );
xor ( n2218 , n1867 , n1837 );
xor ( n2219 , n1815 , n1807 );
and ( n2220 , n76 , n98 );
not ( n2221 , n2220 );
nand ( n2222 , n78 , n96 );
not ( n2223 , n2222 );
and ( n2224 , n83 , n91 );
not ( n2225 , n2224 );
or ( n2226 , n2223 , n2225 );
or ( n2227 , n2224 , n2222 );
nand ( n2228 , n2226 , n2227 );
not ( n2229 , n2228 );
or ( n2230 , n2221 , n2229 );
not ( n2231 , n2224 );
or ( n2232 , n2231 , n2222 );
nand ( n2233 , n2230 , n2232 );
not ( n2234 , n2233 );
not ( n2235 , n11 );
nand ( n2236 , n75 , n99 );
or ( n2237 , n2235 , n2236 );
not ( n2238 , n2237 );
xor ( n2239 , n10 , n1806 );
not ( n2240 , n2239 );
or ( n2241 , n2238 , n2240 );
or ( n2242 , n2237 , n2239 );
nand ( n2243 , n2241 , n2242 );
not ( n2244 , n2243 );
or ( n2245 , n2234 , n2244 );
not ( n2246 , n2237 );
nand ( n2247 , n2246 , n2239 );
nand ( n2248 , n2245 , n2247 );
xor ( n2249 , n2219 , n2248 );
and ( n2250 , n2218 , n2249 );
and ( n2251 , n2219 , n2248 );
nor ( n2252 , n2250 , n2251 );
xor ( n2253 , n2023 , n2010 );
not ( n2254 , n1823 );
not ( n2255 , n1825 );
and ( n2256 , n2254 , n2255 );
and ( n2257 , n1823 , n1825 );
nor ( n2258 , n2256 , n2257 );
and ( n2259 , n2253 , n2258 );
not ( n2260 , n2253 );
not ( n2261 , n2258 );
and ( n2262 , n2260 , n2261 );
nor ( n2263 , n2259 , n2262 );
xor ( n2264 , n2252 , n2263 );
xor ( n2265 , n2233 , n2243 );
and ( n2266 , n1834 , n1831 );
not ( n2267 , n1834 );
not ( n2268 , n1831 );
and ( n2269 , n2267 , n2268 );
nor ( n2270 , n2266 , n2269 );
not ( n2271 , n11 );
not ( n2272 , n2236 );
or ( n2273 , n2271 , n2272 );
or ( n2274 , n11 , n2236 );
nand ( n2275 , n2273 , n2274 );
not ( n2276 , n2275 );
nand ( n2277 , n80 , n94 );
nand ( n2278 , n79 , n95 );
and ( n2279 , n2277 , n2278 );
not ( n2280 , n2277 );
not ( n2281 , n2278 );
and ( n2282 , n2280 , n2281 );
nor ( n2283 , n2279 , n2282 );
not ( n2284 , n2283 );
or ( n2285 , n2276 , n2284 );
not ( n2286 , n2277 );
nand ( n2287 , n2286 , n2281 );
nand ( n2288 , n2285 , n2287 );
xor ( n2289 , n2270 , n2288 );
and ( n2290 , n2265 , n2289 );
and ( n2291 , n2288 , n2270 );
nor ( n2292 , n2290 , n2291 );
not ( n2293 , n2292 );
not ( n2294 , n2293 );
and ( n2295 , n1861 , n1856 );
not ( n2296 , n1861 );
and ( n2297 , n2296 , n1855 );
nor ( n2298 , n2295 , n2297 );
not ( n2299 , n2298 );
not ( n2300 , n1839 );
not ( n2301 , n1849 );
or ( n2302 , n2300 , n2301 );
or ( n2303 , n1839 , n1849 );
nand ( n2304 , n2302 , n2303 );
and ( n2305 , n82 , n92 );
not ( n2306 , n2305 );
nand ( n2307 , n77 , n97 );
not ( n2308 , n2307 );
nand ( n2309 , n81 , n93 );
not ( n2310 , n2309 );
not ( n2311 , n2310 );
or ( n2312 , n2308 , n2311 );
or ( n2313 , n2310 , n2307 );
nand ( n2314 , n2312 , n2313 );
not ( n2315 , n2314 );
or ( n2316 , n2306 , n2315 );
not ( n2317 , n2307 );
nand ( n2318 , n2317 , n2310 );
nand ( n2319 , n2316 , n2318 );
xor ( n2320 , n2304 , n2319 );
not ( n2321 , n2320 );
or ( n2322 , n2299 , n2321 );
nand ( n2323 , n2319 , n2304 );
nand ( n2324 , n2322 , n2323 );
not ( n2325 , n1887 );
and ( n2326 , n1905 , n2325 );
not ( n2327 , n1905 );
and ( n2328 , n2327 , n1887 );
nor ( n2329 , n2326 , n2328 );
not ( n2330 , n2329 );
and ( n2331 , n2324 , n2330 );
not ( n2332 , n2324 );
and ( n2333 , n2332 , n2329 );
nor ( n2334 , n2331 , n2333 );
not ( n2335 , n2334 );
or ( n2336 , n2294 , n2335 );
not ( n2337 , n2324 );
or ( n2338 , n2337 , n2329 );
nand ( n2339 , n2336 , n2338 );
xor ( n2340 , n1913 , n1829 );
and ( n2341 , n2339 , n2340 );
not ( n2342 , n2339 );
not ( n2343 , n2340 );
and ( n2344 , n2342 , n2343 );
nor ( n2345 , n2341 , n2344 );
and ( n2346 , n2264 , n2345 );
and ( n2347 , n2339 , n2340 );
nor ( n2348 , n2346 , n2347 );
not ( n2349 , n1925 );
xor ( n2350 , n2349 , n1920 );
not ( n2351 , n2252 );
not ( n2352 , n2263 );
and ( n2353 , n2351 , n2352 );
and ( n2354 , n2253 , n2261 );
nor ( n2355 , n2353 , n2354 );
xor ( n2356 , n2034 , n2008 );
and ( n2357 , n2355 , n2356 );
not ( n2358 , n2355 );
not ( n2359 , n2356 );
and ( n2360 , n2358 , n2359 );
nor ( n2361 , n2357 , n2360 );
xnor ( n2362 , n2350 , n2361 );
nand ( n2363 , n2348 , n2362 );
not ( n2364 , n2363 );
and ( n2365 , n2334 , n2293 );
not ( n2366 , n2334 );
and ( n2367 , n2366 , n2292 );
nor ( n2368 , n2365 , n2367 );
xnor ( n2369 , n2249 , n2218 );
nand ( n2370 , n81 , n94 );
not ( n2371 , n2370 );
and ( n2372 , n76 , n99 );
xor ( n2373 , n12 , n2372 );
not ( n2374 , n2373 );
not ( n2375 , n2374 );
and ( n2376 , n2371 , n2375 );
nand ( n2377 , n77 , n99 );
not ( n2378 , n2377 );
and ( n2379 , n13 , n2378 );
and ( n2380 , n2370 , n2373 );
not ( n2381 , n2370 );
and ( n2382 , n2381 , n2374 );
or ( n2383 , n2380 , n2382 );
and ( n2384 , n2379 , n2383 );
nor ( n2385 , n2376 , n2384 );
not ( n2386 , n2220 );
and ( n2387 , n2228 , n2386 );
not ( n2388 , n2228 );
and ( n2389 , n2388 , n2220 );
nor ( n2390 , n2387 , n2389 );
and ( n2391 , n2314 , n2305 );
not ( n2392 , n2314 );
not ( n2393 , n2305 );
and ( n2394 , n2392 , n2393 );
nor ( n2395 , n2391 , n2394 );
and ( n2396 , n2390 , n2395 );
not ( n2397 , n2390 );
not ( n2398 , n2395 );
and ( n2399 , n2397 , n2398 );
nor ( n2400 , n2396 , n2399 );
or ( n2401 , n2385 , n2400 );
or ( n2402 , n2390 , n2398 );
nand ( n2403 , n2401 , n2402 );
not ( n2404 , n2403 );
nand ( n2405 , n83 , n92 );
nand ( n2406 , n78 , n97 );
nand ( n2407 , n82 , n93 );
not ( n2408 , n2407 );
and ( n2409 , n2406 , n2408 );
not ( n2410 , n2406 );
and ( n2411 , n2410 , n2407 );
nor ( n2412 , n2409 , n2411 );
or ( n2413 , n2405 , n2412 );
or ( n2414 , n2407 , n2406 );
nand ( n2415 , n2413 , n2414 );
and ( n2416 , n12 , n2372 );
not ( n2417 , n2416 );
and ( n2418 , n80 , n95 );
not ( n2419 , n2418 );
nand ( n2420 , n79 , n96 );
not ( n2421 , n2420 );
nand ( n2422 , n77 , n98 );
not ( n2423 , n2422 );
not ( n2424 , n2423 );
or ( n2425 , n2421 , n2424 );
or ( n2426 , n2423 , n2420 );
nand ( n2427 , n2425 , n2426 );
not ( n2428 , n2427 );
or ( n2429 , n2419 , n2428 );
not ( n2430 , n2420 );
nand ( n2431 , n2430 , n2423 );
nand ( n2432 , n2429 , n2431 );
not ( n2433 , n2432 );
not ( n2434 , n2433 );
or ( n2435 , n2417 , n2434 );
not ( n2436 , n2416 );
nand ( n2437 , n2436 , n2432 );
nand ( n2438 , n2435 , n2437 );
and ( n2439 , n2415 , n2438 );
and ( n2440 , n2416 , n2432 );
nor ( n2441 , n2439 , n2440 );
and ( n2442 , n2320 , n2298 );
not ( n2443 , n2320 );
not ( n2444 , n2298 );
and ( n2445 , n2443 , n2444 );
nor ( n2446 , n2442 , n2445 );
xor ( n2447 , n2441 , n2446 );
not ( n2448 , n2447 );
not ( n2449 , n2448 );
or ( n2450 , n2404 , n2449 );
not ( n2451 , n2441 );
nand ( n2452 , n2451 , n2446 );
nand ( n2453 , n2450 , n2452 );
xnor ( n2454 , n2369 , n2453 );
and ( n2455 , n2368 , n2454 );
not ( n2456 , n2369 );
and ( n2457 , n2456 , n2453 );
nor ( n2458 , n2455 , n2457 );
xor ( n2459 , n2264 , n2345 );
not ( n2460 , n2459 );
nand ( n2461 , n2458 , n2460 );
not ( n2462 , n2461 );
not ( n2463 , n2403 );
not ( n2464 , n2463 );
not ( n2465 , n2448 );
or ( n2466 , n2464 , n2465 );
nand ( n2467 , n2403 , n2447 );
nand ( n2468 , n2466 , n2467 );
xor ( n2469 , n2289 , n2265 );
not ( n2470 , n2469 );
not ( n2471 , n2418 );
and ( n2472 , n2427 , n2471 );
not ( n2473 , n2427 );
and ( n2474 , n2473 , n2418 );
nor ( n2475 , n2472 , n2474 );
not ( n2476 , n2475 );
nand ( n2477 , n82 , n94 );
not ( n2478 , n2477 );
not ( n2479 , n2478 );
nand ( n2480 , n81 , n95 );
not ( n2481 , n2480 );
nand ( n2482 , n78 , n98 );
not ( n2483 , n2482 );
not ( n2484 , n2483 );
or ( n2485 , n2481 , n2484 );
or ( n2486 , n2483 , n2480 );
nand ( n2487 , n2485 , n2486 );
not ( n2488 , n2487 );
or ( n2489 , n2479 , n2488 );
not ( n2490 , n2480 );
nand ( n2491 , n2490 , n2483 );
nand ( n2492 , n2489 , n2491 );
nand ( n2493 , n80 , n96 );
not ( n2494 , n2493 );
not ( n2495 , n2494 );
nand ( n2496 , n79 , n97 );
not ( n2497 , n2496 );
nand ( n2498 , n83 , n93 );
not ( n2499 , n2498 );
not ( n2500 , n2499 );
or ( n2501 , n2497 , n2500 );
or ( n2502 , n2499 , n2496 );
nand ( n2503 , n2501 , n2502 );
not ( n2504 , n2503 );
or ( n2505 , n2495 , n2504 );
not ( n2506 , n2496 );
nand ( n2507 , n2506 , n2499 );
nand ( n2508 , n2505 , n2507 );
xor ( n2509 , n2492 , n2508 );
and ( n2510 , n2476 , n2509 );
and ( n2511 , n2508 , n2492 );
nor ( n2512 , n2510 , n2511 );
not ( n2513 , n2512 );
not ( n2514 , n2513 );
xnor ( n2515 , n2275 , n2283 );
not ( n2516 , n2515 );
not ( n2517 , n2415 );
not ( n2518 , n2517 );
not ( n2519 , n2438 );
or ( n2520 , n2518 , n2519 );
or ( n2521 , n2517 , n2438 );
nand ( n2522 , n2520 , n2521 );
not ( n2523 , n2522 );
or ( n2524 , n2516 , n2523 );
or ( n2525 , n2515 , n2522 );
nand ( n2526 , n2524 , n2525 );
not ( n2527 , n2526 );
or ( n2528 , n2514 , n2527 );
not ( n2529 , n2515 );
nand ( n2530 , n2529 , n2522 );
nand ( n2531 , n2528 , n2530 );
not ( n2532 , n2531 );
not ( n2533 , n2532 );
or ( n2534 , n2470 , n2533 );
not ( n2535 , n2469 );
nand ( n2536 , n2535 , n2531 );
nand ( n2537 , n2534 , n2536 );
and ( n2538 , n2468 , n2537 );
and ( n2539 , n2469 , n2531 );
nor ( n2540 , n2538 , n2539 );
xnor ( n2541 , n2368 , n2454 );
nand ( n2542 , n2540 , n2541 );
not ( n2543 , n2542 );
not ( n2544 , n2512 );
not ( n2545 , n2526 );
or ( n2546 , n2544 , n2545 );
not ( n2547 , n2526 );
nand ( n2548 , n2513 , n2547 );
nand ( n2549 , n2546 , n2548 );
xor ( n2550 , n2383 , n2379 );
not ( n2551 , n2550 );
nand ( n2552 , n79 , n98 );
not ( n2553 , n2552 );
not ( n2554 , n2553 );
nand ( n2555 , n80 , n97 );
not ( n2556 , n2555 );
nand ( n2557 , n81 , n96 );
not ( n2558 , n2557 );
not ( n2559 , n2558 );
or ( n2560 , n2556 , n2559 );
or ( n2561 , n2558 , n2555 );
nand ( n2562 , n2560 , n2561 );
not ( n2563 , n2562 );
or ( n2564 , n2554 , n2563 );
not ( n2565 , n2555 );
nand ( n2566 , n2565 , n2558 );
nand ( n2567 , n2564 , n2566 );
not ( n2568 , n2567 );
nand ( n2569 , n78 , n99 );
not ( n2570 , n2569 );
nand ( n2571 , n14 , n2570 );
not ( n2572 , n2571 );
xor ( n2573 , n13 , n2378 );
not ( n2574 , n2573 );
or ( n2575 , n2572 , n2574 );
or ( n2576 , n2571 , n2573 );
nand ( n2577 , n2575 , n2576 );
not ( n2578 , n2577 );
or ( n2579 , n2568 , n2578 );
not ( n2580 , n2571 );
nand ( n2581 , n2580 , n2573 );
nand ( n2582 , n2579 , n2581 );
not ( n2583 , n2582 );
not ( n2584 , n2405 );
and ( n2585 , n2412 , n2584 );
not ( n2586 , n2412 );
and ( n2587 , n2586 , n2405 );
nor ( n2588 , n2585 , n2587 );
and ( n2589 , n2583 , n2588 );
not ( n2590 , n2583 );
not ( n2591 , n2588 );
and ( n2592 , n2590 , n2591 );
nor ( n2593 , n2589 , n2592 );
not ( n2594 , n2593 );
or ( n2595 , n2551 , n2594 );
nand ( n2596 , n2591 , n2582 );
nand ( n2597 , n2595 , n2596 );
and ( n2598 , n2400 , n2385 );
not ( n2599 , n2400 );
not ( n2600 , n2385 );
and ( n2601 , n2599 , n2600 );
nor ( n2602 , n2598 , n2601 );
xor ( n2603 , n2597 , n2602 );
and ( n2604 , n2549 , n2603 );
and ( n2605 , n2602 , n2597 );
nor ( n2606 , n2604 , n2605 );
xor ( n2607 , n2537 , n2468 );
not ( n2608 , n2607 );
nand ( n2609 , n2606 , n2608 );
not ( n2610 , n2609 );
xor ( n2611 , n2549 , n2603 );
not ( n2612 , n2611 );
xor ( n2613 , n2550 , n2593 );
not ( n2614 , n2613 );
and ( n2615 , n83 , n94 );
not ( n2616 , n2615 );
nand ( n2617 , n82 , n95 );
or ( n2618 , n2616 , n2617 );
nand ( n2619 , n79 , n99 );
not ( n2620 , n2619 );
and ( n2621 , n15 , n2620 );
xnor ( n2622 , n2617 , n2615 );
nand ( n2623 , n2621 , n2622 );
nand ( n2624 , n2618 , n2623 );
not ( n2625 , n2624 );
xor ( n2626 , n2493 , n2503 );
not ( n2627 , n2626 );
not ( n2628 , n2627 );
xnor ( n2629 , n2477 , n2487 );
not ( n2630 , n2629 );
not ( n2631 , n2630 );
or ( n2632 , n2628 , n2631 );
nand ( n2633 , n2629 , n2626 );
nand ( n2634 , n2632 , n2633 );
not ( n2635 , n2634 );
or ( n2636 , n2625 , n2635 );
nand ( n2637 , n2627 , n2629 );
nand ( n2638 , n2636 , n2637 );
not ( n2639 , n2638 );
not ( n2640 , n2639 );
not ( n2641 , n2475 );
not ( n2642 , n2509 );
and ( n2643 , n2641 , n2642 );
and ( n2644 , n2475 , n2509 );
nor ( n2645 , n2643 , n2644 );
not ( n2646 , n2645 );
not ( n2647 , n2646 );
or ( n2648 , n2640 , n2647 );
nand ( n2649 , n2638 , n2645 );
nand ( n2650 , n2648 , n2649 );
not ( n2651 , n2650 );
or ( n2652 , n2614 , n2651 );
or ( n2653 , n2639 , n2645 );
nand ( n2654 , n2652 , n2653 );
not ( n2655 , n2654 );
nand ( n2656 , n2612 , n2655 );
not ( n2657 , n2656 );
xnor ( n2658 , n2634 , n2624 );
not ( n2659 , n2552 );
not ( n2660 , n2562 );
or ( n2661 , n2659 , n2660 );
or ( n2662 , n2552 , n2562 );
nand ( n2663 , n2661 , n2662 );
not ( n2664 , n2663 );
xor ( n2665 , n14 , n2569 );
not ( n2666 , n2665 );
and ( n2667 , n80 , n98 );
not ( n2668 , n2667 );
nand ( n2669 , n81 , n97 );
not ( n2670 , n2669 );
nand ( n2671 , n82 , n96 );
not ( n2672 , n2671 );
not ( n2673 , n2672 );
or ( n2674 , n2670 , n2673 );
not ( n2675 , n2671 );
nand ( n2676 , n81 , n97 );
or ( n2677 , n2675 , n2676 );
nand ( n2678 , n2674 , n2677 );
not ( n2679 , n2678 );
or ( n2680 , n2668 , n2679 );
not ( n2681 , n2676 );
nand ( n2682 , n2675 , n2681 );
nand ( n2683 , n2680 , n2682 );
not ( n2684 , n2683 );
or ( n2685 , n2666 , n2684 );
or ( n2686 , n2665 , n2683 );
nand ( n2687 , n2685 , n2686 );
not ( n2688 , n2687 );
or ( n2689 , n2664 , n2688 );
not ( n2690 , n2665 );
nand ( n2691 , n2690 , n2683 );
nand ( n2692 , n2689 , n2691 );
not ( n2693 , n2692 );
xor ( n2694 , n2567 , n2577 );
not ( n2695 , n2694 );
and ( n2696 , n2693 , n2695 );
not ( n2697 , n2693 );
and ( n2698 , n2697 , n2694 );
nor ( n2699 , n2696 , n2698 );
not ( n2700 , n2699 );
or ( n2701 , n2658 , n2700 );
or ( n2702 , n2695 , n2693 );
nand ( n2703 , n2701 , n2702 );
not ( n2704 , n2703 );
and ( n2705 , n2650 , n2613 );
not ( n2706 , n2650 );
not ( n2707 , n2613 );
and ( n2708 , n2706 , n2707 );
nor ( n2709 , n2705 , n2708 );
not ( n2710 , n2709 );
nand ( n2711 , n2704 , n2710 );
not ( n2712 , n2711 );
xnor ( n2713 , n2622 , n2621 );
not ( n2714 , n2713 );
nand ( n2715 , n81 , n98 );
not ( n2716 , n2715 );
not ( n2717 , n2716 );
nand ( n2718 , n82 , n97 );
not ( n2719 , n2718 );
nand ( n2720 , n83 , n96 );
not ( n2721 , n2720 );
not ( n2722 , n2721 );
or ( n2723 , n2719 , n2722 );
or ( n2724 , n2721 , n2718 );
nand ( n2725 , n2723 , n2724 );
not ( n2726 , n2725 );
or ( n2727 , n2717 , n2726 );
not ( n2728 , n2718 );
nand ( n2729 , n2728 , n2721 );
nand ( n2730 , n2727 , n2729 );
not ( n2731 , n2730 );
nand ( n2732 , n83 , n95 );
xor ( n2733 , n15 , n2620 );
xnor ( n2734 , n2732 , n2733 );
not ( n2735 , n2734 );
or ( n2736 , n2731 , n2735 );
not ( n2737 , n2732 );
nand ( n2738 , n2737 , n2733 );
nand ( n2739 , n2736 , n2738 );
not ( n2740 , n2739 );
or ( n2741 , n2714 , n2740 );
or ( n2742 , n2713 , n2739 );
nand ( n2743 , n2741 , n2742 );
not ( n2744 , n2743 );
not ( n2745 , n2687 );
and ( n2746 , n2663 , n2745 );
not ( n2747 , n2663 );
and ( n2748 , n2747 , n2687 );
nor ( n2749 , n2746 , n2748 );
not ( n2750 , n2749 );
not ( n2751 , n2750 );
or ( n2752 , n2744 , n2751 );
not ( n2753 , n2739 );
or ( n2754 , n2713 , n2753 );
nand ( n2755 , n2752 , n2754 );
and ( n2756 , n2658 , n2699 );
not ( n2757 , n2658 );
and ( n2758 , n2757 , n2700 );
nor ( n2759 , n2756 , n2758 );
not ( n2760 , n2759 );
nand ( n2761 , n2755 , n2760 );
not ( n2762 , n2755 );
nand ( n2763 , n2762 , n2759 );
not ( n2764 , n16 );
nand ( n2765 , n80 , n99 );
and ( n2766 , n2764 , n2765 );
not ( n2767 , n2667 );
not ( n2768 , n2678 );
not ( n2769 , n2768 );
or ( n2770 , n2767 , n2769 );
not ( n2771 , n2667 );
nand ( n2772 , n2771 , n2678 );
nand ( n2773 , n2770 , n2772 );
and ( n2774 , n2766 , n2773 );
not ( n2775 , n2766 );
not ( n2776 , n2773 );
and ( n2777 , n2775 , n2776 );
nor ( n2778 , n2774 , n2777 );
not ( n2779 , n2778 );
not ( n2780 , n2779 );
not ( n2781 , n2730 );
not ( n2782 , n2734 );
not ( n2783 , n2782 );
or ( n2784 , n2781 , n2783 );
or ( n2785 , n2730 , n2782 );
nand ( n2786 , n2784 , n2785 );
not ( n2787 , n2786 );
or ( n2788 , n2780 , n2787 );
or ( n2789 , n2766 , n2776 );
nand ( n2790 , n2788 , n2789 );
not ( n2791 , n2750 );
not ( n2792 , n2743 );
not ( n2793 , n2792 );
or ( n2794 , n2791 , n2793 );
nand ( n2795 , n2743 , n2749 );
nand ( n2796 , n2794 , n2795 );
and ( n2797 , n2790 , n2796 );
not ( n2798 , n2797 );
or ( n2799 , n2790 , n2796 );
xor ( n2800 , n2764 , n2765 );
not ( n2801 , n17 );
nand ( n2802 , n81 , n99 );
nor ( n2803 , n2801 , n2802 );
and ( n2804 , n2800 , n2803 );
not ( n2805 , n2800 );
not ( n2806 , n2803 );
and ( n2807 , n2805 , n2806 );
nor ( n2808 , n2804 , n2807 );
xor ( n2809 , n2715 , n2725 );
or ( n2810 , n2808 , n2809 );
or ( n2811 , n2806 , n2800 );
nand ( n2812 , n2810 , n2811 );
not ( n2813 , n2779 );
not ( n2814 , n2786 );
not ( n2815 , n2814 );
or ( n2816 , n2813 , n2815 );
nand ( n2817 , n2778 , n2786 );
nand ( n2818 , n2816 , n2817 );
nand ( n2819 , n2812 , n2818 );
or ( n2820 , n2812 , n2818 );
xor ( n2821 , n2809 , n2808 );
not ( n2822 , n2821 );
and ( n2823 , n2802 , n2801 );
not ( n2824 , n2802 );
and ( n2825 , n2824 , n17 );
nor ( n2826 , n2823 , n2825 );
not ( n2827 , n2826 );
nand ( n2828 , n83 , n97 );
nand ( n2829 , n82 , n98 );
and ( n2830 , n2828 , n2829 );
not ( n2831 , n2828 );
not ( n2832 , n2829 );
and ( n2833 , n2831 , n2832 );
nor ( n2834 , n2830 , n2833 );
not ( n2835 , n2834 );
or ( n2836 , n2827 , n2835 );
or ( n2837 , n2828 , n2829 );
nand ( n2838 , n2836 , n2837 );
not ( n2839 , n2838 );
nand ( n2840 , n2822 , n2839 );
not ( n2841 , n2840 );
xor ( n2842 , n2834 , n2826 );
not ( n2843 , n2842 );
and ( n2844 , n83 , n98 );
xor ( n2845 , n18 , n2844 );
not ( n2846 , n2845 );
nand ( n2847 , n83 , n99 );
not ( n2848 , n2847 );
nand ( n2849 , n2848 , n19 );
nand ( n2850 , n82 , n99 );
and ( n2851 , n2849 , n2850 );
not ( n2852 , n2849 );
not ( n2853 , n2850 );
and ( n2854 , n2852 , n2853 );
nor ( n2855 , n2851 , n2854 );
not ( n2856 , n2855 );
or ( n2857 , n2846 , n2856 );
not ( n2858 , n2849 );
nand ( n2859 , n2853 , n2858 );
nand ( n2860 , n2857 , n2859 );
and ( n2861 , n18 , n2844 );
and ( n2862 , n2860 , n2861 );
not ( n2863 , n2860 );
not ( n2864 , n2861 );
and ( n2865 , n2863 , n2864 );
nor ( n2866 , n2862 , n2865 );
not ( n2867 , n2866 );
or ( n2868 , n2843 , n2867 );
nand ( n2869 , n2861 , n2860 );
nand ( n2870 , n2868 , n2869 );
not ( n2871 , n2870 );
or ( n2872 , n2841 , n2871 );
nand ( n2873 , n2838 , n2821 );
nand ( n2874 , n2872 , n2873 );
nand ( n2875 , n2820 , n2874 );
nand ( n2876 , n2819 , n2875 );
nand ( n2877 , n2799 , n2876 );
nand ( n2878 , n2798 , n2877 );
nand ( n2879 , n2763 , n2878 );
nand ( n2880 , n2761 , n2879 );
not ( n2881 , n2880 );
or ( n2882 , n2712 , n2881 );
nand ( n2883 , n2703 , n2709 );
nand ( n2884 , n2882 , n2883 );
not ( n2885 , n2884 );
or ( n2886 , n2657 , n2885 );
nand ( n2887 , n2654 , n2611 );
nand ( n2888 , n2886 , n2887 );
not ( n2889 , n2888 );
or ( n2890 , n2610 , n2889 );
not ( n2891 , n2606 );
nand ( n2892 , n2891 , n2607 );
nand ( n2893 , n2890 , n2892 );
not ( n2894 , n2893 );
or ( n2895 , n2543 , n2894 );
not ( n2896 , n2540 );
not ( n2897 , n2541 );
nand ( n2898 , n2896 , n2897 );
nand ( n2899 , n2895 , n2898 );
not ( n2900 , n2899 );
or ( n2901 , n2462 , n2900 );
not ( n2902 , n2458 );
nand ( n2903 , n2902 , n2459 );
nand ( n2904 , n2901 , n2903 );
not ( n2905 , n2904 );
or ( n2906 , n2364 , n2905 );
not ( n2907 , n2348 );
not ( n2908 , n2362 );
nand ( n2909 , n2907 , n2908 );
nand ( n2910 , n2906 , n2909 );
not ( n2911 , n2910 );
not ( n2912 , n2067 );
and ( n2913 , n2912 , n2063 );
not ( n2914 , n2912 );
not ( n2915 , n2063 );
and ( n2916 , n2914 , n2915 );
nor ( n2917 , n2913 , n2916 );
or ( n2918 , n2350 , n2361 );
or ( n2919 , n2359 , n2355 );
nand ( n2920 , n2918 , n2919 );
xnor ( n2921 , n2917 , n2920 );
not ( n2922 , n2921 );
or ( n2923 , n2911 , n2922 );
not ( n2924 , n2917 );
nand ( n2925 , n2920 , n2924 );
nand ( n2926 , n2923 , n2925 );
nand ( n2927 , n2217 , n2926 );
nor ( n2928 , n2927 , n2154 );
nand ( n2929 , n2214 , n2928 , n1405 );
nand ( n2930 , n2213 , n2929 );
and ( n2931 , n843 , n1304 , n2930 );
nand ( n2932 , n667 , n2931 );
not ( n2933 , n843 );
nand ( n2934 , n1285 , n1295 );
or ( n2935 , n2934 , n1303 );
nand ( n2936 , n1299 , n1302 );
nand ( n2937 , n2935 , n2936 );
not ( n2938 , n2937 );
or ( n2939 , n2933 , n2938 );
not ( n2940 , n668 );
nand ( n2941 , n2940 , n841 );
nand ( n2942 , n2939 , n2941 );
and ( n2943 , n2942 , n667 );
nor ( n2944 , n581 , n666 );
nor ( n2945 , n2943 , n2944 );
nand ( n2946 , n2932 , n2945 );
buf ( n2947 , n2946 );
or ( n2948 , n523 , n526 );
or ( n2949 , n524 , n525 );
nand ( n2950 , n2948 , n2949 );
nand ( n2951 , n74 , n84 );
not ( n2952 , n2951 );
or ( n2953 , n551 , n550 );
or ( n2954 , n548 , n549 );
nand ( n2955 , n2953 , n2954 );
not ( n2956 , n2955 );
or ( n2957 , n2952 , n2956 );
or ( n2958 , n2951 , n2955 );
nand ( n2959 , n2957 , n2958 );
xnor ( n2960 , n2950 , n2959 );
and ( n2961 , n552 , n559 );
and ( n2962 , n555 , n558 );
nor ( n2963 , n2961 , n2962 );
xor ( n2964 , n2960 , n2963 );
or ( n2965 , n541 , n528 );
or ( n2966 , n527 , n522 );
nand ( n2967 , n2965 , n2966 );
xor ( n2968 , n2964 , n2967 );
nand ( n2969 , n71 , n87 );
nand ( n2970 , n69 , n89 );
nand ( n2971 , n68 , n90 );
xnor ( n2972 , n2970 , n2971 );
xnor ( n2973 , n2969 , n2972 );
nand ( n2974 , n73 , n85 );
nand ( n2975 , n72 , n86 );
nand ( n2976 , n70 , n88 );
xnor ( n2977 , n2975 , n2976 );
xnor ( n2978 , n2974 , n2977 );
xnor ( n2979 , n2973 , n2978 );
and ( n2980 , n521 , n518 );
and ( n2981 , n520 , n519 );
nor ( n2982 , n2980 , n2981 );
xor ( n2983 , n2979 , n2982 );
xor ( n2984 , n2968 , n2983 );
or ( n2985 , n561 , n578 );
or ( n2986 , n547 , n560 );
nand ( n2987 , n2985 , n2986 );
xor ( n2988 , n2984 , n2987 );
not ( n2989 , n2988 );
or ( n2990 , n514 , n580 );
or ( n2991 , n542 , n579 );
nand ( n2992 , n2990 , n2991 );
not ( n2993 , n2992 );
nand ( n2994 , n2989 , n2993 );
not ( n2995 , n2994 );
xor ( n2996 , n303 , n300 );
or ( n2997 , n2974 , n2977 );
or ( n2998 , n2975 , n2976 );
nand ( n2999 , n2997 , n2998 );
or ( n3000 , n2969 , n2972 );
or ( n3001 , n2970 , n2971 );
nand ( n3002 , n3000 , n3001 );
xor ( n3003 , n2999 , n3002 );
xnor ( n3004 , n2996 , n3003 );
xnor ( n3005 , n286 , n289 );
and ( n3006 , n2950 , n2959 );
not ( n3007 , n2951 );
and ( n3008 , n3007 , n2955 );
nor ( n3009 , n3006 , n3008 );
xnor ( n3010 , n3005 , n3009 );
or ( n3011 , n3004 , n3010 );
or ( n3012 , n3005 , n3009 );
nand ( n3013 , n3011 , n3012 );
xnor ( n3014 , n298 , n307 );
and ( n3015 , n2996 , n3003 );
and ( n3016 , n2999 , n3002 );
nor ( n3017 , n3015 , n3016 );
xor ( n3018 , n3014 , n3017 );
xnor ( n3019 , n3013 , n3018 );
not ( n3020 , n2967 );
not ( n3021 , n2964 );
or ( n3022 , n3020 , n3021 );
or ( n3023 , n2960 , n2963 );
nand ( n3024 , n3022 , n3023 );
xor ( n3025 , n3010 , n3004 );
or ( n3026 , n2982 , n2979 );
or ( n3027 , n2978 , n2973 );
nand ( n3028 , n3026 , n3027 );
xor ( n3029 , n3025 , n3028 );
and ( n3030 , n3024 , n3029 );
and ( n3031 , n3028 , n3025 );
nor ( n3032 , n3030 , n3031 );
nand ( n3033 , n3019 , n3032 );
xnor ( n3034 , n3029 , n3024 );
and ( n3035 , n2987 , n2984 );
and ( n3036 , n2983 , n2968 );
nor ( n3037 , n3035 , n3036 );
nand ( n3038 , n3034 , n3037 );
nand ( n3039 , n3033 , n3038 );
nor ( n3040 , n2995 , n3039 );
nand ( n3041 , n2947 , n3040 );
not ( n3042 , n3041 );
xor ( n3043 , n315 , n310 );
not ( n3044 , n3013 );
not ( n3045 , n3018 );
or ( n3046 , n3044 , n3045 );
or ( n3047 , n3017 , n3014 );
nand ( n3048 , n3046 , n3047 );
nor ( n3049 , n3043 , n3048 );
not ( n3050 , n3049 );
nand ( n3051 , n320 , n3042 , n3050 );
not ( n3052 , n281 );
nand ( n3053 , n285 , n318 );
not ( n3054 , n3053 );
and ( n3055 , n3052 , n3054 );
not ( n3056 , n251 );
nor ( n3057 , n3056 , n279 );
nor ( n3058 , n3055 , n3057 );
nand ( n3059 , n3043 , n3048 );
not ( n3060 , n3059 );
nand ( n3061 , n2988 , n2992 );
or ( n3062 , n3039 , n3061 );
nor ( n3063 , n3034 , n3037 );
and ( n3064 , n3033 , n3063 );
nor ( n3065 , n3019 , n3032 );
nor ( n3066 , n3064 , n3065 );
nand ( n3067 , n3062 , n3066 );
nand ( n3068 , n3050 , n3067 );
not ( n3069 , n3068 );
or ( n3070 , n3060 , n3069 );
nand ( n3071 , n3070 , n320 );
nand ( n3072 , n3051 , n3058 , n3071 );
nand ( n3073 , n68 , n84 );
and ( n3074 , n250 , n245 );
and ( n3075 , n249 , n246 );
nor ( n3076 , n3074 , n3075 );
or ( n3077 , n3073 , n3076 );
nand ( n3078 , n3073 , n3076 );
nand ( n3079 , n3077 , n3078 );
not ( n3080 , n3079 );
and ( n3081 , n3072 , n3080 );
not ( n3082 , n3072 );
and ( n3083 , n3082 , n3079 );
nor ( n3084 , n3081 , n3083 );
not ( n3085 , n3084 );
or ( n3086 , n238 , n3085 );
xor ( n3087 , n39 , n40 );
not ( n3088 , n3087 );
xor ( n3089 , n38 , n39 );
and ( n3090 , n3088 , n3089 );
buf ( n3091 , n3090 );
buf ( n3092 , n3091 );
not ( n3093 , n3092 );
not ( n3094 , n3093 );
not ( n3095 , n3094 );
not ( n3096 , n38 );
and ( n3097 , n3 , n4 );
not ( n3098 , n3 );
and ( n3099 , n3098 , n20 );
nor ( n3100 , n3097 , n3099 );
not ( n3101 , n3100 );
buf ( n3102 , n3101 );
buf ( n3103 , n3102 );
not ( n3104 , n3103 );
nand ( n3105 , n3096 , n3104 );
buf ( n3106 , n3102 );
nand ( n3107 , n38 , n3106 );
and ( n3108 , n3105 , n3107 );
not ( n3109 , n3108 );
or ( n3110 , n3095 , n3109 );
buf ( n3111 , n3087 );
buf ( n3112 , n3111 );
buf ( n3113 , n3112 );
not ( n3114 , n3113 );
not ( n3115 , n3114 );
nand ( n3116 , n38 , n3115 );
nand ( n3117 , n3110 , n3116 );
nand ( n3118 , n36 , n37 );
nor ( n3119 , n36 , n37 );
not ( n3120 , n3119 );
xor ( n3121 , n37 , n38 );
not ( n3122 , n3121 );
and ( n3123 , n3118 , n3120 , n3122 );
buf ( n3124 , n3123 );
not ( n3125 , n3124 );
not ( n3126 , n36 );
and ( n3127 , n3 , n6 );
not ( n3128 , n3 );
and ( n3129 , n3128 , n22 );
nor ( n3130 , n3127 , n3129 );
not ( n3131 , n3130 );
buf ( n3132 , n3131 );
not ( n3133 , n3132 );
not ( n3134 , n3133 );
not ( n3135 , n3134 );
not ( n3136 , n3135 );
and ( n3137 , n3126 , n3136 );
and ( n3138 , n36 , n3135 );
nor ( n3139 , n3137 , n3138 );
or ( n3140 , n3125 , n3139 );
not ( n3141 , n3122 );
buf ( n3142 , n3141 );
not ( n3143 , n3142 );
not ( n3144 , n3143 );
not ( n3145 , n3144 );
not ( n3146 , n3145 );
not ( n3147 , n3146 );
not ( n3148 , n3147 );
not ( n3149 , n3148 );
and ( n3150 , n3 , n5 );
not ( n3151 , n3 );
and ( n3152 , n3151 , n21 );
nor ( n3153 , n3150 , n3152 );
buf ( n3154 , n3153 );
not ( n3155 , n3154 );
not ( n3156 , n3155 );
not ( n3157 , n3156 );
not ( n3158 , n3157 );
buf ( n3159 , n3158 );
not ( n3160 , n3159 );
or ( n3161 , n36 , n3160 );
or ( n3162 , n3126 , n3159 );
nand ( n3163 , n3161 , n3162 );
or ( n3164 , n3149 , n3163 );
nand ( n3165 , n3140 , n3164 );
not ( n3166 , n7 );
and ( n3167 , n3 , n3166 );
not ( n3168 , n3 );
not ( n3169 , n23 );
and ( n3170 , n3168 , n3169 );
nor ( n3171 , n3167 , n3170 );
buf ( n3172 , n3171 );
not ( n3173 , n3172 );
not ( n3174 , n3173 );
and ( n3175 , n36 , n3174 );
not ( n3176 , n3175 );
not ( n3177 , n3117 );
or ( n3178 , n3176 , n3177 );
or ( n3179 , n3175 , n3117 );
nand ( n3180 , n3178 , n3179 );
and ( n3181 , n3165 , n3180 );
not ( n3182 , n3117 );
and ( n3183 , n3175 , n3182 );
nor ( n3184 , n3181 , n3183 );
and ( n3185 , n3117 , n3184 );
nor ( n3186 , n3117 , n3184 );
nor ( n3187 , n3185 , n3186 );
not ( n3188 , n3125 );
not ( n3189 , n3163 );
and ( n3190 , n3188 , n3189 );
not ( n3191 , n3149 );
not ( n3192 , n3102 );
not ( n3193 , n3192 );
not ( n3194 , n3193 );
not ( n3195 , n3194 );
not ( n3196 , n3195 );
not ( n3197 , n3196 );
not ( n3198 , n3197 );
and ( n3199 , n3126 , n3198 );
and ( n3200 , n36 , n3197 );
nor ( n3201 , n3199 , n3200 );
and ( n3202 , n3191 , n3201 );
nor ( n3203 , n3190 , n3202 );
not ( n3204 , n3136 );
not ( n3205 , n3204 );
not ( n3206 , n3205 );
not ( n3207 , n3206 );
nand ( n3208 , n36 , n3207 );
buf ( n3209 , n3115 );
buf ( n3210 , n3209 );
not ( n3211 , n3210 );
not ( n3212 , n3094 );
and ( n3213 , n3211 , n3212 );
nor ( n3214 , n3213 , n3096 );
xnor ( n3215 , n3208 , n3214 );
xnor ( n3216 , n3203 , n3215 );
xor ( n3217 , n3187 , n3216 );
xor ( n3218 , n40 , n41 );
not ( n3219 , n3218 );
xor ( n3220 , n41 , n42 );
nor ( n3221 , n3219 , n3220 );
buf ( n3222 , n3221 );
not ( n3223 , n3222 );
not ( n3224 , n3223 );
buf ( n3225 , n3224 );
not ( n3226 , n40 );
not ( n3227 , n3192 );
or ( n3228 , n3226 , n3227 );
not ( n3229 , n40 );
nand ( n3230 , n3229 , n3106 );
nand ( n3231 , n3228 , n3230 );
and ( n3232 , n3225 , n3231 );
xor ( n3233 , n41 , n42 );
buf ( n3234 , n3233 );
buf ( n3235 , n3234 );
buf ( n3236 , n3235 );
not ( n3237 , n3236 );
not ( n3238 , n3237 );
and ( n3239 , n3238 , n40 );
nor ( n3240 , n3232 , n3239 );
not ( n3241 , n3240 );
xor ( n3242 , n36 , n3174 );
not ( n3243 , n3242 );
or ( n3244 , n3125 , n3243 );
not ( n3245 , n3148 );
or ( n3246 , n3245 , n3139 );
nand ( n3247 , n3244 , n3246 );
and ( n3248 , n3241 , n3247 );
and ( n3249 , n3247 , n3241 );
not ( n3250 , n3247 );
and ( n3251 , n3250 , n3240 );
nor ( n3252 , n3249 , n3251 );
and ( n3253 , n3 , n9 );
not ( n3254 , n3 );
and ( n3255 , n3254 , n25 );
nor ( n3256 , n3253 , n3255 );
not ( n3257 , n3256 );
buf ( n3258 , n3257 );
not ( n3259 , n3258 );
not ( n3260 , n3259 );
nand ( n3261 , n36 , n3260 );
not ( n3262 , n3261 );
not ( n3263 , n3262 );
not ( n3264 , n3124 );
and ( n3265 , n3 , n8 );
not ( n3266 , n3 );
and ( n3267 , n3266 , n24 );
nor ( n3268 , n3265 , n3267 );
not ( n3269 , n3268 );
buf ( n3270 , n3269 );
buf ( n3271 , n3270 );
buf ( n3272 , n3271 );
and ( n3273 , n36 , n3272 );
not ( n3274 , n36 );
not ( n3275 , n3271 );
and ( n3276 , n3274 , n3275 );
nor ( n3277 , n3273 , n3276 );
not ( n3278 , n3277 );
or ( n3279 , n3264 , n3278 );
not ( n3280 , n3143 );
nand ( n3281 , n3280 , n3242 );
nand ( n3282 , n3279 , n3281 );
not ( n3283 , n3282 );
or ( n3284 , n3263 , n3283 );
and ( n3285 , n3096 , n3134 );
buf ( n3286 , n3132 );
not ( n3287 , n3286 );
and ( n3288 , n3287 , n38 );
nor ( n3289 , n3285 , n3288 );
buf ( n3290 , n3289 );
or ( n3291 , n3093 , n3290 );
not ( n3292 , n3157 );
not ( n3293 , n3292 );
and ( n3294 , n3096 , n3293 );
and ( n3295 , n38 , n3158 );
nor ( n3296 , n3294 , n3295 );
or ( n3297 , n3114 , n3296 );
nand ( n3298 , n3291 , n3297 );
and ( n3299 , n3282 , n3261 );
not ( n3300 , n3282 );
and ( n3301 , n3300 , n3262 );
nor ( n3302 , n3299 , n3301 );
not ( n3303 , n3302 );
nand ( n3304 , n3298 , n3303 );
nand ( n3305 , n3284 , n3304 );
and ( n3306 , n3252 , n3305 );
nor ( n3307 , n3248 , n3306 );
not ( n3308 , n3209 );
not ( n3309 , n3108 );
or ( n3310 , n3308 , n3309 );
or ( n3311 , n3212 , n3296 );
nand ( n3312 , n3310 , n3311 );
not ( n3313 , n3275 );
not ( n3314 , n3313 );
not ( n3315 , n3314 );
and ( n3316 , n36 , n3315 );
buf ( n3317 , n3235 );
not ( n3318 , n3317 );
not ( n3319 , n3318 );
not ( n3320 , n3225 );
not ( n3321 , n3320 );
or ( n3322 , n3319 , n3321 );
nand ( n3323 , n3322 , n40 );
xor ( n3324 , n3316 , n3323 );
and ( n3325 , n3312 , n3324 );
and ( n3326 , n3316 , n3323 );
nor ( n3327 , n3325 , n3326 );
xnor ( n3328 , n3165 , n3180 );
xnor ( n3329 , n3327 , n3328 );
or ( n3330 , n3307 , n3329 );
or ( n3331 , n3327 , n3328 );
nand ( n3332 , n3330 , n3331 );
nand ( n3333 , n3217 , n3332 );
not ( n3334 , n3217 );
not ( n3335 , n3332 );
nand ( n3336 , n3334 , n3335 );
nand ( n3337 , n3333 , n3336 );
xnor ( n3338 , n3307 , n3329 );
xor ( n3339 , n3312 , n3324 );
xor ( n3340 , n3252 , n3305 );
xor ( n3341 , n3339 , n3340 );
not ( n3342 , n3298 );
not ( n3343 , n3302 );
and ( n3344 , n3342 , n3343 );
and ( n3345 , n3298 , n3302 );
nor ( n3346 , n3344 , n3345 );
xor ( n3347 , n43 , n44 );
buf ( n3348 , n3347 );
buf ( n3349 , n3348 );
buf ( n3350 , n3349 );
not ( n3351 , n3350 );
not ( n3352 , n3351 );
xor ( n3353 , n42 , n43 );
not ( n3354 , n3353 );
xor ( n3355 , n43 , n44 );
nor ( n3356 , n3354 , n3355 );
not ( n3357 , n3356 );
buf ( n3358 , n3357 );
not ( n3359 , n3358 );
or ( n3360 , n3352 , n3359 );
nand ( n3361 , n3360 , n42 );
not ( n3362 , n3280 );
not ( n3363 , n3277 );
or ( n3364 , n3362 , n3363 );
not ( n3365 , n3126 );
not ( n3366 , n3258 );
or ( n3367 , n3365 , n3366 );
buf ( n3368 , n3256 );
not ( n3369 , n3368 );
or ( n3370 , n3126 , n3369 );
nand ( n3371 , n3367 , n3370 );
nand ( n3372 , n3124 , n3371 );
nand ( n3373 , n3364 , n3372 );
nand ( n3374 , n3361 , n3373 );
not ( n3375 , n40 );
not ( n3376 , n3156 );
or ( n3377 , n3375 , n3376 );
not ( n3378 , n3155 );
or ( n3379 , n40 , n3378 );
nand ( n3380 , n3377 , n3379 );
not ( n3381 , n3380 );
or ( n3382 , n3320 , n3381 );
not ( n3383 , n3231 );
or ( n3384 , n3383 , n3318 );
nand ( n3385 , n3382 , n3384 );
not ( n3386 , n3361 );
not ( n3387 , n3373 );
not ( n3388 , n3387 );
or ( n3389 , n3386 , n3388 );
not ( n3390 , n3361 );
nand ( n3391 , n3390 , n3373 );
nand ( n3392 , n3389 , n3391 );
nand ( n3393 , n3385 , n3392 );
and ( n3394 , n3374 , n3393 );
and ( n3395 , n3394 , n3240 );
not ( n3396 , n3394 );
and ( n3397 , n3396 , n3241 );
nor ( n3398 , n3395 , n3397 );
or ( n3399 , n3346 , n3398 );
or ( n3400 , n3241 , n3394 );
nand ( n3401 , n3399 , n3400 );
and ( n3402 , n3341 , n3401 );
and ( n3403 , n3339 , n3340 );
nor ( n3404 , n3402 , n3403 );
nor ( n3405 , n3338 , n3404 );
not ( n3406 , n3405 );
not ( n3407 , n3091 );
and ( n3408 , n3 , n12 );
not ( n3409 , n3 );
and ( n3410 , n3409 , n28 );
nor ( n3411 , n3408 , n3410 );
buf ( n3412 , n3411 );
not ( n3413 , n3412 );
buf ( n3414 , n3413 );
not ( n3415 , n3414 );
and ( n3416 , n3415 , n3096 );
not ( n3417 , n3415 );
and ( n3418 , n3417 , n38 );
nor ( n3419 , n3416 , n3418 );
not ( n3420 , n3419 );
or ( n3421 , n3407 , n3420 );
buf ( n3422 , n3112 );
not ( n3423 , n3096 );
not ( n3424 , n11 );
and ( n3425 , n3 , n3424 );
not ( n3426 , n3 );
not ( n3427 , n27 );
and ( n3428 , n3426 , n3427 );
nor ( n3429 , n3425 , n3428 );
not ( n3430 , n3429 );
buf ( n3431 , n3430 );
not ( n3432 , n3431 );
buf ( n3433 , n3432 );
not ( n3434 , n3433 );
or ( n3435 , n3423 , n3434 );
and ( n3436 , n3 , n11 );
not ( n3437 , n3 );
and ( n3438 , n3437 , n27 );
nor ( n3439 , n3436 , n3438 );
nand ( n3440 , n38 , n3439 );
nand ( n3441 , n3435 , n3440 );
nand ( n3442 , n3422 , n3441 );
nand ( n3443 , n3421 , n3442 );
not ( n3444 , n3443 );
xor ( n3445 , n45 , n46 );
not ( n3446 , n3445 );
not ( n3447 , n44 );
not ( n3448 , n45 );
and ( n3449 , n3447 , n3448 );
and ( n3450 , n44 , n45 );
nor ( n3451 , n3449 , n3450 );
and ( n3452 , n3446 , n3451 );
buf ( n3453 , n3452 );
buf ( n3454 , n3453 );
not ( n3455 , n3454 );
xor ( n3456 , n44 , n3132 );
not ( n3457 , n3456 );
or ( n3458 , n3455 , n3457 );
not ( n3459 , n45 );
not ( n3460 , n46 );
or ( n3461 , n3459 , n3460 );
or ( n3462 , n45 , n46 );
nand ( n3463 , n3461 , n3462 );
buf ( n3464 , n3463 );
not ( n3465 , n3464 );
buf ( n3466 , n3465 );
not ( n3467 , n3466 );
not ( n3468 , n3467 );
xor ( n3469 , n44 , n3155 );
nand ( n3470 , n3468 , n3469 );
nand ( n3471 , n3458 , n3470 );
xor ( n3472 , n3444 , n3471 );
not ( n3473 , n3224 );
not ( n3474 , n3229 );
not ( n3475 , n10 );
and ( n3476 , n3 , n3475 );
not ( n3477 , n3 );
not ( n3478 , n26 );
and ( n3479 , n3477 , n3478 );
nor ( n3480 , n3476 , n3479 );
buf ( n3481 , n3480 );
buf ( n3482 , n3481 );
not ( n3483 , n3482 );
or ( n3484 , n3474 , n3483 );
or ( n3485 , n3229 , n3482 );
nand ( n3486 , n3484 , n3485 );
not ( n3487 , n3486 );
or ( n3488 , n3473 , n3487 );
not ( n3489 , n3229 );
not ( n3490 , n3258 );
or ( n3491 , n3489 , n3490 );
or ( n3492 , n3229 , n3369 );
nand ( n3493 , n3491 , n3492 );
nand ( n3494 , n3317 , n3493 );
nand ( n3495 , n3488 , n3494 );
not ( n3496 , n3495 );
xor ( n3497 , n3472 , n3496 );
not ( n3498 , n3358 );
not ( n3499 , n3498 );
and ( n3500 , n3270 , n42 );
not ( n3501 , n3270 );
not ( n3502 , n42 );
and ( n3503 , n3501 , n3502 );
nor ( n3504 , n3500 , n3503 );
not ( n3505 , n3504 );
or ( n3506 , n3499 , n3505 );
not ( n3507 , n3172 );
xnor ( n3508 , n42 , n3507 );
nand ( n3509 , n3350 , n3508 );
nand ( n3510 , n3506 , n3509 );
and ( n3511 , n3 , n15 );
not ( n3512 , n3 );
and ( n3513 , n3512 , n31 );
nor ( n3514 , n3511 , n3513 );
buf ( n3515 , n3514 );
not ( n3516 , n3515 );
not ( n3517 , n3516 );
not ( n3518 , n3517 );
and ( n3519 , n36 , n3518 );
not ( n3520 , n3519 );
buf ( n3521 , n3141 );
not ( n3522 , n3521 );
and ( n3523 , n3 , n13 );
not ( n3524 , n3 );
and ( n3525 , n3524 , n29 );
nor ( n3526 , n3523 , n3525 );
not ( n3527 , n3526 );
not ( n3528 , n3527 );
and ( n3529 , n36 , n3528 );
not ( n3530 , n36 );
buf ( n3531 , n3526 );
not ( n3532 , n3531 );
and ( n3533 , n3530 , n3532 );
or ( n3534 , n3529 , n3533 );
not ( n3535 , n3534 );
or ( n3536 , n3522 , n3535 );
not ( n3537 , n36 );
and ( n3538 , n3 , n14 );
not ( n3539 , n3 );
and ( n3540 , n3539 , n30 );
nor ( n3541 , n3538 , n3540 );
not ( n3542 , n3541 );
buf ( n3543 , n3542 );
not ( n3544 , n3543 );
not ( n3545 , n3544 );
or ( n3546 , n3537 , n3545 );
not ( n3547 , n3543 );
or ( n3548 , n3547 , n36 );
nand ( n3549 , n3546 , n3548 );
nand ( n3550 , n3123 , n3549 );
nand ( n3551 , n3536 , n3550 );
not ( n3552 , n3551 );
not ( n3553 , n3552 );
or ( n3554 , n3520 , n3553 );
not ( n3555 , n3519 );
nand ( n3556 , n3555 , n3551 );
nand ( n3557 , n3554 , n3556 );
xor ( n3558 , n3510 , n3557 );
xor ( n3559 , n3101 , n48 );
not ( n3560 , n3559 );
xor ( n3561 , n48 , n49 );
xor ( n3562 , n49 , n50 );
not ( n3563 , n3562 );
nand ( n3564 , n3561 , n3563 );
buf ( n3565 , n3564 );
not ( n3566 , n3565 );
not ( n3567 , n3566 );
or ( n3568 , n3560 , n3567 );
buf ( n3569 , n3562 );
not ( n3570 , n3569 );
buf ( n3571 , n3570 );
not ( n3572 , n3571 );
nand ( n3573 , n48 , n3572 );
nand ( n3574 , n3568 , n3573 );
not ( n3575 , n3574 );
not ( n3576 , n3575 );
not ( n3577 , n3576 );
not ( n3578 , n3123 );
xor ( n3579 , n36 , n3518 );
not ( n3580 , n3579 );
or ( n3581 , n3578 , n3580 );
not ( n3582 , n3141 );
not ( n3583 , n3582 );
nand ( n3584 , n3583 , n3549 );
nand ( n3585 , n3581 , n3584 );
not ( n3586 , n3585 );
or ( n3587 , n3577 , n3586 );
or ( n3588 , n3576 , n3585 );
not ( n3589 , n3091 );
not ( n3590 , n3096 );
not ( n3591 , n3528 );
and ( n3592 , n3590 , n3591 );
and ( n3593 , n3096 , n3528 );
nor ( n3594 , n3592 , n3593 );
not ( n3595 , n3594 );
or ( n3596 , n3589 , n3595 );
nand ( n3597 , n3422 , n3419 );
nand ( n3598 , n3596 , n3597 );
nand ( n3599 , n3588 , n3598 );
nand ( n3600 , n3587 , n3599 );
not ( n3601 , n3600 );
xnor ( n3602 , n3558 , n3601 );
xor ( n3603 , n3497 , n3602 );
not ( n3604 , n3603 );
nor ( n3605 , n46 , n47 );
not ( n3606 , n3605 );
nand ( n3607 , n46 , n47 );
xor ( n3608 , n47 , n48 );
not ( n3609 , n3608 );
nand ( n3610 , n3606 , n3607 , n3609 );
not ( n3611 , n3610 );
not ( n3612 , n3611 );
not ( n3613 , n3612 );
not ( n3614 , n3613 );
and ( n3615 , n46 , n3100 );
not ( n3616 , n46 );
and ( n3617 , n3 , n4 );
not ( n3618 , n3 );
and ( n3619 , n3618 , n20 );
nor ( n3620 , n3617 , n3619 );
not ( n3621 , n3620 );
and ( n3622 , n3616 , n3621 );
or ( n3623 , n3615 , n3622 );
not ( n3624 , n3623 );
or ( n3625 , n3614 , n3624 );
xor ( n3626 , n47 , n48 );
not ( n3627 , n3626 );
not ( n3628 , n3627 );
not ( n3629 , n3628 );
not ( n3630 , n3629 );
nand ( n3631 , n46 , n3630 );
nand ( n3632 , n3625 , n3631 );
not ( n3633 , n3632 );
buf ( n3634 , n3348 );
not ( n3635 , n3634 );
not ( n3636 , n3504 );
or ( n3637 , n3635 , n3636 );
not ( n3638 , n42 );
not ( n3639 , n3256 );
or ( n3640 , n3638 , n3639 );
or ( n3641 , n42 , n3256 );
nand ( n3642 , n3640 , n3641 );
nand ( n3643 , n3356 , n3642 );
nand ( n3644 , n3637 , n3643 );
not ( n3645 , n3644 );
not ( n3646 , n3561 );
not ( n3647 , n3646 );
not ( n3648 , n3570 );
or ( n3649 , n3647 , n3648 );
nand ( n3650 , n3649 , n48 );
not ( n3651 , n3650 );
not ( n3652 , n3651 );
not ( n3653 , n3628 );
not ( n3654 , n3623 );
or ( n3655 , n3653 , n3654 );
xnor ( n3656 , n3153 , n46 );
nand ( n3657 , n3611 , n3656 );
nand ( n3658 , n3655 , n3657 );
not ( n3659 , n3658 );
or ( n3660 , n3652 , n3659 );
or ( n3661 , n3651 , n3658 );
nand ( n3662 , n3660 , n3661 );
not ( n3663 , n3662 );
or ( n3664 , n3645 , n3663 );
not ( n3665 , n3651 );
not ( n3666 , n3658 );
not ( n3667 , n3666 );
nand ( n3668 , n3665 , n3667 );
nand ( n3669 , n3664 , n3668 );
xor ( n3670 , n3633 , n3669 );
not ( n3671 , n3468 );
not ( n3672 , n3456 );
or ( n3673 , n3671 , n3672 );
buf ( n3674 , n3452 );
buf ( n3675 , n3674 );
not ( n3676 , n44 );
not ( n3677 , n3173 );
or ( n3678 , n3676 , n3677 );
or ( n3679 , n44 , n3173 );
nand ( n3680 , n3678 , n3679 );
nand ( n3681 , n3675 , n3680 );
nand ( n3682 , n3673 , n3681 );
not ( n3683 , n3682 );
not ( n3684 , n16 );
and ( n3685 , n3 , n3684 );
not ( n3686 , n3 );
not ( n3687 , n32 );
and ( n3688 , n3686 , n3687 );
nor ( n3689 , n3685 , n3688 );
buf ( n3690 , n3689 );
not ( n3691 , n3690 );
not ( n3692 , n3691 );
buf ( n3693 , n3692 );
nand ( n3694 , n36 , n3693 );
not ( n3695 , n3694 );
not ( n3696 , n3235 );
not ( n3697 , n3486 );
or ( n3698 , n3696 , n3697 );
not ( n3699 , n3229 );
not ( n3700 , n3432 );
or ( n3701 , n3699 , n3700 );
nand ( n3702 , n40 , n3439 );
nand ( n3703 , n3701 , n3702 );
nand ( n3704 , n3222 , n3703 );
nand ( n3705 , n3698 , n3704 );
not ( n3706 , n3705 );
or ( n3707 , n3695 , n3706 );
or ( n3708 , n3694 , n3705 );
nand ( n3709 , n3707 , n3708 );
not ( n3710 , n3709 );
or ( n3711 , n3683 , n3710 );
not ( n3712 , n3694 );
nand ( n3713 , n3712 , n3705 );
nand ( n3714 , n3711 , n3713 );
not ( n3715 , n3714 );
and ( n3716 , n3670 , n3715 );
not ( n3717 , n3670 );
and ( n3718 , n3717 , n3714 );
nor ( n3719 , n3716 , n3718 );
not ( n3720 , n3719 );
not ( n3721 , n3454 );
xor ( n3722 , n44 , n3271 );
not ( n3723 , n3722 );
or ( n3724 , n3721 , n3723 );
not ( n3725 , n3464 );
not ( n3726 , n3725 );
not ( n3727 , n3726 );
buf ( n3728 , n3727 );
nand ( n3729 , n3728 , n3680 );
nand ( n3730 , n3724 , n3729 );
not ( n3731 , n3730 );
not ( n3732 , n3222 );
xnor ( n3733 , n3229 , n3413 );
not ( n3734 , n3733 );
or ( n3735 , n3732 , n3734 );
buf ( n3736 , n3234 );
nand ( n3737 , n3736 , n3703 );
nand ( n3738 , n3735 , n3737 );
not ( n3739 , n3112 );
not ( n3740 , n3594 );
or ( n3741 , n3739 , n3740 );
not ( n3742 , n38 );
and ( n3743 , n3 , n14 );
not ( n3744 , n3 );
and ( n3745 , n3744 , n30 );
nor ( n3746 , n3743 , n3745 );
not ( n3747 , n3746 );
not ( n3748 , n3747 );
not ( n3749 , n3748 );
or ( n3750 , n3742 , n3749 );
or ( n3751 , n38 , n3748 );
nand ( n3752 , n3750 , n3751 );
nand ( n3753 , n3090 , n3752 );
nand ( n3754 , n3741 , n3753 );
and ( n3755 , n3738 , n3754 );
not ( n3756 , n3738 );
not ( n3757 , n3754 );
and ( n3758 , n3756 , n3757 );
nor ( n3759 , n3755 , n3758 );
not ( n3760 , n3759 );
or ( n3761 , n3731 , n3760 );
not ( n3762 , n3757 );
nand ( n3763 , n3738 , n3762 );
nand ( n3764 , n3761 , n3763 );
not ( n3765 , n3764 );
and ( n3766 , n3 , n17 );
not ( n3767 , n3 );
and ( n3768 , n3767 , n33 );
nor ( n3769 , n3766 , n3768 );
not ( n3770 , n3769 );
not ( n3771 , n3770 );
not ( n3772 , n3771 );
not ( n3773 , n3772 );
not ( n3774 , n3773 );
and ( n3775 , n36 , n3774 );
not ( n3776 , n3775 );
xor ( n3777 , n46 , n3131 );
not ( n3778 , n3777 );
buf ( n3779 , n3611 );
not ( n3780 , n3779 );
or ( n3781 , n3778 , n3780 );
not ( n3782 , n3629 );
nand ( n3783 , n3782 , n3656 );
nand ( n3784 , n3781 , n3783 );
not ( n3785 , n3784 );
or ( n3786 , n3776 , n3785 );
or ( n3787 , n3775 , n3784 );
buf ( n3788 , n3356 );
not ( n3789 , n3788 );
not ( n3790 , n3481 );
xnor ( n3791 , n42 , n3790 );
not ( n3792 , n3791 );
or ( n3793 , n3789 , n3792 );
nand ( n3794 , n3634 , n3642 );
nand ( n3795 , n3793 , n3794 );
nand ( n3796 , n3787 , n3795 );
nand ( n3797 , n3786 , n3796 );
buf ( n3798 , n3797 );
xor ( n3799 , n3650 , n3666 );
xnor ( n3800 , n3799 , n3644 );
and ( n3801 , n3798 , n3800 );
not ( n3802 , n3798 );
not ( n3803 , n3800 );
and ( n3804 , n3802 , n3803 );
nor ( n3805 , n3801 , n3804 );
not ( n3806 , n3805 );
or ( n3807 , n3765 , n3806 );
nand ( n3808 , n3798 , n3800 );
nand ( n3809 , n3807 , n3808 );
not ( n3810 , n3809 );
or ( n3811 , n3720 , n3810 );
or ( n3812 , n3719 , n3809 );
nand ( n3813 , n3811 , n3812 );
not ( n3814 , n3813 );
not ( n3815 , n3814 );
or ( n3816 , n3604 , n3815 );
not ( n3817 , n3603 );
nand ( n3818 , n3817 , n3813 );
nand ( n3819 , n3816 , n3818 );
xor ( n3820 , n3585 , n3598 );
not ( n3821 , n3576 );
xor ( n3822 , n3820 , n3821 );
not ( n3823 , n3822 );
not ( n3824 , n3823 );
not ( n3825 , n3728 );
not ( n3826 , n3722 );
or ( n3827 , n3825 , n3826 );
and ( n3828 , n44 , n3256 );
not ( n3829 , n44 );
and ( n3830 , n3 , n9 );
not ( n3831 , n3 );
and ( n3832 , n3831 , n25 );
nor ( n3833 , n3830 , n3832 );
not ( n3834 , n3833 );
and ( n3835 , n3829 , n3834 );
or ( n3836 , n3828 , n3835 );
nand ( n3837 , n3674 , n3836 );
nand ( n3838 , n3827 , n3837 );
buf ( n3839 , n3838 );
not ( n3840 , n3839 );
not ( n3841 , n3575 );
not ( n3842 , n3521 );
not ( n3843 , n3579 );
or ( n3844 , n3842 , n3843 );
nand ( n3845 , n3120 , n3122 );
not ( n3846 , n3118 );
nor ( n3847 , n3845 , n3846 );
not ( n3848 , n36 );
not ( n3849 , n3691 );
or ( n3850 , n3848 , n3849 );
not ( n3851 , n3690 );
not ( n3852 , n3851 );
nand ( n3853 , n3126 , n3852 );
nand ( n3854 , n3850 , n3853 );
nand ( n3855 , n3847 , n3854 );
nand ( n3856 , n3844 , n3855 );
not ( n3857 , n3856 );
not ( n3858 , n3857 );
or ( n3859 , n3841 , n3858 );
nand ( n3860 , n3574 , n3856 );
nand ( n3861 , n3859 , n3860 );
not ( n3862 , n3861 );
or ( n3863 , n3840 , n3862 );
nand ( n3864 , n3821 , n3856 );
nand ( n3865 , n3863 , n3864 );
xor ( n3866 , n3682 , n3709 );
xor ( n3867 , n3865 , n3866 );
not ( n3868 , n3867 );
or ( n3869 , n3824 , n3868 );
nand ( n3870 , n3865 , n3866 );
nand ( n3871 , n3869 , n3870 );
not ( n3872 , n3871 );
xor ( n3873 , n3775 , n3784 );
buf ( n3874 , n3795 );
xnor ( n3875 , n3873 , n3874 );
not ( n3876 , n3839 );
not ( n3877 , n3876 );
not ( n3878 , n3861 );
or ( n3879 , n3877 , n3878 );
not ( n3880 , n3839 );
or ( n3881 , n3880 , n3861 );
nand ( n3882 , n3879 , n3881 );
xnor ( n3883 , n3875 , n3882 );
not ( n3884 , n3883 );
not ( n3885 , n3357 );
not ( n3886 , n3885 );
not ( n3887 , n3412 );
and ( n3888 , n3887 , n42 );
not ( n3889 , n3887 );
and ( n3890 , n3889 , n3502 );
nor ( n3891 , n3888 , n3890 );
not ( n3892 , n3891 );
or ( n3893 , n3886 , n3892 );
buf ( n3894 , n3348 );
not ( n3895 , n3502 );
not ( n3896 , n3430 );
not ( n3897 , n3896 );
or ( n3898 , n3895 , n3897 );
not ( n3899 , n3431 );
or ( n3900 , n3502 , n3899 );
nand ( n3901 , n3898 , n3900 );
nand ( n3902 , n3894 , n3901 );
nand ( n3903 , n3893 , n3902 );
not ( n3904 , n3453 );
not ( n3905 , n44 );
not ( n3906 , n3481 );
not ( n3907 , n3906 );
or ( n3908 , n3905 , n3907 );
not ( n3909 , n44 );
nand ( n3910 , n3909 , n3481 );
nand ( n3911 , n3908 , n3910 );
not ( n3912 , n3911 );
or ( n3913 , n3904 , n3912 );
not ( n3914 , n3446 );
nand ( n3915 , n3914 , n3836 );
nand ( n3916 , n3913 , n3915 );
xor ( n3917 , n3903 , n3916 );
not ( n3918 , n3917 );
not ( n3919 , n3142 );
not ( n3920 , n36 );
not ( n3921 , n3772 );
not ( n3922 , n3921 );
or ( n3923 , n3920 , n3922 );
or ( n3924 , n36 , n3921 );
nand ( n3925 , n3923 , n3924 );
not ( n3926 , n3925 );
or ( n3927 , n3919 , n3926 );
and ( n3928 , n3 , n18 );
not ( n3929 , n3 );
and ( n3930 , n3929 , n34 );
nor ( n3931 , n3928 , n3930 );
not ( n3932 , n3931 );
not ( n3933 , n3932 );
and ( n3934 , n3126 , n3933 );
not ( n3935 , n3126 );
not ( n3936 , n3931 );
and ( n3937 , n3935 , n3936 );
nor ( n3938 , n3934 , n3937 );
nand ( n3939 , n3123 , n3938 );
nand ( n3940 , n3927 , n3939 );
not ( n3941 , n3940 );
not ( n3942 , n3941 );
not ( n3943 , n3942 );
or ( n3944 , n3918 , n3943 );
nand ( n3945 , n3903 , n3916 );
nand ( n3946 , n3944 , n3945 );
not ( n3947 , n3946 );
nand ( n3948 , n3229 , n3542 );
not ( n3949 , n3747 );
nand ( n3950 , n40 , n3949 );
nand ( n3951 , n3948 , n3950 );
not ( n3952 , n3951 );
not ( n3953 , n3222 );
or ( n3954 , n3952 , n3953 );
not ( n3955 , n40 );
not ( n3956 , n3528 );
or ( n3957 , n3955 , n3956 );
or ( n3958 , n40 , n3528 );
nand ( n3959 , n3957 , n3958 );
nand ( n3960 , n3234 , n3959 );
nand ( n3961 , n3954 , n3960 );
not ( n3962 , n3961 );
not ( n3963 , n3089 );
nor ( n3964 , n3111 , n3963 );
not ( n3965 , n3964 );
and ( n3966 , n3690 , n38 );
not ( n3967 , n3690 );
and ( n3968 , n3967 , n3096 );
nor ( n3969 , n3966 , n3968 );
not ( n3970 , n3969 );
or ( n3971 , n3965 , n3970 );
buf ( n3972 , n3087 );
not ( n3973 , n3972 );
not ( n3974 , n3973 );
and ( n3975 , n3515 , n3096 );
not ( n3976 , n3515 );
and ( n3977 , n3976 , n38 );
nor ( n3978 , n3975 , n3977 );
nand ( n3979 , n3974 , n3978 );
nand ( n3980 , n3971 , n3979 );
not ( n3981 , n3605 );
nand ( n3982 , n3609 , n3981 , n3607 );
not ( n3983 , n3982 );
not ( n3984 , n3983 );
and ( n3985 , n3 , n8 );
not ( n3986 , n3 );
and ( n3987 , n3986 , n24 );
or ( n3988 , n3985 , n3987 );
and ( n3989 , n46 , n3988 );
not ( n3990 , n46 );
and ( n3991 , n3990 , n3268 );
or ( n3992 , n3989 , n3991 );
not ( n3993 , n3992 );
not ( n3994 , n3993 );
or ( n3995 , n3984 , n3994 );
not ( n3996 , n3627 );
not ( n3997 , n7 );
and ( n3998 , n3 , n3997 );
not ( n3999 , n3 );
not ( n4000 , n23 );
and ( n4001 , n3999 , n4000 );
nor ( n4002 , n3998 , n4001 );
xor ( n4003 , n46 , n4002 );
nand ( n4004 , n3996 , n4003 );
nand ( n4005 , n3995 , n4004 );
and ( n4006 , n3980 , n4005 );
not ( n4007 , n3980 );
not ( n4008 , n4005 );
and ( n4009 , n4007 , n4008 );
nor ( n4010 , n4006 , n4009 );
not ( n4011 , n4010 );
or ( n4012 , n3962 , n4011 );
not ( n4013 , n4008 );
nand ( n4014 , n4013 , n3980 );
nand ( n4015 , n4012 , n4014 );
not ( n4016 , n3565 );
buf ( n4017 , n4016 );
not ( n4018 , n4017 );
xor ( n4019 , n48 , n3131 );
not ( n4020 , n4019 );
or ( n4021 , n4018 , n4020 );
buf ( n4022 , n3569 );
buf ( n4023 , n4022 );
not ( n4024 , n3154 );
xor ( n4025 , n48 , n4024 );
nand ( n4026 , n4023 , n4025 );
nand ( n4027 , n4021 , n4026 );
not ( n4028 , n4027 );
not ( n4029 , n51 );
nand ( n4030 , n50 , n4029 );
buf ( n4031 , n4030 );
not ( n4032 , n4031 );
not ( n4033 , n4032 );
not ( n4034 , n50 );
not ( n4035 , n4034 );
not ( n4036 , n3621 );
or ( n4037 , n4035 , n4036 );
nand ( n4038 , n50 , n3620 );
nand ( n4039 , n4037 , n4038 );
not ( n4040 , n4039 );
or ( n4041 , n4033 , n4040 );
nand ( n4042 , n50 , n51 );
nand ( n4043 , n4041 , n4042 );
not ( n4044 , n4043 );
not ( n4045 , n35 );
or ( n4046 , n4045 , n3 );
not ( n4047 , n35 );
or ( n4048 , n4047 , n19 );
nand ( n4049 , n4048 , n3 );
nand ( n4050 , n4046 , n4049 );
buf ( n4051 , n4050 );
not ( n4052 , n4051 );
not ( n4053 , n4052 );
nand ( n4054 , n4053 , n36 );
not ( n4055 , n4054 );
or ( n4056 , n4044 , n4055 );
or ( n4057 , n4054 , n4043 );
nand ( n4058 , n4056 , n4057 );
not ( n4059 , n4058 );
or ( n4060 , n4028 , n4059 );
not ( n4061 , n4054 );
nand ( n4062 , n4061 , n4043 );
nand ( n4063 , n4060 , n4062 );
not ( n4064 , n4063 );
and ( n4065 , n4015 , n4064 );
not ( n4066 , n4015 );
and ( n4067 , n4066 , n4063 );
or ( n4068 , n4065 , n4067 );
not ( n4069 , n4068 );
or ( n4070 , n3947 , n4069 );
nand ( n4071 , n4063 , n4015 );
nand ( n4072 , n4070 , n4071 );
not ( n4073 , n4072 );
or ( n4074 , n3884 , n4073 );
not ( n4075 , n3875 );
nand ( n4076 , n4075 , n3882 );
nand ( n4077 , n4074 , n4076 );
not ( n4078 , n4077 );
not ( n4079 , n3349 );
not ( n4080 , n3791 );
or ( n4081 , n4079 , n4080 );
buf ( n4082 , n3356 );
nand ( n4083 , n4082 , n3901 );
nand ( n4084 , n4081 , n4083 );
not ( n4085 , n4084 );
not ( n4086 , n3782 );
not ( n4087 , n3777 );
or ( n4088 , n4086 , n4087 );
nand ( n4089 , n3779 , n4003 );
nand ( n4090 , n4088 , n4089 );
not ( n4091 , n4090 );
or ( n4092 , n4085 , n4091 );
or ( n4093 , n4084 , n4090 );
not ( n4094 , n4025 );
not ( n4095 , n3566 );
or ( n4096 , n4094 , n4095 );
nand ( n4097 , n4023 , n3559 );
nand ( n4098 , n4096 , n4097 );
nand ( n4099 , n4093 , n4098 );
nand ( n4100 , n4092 , n4099 );
not ( n4101 , n3933 );
nand ( n4102 , n36 , n4101 );
nand ( n4103 , n50 , n4102 );
not ( n4104 , n4103 );
not ( n4105 , n3521 );
not ( n4106 , n3854 );
or ( n4107 , n4105 , n4106 );
nand ( n4108 , n3847 , n3925 );
nand ( n4109 , n4107 , n4108 );
not ( n4110 , n4109 );
or ( n4111 , n4104 , n4110 );
not ( n4112 , n50 );
not ( n4113 , n4102 );
nand ( n4114 , n4112 , n4113 );
nand ( n4115 , n4111 , n4114 );
and ( n4116 , n4100 , n4115 );
not ( n4117 , n4100 );
not ( n4118 , n4115 );
and ( n4119 , n4117 , n4118 );
nor ( n4120 , n4116 , n4119 );
not ( n4121 , n4120 );
not ( n4122 , n3730 );
not ( n4123 , n4122 );
not ( n4124 , n3759 );
and ( n4125 , n4123 , n4124 );
and ( n4126 , n4122 , n3759 );
nor ( n4127 , n4125 , n4126 );
not ( n4128 , n4127 );
not ( n4129 , n4128 );
or ( n4130 , n4121 , n4129 );
not ( n4131 , n4118 );
nand ( n4132 , n4131 , n4100 );
nand ( n4133 , n4130 , n4132 );
not ( n4134 , n4133 );
not ( n4135 , n4134 );
xor ( n4136 , n3797 , n3800 );
xnor ( n4137 , n4136 , n3764 );
not ( n4138 , n4137 );
not ( n4139 , n4138 );
or ( n4140 , n4135 , n4139 );
nand ( n4141 , n4133 , n4137 );
nand ( n4142 , n4140 , n4141 );
not ( n4143 , n4142 );
or ( n4144 , n4078 , n4143 );
not ( n4145 , n4134 );
not ( n4146 , n4137 );
nand ( n4147 , n4145 , n4146 );
nand ( n4148 , n4144 , n4147 );
not ( n4149 , n4148 );
not ( n4150 , n4149 );
or ( n4151 , n3872 , n4150 );
not ( n4152 , n3871 );
nand ( n4153 , n4152 , n4148 );
nand ( n4154 , n4151 , n4153 );
xnor ( n4155 , n3819 , n4154 );
xor ( n4156 , n4142 , n4077 );
not ( n4157 , n4156 );
not ( n4158 , n3865 );
xor ( n4159 , n3866 , n4158 );
xnor ( n4160 , n4159 , n3822 );
not ( n4161 , n46 );
not ( n4162 , n4161 );
not ( n4163 , n3257 );
or ( n4164 , n4162 , n4163 );
not ( n4165 , n46 );
not ( n4166 , n3368 );
or ( n4167 , n4165 , n4166 );
nand ( n4168 , n4164 , n4167 );
not ( n4169 , n4168 );
not ( n4170 , n3612 );
not ( n4171 , n4170 );
or ( n4172 , n4169 , n4171 );
not ( n4173 , n3992 );
nand ( n4174 , n3630 , n4173 );
nand ( n4175 , n4172 , n4174 );
not ( n4176 , n4175 );
nor ( n4177 , n3219 , n3233 );
not ( n4178 , n4177 );
and ( n4179 , n3515 , n40 );
not ( n4180 , n3515 );
and ( n4181 , n4180 , n3229 );
or ( n4182 , n4179 , n4181 );
not ( n4183 , n4182 );
or ( n4184 , n4178 , n4183 );
not ( n4185 , n3948 );
not ( n4186 , n3950 );
or ( n4187 , n4185 , n4186 );
nand ( n4188 , n4187 , n3234 );
nand ( n4189 , n4184 , n4188 );
not ( n4190 , n4189 );
not ( n4191 , n4190 );
not ( n4192 , n3348 );
not ( n4193 , n3891 );
or ( n4194 , n4192 , n4193 );
nor ( n4195 , n3354 , n3355 );
xnor ( n4196 , n42 , n3526 );
nand ( n4197 , n4195 , n4196 );
nand ( n4198 , n4194 , n4197 );
not ( n4199 , n4198 );
or ( n4200 , n4191 , n4199 );
not ( n4201 , n4189 );
or ( n4202 , n4201 , n4198 );
nand ( n4203 , n4200 , n4202 );
not ( n4204 , n4203 );
or ( n4205 , n4176 , n4204 );
not ( n4206 , n4201 );
nand ( n4207 , n4206 , n4198 );
nand ( n4208 , n4205 , n4207 );
not ( n4209 , n4208 );
not ( n4210 , n51 );
not ( n4211 , n4039 );
or ( n4212 , n4210 , n4211 );
not ( n4213 , n4031 );
and ( n4214 , n3 , n5 );
not ( n4215 , n3 );
and ( n4216 , n4215 , n21 );
nor ( n4217 , n4214 , n4216 );
xnor ( n4218 , n50 , n4217 );
nand ( n4219 , n4213 , n4218 );
nand ( n4220 , n4212 , n4219 );
not ( n4221 , n4220 );
not ( n4222 , n4221 );
nor ( n4223 , n37 , n38 );
not ( n4224 , n4223 );
not ( n4225 , n4224 );
not ( n4226 , n4050 );
not ( n4227 , n4226 );
not ( n4228 , n4227 );
or ( n4229 , n4225 , n4228 );
nand ( n4230 , n37 , n38 );
not ( n4231 , n4230 );
nor ( n4232 , n4231 , n3126 );
nand ( n4233 , n4229 , n4232 );
not ( n4234 , n4233 );
nand ( n4235 , n4222 , n4234 );
not ( n4236 , n4235 );
not ( n4237 , n4236 );
not ( n4238 , n3674 );
not ( n4239 , n3896 );
not ( n4240 , n44 );
and ( n4241 , n4239 , n4240 );
not ( n4242 , n4239 );
and ( n4243 , n4242 , n44 );
nor ( n4244 , n4241 , n4243 );
not ( n4245 , n4244 );
or ( n4246 , n4238 , n4245 );
buf ( n4247 , n3463 );
buf ( n4248 , n4247 );
not ( n4249 , n4248 );
nand ( n4250 , n4249 , n3911 );
nand ( n4251 , n4246 , n4250 );
not ( n4252 , n3847 );
not ( n4253 , n36 );
not ( n4254 , n4050 );
buf ( n4255 , n4254 );
not ( n4256 , n4255 );
or ( n4257 , n4253 , n4256 );
or ( n4258 , n36 , n4255 );
nand ( n4259 , n4257 , n4258 );
not ( n4260 , n4259 );
or ( n4261 , n4252 , n4260 );
not ( n4262 , n3582 );
nand ( n4263 , n4262 , n3938 );
nand ( n4264 , n4261 , n4263 );
nand ( n4265 , n4251 , n4264 );
or ( n4266 , n4264 , n4251 );
not ( n4267 , n3571 );
not ( n4268 , n4267 );
not ( n4269 , n4019 );
or ( n4270 , n4268 , n4269 );
xor ( n4271 , n48 , n3172 );
nand ( n4272 , n3566 , n4271 );
nand ( n4273 , n4270 , n4272 );
nand ( n4274 , n4266 , n4273 );
nand ( n4275 , n4265 , n4274 );
not ( n4276 , n4275 );
not ( n4277 , n4276 );
or ( n4278 , n4237 , n4277 );
not ( n4279 , n4265 );
not ( n4280 , n4274 );
or ( n4281 , n4279 , n4280 );
nand ( n4282 , n4281 , n4235 );
nand ( n4283 , n4278 , n4282 );
not ( n4284 , n4283 );
or ( n4285 , n4209 , n4284 );
nand ( n4286 , n4236 , n4275 );
nand ( n4287 , n4285 , n4286 );
not ( n4288 , n4287 );
xor ( n4289 , n4113 , n50 );
xor ( n4290 , n4109 , n4289 );
not ( n4291 , n4290 );
not ( n4292 , n4084 );
not ( n4293 , n4098 );
not ( n4294 , n4293 );
or ( n4295 , n4292 , n4294 );
not ( n4296 , n4098 );
or ( n4297 , n4084 , n4296 );
nand ( n4298 , n4295 , n4297 );
and ( n4299 , n4298 , n4090 );
not ( n4300 , n4298 );
not ( n4301 , n4090 );
and ( n4302 , n4300 , n4301 );
nor ( n4303 , n4299 , n4302 );
not ( n4304 , n4303 );
or ( n4305 , n4291 , n4304 );
or ( n4306 , n4290 , n4303 );
nand ( n4307 , n4305 , n4306 );
not ( n4308 , n4307 );
or ( n4309 , n4288 , n4308 );
not ( n4310 , n4290 );
nand ( n4311 , n4310 , n4303 );
nand ( n4312 , n4309 , n4311 );
not ( n4313 , n4312 );
not ( n4314 , n3839 );
not ( n4315 , n4314 );
not ( n4316 , n3222 );
not ( n4317 , n3959 );
or ( n4318 , n4316 , n4317 );
nand ( n4319 , n3235 , n3733 );
nand ( n4320 , n4318 , n4319 );
buf ( n4321 , n3972 );
not ( n4322 , n4321 );
not ( n4323 , n3752 );
or ( n4324 , n4322 , n4323 );
nand ( n4325 , n3090 , n3978 );
nand ( n4326 , n4324 , n4325 );
xor ( n4327 , n4320 , n4326 );
not ( n4328 , n4327 );
or ( n4329 , n4315 , n4328 );
nand ( n4330 , n4320 , n4326 );
nand ( n4331 , n4329 , n4330 );
not ( n4332 , n4331 );
not ( n4333 , n4332 );
not ( n4334 , n4128 );
not ( n4335 , n4120 );
not ( n4336 , n4335 );
or ( n4337 , n4334 , n4336 );
nand ( n4338 , n4127 , n4120 );
nand ( n4339 , n4337 , n4338 );
not ( n4340 , n4339 );
or ( n4341 , n4333 , n4340 );
or ( n4342 , n4332 , n4339 );
nand ( n4343 , n4341 , n4342 );
not ( n4344 , n4343 );
or ( n4345 , n4313 , n4344 );
not ( n4346 , n4332 );
nand ( n4347 , n4346 , n4339 );
nand ( n4348 , n4345 , n4347 );
not ( n4349 , n4348 );
and ( n4350 , n4160 , n4349 );
not ( n4351 , n4160 );
not ( n4352 , n4349 );
and ( n4353 , n4351 , n4352 );
nor ( n4354 , n4350 , n4353 );
not ( n4355 , n4354 );
or ( n4356 , n4157 , n4355 );
not ( n4357 , n4160 );
nand ( n4358 , n4357 , n4352 );
nand ( n4359 , n4356 , n4358 );
not ( n4360 , n4359 );
nor ( n4361 , n4155 , n4360 );
not ( n4362 , n3510 );
not ( n4363 , n3557 );
or ( n4364 , n4362 , n4363 );
nand ( n4365 , n3519 , n3551 );
nand ( n4366 , n4364 , n4365 );
not ( n4367 , n4366 );
not ( n4368 , n4367 );
not ( n4369 , n3238 );
not ( n4370 , n40 );
not ( n4371 , n3275 );
or ( n4372 , n4370 , n4371 );
not ( n4373 , n3272 );
or ( n4374 , n40 , n4373 );
nand ( n4375 , n4372 , n4374 );
not ( n4376 , n4375 );
or ( n4377 , n4369 , n4376 );
nand ( n4378 , n3225 , n3493 );
nand ( n4379 , n4377 , n4378 );
not ( n4380 , n3629 );
not ( n4381 , n4380 );
not ( n4382 , n4381 );
not ( n4383 , n3612 );
or ( n4384 , n4382 , n4383 );
nand ( n4385 , n4384 , n46 );
not ( n4386 , n4385 );
not ( n4387 , n4386 );
not ( n4388 , n3468 );
xor ( n4389 , n3102 , n44 );
not ( n4390 , n4389 );
or ( n4391 , n4388 , n4390 );
nand ( n4392 , n3674 , n3469 );
nand ( n4393 , n4391 , n4392 );
not ( n4394 , n4393 );
or ( n4395 , n4387 , n4394 );
or ( n4396 , n4386 , n4393 );
nand ( n4397 , n4395 , n4396 );
xnor ( n4398 , n4379 , n4397 );
not ( n4399 , n4398 );
not ( n4400 , n4399 );
or ( n4401 , n4368 , n4400 );
nand ( n4402 , n4366 , n4398 );
nand ( n4403 , n4401 , n4402 );
not ( n4404 , n3350 );
not ( n4405 , n42 );
not ( n4406 , n3133 );
or ( n4407 , n4405 , n4406 );
nand ( n4408 , n3502 , n3286 );
nand ( n4409 , n4407 , n4408 );
not ( n4410 , n4409 );
or ( n4411 , n4404 , n4410 );
not ( n4412 , n3358 );
nand ( n4413 , n4412 , n3508 );
nand ( n4414 , n4411 , n4413 );
not ( n4415 , n3422 );
not ( n4416 , n4415 );
not ( n4417 , n4416 );
not ( n4418 , n38 );
buf ( n4419 , n3481 );
not ( n4420 , n4419 );
not ( n4421 , n4420 );
or ( n4422 , n4418 , n4421 );
nand ( n4423 , n3096 , n4419 );
nand ( n4424 , n4422 , n4423 );
not ( n4425 , n4424 );
or ( n4426 , n4417 , n4425 );
nand ( n4427 , n3092 , n3441 );
nand ( n4428 , n4426 , n4427 );
and ( n4429 , n4414 , n4428 );
not ( n4430 , n4414 );
not ( n4431 , n4428 );
and ( n4432 , n4430 , n4431 );
nor ( n4433 , n4429 , n4432 );
not ( n4434 , n3124 );
not ( n4435 , n3534 );
or ( n4436 , n4434 , n4435 );
buf ( n4437 , n3414 );
and ( n4438 , n36 , n4437 );
not ( n4439 , n36 );
not ( n4440 , n4437 );
and ( n4441 , n4439 , n4440 );
nor ( n4442 , n4438 , n4441 );
not ( n4443 , n4442 );
or ( n4444 , n3145 , n4443 );
nand ( n4445 , n4436 , n4444 );
buf ( n4446 , n4445 );
xor ( n4447 , n4433 , n4446 );
xnor ( n4448 , n4403 , n4447 );
not ( n4449 , n4448 );
not ( n4450 , n3497 );
not ( n4451 , n3602 );
or ( n4452 , n4450 , n4451 );
not ( n4453 , n3601 );
not ( n4454 , n3557 );
xnor ( n4455 , n3510 , n4454 );
nand ( n4456 , n4453 , n4455 );
nand ( n4457 , n4452 , n4456 );
not ( n4458 , n4457 );
not ( n4459 , n4458 );
not ( n4460 , n3547 );
buf ( n4461 , n4460 );
nand ( n4462 , n36 , n4461 );
xor ( n4463 , n4462 , n3632 );
not ( n4464 , n4463 );
not ( n4465 , n3443 );
not ( n4466 , n3471 );
or ( n4467 , n4465 , n4466 );
not ( n4468 , n3443 );
not ( n4469 , n4468 );
not ( n4470 , n3471 );
not ( n4471 , n4470 );
or ( n4472 , n4469 , n4471 );
nand ( n4473 , n4472 , n3495 );
nand ( n4474 , n4467 , n4473 );
not ( n4475 , n4474 );
or ( n4476 , n4464 , n4475 );
or ( n4477 , n4463 , n4474 );
nand ( n4478 , n4476 , n4477 );
not ( n4479 , n3670 );
not ( n4480 , n3714 );
or ( n4481 , n4479 , n4480 );
nand ( n4482 , n3633 , n3669 );
nand ( n4483 , n4481 , n4482 );
and ( n4484 , n4478 , n4483 );
not ( n4485 , n4478 );
not ( n4486 , n4483 );
and ( n4487 , n4485 , n4486 );
nor ( n4488 , n4484 , n4487 );
not ( n4489 , n4488 );
or ( n4490 , n4459 , n4489 );
or ( n4491 , n4458 , n4488 );
nand ( n4492 , n4490 , n4491 );
not ( n4493 , n4492 );
or ( n4494 , n4449 , n4493 );
or ( n4495 , n4448 , n4492 );
nand ( n4496 , n4494 , n4495 );
not ( n4497 , n4496 );
not ( n4498 , n3603 );
not ( n4499 , n3813 );
or ( n4500 , n4498 , n4499 );
not ( n4501 , n3719 );
nand ( n4502 , n4501 , n3809 );
nand ( n4503 , n4500 , n4502 );
not ( n4504 , n4503 );
not ( n4505 , n4504 );
and ( n4506 , n4497 , n4505 );
and ( n4507 , n4504 , n4496 );
nor ( n4508 , n4506 , n4507 );
not ( n4509 , n3819 );
not ( n4510 , n4154 );
or ( n4511 , n4509 , n4510 );
nand ( n4512 , n3871 , n4148 );
nand ( n4513 , n4511 , n4512 );
not ( n4514 , n4513 );
nand ( n4515 , n4508 , n4514 );
nand ( n4516 , n4361 , n4515 );
not ( n4517 , n4514 );
not ( n4518 , n4508 );
nand ( n4519 , n4517 , n4518 );
nand ( n4520 , n4516 , n4519 );
not ( n4521 , n4520 );
not ( n4522 , n3092 );
not ( n4523 , n4424 );
or ( n4524 , n4522 , n4523 );
buf ( n4525 , n4321 );
not ( n4526 , n3096 );
not ( n4527 , n3368 );
not ( n4528 , n4527 );
or ( n4529 , n4526 , n4528 );
buf ( n4530 , n3257 );
or ( n4531 , n3096 , n4530 );
nand ( n4532 , n4529 , n4531 );
nand ( n4533 , n4525 , n4532 );
nand ( n4534 , n4524 , n4533 );
not ( n4535 , n3675 );
not ( n4536 , n4389 );
or ( n4537 , n4535 , n4536 );
nand ( n4538 , n44 , n3728 );
nand ( n4539 , n4537 , n4538 );
xor ( n4540 , n4534 , n4539 );
not ( n4541 , n3124 );
not ( n4542 , n4442 );
or ( n4543 , n4541 , n4542 );
not ( n4544 , n3126 );
buf ( n4545 , n3431 );
not ( n4546 , n4545 );
not ( n4547 , n4546 );
or ( n4548 , n4544 , n4547 );
not ( n4549 , n4545 );
or ( n4550 , n3126 , n4549 );
nand ( n4551 , n4548 , n4550 );
nand ( n4552 , n3280 , n4551 );
nand ( n4553 , n4543 , n4552 );
xor ( n4554 , n4540 , n4553 );
not ( n4555 , n4379 );
not ( n4556 , n4397 );
or ( n4557 , n4555 , n4556 );
not ( n4558 , n4386 );
nand ( n4559 , n4558 , n4393 );
nand ( n4560 , n4557 , n4559 );
not ( n4561 , n4560 );
not ( n4562 , n4561 );
not ( n4563 , n4445 );
not ( n4564 , n4433 );
or ( n4565 , n4563 , n4564 );
not ( n4566 , n4431 );
nand ( n4567 , n4566 , n4414 );
nand ( n4568 , n4565 , n4567 );
not ( n4569 , n4568 );
or ( n4570 , n4562 , n4569 );
or ( n4571 , n4561 , n4568 );
nand ( n4572 , n4570 , n4571 );
and ( n4573 , n4554 , n4572 );
not ( n4574 , n4554 );
not ( n4575 , n4572 );
and ( n4576 , n4574 , n4575 );
or ( n4577 , n4573 , n4576 );
not ( n4578 , n4457 );
not ( n4579 , n4488 );
or ( n4580 , n4578 , n4579 );
not ( n4581 , n4486 );
nand ( n4582 , n4478 , n4581 );
nand ( n4583 , n4580 , n4582 );
not ( n4584 , n4583 );
xor ( n4585 , n4577 , n4584 );
not ( n4586 , n4463 );
not ( n4587 , n4586 );
not ( n4588 , n4474 );
or ( n4589 , n4587 , n4588 );
not ( n4590 , n4462 );
nand ( n4591 , n4590 , n3632 );
nand ( n4592 , n4589 , n4591 );
not ( n4593 , n3532 );
not ( n4594 , n4593 );
and ( n4595 , n36 , n4594 );
not ( n4596 , n4595 );
not ( n4597 , n3358 );
not ( n4598 , n4597 );
not ( n4599 , n4409 );
or ( n4600 , n4598 , n4599 );
buf ( n4601 , n3350 );
not ( n4602 , n3502 );
not ( n4603 , n3155 );
or ( n4604 , n4602 , n4603 );
or ( n4605 , n3502 , n3155 );
nand ( n4606 , n4604 , n4605 );
nand ( n4607 , n4601 , n4606 );
nand ( n4608 , n4600 , n4607 );
not ( n4609 , n4608 );
or ( n4610 , n4596 , n4609 );
or ( n4611 , n4595 , n4608 );
nand ( n4612 , n4610 , n4611 );
not ( n4613 , n3225 );
not ( n4614 , n4375 );
or ( n4615 , n4613 , n4614 );
not ( n4616 , n40 );
not ( n4617 , n3172 );
not ( n4618 , n4617 );
or ( n4619 , n4616 , n4618 );
or ( n4620 , n40 , n4617 );
nand ( n4621 , n4619 , n4620 );
nand ( n4622 , n3317 , n4621 );
nand ( n4623 , n4615 , n4622 );
and ( n4624 , n4612 , n4623 );
not ( n4625 , n4612 );
not ( n4626 , n4623 );
and ( n4627 , n4625 , n4626 );
nor ( n4628 , n4624 , n4627 );
xor ( n4629 , n4592 , n4628 );
not ( n4630 , n4447 );
not ( n4631 , n4403 );
or ( n4632 , n4630 , n4631 );
nand ( n4633 , n4366 , n4399 );
nand ( n4634 , n4632 , n4633 );
xor ( n4635 , n4629 , n4634 );
xnor ( n4636 , n4585 , n4635 );
not ( n4637 , n4636 );
not ( n4638 , n4503 );
not ( n4639 , n4496 );
or ( n4640 , n4638 , n4639 );
not ( n4641 , n4448 );
nand ( n4642 , n4641 , n4492 );
nand ( n4643 , n4640 , n4642 );
not ( n4644 , n4643 );
not ( n4645 , n4644 );
nand ( n4646 , n4637 , n4645 );
nand ( n4647 , n4521 , n4646 );
not ( n4648 , n4636 );
not ( n4649 , n4643 );
not ( n4650 , n4649 );
or ( n4651 , n4648 , n4650 );
not ( n4652 , n4629 );
not ( n4653 , n4634 );
or ( n4654 , n4652 , n4653 );
nand ( n4655 , n4628 , n4592 );
nand ( n4656 , n4654 , n4655 );
not ( n4657 , n4554 );
not ( n4658 , n4572 );
or ( n4659 , n4657 , n4658 );
not ( n4660 , n4568 );
or ( n4661 , n4561 , n4660 );
nand ( n4662 , n4659 , n4661 );
not ( n4663 , n4662 );
not ( n4664 , n3126 );
buf ( n4665 , n4419 );
not ( n4666 , n4665 );
not ( n4667 , n4666 );
or ( n4668 , n4664 , n4667 );
not ( n4669 , n4420 );
nand ( n4670 , n36 , n4669 );
nand ( n4671 , n4668 , n4670 );
not ( n4672 , n4671 );
and ( n4673 , n4672 , n3146 );
not ( n4674 , n4551 );
nor ( n4675 , n4434 , n4674 );
nor ( n4676 , n4673 , n4675 );
not ( n4677 , n4676 );
not ( n4678 , n3415 );
and ( n4679 , n36 , n4678 );
not ( n4680 , n3236 );
not ( n4681 , n40 );
not ( n4682 , n3133 );
or ( n4683 , n4681 , n4682 );
nand ( n4684 , n3229 , n3132 );
nand ( n4685 , n4683 , n4684 );
not ( n4686 , n4685 );
or ( n4687 , n4680 , n4686 );
nand ( n4688 , n3224 , n4621 );
nand ( n4689 , n4687 , n4688 );
xor ( n4690 , n4679 , n4689 );
not ( n4691 , n4690 );
or ( n4692 , n4677 , n4691 );
or ( n4693 , n4676 , n4690 );
nand ( n4694 , n4692 , n4693 );
not ( n4695 , n4694 );
not ( n4696 , n4608 );
not ( n4697 , n4696 );
not ( n4698 , n4539 );
not ( n4699 , n4553 );
or ( n4700 , n4698 , n4699 );
or ( n4701 , n4553 , n4539 );
nand ( n4702 , n4701 , n4534 );
nand ( n4703 , n4700 , n4702 );
not ( n4704 , n4703 );
or ( n4705 , n4697 , n4704 );
or ( n4706 , n4696 , n4703 );
nand ( n4707 , n4705 , n4706 );
nand ( n4708 , n4695 , n4707 );
not ( n4709 , n4708 );
not ( n4710 , n4694 );
nor ( n4711 , n4710 , n4707 );
nor ( n4712 , n4709 , n4711 );
not ( n4713 , n4712 );
not ( n4714 , n4623 );
not ( n4715 , n4612 );
or ( n4716 , n4714 , n4715 );
nand ( n4717 , n4595 , n4696 );
nand ( n4718 , n4716 , n4717 );
not ( n4719 , n4718 );
not ( n4720 , n4597 );
not ( n4721 , n4606 );
or ( n4722 , n4720 , n4721 );
not ( n4723 , n42 );
not ( n4724 , n3102 );
not ( n4725 , n4724 );
or ( n4726 , n4723 , n4725 );
nand ( n4727 , n3502 , n3102 );
nand ( n4728 , n4726 , n4727 );
nand ( n4729 , n4601 , n4728 );
nand ( n4730 , n4722 , n4729 );
not ( n4731 , n4248 );
not ( n4732 , n4731 );
not ( n4733 , n4732 );
not ( n4734 , n3675 );
not ( n4735 , n4734 );
or ( n4736 , n4733 , n4735 );
nand ( n4737 , n4736 , n44 );
not ( n4738 , n38 );
not ( n4739 , n3271 );
not ( n4740 , n4739 );
or ( n4741 , n4738 , n4740 );
nand ( n4742 , n3096 , n3271 );
nand ( n4743 , n4741 , n4742 );
nand ( n4744 , n3113 , n4743 );
nand ( n4745 , n3092 , n4532 );
nand ( n4746 , n4744 , n4745 );
xor ( n4747 , n4737 , n4746 );
xnor ( n4748 , n4730 , n4747 );
not ( n4749 , n4748 );
or ( n4750 , n4719 , n4749 );
or ( n4751 , n4718 , n4748 );
nand ( n4752 , n4750 , n4751 );
not ( n4753 , n4752 );
and ( n4754 , n4713 , n4753 );
and ( n4755 , n4752 , n4712 );
nor ( n4756 , n4754 , n4755 );
not ( n4757 , n4756 );
or ( n4758 , n4663 , n4757 );
or ( n4759 , n4662 , n4756 );
nand ( n4760 , n4758 , n4759 );
xnor ( n4761 , n4656 , n4760 );
not ( n4762 , t_0 );
nand ( n4763 , n4761 , n4762 );
nand ( n4764 , n4651 , n4763 );
not ( n4765 , n4764 );
nand ( n4766 , n4647 , n4765 );
xor ( n4767 , n4343 , n4312 );
not ( n4768 , n4767 );
not ( n4769 , n3883 );
xnor ( n4770 , n4769 , n4072 );
not ( n4771 , n4770 );
and ( n4772 , n4068 , n3946 );
not ( n4773 , n4068 );
not ( n4774 , n3946 );
and ( n4775 , n4773 , n4774 );
nor ( n4776 , n4772 , n4775 );
not ( n4777 , n4776 );
xor ( n4778 , n3839 , n4327 );
and ( n4779 , n3917 , n3940 );
not ( n4780 , n3917 );
and ( n4781 , n4780 , n3941 );
or ( n4782 , n4779 , n4781 );
xor ( n4783 , n4005 , n3980 );
not ( n4784 , n3961 );
xnor ( n4785 , n4783 , n4784 );
xor ( n4786 , n4027 , n4058 );
nor ( n4787 , n4785 , n4786 );
or ( n4788 , n4782 , n4787 );
nand ( n4789 , n4786 , n4785 );
nand ( n4790 , n4788 , n4789 );
not ( n4791 , n4790 );
and ( n4792 , n4778 , n4791 );
not ( n4793 , n4778 );
not ( n4794 , n4791 );
and ( n4795 , n4793 , n4794 );
nor ( n4796 , n4792 , n4795 );
not ( n4797 , n4796 );
or ( n4798 , n4777 , n4797 );
not ( n4799 , n4778 );
nand ( n4800 , n4799 , n4794 );
nand ( n4801 , n4798 , n4800 );
not ( n4802 , n4801 );
not ( n4803 , n4802 );
or ( n4804 , n4771 , n4803 );
not ( n4805 , n4770 );
nand ( n4806 , n4805 , n4801 );
nand ( n4807 , n4804 , n4806 );
not ( n4808 , n4807 );
or ( n4809 , n4768 , n4808 );
nand ( n4810 , n4770 , n4801 );
nand ( n4811 , n4809 , n4810 );
not ( n4812 , n4811 );
xor ( n4813 , n4160 , n4349 );
xnor ( n4814 , n4813 , n4156 );
nand ( n4815 , n4812 , n4814 );
not ( n4816 , n4815 );
nor ( n4817 , n4816 , n4764 );
and ( n4818 , n4264 , n4251 );
not ( n4819 , n4264 );
not ( n4820 , n4251 );
and ( n4821 , n4819 , n4820 );
nor ( n4822 , n4818 , n4821 );
and ( n4823 , n4822 , n4273 );
not ( n4824 , n4822 );
not ( n4825 , n4273 );
and ( n4826 , n4824 , n4825 );
nor ( n4827 , n4823 , n4826 );
not ( n4828 , n4827 );
not ( n4829 , n3356 );
not ( n4830 , n42 );
not ( n4831 , n3748 );
or ( n4832 , n4830 , n4831 );
nand ( n4833 , n3502 , n3543 );
nand ( n4834 , n4832 , n4833 );
not ( n4835 , n4834 );
or ( n4836 , n4829 , n4835 );
nand ( n4837 , n3894 , n4196 );
nand ( n4838 , n4836 , n4837 );
not ( n4839 , n4838 );
not ( n4840 , n4839 );
not ( n4841 , n3674 );
xor ( n4842 , n44 , n3413 );
not ( n4843 , n4842 );
or ( n4844 , n4841 , n4843 );
nand ( n4845 , n4249 , n4244 );
nand ( n4846 , n4844 , n4845 );
nand ( n4847 , n4840 , n4846 );
not ( n4848 , n4839 );
not ( n4849 , n4846 );
not ( n4850 , n4849 );
or ( n4851 , n4848 , n4850 );
not ( n4852 , n4380 );
not ( n4853 , n4168 );
or ( n4854 , n4852 , n4853 );
xor ( n4855 , n3480 , n46 );
buf ( n4856 , n4855 );
nand ( n4857 , n3779 , n4856 );
nand ( n4858 , n4854 , n4857 );
nand ( n4859 , n4851 , n4858 );
nand ( n4860 , n4847 , n4859 );
not ( n4861 , n4860 );
not ( n4862 , n4175 );
and ( n4863 , n4203 , n4862 );
not ( n4864 , n4203 );
and ( n4865 , n4864 , n4175 );
nor ( n4866 , n4863 , n4865 );
not ( n4867 , n4866 );
or ( n4868 , n4861 , n4867 );
buf ( n4869 , n4860 );
or ( n4870 , n4869 , n4866 );
nand ( n4871 , n4868 , n4870 );
not ( n4872 , n4871 );
or ( n4873 , n4828 , n4872 );
not ( n4874 , n4866 );
nand ( n4875 , n4869 , n4874 );
nand ( n4876 , n4873 , n4875 );
not ( n4877 , n4876 );
not ( n4878 , n3566 );
xor ( n4879 , n48 , n3270 );
not ( n4880 , n4879 );
or ( n4881 , n4878 , n4880 );
nand ( n4882 , n4267 , n4271 );
nand ( n4883 , n4881 , n4882 );
not ( n4884 , n4883 );
not ( n4885 , n4255 );
nand ( n4886 , n4885 , n3141 );
not ( n4887 , n4886 );
not ( n4888 , n4030 );
not ( n4889 , n4888 );
not ( n4890 , n50 );
not ( n4891 , n4890 );
and ( n4892 , n3 , n6 );
not ( n4893 , n3 );
and ( n4894 , n4893 , n22 );
nor ( n4895 , n4892 , n4894 );
not ( n4896 , n4895 );
not ( n4897 , n4896 );
or ( n4898 , n4891 , n4897 );
not ( n4899 , n50 );
not ( n4900 , n3130 );
or ( n4901 , n4899 , n4900 );
nand ( n4902 , n4898 , n4901 );
not ( n4903 , n4902 );
or ( n4904 , n4889 , n4903 );
nand ( n4905 , n51 , n4218 );
nand ( n4906 , n4904 , n4905 );
not ( n4907 , n4906 );
and ( n4908 , n4887 , n4907 );
and ( n4909 , n4886 , n4906 );
nor ( n4910 , n4908 , n4909 );
or ( n4911 , n4884 , n4910 );
not ( n4912 , n4886 );
nand ( n4913 , n4912 , n4906 );
nand ( n4914 , n4911 , n4913 );
not ( n4915 , n4914 );
not ( n4916 , n4233 );
not ( n4917 , n4916 );
not ( n4918 , n4221 );
or ( n4919 , n4917 , n4918 );
nand ( n4920 , n4233 , n4220 );
nand ( n4921 , n4919 , n4920 );
not ( n4922 , n3422 );
not ( n4923 , n3969 );
or ( n4924 , n4922 , n4923 );
not ( n4925 , n38 );
not ( n4926 , n3772 );
not ( n4927 , n4926 );
or ( n4928 , n4925 , n4927 );
not ( n4929 , n3772 );
or ( n4930 , n38 , n4929 );
nand ( n4931 , n4928 , n4930 );
nand ( n4932 , n3091 , n4931 );
nand ( n4933 , n4924 , n4932 );
xnor ( n4934 , n4921 , n4933 );
not ( n4935 , n4934 );
not ( n4936 , n4935 );
or ( n4937 , n4915 , n4936 );
nand ( n4938 , n4933 , n4921 );
nand ( n4939 , n4937 , n4938 );
not ( n4940 , n4939 );
not ( n4941 , n4208 );
and ( n4942 , n4283 , n4941 );
not ( n4943 , n4283 );
and ( n4944 , n4943 , n4208 );
nor ( n4945 , n4942 , n4944 );
not ( n4946 , n4945 );
and ( n4947 , n4940 , n4946 );
not ( n4948 , n4940 );
and ( n4949 , n4948 , n4945 );
nor ( n4950 , n4947 , n4949 );
not ( n4951 , n4950 );
not ( n4952 , n4951 );
or ( n4953 , n4877 , n4952 );
nand ( n4954 , n4939 , n4946 );
nand ( n4955 , n4953 , n4954 );
not ( n4956 , n4955 );
and ( n4957 , n4287 , n4307 );
not ( n4958 , n4287 );
not ( n4959 , n4307 );
and ( n4960 , n4958 , n4959 );
nor ( n4961 , n4957 , n4960 );
xor ( n4962 , n4778 , n4791 );
xnor ( n4963 , n4962 , n4776 );
not ( n4964 , n4963 );
and ( n4965 , n4961 , n4964 );
not ( n4966 , n4961 );
not ( n4967 , n4964 );
and ( n4968 , n4966 , n4967 );
nor ( n4969 , n4965 , n4968 );
not ( n4970 , n4969 );
or ( n4971 , n4956 , n4970 );
not ( n4972 , n4967 );
nand ( n4973 , n4961 , n4972 );
nand ( n4974 , n4971 , n4973 );
not ( n4975 , n4974 );
not ( n4976 , n4767 );
and ( n4977 , n4807 , n4976 );
not ( n4978 , n4807 );
and ( n4979 , n4978 , n4767 );
nor ( n4980 , n4977 , n4979 );
nand ( n4981 , n4975 , n4980 );
not ( n4982 , n4981 );
not ( n4983 , n4876 );
not ( n4984 , n4983 );
not ( n4985 , n4951 );
or ( n4986 , n4984 , n4985 );
nand ( n4987 , n4876 , n4950 );
nand ( n4988 , n4986 , n4987 );
not ( n4989 , n4988 );
buf ( n4990 , n4782 );
not ( n4991 , n4990 );
buf ( n4992 , n4786 );
not ( n4993 , n4785 );
not ( n4994 , n4993 );
nand ( n4995 , n4991 , n4992 , n4994 );
not ( n4996 , n4990 );
not ( n4997 , n4992 );
nand ( n4998 , n4996 , n4997 , n4993 );
not ( n4999 , n4992 );
not ( n5000 , n4993 );
nand ( n5001 , n4999 , n4990 , n5000 );
nand ( n5002 , n4992 , n4990 , n4993 );
nand ( n5003 , n4995 , n4998 , n5001 , n5002 );
not ( n5004 , n5003 );
and ( n5005 , n4910 , n4884 );
not ( n5006 , n4910 );
and ( n5007 , n5006 , n4883 );
nor ( n5008 , n5005 , n5007 );
not ( n5009 , n3235 );
and ( n5010 , n3229 , n3851 );
not ( n5011 , n3229 );
and ( n5012 , n5011 , n3852 );
nor ( n5013 , n5010 , n5012 );
not ( n5014 , n5013 );
or ( n5015 , n5009 , n5014 );
not ( n5016 , n40 );
not ( n5017 , n3773 );
or ( n5018 , n5016 , n5017 );
or ( n5019 , n40 , n3921 );
nand ( n5020 , n5018 , n5019 );
nand ( n5021 , n3222 , n5020 );
nand ( n5022 , n5015 , n5021 );
not ( n5023 , n5022 );
not ( n5024 , n3628 );
not ( n5025 , n4855 );
or ( n5026 , n5024 , n5025 );
not ( n5027 , n46 );
not ( n5028 , n3431 );
or ( n5029 , n5027 , n5028 );
or ( n5030 , n46 , n3431 );
nand ( n5031 , n5029 , n5030 );
nand ( n5032 , n3611 , n5031 );
nand ( n5033 , n5026 , n5032 );
not ( n5034 , n5033 );
nand ( n5035 , n5023 , n5034 );
not ( n5036 , n5033 );
not ( n5037 , n5022 );
or ( n5038 , n5036 , n5037 );
not ( n5039 , n3964 );
not ( n5040 , n38 );
not ( n5041 , n4226 );
or ( n5042 , n5040 , n5041 );
or ( n5043 , n4052 , n38 );
nand ( n5044 , n5042 , n5043 );
not ( n5045 , n5044 );
or ( n5046 , n5039 , n5045 );
not ( n5047 , n3973 );
and ( n5048 , n38 , n3936 );
not ( n5049 , n38 );
not ( n5050 , n3932 );
and ( n5051 , n5049 , n5050 );
nor ( n5052 , n5048 , n5051 );
nand ( n5053 , n5047 , n5052 );
nand ( n5054 , n5046 , n5053 );
not ( n5055 , n5054 );
nand ( n5056 , n5038 , n5055 );
nand ( n5057 , n5035 , n5056 );
not ( n5058 , n5057 );
xor ( n5059 , n5008 , n5058 );
not ( n5060 , n3727 );
not ( n5061 , n4842 );
or ( n5062 , n5060 , n5061 );
and ( n5063 , n3 , n13 );
not ( n5064 , n3 );
and ( n5065 , n5064 , n29 );
nor ( n5066 , n5063 , n5065 );
xnor ( n5067 , n44 , n5066 );
nand ( n5068 , n3674 , n5067 );
nand ( n5069 , n5062 , n5068 );
not ( n5070 , n3349 );
not ( n5071 , n4834 );
or ( n5072 , n5070 , n5071 );
not ( n5073 , n42 );
not ( n5074 , n3516 );
and ( n5075 , n5073 , n5074 );
not ( n5076 , n3517 );
and ( n5077 , n42 , n5076 );
nor ( n5078 , n5075 , n5077 );
nand ( n5079 , n3788 , n5078 );
nand ( n5080 , n5072 , n5079 );
xor ( n5081 , n5069 , n5080 );
not ( n5082 , n4267 );
not ( n5083 , n4879 );
or ( n5084 , n5082 , n5083 );
not ( n5085 , n3565 );
not ( n5086 , n48 );
not ( n5087 , n3256 );
or ( n5088 , n5086 , n5087 );
or ( n5089 , n48 , n3256 );
nand ( n5090 , n5088 , n5089 );
nand ( n5091 , n5085 , n5090 );
nand ( n5092 , n5084 , n5091 );
and ( n5093 , n5081 , n5092 );
and ( n5094 , n5069 , n5080 );
or ( n5095 , n5093 , n5094 );
and ( n5096 , n5059 , n5095 );
and ( n5097 , n5008 , n5058 );
or ( n5098 , n5096 , n5097 );
not ( n5099 , n5098 );
not ( n5100 , n4914 );
not ( n5101 , n4934 );
or ( n5102 , n5100 , n5101 );
or ( n5103 , n4914 , n4934 );
nand ( n5104 , n5102 , n5103 );
nand ( n5105 , n39 , n40 );
not ( n5106 , n5105 );
not ( n5107 , n4052 );
or ( n5108 , n5106 , n5107 );
nor ( n5109 , n39 , n40 );
not ( n5110 , n5109 );
nand ( n5111 , n5108 , n5110 );
nand ( n5112 , n38 , n5111 );
not ( n5113 , n5112 );
not ( n5114 , n51 );
not ( n5115 , n4902 );
or ( n5116 , n5114 , n5115 );
not ( n5117 , n50 );
not ( n5118 , n5117 );
not ( n5119 , n3171 );
or ( n5120 , n5118 , n5119 );
not ( n5121 , n50 );
or ( n5122 , n5121 , n3171 );
nand ( n5123 , n5120 , n5122 );
nand ( n5124 , n4032 , n5123 );
nand ( n5125 , n5116 , n5124 );
nand ( n5126 , n5113 , n5125 );
not ( n5127 , n5126 );
not ( n5128 , n5127 );
not ( n5129 , n3090 );
not ( n5130 , n5052 );
or ( n5131 , n5129 , n5130 );
buf ( n5132 , n5047 );
nand ( n5133 , n5132 , n4931 );
nand ( n5134 , n5131 , n5133 );
not ( n5135 , n5134 );
not ( n5136 , n5135 );
not ( n5137 , n3222 );
not ( n5138 , n5013 );
or ( n5139 , n5137 , n5138 );
nand ( n5140 , n3736 , n4182 );
nand ( n5141 , n5139 , n5140 );
not ( n5142 , n5141 );
or ( n5143 , n5136 , n5142 );
not ( n5144 , n5134 );
or ( n5145 , n5141 , n5144 );
nand ( n5146 , n5143 , n5145 );
not ( n5147 , n5146 );
or ( n5148 , n5128 , n5147 );
not ( n5149 , n5144 );
nand ( n5150 , n5141 , n5149 );
nand ( n5151 , n5148 , n5150 );
not ( n5152 , n5151 );
and ( n5153 , n5104 , n5152 );
not ( n5154 , n5104 );
and ( n5155 , n5154 , n5151 );
nor ( n5156 , n5153 , n5155 );
nor ( n5157 , n5099 , n5156 );
not ( n5158 , n5152 );
and ( n5159 , n5104 , n5158 );
nor ( n5160 , n5157 , n5159 );
not ( n5161 , n5160 );
or ( n5162 , n5004 , n5161 );
not ( n5163 , n5159 );
not ( n5164 , n5163 );
not ( n5165 , n5157 );
not ( n5166 , n5165 );
or ( n5167 , n5164 , n5166 );
not ( n5168 , n4996 );
not ( n5169 , n4787 );
or ( n5170 , n5168 , n5169 );
nand ( n5171 , n5170 , n4995 );
not ( n5172 , n4997 );
nand ( n5173 , n4990 , n5000 );
or ( n5174 , n5172 , n5173 );
nand ( n5175 , n5174 , n5002 );
nor ( n5176 , n5171 , n5175 );
nand ( n5177 , n5167 , n5176 );
nand ( n5178 , n5162 , n5177 );
not ( n5179 , n5178 );
or ( n5180 , n4989 , n5179 );
not ( n5181 , n5160 );
nand ( n5182 , n5003 , n5181 );
nand ( n5183 , n5180 , n5182 );
not ( n5184 , n5183 );
not ( n5185 , n5184 );
xor ( n5186 , n4961 , n4964 );
xnor ( n5187 , n5186 , n4955 );
not ( n5188 , n5187 );
nor ( n5189 , n5185 , n5188 );
xor ( n5190 , n5156 , n5099 );
not ( n5191 , n5190 );
xor ( n5192 , n4860 , n4866 );
xor ( n5193 , n5192 , n4827 );
buf ( n5194 , n5193 );
not ( n5195 , n5194 );
not ( n5196 , n4213 );
xor ( n5197 , n3269 , n50 );
not ( n5198 , n5197 );
or ( n5199 , n5196 , n5198 );
nand ( n5200 , n51 , n5123 );
nand ( n5201 , n5199 , n5200 );
not ( n5202 , n3634 );
not ( n5203 , n5078 );
or ( n5204 , n5202 , n5203 );
not ( n5205 , n42 );
not ( n5206 , n3691 );
or ( n5207 , n5205 , n5206 );
or ( n5208 , n42 , n3691 );
nand ( n5209 , n5207 , n5208 );
nand ( n5210 , n3885 , n5209 );
nand ( n5211 , n5204 , n5210 );
xor ( n5212 , n5201 , n5211 );
not ( n5213 , n3223 );
not ( n5214 , n5213 );
not ( n5215 , n40 );
not ( n5216 , n3933 );
or ( n5217 , n5215 , n5216 );
or ( n5218 , n40 , n3933 );
nand ( n5219 , n5217 , n5218 );
not ( n5220 , n5219 );
or ( n5221 , n5214 , n5220 );
nand ( n5222 , n3235 , n5020 );
nand ( n5223 , n5221 , n5222 );
and ( n5224 , n5212 , n5223 );
and ( n5225 , n5201 , n5211 );
or ( n5226 , n5224 , n5225 );
not ( n5227 , n5226 );
not ( n5228 , n3570 );
not ( n5229 , n5228 );
not ( n5230 , n5090 );
or ( n5231 , n5229 , n5230 );
not ( n5232 , n3565 );
not ( n5233 , n10 );
and ( n5234 , n3 , n5233 );
not ( n5235 , n3 );
not ( n5236 , n26 );
and ( n5237 , n5235 , n5236 );
nor ( n5238 , n5234 , n5237 );
xor ( n5239 , n5238 , n48 );
nand ( n5240 , n5232 , n5239 );
nand ( n5241 , n5231 , n5240 );
not ( n5242 , n5241 );
not ( n5243 , n3452 );
and ( n5244 , n3 , n14 );
not ( n5245 , n3 );
and ( n5246 , n5245 , n30 );
nor ( n5247 , n5244 , n5246 );
and ( n5248 , n44 , n5247 );
not ( n5249 , n44 );
and ( n5250 , n5249 , n3542 );
or ( n5251 , n5248 , n5250 );
not ( n5252 , n5251 );
or ( n5253 , n5243 , n5252 );
nand ( n5254 , n3725 , n5067 );
nand ( n5255 , n5253 , n5254 );
nand ( n5256 , n3111 , n4051 );
not ( n5257 , n5256 );
and ( n5258 , n5255 , n5257 );
not ( n5259 , n5255 );
not ( n5260 , n5257 );
and ( n5261 , n5259 , n5260 );
nor ( n5262 , n5258 , n5261 );
not ( n5263 , n5262 );
or ( n5264 , n5242 , n5263 );
not ( n5265 , n5260 );
nand ( n5266 , n5265 , n5255 );
nand ( n5267 , n5264 , n5266 );
not ( n5268 , n5267 );
not ( n5269 , n5268 );
not ( n5270 , n5112 );
not ( n5271 , n5270 );
not ( n5272 , n5125 );
not ( n5273 , n5272 );
or ( n5274 , n5271 , n5273 );
not ( n5275 , n38 );
not ( n5276 , n5111 );
or ( n5277 , n5275 , n5276 );
nand ( n5278 , n5277 , n5125 );
nand ( n5279 , n5274 , n5278 );
buf ( n5280 , n5279 );
and ( n5281 , n5269 , n5280 );
not ( n5282 , n5269 );
not ( n5283 , n5280 );
and ( n5284 , n5282 , n5283 );
nor ( n5285 , n5281 , n5284 );
not ( n5286 , n5285 );
or ( n5287 , n5227 , n5286 );
not ( n5288 , n5283 );
nand ( n5289 , n5288 , n5269 );
nand ( n5290 , n5287 , n5289 );
not ( n5291 , n5290 );
xor ( n5292 , n5126 , n5146 );
not ( n5293 , n5292 );
not ( n5294 , n5293 );
not ( n5295 , n4858 );
not ( n5296 , n4839 );
nor ( n5297 , n5296 , n4846 );
not ( n5298 , n5297 );
or ( n5299 , n5295 , n5298 );
not ( n5300 , n4839 );
nand ( n5301 , n4858 , n5300 , n4846 );
nand ( n5302 , n5299 , n5301 );
not ( n5303 , n4858 );
not ( n5304 , n5303 );
and ( n5305 , n4846 , n4839 );
not ( n5306 , n4846 );
and ( n5307 , n5306 , n5300 );
nor ( n5308 , n5305 , n5307 );
nor ( n5309 , n5304 , n5308 );
nor ( n5310 , n5302 , n5309 );
not ( n5311 , n5310 );
or ( n5312 , n5294 , n5311 );
not ( n5313 , n5309 );
not ( n5314 , n5302 );
nand ( n5315 , n5313 , n5314 );
nand ( n5316 , n5292 , n5315 );
nand ( n5317 , n5312 , n5316 );
not ( n5318 , n5317 );
or ( n5319 , n5291 , n5318 );
not ( n5320 , n5292 );
nand ( n5321 , n5320 , n5315 );
nand ( n5322 , n5319 , n5321 );
not ( n5323 , n5322 );
not ( n5324 , n5323 );
not ( n5325 , n5324 );
or ( n5326 , n5195 , n5325 );
not ( n5327 , n5323 );
or ( n5328 , n5194 , n5327 );
nand ( n5329 , n5326 , n5328 );
not ( n5330 , n5329 );
or ( n5331 , n5191 , n5330 );
not ( n5332 , n5194 );
not ( n5333 , n5323 );
nand ( n5334 , n5332 , n5333 );
nand ( n5335 , n5331 , n5334 );
not ( n5336 , n4988 );
not ( n5337 , n5336 );
not ( n5338 , n5178 );
or ( n5339 , n5337 , n5338 );
or ( n5340 , n5336 , n5178 );
nand ( n5341 , n5339 , n5340 );
nand ( n5342 , n5335 , n5341 );
or ( n5343 , n5189 , n5342 );
not ( n5344 , n5184 );
nand ( n5345 , n5344 , n5188 );
nand ( n5346 , n5343 , n5345 );
not ( n5347 , n5346 );
or ( n5348 , n4982 , n5347 );
not ( n5349 , n4975 );
not ( n5350 , n4980 );
nand ( n5351 , n5349 , n5350 );
not ( n5352 , n4814 );
nand ( n5353 , n5352 , n4811 );
nand ( n5354 , n5351 , n5353 );
not ( n5355 , n5354 );
nand ( n5356 , n5348 , n5355 );
nand ( n5357 , n4155 , n4360 );
not ( n5358 , n5357 );
not ( n5359 , n4515 );
nor ( n5360 , n5358 , n5359 );
and ( n5361 , n4817 , n5356 , n5360 );
not ( n5362 , n4761 );
nand ( n5363 , t_1 , n5362 );
not ( n5364 , n5363 );
nor ( n5365 , n5361 , n5364 );
xor ( n5366 , n5008 , n5058 );
xor ( n5367 , n5366 , n5095 );
nor ( n5368 , n41 , n42 );
not ( n5369 , n5368 );
not ( n5370 , n5369 );
not ( n5371 , n3 );
nand ( n5372 , n5371 , n35 );
nand ( n5373 , n5372 , n4049 );
not ( n5374 , n5373 );
not ( n5375 , n5374 );
not ( n5376 , n5375 );
or ( n5377 , n5370 , n5376 );
nand ( n5378 , n41 , n42 );
nand ( n5379 , n40 , n5378 );
not ( n5380 , n5379 );
nand ( n5381 , n5377 , n5380 );
not ( n5382 , n5381 );
not ( n5383 , n3429 );
not ( n5384 , n48 );
not ( n5385 , n5384 );
and ( n5386 , n5383 , n5385 );
not ( n5387 , n48 );
and ( n5388 , n5387 , n3429 );
nor ( n5389 , n5386 , n5388 );
not ( n5390 , n5389 );
not ( n5391 , n3564 );
and ( n5392 , n5390 , n5391 );
and ( n5393 , n3569 , n5239 );
nor ( n5394 , n5392 , n5393 );
not ( n5395 , n5394 );
nand ( n5396 , n5382 , n5395 );
not ( n5397 , n5396 );
not ( n5398 , n4381 );
nand ( n5399 , n5398 , n5031 );
not ( n5400 , n46 );
not ( n5401 , n5400 );
not ( n5402 , n3887 );
or ( n5403 , n5401 , n5402 );
not ( n5404 , n46 );
or ( n5405 , n5404 , n3413 );
nand ( n5406 , n5403 , n5405 );
nand ( n5407 , n3613 , n5406 );
nand ( n5408 , n5399 , n5407 );
not ( n5409 , n5408 );
or ( n5410 , n5397 , n5409 );
nand ( n5411 , n5399 , n5407 , n5382 , n5395 );
nand ( n5412 , n5410 , n5411 );
not ( n5413 , n5412 );
not ( n5414 , n51 );
not ( n5415 , n5197 );
or ( n5416 , n5414 , n5415 );
and ( n5417 , n50 , n3834 );
not ( n5418 , n50 );
and ( n5419 , n5418 , n3833 );
nor ( n5420 , n5417 , n5419 );
nand ( n5421 , n4213 , n5420 );
nand ( n5422 , n5416 , n5421 );
not ( n5423 , n5422 );
not ( n5424 , n3894 );
not ( n5425 , n5209 );
or ( n5426 , n5424 , n5425 );
not ( n5427 , n3769 );
buf ( n5428 , n5427 );
not ( n5429 , n5428 );
and ( n5430 , n5429 , n3502 );
not ( n5431 , n5429 );
and ( n5432 , n5431 , n42 );
nor ( n5433 , n5430 , n5432 );
nand ( n5434 , n4082 , n5433 );
nand ( n5435 , n5426 , n5434 );
not ( n5436 , n5435 );
or ( n5437 , n5423 , n5436 );
not ( n5438 , n3728 );
not ( n5439 , n5251 );
or ( n5440 , n5438 , n5439 );
xnor ( n5441 , n44 , n3515 );
nand ( n5442 , n3454 , n5441 );
nand ( n5443 , n5440 , n5442 );
not ( n5444 , n5422 );
not ( n5445 , n5435 );
not ( n5446 , n5445 );
or ( n5447 , n5444 , n5446 );
not ( n5448 , n5422 );
nand ( n5449 , n5448 , n5435 );
nand ( n5450 , n5447 , n5449 );
nand ( n5451 , n5443 , n5450 );
nand ( n5452 , n5437 , n5451 );
not ( n5453 , n5452 );
or ( n5454 , n5413 , n5453 );
not ( n5455 , n5396 );
nand ( n5456 , n5408 , n5455 );
nand ( n5457 , n5454 , n5456 );
not ( n5458 , n5457 );
xor ( n5459 , n5069 , n5080 );
xor ( n5460 , n5459 , n5092 );
not ( n5461 , n5460 );
xor ( n5462 , n5033 , n5055 );
xor ( n5463 , n5462 , n5022 );
not ( n5464 , n5463 );
or ( n5465 , n5461 , n5464 );
or ( n5466 , n5463 , n5460 );
nand ( n5467 , n5465 , n5466 );
not ( n5468 , n5467 );
or ( n5469 , n5458 , n5468 );
not ( n5470 , n5463 );
nand ( n5471 , n5460 , n5470 );
nand ( n5472 , n5469 , n5471 );
xor ( n5473 , n5367 , n5472 );
xor ( n5474 , n5290 , n5317 );
xnor ( n5475 , n5473 , n5474 );
and ( n5476 , n5467 , n5457 );
not ( n5477 , n5467 );
not ( n5478 , n5457 );
and ( n5479 , n5477 , n5478 );
nor ( n5480 , n5476 , n5479 );
not ( n5481 , n5480 );
not ( n5482 , n5481 );
not ( n5483 , n5482 );
xor ( n5484 , n5279 , n5268 );
xnor ( n5485 , n5484 , n5226 );
not ( n5486 , n5485 );
xor ( n5487 , n5201 , n5211 );
xor ( n5488 , n5487 , n5223 );
not ( n5489 , n5488 );
not ( n5490 , n5255 );
xor ( n5491 , n5257 , n5490 );
xnor ( n5492 , n5491 , n5241 );
not ( n5493 , n3611 );
not ( n5494 , n46 );
not ( n5495 , n3531 );
or ( n5496 , n5494 , n5495 );
or ( n5497 , n46 , n3531 );
nand ( n5498 , n5496 , n5497 );
not ( n5499 , n5498 );
or ( n5500 , n5493 , n5499 );
nand ( n5501 , n3628 , n5406 );
nand ( n5502 , n5500 , n5501 );
not ( n5503 , n5502 );
not ( n5504 , n5381 );
not ( n5505 , n5394 );
not ( n5506 , n5505 );
or ( n5507 , n5504 , n5506 );
nand ( n5508 , n5382 , n5394 );
nand ( n5509 , n5507 , n5508 );
not ( n5510 , n5509 );
or ( n5511 , n5503 , n5510 );
or ( n5512 , n5502 , n5509 );
not ( n5513 , n3234 );
not ( n5514 , n5219 );
or ( n5515 , n5513 , n5514 );
not ( n5516 , n3229 );
not ( n5517 , n4052 );
or ( n5518 , n5516 , n5517 );
nand ( n5519 , n5518 , n4177 );
not ( n5520 , n5519 );
nand ( n5521 , n40 , n4053 );
nand ( n5522 , n5520 , n5521 );
nand ( n5523 , n5515 , n5522 );
nand ( n5524 , n5512 , n5523 );
nand ( n5525 , n5511 , n5524 );
xor ( n5526 , n5492 , n5525 );
not ( n5527 , n5526 );
or ( n5528 , n5489 , n5527 );
nand ( n5529 , n5492 , n5525 );
nand ( n5530 , n5528 , n5529 );
not ( n5531 , n5530 );
not ( n5532 , n5531 );
or ( n5533 , n5486 , n5532 );
not ( n5534 , n5485 );
nand ( n5535 , n5534 , n5530 );
nand ( n5536 , n5533 , n5535 );
not ( n5537 , n5536 );
or ( n5538 , n5483 , n5537 );
nand ( n5539 , n5485 , n5530 );
nand ( n5540 , n5538 , n5539 );
not ( n5541 , n5540 );
nand ( n5542 , n5475 , n5541 );
not ( n5543 , n3356 );
not ( n5544 , n42 );
and ( n5545 , n3 , n18 );
not ( n5546 , n3 );
and ( n5547 , n5546 , n34 );
nor ( n5548 , n5545 , n5547 );
not ( n5549 , n5548 );
or ( n5550 , n5544 , n5549 );
or ( n5551 , n42 , n3931 );
nand ( n5552 , n5550 , n5551 );
not ( n5553 , n5552 );
or ( n5554 , n5543 , n5553 );
not ( n5555 , n3348 );
not ( n5556 , n5555 );
nand ( n5557 , n5556 , n5433 );
nand ( n5558 , n5554 , n5557 );
not ( n5559 , n4213 );
not ( n5560 , n50 );
not ( n5561 , n3480 );
and ( n5562 , n5560 , n5561 );
and ( n5563 , n50 , n3480 );
nor ( n5564 , n5562 , n5563 );
not ( n5565 , n5564 );
or ( n5566 , n5559 , n5565 );
nand ( n5567 , n51 , n5420 );
nand ( n5568 , n5566 , n5567 );
not ( n5569 , n5568 );
not ( n5570 , n5569 );
nand ( n5571 , n5558 , n5570 );
not ( n5572 , n5569 );
not ( n5573 , n5558 );
not ( n5574 , n5573 );
or ( n5575 , n5572 , n5574 );
not ( n5576 , n3630 );
not ( n5577 , n5498 );
or ( n5578 , n5576 , n5577 );
xnor ( n5579 , n46 , n3748 );
nand ( n5580 , n4170 , n5579 );
nand ( n5581 , n5578 , n5580 );
nand ( n5582 , n5575 , n5581 );
nand ( n5583 , n5571 , n5582 );
not ( n5584 , n3453 );
xor ( n5585 , n44 , n3690 );
not ( n5586 , n5585 );
or ( n5587 , n5584 , n5586 );
not ( n5588 , n3725 );
not ( n5589 , n5588 );
nand ( n5590 , n5441 , n5589 );
nand ( n5591 , n5587 , n5590 );
not ( n5592 , n5591 );
nand ( n5593 , n3233 , n4051 );
not ( n5594 , n3564 );
not ( n5595 , n5594 );
and ( n5596 , n3 , n12 );
not ( n5597 , n3 );
and ( n5598 , n5597 , n28 );
nor ( n5599 , n5596 , n5598 );
not ( n5600 , n5599 );
not ( n5601 , n5600 );
not ( n5602 , n48 );
not ( n5603 , n5602 );
and ( n5604 , n5601 , n5603 );
not ( n5605 , n48 );
not ( n5606 , n3411 );
and ( n5607 , n5605 , n5606 );
nor ( n5608 , n5604 , n5607 );
not ( n5609 , n5608 );
not ( n5610 , n5609 );
or ( n5611 , n5595 , n5610 );
not ( n5612 , n5389 );
nand ( n5613 , n5612 , n3569 );
nand ( n5614 , n5611 , n5613 );
not ( n5615 , n5614 );
and ( n5616 , n5593 , n5615 );
not ( n5617 , n5593 );
and ( n5618 , n5617 , n5614 );
or ( n5619 , n5616 , n5618 );
not ( n5620 , n5619 );
not ( n5621 , n5620 );
or ( n5622 , n5592 , n5621 );
not ( n5623 , n5593 );
nand ( n5624 , n5623 , n5614 );
nand ( n5625 , n5622 , n5624 );
xor ( n5626 , n5583 , n5625 );
xor ( n5627 , n5450 , n5443 );
not ( n5628 , n5627 );
xor ( n5629 , n5626 , n5628 );
not ( n5630 , n5629 );
not ( n5631 , n5630 );
not ( n5632 , n5509 );
not ( n5633 , n5502 );
and ( n5634 , n5523 , n5633 );
not ( n5635 , n5523 );
and ( n5636 , n5635 , n5502 );
nor ( n5637 , n5634 , n5636 );
not ( n5638 , n5637 );
or ( n5639 , n5632 , n5638 );
or ( n5640 , n5637 , n5509 );
nand ( n5641 , n5639 , n5640 );
not ( n5642 , n5641 );
not ( n5643 , n4731 );
not ( n5644 , n5585 );
or ( n5645 , n5643 , n5644 );
xnor ( n5646 , n44 , n5429 );
nand ( n5647 , n3674 , n5646 );
nand ( n5648 , n5645 , n5647 );
not ( n5649 , n5648 );
not ( n5650 , n51 );
not ( n5651 , n5564 );
or ( n5652 , n5650 , n5651 );
not ( n5653 , n51 );
nand ( n5654 , n5653 , n50 );
not ( n5655 , n5654 );
not ( n5656 , n50 );
not ( n5657 , n5656 );
not ( n5658 , n3896 );
or ( n5659 , n5657 , n5658 );
nand ( n5660 , n50 , n3439 );
nand ( n5661 , n5659 , n5660 );
nand ( n5662 , n5655 , n5661 );
nand ( n5663 , n5652 , n5662 );
not ( n5664 , n5663 );
not ( n5665 , n4195 );
not ( n5666 , n42 );
not ( n5667 , n5374 );
or ( n5668 , n5666 , n5667 );
or ( n5669 , n42 , n5374 );
nand ( n5670 , n5668 , n5669 );
not ( n5671 , n5670 );
or ( n5672 , n5665 , n5671 );
nand ( n5673 , n3348 , n5552 );
nand ( n5674 , n5672 , n5673 );
not ( n5675 , n5674 );
not ( n5676 , n5675 );
or ( n5677 , n5664 , n5676 );
not ( n5678 , n5674 );
or ( n5679 , n5678 , n5663 );
nand ( n5680 , n5677 , n5679 );
not ( n5681 , n5680 );
or ( n5682 , n5649 , n5681 );
not ( n5683 , n5678 );
nand ( n5684 , n5663 , n5683 );
nand ( n5685 , n5682 , n5684 );
not ( n5686 , n5685 );
xor ( n5687 , n5591 , n5619 );
nand ( n5688 , n43 , n44 );
not ( n5689 , n5688 );
not ( n5690 , n4254 );
or ( n5691 , n5689 , n5690 );
nor ( n5692 , n43 , n44 );
not ( n5693 , n5692 );
nand ( n5694 , n5691 , n5693 );
nand ( n5695 , n5694 , n42 );
not ( n5696 , n5695 );
not ( n5697 , n5232 );
and ( n5698 , n48 , n3527 );
not ( n5699 , n48 );
and ( n5700 , n5699 , n3526 );
nor ( n5701 , n5698 , n5700 );
not ( n5702 , n5701 );
or ( n5703 , n5697 , n5702 );
not ( n5704 , n5608 );
nand ( n5705 , n4022 , n5704 );
nand ( n5706 , n5703 , n5705 );
and ( n5707 , n5696 , n5706 );
xnor ( n5708 , n5687 , n5707 );
not ( n5709 , n5708 );
or ( n5710 , n5686 , n5709 );
not ( n5711 , n5591 );
nand ( n5712 , n5711 , n5620 );
not ( n5713 , n5712 );
not ( n5714 , n5620 );
nand ( n5715 , n5591 , n5714 );
not ( n5716 , n5715 );
or ( n5717 , n5713 , n5716 );
nand ( n5718 , n5717 , n5707 );
nand ( n5719 , n5710 , n5718 );
not ( n5720 , n5719 );
not ( n5721 , n5720 );
or ( n5722 , n5642 , n5721 );
not ( n5723 , n5719 );
or ( n5724 , n5641 , n5723 );
nand ( n5725 , n5722 , n5724 );
not ( n5726 , n5725 );
or ( n5727 , n5631 , n5726 );
not ( n5728 , n5723 );
nand ( n5729 , n5641 , n5728 );
nand ( n5730 , n5727 , n5729 );
not ( n5731 , n5730 );
and ( n5732 , n5452 , n5412 );
not ( n5733 , n5452 );
not ( n5734 , n5412 );
and ( n5735 , n5733 , n5734 );
nor ( n5736 , n5732 , n5735 );
not ( n5737 , n5627 );
not ( n5738 , n5626 );
or ( n5739 , n5737 , n5738 );
nand ( n5740 , n5583 , n5625 );
nand ( n5741 , n5739 , n5740 );
not ( n5742 , n5741 );
xor ( n5743 , n5736 , n5742 );
xor ( n5744 , n5526 , n5488 );
xnor ( n5745 , n5743 , n5744 );
not ( n5746 , n5745 );
nand ( n5747 , n5731 , n5746 );
and ( n5748 , n5536 , n5480 );
not ( n5749 , n5536 );
and ( n5750 , n5749 , n5481 );
nor ( n5751 , n5748 , n5750 );
not ( n5752 , n5744 );
not ( n5753 , n5736 );
not ( n5754 , n5753 );
not ( n5755 , n5741 );
or ( n5756 , n5754 , n5755 );
or ( n5757 , n5753 , n5741 );
nand ( n5758 , n5756 , n5757 );
not ( n5759 , n5758 );
or ( n5760 , n5752 , n5759 );
not ( n5761 , n5753 );
nand ( n5762 , n5761 , n5741 );
nand ( n5763 , n5760 , n5762 );
nor ( n5764 , n5751 , n5763 );
not ( n5765 , n5764 );
and ( n5766 , n5542 , n5747 , n5765 );
not ( n5767 , n5570 );
not ( n5768 , n5558 );
not ( n5769 , n5768 );
or ( n5770 , n5767 , n5769 );
or ( n5771 , n5570 , n5768 );
nand ( n5772 , n5770 , n5771 );
xor ( n5773 , n5581 , n5772 );
not ( n5774 , n5773 );
not ( n5775 , n4254 );
nand ( n5776 , n5775 , n3348 );
buf ( n5777 , n5776 );
not ( n5778 , n5777 );
not ( n5779 , n5778 );
not ( n5780 , n4248 );
not ( n5781 , n5780 );
not ( n5782 , n5646 );
or ( n5783 , n5781 , n5782 );
not ( n5784 , n44 );
not ( n5785 , n5784 );
not ( n5786 , n5548 );
not ( n5787 , n5786 );
or ( n5788 , n5785 , n5787 );
not ( n5789 , n44 );
not ( n5790 , n5548 );
or ( n5791 , n5789 , n5790 );
nand ( n5792 , n5788 , n5791 );
nand ( n5793 , n3674 , n5792 );
nand ( n5794 , n5783 , n5793 );
not ( n5795 , n5794 );
or ( n5796 , n5779 , n5795 );
not ( n5797 , n5777 );
not ( n5798 , n5794 );
not ( n5799 , n5798 );
or ( n5800 , n5797 , n5799 );
not ( n5801 , n4030 );
not ( n5802 , n5801 );
xnor ( n5803 , n3412 , n50 );
not ( n5804 , n5803 );
or ( n5805 , n5802 , n5804 );
nand ( n5806 , n51 , n5661 );
nand ( n5807 , n5805 , n5806 );
nand ( n5808 , n5800 , n5807 );
nand ( n5809 , n5796 , n5808 );
not ( n5810 , n5809 );
not ( n5811 , n3611 );
xnor ( n5812 , n46 , n3515 );
not ( n5813 , n5812 );
or ( n5814 , n5811 , n5813 );
nand ( n5815 , n3628 , n5579 );
nand ( n5816 , n5814 , n5815 );
not ( n5817 , n5816 );
xor ( n5818 , n5696 , n5706 );
not ( n5819 , n5818 );
not ( n5820 , n5819 );
or ( n5821 , n5817 , n5820 );
not ( n5822 , n5816 );
nand ( n5823 , n5822 , n5818 );
nand ( n5824 , n5821 , n5823 );
not ( n5825 , n5824 );
or ( n5826 , n5810 , n5825 );
nand ( n5827 , n5816 , n5818 );
nand ( n5828 , n5826 , n5827 );
not ( n5829 , n5828 );
not ( n5830 , n5829 );
or ( n5831 , n5774 , n5830 );
not ( n5832 , n5828 );
or ( n5833 , n5773 , n5832 );
nand ( n5834 , n5831 , n5833 );
not ( n5835 , n5834 );
not ( n5836 , n5685 );
and ( n5837 , n5708 , n5836 );
not ( n5838 , n5708 );
and ( n5839 , n5838 , n5685 );
nor ( n5840 , n5837 , n5839 );
not ( n5841 , n5840 );
not ( n5842 , n5841 );
or ( n5843 , n5835 , n5842 );
not ( n5844 , n5832 );
nand ( n5845 , n5773 , n5844 );
nand ( n5846 , n5843 , n5845 );
not ( n5847 , n5846 );
not ( n5848 , n5629 );
not ( n5849 , n5725 );
or ( n5850 , n5848 , n5849 );
or ( n5851 , n5629 , n5725 );
nand ( n5852 , n5850 , n5851 );
not ( n5853 , n5852 );
nand ( n5854 , n5847 , n5853 );
not ( n5855 , n5854 );
not ( n5856 , n5834 );
not ( n5857 , n5840 );
and ( n5858 , n5856 , n5857 );
and ( n5859 , n5834 , n5840 );
nor ( n5860 , n5858 , n5859 );
not ( n5861 , n5860 );
not ( n5862 , n5824 );
xnor ( n5863 , n5862 , n5809 );
not ( n5864 , n5863 );
nand ( n5865 , n45 , n46 );
not ( n5866 , n5865 );
nor ( n5867 , n45 , n46 );
not ( n5868 , n5867 );
not ( n5869 , n5868 );
not ( n5870 , n4227 );
or ( n5871 , n5869 , n5870 );
nand ( n5872 , n5871 , n44 );
nor ( n5873 , n5866 , n5872 );
not ( n5874 , n51 );
not ( n5875 , n5803 );
or ( n5876 , n5874 , n5875 );
xnor ( n5877 , n50 , n5066 );
nand ( n5878 , n4213 , n5877 );
nand ( n5879 , n5876 , n5878 );
nand ( n5880 , n5873 , n5879 );
not ( n5881 , n5880 );
not ( n5882 , n5881 );
not ( n5883 , n4016 );
not ( n5884 , n48 );
not ( n5885 , n5884 );
not ( n5886 , n5247 );
not ( n5887 , n5886 );
or ( n5888 , n5885 , n5887 );
not ( n5889 , n48 );
or ( n5890 , n5889 , n3747 );
nand ( n5891 , n5888 , n5890 );
not ( n5892 , n5891 );
or ( n5893 , n5883 , n5892 );
nand ( n5894 , n4022 , n5701 );
nand ( n5895 , n5893 , n5894 );
not ( n5896 , n3982 );
not ( n5897 , n5896 );
xor ( n5898 , n46 , n3690 );
not ( n5899 , n5898 );
or ( n5900 , n5897 , n5899 );
not ( n5901 , n3627 );
nand ( n5902 , n5812 , n5901 );
nand ( n5903 , n5900 , n5902 );
and ( n5904 , n5895 , n5903 );
not ( n5905 , n5895 );
not ( n5906 , n5903 );
and ( n5907 , n5905 , n5906 );
nor ( n5908 , n5904 , n5907 );
not ( n5909 , n5908 );
or ( n5910 , n5882 , n5909 );
not ( n5911 , n5906 );
nand ( n5912 , n5895 , n5911 );
nand ( n5913 , n5910 , n5912 );
not ( n5914 , n5913 );
not ( n5915 , n5914 );
not ( n5916 , n5648 );
not ( n5917 , n5916 );
not ( n5918 , n5680 );
or ( n5919 , n5917 , n5918 );
not ( n5920 , n5648 );
or ( n5921 , n5920 , n5680 );
nand ( n5922 , n5919 , n5921 );
not ( n5923 , n5922 );
and ( n5924 , n5915 , n5923 );
not ( n5925 , n5913 );
and ( n5926 , n5925 , n5922 );
nor ( n5927 , n5924 , n5926 );
not ( n5928 , n5927 );
not ( n5929 , n5928 );
or ( n5930 , n5864 , n5929 );
not ( n5931 , n5925 );
nand ( n5932 , n5931 , n5922 );
nand ( n5933 , n5930 , n5932 );
nand ( n5934 , n5861 , n5933 );
nand ( n5935 , n5852 , n5846 );
xor ( n5936 , n5908 , n5881 );
not ( n5937 , n5936 );
not ( n5938 , n4017 );
and ( n5939 , n48 , n3517 );
not ( n5940 , n48 );
and ( n5941 , n5940 , n3516 );
or ( n5942 , n5939 , n5941 );
not ( n5943 , n5942 );
or ( n5944 , n5938 , n5943 );
nand ( n5945 , n4023 , n5891 );
nand ( n5946 , n5944 , n5945 );
not ( n5947 , n5946 );
not ( n5948 , n5901 );
not ( n5949 , n5898 );
or ( n5950 , n5948 , n5949 );
not ( n5951 , n46 );
not ( n5952 , n5951 );
not ( n5953 , n3770 );
or ( n5954 , n5952 , n5953 );
not ( n5955 , n46 );
or ( n5956 , n5955 , n5428 );
nand ( n5957 , n5954 , n5956 );
nand ( n5958 , n5896 , n5957 );
nand ( n5959 , n5950 , n5958 );
not ( n5960 , n5959 );
not ( n5961 , n3452 );
and ( n5962 , n5373 , n44 );
not ( n5963 , n5373 );
not ( n5964 , n44 );
and ( n5965 , n5963 , n5964 );
nor ( n5966 , n5962 , n5965 );
not ( n5967 , n5966 );
or ( n5968 , n5961 , n5967 );
nand ( n5969 , n3465 , n5792 );
nand ( n5970 , n5968 , n5969 );
not ( n5971 , n5970 );
not ( n5972 , n5971 );
or ( n5973 , n5960 , n5972 );
not ( n5974 , n5970 );
or ( n5975 , n5959 , n5974 );
nand ( n5976 , n5973 , n5975 );
not ( n5977 , n5976 );
or ( n5978 , n5947 , n5977 );
not ( n5979 , n5974 );
nand ( n5980 , n5959 , n5979 );
nand ( n5981 , n5978 , n5980 );
not ( n5982 , n5981 );
xor ( n5983 , n5776 , n5807 );
xnor ( n5984 , n5983 , n5794 );
and ( n5985 , n5982 , n5984 );
not ( n5986 , n5982 );
not ( n5987 , n5984 );
and ( n5988 , n5986 , n5987 );
nor ( n5989 , n5985 , n5988 );
not ( n5990 , n5989 );
not ( n5991 , n5990 );
or ( n5992 , n5937 , n5991 );
nand ( n5993 , n5984 , n5981 );
nand ( n5994 , n5992 , n5993 );
not ( n5995 , n5994 );
not ( n5996 , n5863 );
not ( n5997 , n5927 );
or ( n5998 , n5996 , n5997 );
or ( n5999 , n5863 , n5927 );
nand ( n6000 , n5998 , n5999 );
not ( n6001 , n6000 );
or ( n6002 , n5995 , n6001 );
xor ( n6003 , n5976 , n5946 );
not ( n6004 , n6003 );
not ( n6005 , n5228 );
not ( n6006 , n5942 );
or ( n6007 , n6005 , n6006 );
not ( n6008 , n48 );
not ( n6009 , n3851 );
or ( n6010 , n6008 , n6009 );
not ( n6011 , n48 );
nand ( n6012 , n6011 , n3690 );
nand ( n6013 , n6010 , n6012 );
buf ( n6014 , n6013 );
nand ( n6015 , n3566 , n6014 );
nand ( n6016 , n6007 , n6015 );
not ( n6017 , n6016 );
and ( n6018 , n3466 , n4227 );
not ( n6019 , n6018 );
not ( n6020 , n51 );
not ( n6021 , n5877 );
or ( n6022 , n6020 , n6021 );
not ( n6023 , n50 );
not ( n6024 , n6023 );
not ( n6025 , n5886 );
or ( n6026 , n6024 , n6025 );
not ( n6027 , n50 );
or ( n6028 , n6027 , n3747 );
nand ( n6029 , n6026 , n6028 );
nand ( n6030 , n4888 , n6029 );
nand ( n6031 , n6022 , n6030 );
not ( n6032 , n6031 );
not ( n6033 , n6032 );
or ( n6034 , n6019 , n6033 );
nor ( n6035 , n3726 , n4052 );
not ( n6036 , n6035 );
nand ( n6037 , n6036 , n6031 );
nand ( n6038 , n6034 , n6037 );
not ( n6039 , n6038 );
or ( n6040 , n6017 , n6039 );
nand ( n6041 , n6018 , n6031 );
nand ( n6042 , n6040 , n6041 );
not ( n6043 , n6042 );
not ( n6044 , n6043 );
nand ( n6045 , n5868 , n4227 );
nand ( n6046 , n5865 , n44 , n6045 );
not ( n6047 , n6046 );
not ( n6048 , n5879 );
and ( n6049 , n6047 , n6048 );
and ( n6050 , n6046 , n5879 );
nor ( n6051 , n6049 , n6050 );
not ( n6052 , n6051 );
and ( n6053 , n6044 , n6052 );
not ( n6054 , n6044 );
and ( n6055 , n6054 , n6051 );
nor ( n6056 , n6053 , n6055 );
not ( n6057 , n6056 );
or ( n6058 , n6004 , n6057 );
not ( n6059 , n6051 );
nand ( n6060 , n6059 , n6044 );
nand ( n6061 , n6058 , n6060 );
not ( n6062 , n6061 );
not ( n6063 , n5989 );
not ( n6064 , n5936 );
and ( n6065 , n6063 , n6064 );
and ( n6066 , n5936 , n5989 );
nor ( n6067 , n6065 , n6066 );
nor ( n6068 , n6062 , n6067 );
not ( n6069 , n6068 );
nand ( n6070 , n6002 , n6069 );
nor ( n6071 , n6000 , n5994 );
not ( n6072 , n6071 );
not ( n6073 , n5933 );
nand ( n6074 , n6073 , n5860 );
nand ( n6075 , n6070 , n6072 , n6074 );
nand ( n6076 , n5934 , n5935 , n6075 );
not ( n6077 , n6076 );
or ( n6078 , n5855 , n6077 );
not ( n6079 , n6074 );
not ( n6080 , n6079 );
not ( n6081 , n3779 );
not ( n6082 , n46 );
not ( n6083 , n6082 );
not ( n6084 , n3932 );
or ( n6085 , n6083 , n6084 );
not ( n6086 , n46 );
not ( n6087 , n3931 );
or ( n6088 , n6086 , n6087 );
nand ( n6089 , n6085 , n6088 );
not ( n6090 , n6089 );
or ( n6091 , n6081 , n6090 );
nand ( n6092 , n3782 , n5957 );
nand ( n6093 , n6091 , n6092 );
not ( n6094 , n6093 );
not ( n6095 , n6094 );
nand ( n6096 , n47 , n48 );
not ( n6097 , n6096 );
nor ( n6098 , n47 , n48 );
not ( n6099 , n6098 );
not ( n6100 , n6099 );
not ( n6101 , n4051 );
or ( n6102 , n6100 , n6101 );
nand ( n6103 , n6102 , n46 );
nor ( n6104 , n6097 , n6103 );
not ( n6105 , n51 );
not ( n6106 , n6029 );
or ( n6107 , n6105 , n6106 );
xnor ( n6108 , n50 , n3514 );
nand ( n6109 , n5801 , n6108 );
nand ( n6110 , n6107 , n6109 );
nand ( n6111 , n6104 , n6110 );
not ( n6112 , n6111 );
not ( n6113 , n6112 );
and ( n6114 , n6095 , n6113 );
not ( n6115 , n6093 );
not ( n6116 , n6111 );
and ( n6117 , n6115 , n6116 );
nor ( n6118 , n6114 , n6117 );
not ( n6119 , n6118 );
not ( n6120 , n6119 );
not ( n6121 , n6016 );
not ( n6122 , n6121 );
not ( n6123 , n6038 );
or ( n6124 , n6122 , n6123 );
or ( n6125 , n6121 , n6038 );
nand ( n6126 , n6124 , n6125 );
not ( n6127 , n6126 );
or ( n6128 , n6120 , n6127 );
not ( n6129 , n6115 );
nand ( n6130 , n6129 , n6116 );
nand ( n6131 , n6128 , n6130 );
not ( n6132 , n6131 );
xor ( n6133 , n6051 , n6043 );
xnor ( n6134 , n6133 , n6003 );
nand ( n6135 , n6132 , n6134 );
not ( n6136 , n6135 );
not ( n6137 , n6104 );
not ( n6138 , n6110 );
not ( n6139 , n6138 );
and ( n6140 , n6137 , n6139 );
and ( n6141 , n6104 , n6138 );
nor ( n6142 , n6140 , n6141 );
not ( n6143 , n6142 );
not ( n6144 , n6143 );
not ( n6145 , n3611 );
not ( n6146 , n46 );
not ( n6147 , n4254 );
or ( n6148 , n6146 , n6147 );
or ( n6149 , n46 , n4226 );
nand ( n6150 , n6148 , n6149 );
not ( n6151 , n6150 );
or ( n6152 , n6145 , n6151 );
nand ( n6153 , n3628 , n6089 );
nand ( n6154 , n6152 , n6153 );
not ( n6155 , n4016 );
not ( n6156 , n48 );
not ( n6157 , n3771 );
or ( n6158 , n6156 , n6157 );
not ( n6159 , n48 );
nand ( n6160 , n6159 , n5428 );
nand ( n6161 , n6158 , n6160 );
not ( n6162 , n6161 );
or ( n6163 , n6155 , n6162 );
not ( n6164 , n3570 );
nand ( n6165 , n6164 , n6013 );
nand ( n6166 , n6163 , n6165 );
and ( n6167 , n6154 , n6166 );
not ( n6168 , n6154 );
not ( n6169 , n6166 );
and ( n6170 , n6168 , n6169 );
nor ( n6171 , n6167 , n6170 );
not ( n6172 , n6171 );
or ( n6173 , n6144 , n6172 );
not ( n6174 , n6169 );
nand ( n6175 , n6174 , n6154 );
nand ( n6176 , n6173 , n6175 );
not ( n6177 , n6176 );
not ( n6178 , n6118 );
not ( n6179 , n6126 );
and ( n6180 , n6178 , n6179 );
and ( n6181 , n6118 , n6126 );
nor ( n6182 , n6180 , n6181 );
nand ( n6183 , n6177 , n6182 );
not ( n6184 , n6183 );
not ( n6185 , n5085 );
and ( n6186 , n48 , n3931 );
not ( n6187 , n48 );
and ( n6188 , n6187 , n3932 );
or ( n6189 , n6186 , n6188 );
not ( n6190 , n6189 );
or ( n6191 , n6185 , n6190 );
not ( n6192 , n6161 );
or ( n6193 , n3571 , n6192 );
nand ( n6194 , n6191 , n6193 );
not ( n6195 , n6194 );
not ( n6196 , n5654 );
not ( n6197 , n6196 );
not ( n6198 , n50 );
not ( n6199 , n6198 );
not ( n6200 , n16 );
and ( n6201 , n3 , n6200 );
not ( n6202 , n3 );
not ( n6203 , n32 );
and ( n6204 , n6202 , n6203 );
nor ( n6205 , n6201 , n6204 );
not ( n6206 , n6205 );
or ( n6207 , n6199 , n6206 );
not ( n6208 , n50 );
or ( n6209 , n6208 , n6205 );
nand ( n6210 , n6207 , n6209 );
not ( n6211 , n6210 );
or ( n6212 , n6197 , n6211 );
nand ( n6213 , n51 , n6108 );
nand ( n6214 , n6212 , n6213 );
not ( n6215 , n5373 );
nor ( n6216 , n6215 , n3627 );
xnor ( n6217 , n6214 , n6216 );
not ( n6218 , n6217 );
not ( n6219 , n6218 );
or ( n6220 , n6195 , n6219 );
nand ( n6221 , n6216 , n6214 );
nand ( n6222 , n6220 , n6221 );
not ( n6223 , n6222 );
not ( n6224 , n6142 );
not ( n6225 , n6171 );
and ( n6226 , n6224 , n6225 );
and ( n6227 , n6142 , n6171 );
nor ( n6228 , n6226 , n6227 );
nand ( n6229 , n6223 , n6228 );
not ( n6230 , n6229 );
nand ( n6231 , n49 , n50 );
not ( n6232 , n6231 );
not ( n6233 , n5374 );
or ( n6234 , n6232 , n6233 );
nor ( n6235 , n49 , n50 );
not ( n6236 , n6235 );
nand ( n6237 , n6234 , n6236 );
nand ( n6238 , n6237 , n48 );
not ( n6239 , n6238 );
not ( n6240 , n51 );
not ( n6241 , n6210 );
or ( n6242 , n6240 , n6241 );
not ( n6243 , n50 );
not ( n6244 , n6243 );
not ( n6245 , n5427 );
or ( n6246 , n6244 , n6245 );
not ( n6247 , n50 );
or ( n6248 , n3770 , n6247 );
nand ( n6249 , n6246 , n6248 );
nand ( n6250 , n6196 , n6249 );
nand ( n6251 , n6242 , n6250 );
nand ( n6252 , n6239 , n6251 );
not ( n6253 , n6252 );
not ( n6254 , n6217 );
not ( n6255 , n6194 );
and ( n6256 , n6254 , n6255 );
and ( n6257 , n6194 , n6217 );
nor ( n6258 , n6256 , n6257 );
not ( n6259 , n6258 );
nand ( n6260 , n6253 , n6259 );
nand ( n6261 , n6258 , n6252 );
nand ( n6262 , n5228 , n4053 );
not ( n6263 , n6262 );
not ( n6264 , n4030 );
not ( n6265 , n6264 );
not ( n6266 , n5786 );
not ( n6267 , n50 );
not ( n6268 , n6267 );
and ( n6269 , n6266 , n6268 );
not ( n6270 , n50 );
and ( n6271 , n6270 , n5790 );
nor ( n6272 , n6269 , n6271 );
nand ( n6273 , n6265 , n6272 );
nand ( n6274 , n50 , n4255 , n6273 );
not ( n6275 , n6274 );
or ( n6276 , n6263 , n6275 );
not ( n6277 , n5801 );
or ( n6278 , n6277 , n6272 );
not ( n6279 , n51 );
not ( n6280 , n6249 );
or ( n6281 , n6279 , n6280 );
nand ( n6282 , n6278 , n6281 );
nand ( n6283 , n6276 , n6282 );
not ( n6284 , n6283 );
not ( n6285 , n4016 );
not ( n6286 , n48 );
not ( n6287 , n4254 );
or ( n6288 , n6286 , n6287 );
or ( n6289 , n48 , n4226 );
nand ( n6290 , n6288 , n6289 );
not ( n6291 , n6290 );
or ( n6292 , n6285 , n6291 );
not ( n6293 , n3570 );
nand ( n6294 , n6293 , n6189 );
nand ( n6295 , n6292 , n6294 );
not ( n6296 , n6295 );
not ( n6297 , n6238 );
not ( n6298 , n6251 );
and ( n6299 , n6297 , n6298 );
and ( n6300 , n6238 , n6251 );
nor ( n6301 , n6299 , n6300 );
nand ( n6302 , n6296 , n6301 );
nand ( n6303 , n6284 , n6302 );
not ( n6304 , n6301 );
nand ( n6305 , n6295 , n6304 );
nand ( n6306 , n6303 , n6305 );
nand ( n6307 , n6261 , n6306 );
nand ( n6308 , n6260 , n6307 );
not ( n6309 , n6308 );
or ( n6310 , n6230 , n6309 );
not ( n6311 , n6223 );
not ( n6312 , n6228 );
nand ( n6313 , n6311 , n6312 );
nand ( n6314 , n6310 , n6313 );
not ( n6315 , n6314 );
or ( n6316 , n6184 , n6315 );
not ( n6317 , n6177 );
not ( n6318 , n6182 );
nand ( n6319 , n6317 , n6318 );
nand ( n6320 , n6316 , n6319 );
not ( n6321 , n6320 );
or ( n6322 , n6136 , n6321 );
not ( n6323 , n6132 );
not ( n6324 , n6134 );
nand ( n6325 , n6323 , n6324 );
nand ( n6326 , n6322 , n6325 );
not ( n6327 , n6067 );
nor ( n6328 , n6061 , n6327 );
nor ( n6329 , n6071 , n6328 );
nand ( n6330 , n6326 , n6329 );
not ( n6331 , n6330 );
nand ( n6332 , n5854 , n6080 , n6331 );
nand ( n6333 , n6078 , n6332 );
xor ( n6334 , n5193 , n5323 );
xnor ( n6335 , n6334 , n5190 );
not ( n6336 , n5474 );
and ( n6337 , n5472 , n5367 );
not ( n6338 , n5472 );
not ( n6339 , n5367 );
and ( n6340 , n6338 , n6339 );
nor ( n6341 , n6337 , n6340 );
not ( n6342 , n6341 );
or ( n6343 , n6336 , n6342 );
not ( n6344 , n6339 );
nand ( n6345 , n6344 , n5472 );
nand ( n6346 , n6343 , n6345 );
not ( n6347 , n6346 );
nand ( n6348 , n6335 , n6347 );
nand ( n6349 , n5766 , n6333 , n6348 );
not ( n6350 , n5541 );
not ( n6351 , n5475 );
nand ( n6352 , n6350 , n6351 );
not ( n6353 , n6352 );
nand ( n6354 , n5745 , n5730 );
or ( n6355 , n6354 , n5764 );
not ( n6356 , n5763 );
not ( n6357 , n6356 );
nand ( n6358 , n6357 , n5751 );
nand ( n6359 , n6355 , n6358 );
nand ( n6360 , n6359 , n5542 );
not ( n6361 , n6360 );
or ( n6362 , n6353 , n6361 );
nand ( n6363 , n6362 , n6348 );
not ( n6364 , n6347 );
not ( n6365 , n6335 );
nand ( n6366 , n6364 , n6365 );
nand ( n6367 , n6349 , n6363 , n6366 );
nand ( n6368 , n4981 , n4815 );
nor ( n6369 , n5341 , n5335 );
not ( n6370 , n6369 );
nand ( n6371 , n5184 , n5187 );
nand ( n6372 , n6370 , n6371 );
nor ( n6373 , n6368 , n6372 );
and ( n6374 , n6367 , n6373 );
nand ( n6375 , n4644 , n4636 );
and ( n6376 , n4515 , n6375 , n5357 );
nand ( n6377 , n6374 , n6376 , n4763 );
nand ( n6378 , n4766 , n5365 , n6377 );
not ( n6379 , n6378 );
not ( n6380 , n6379 );
nand ( n6381 , n3338 , n3404 );
buf ( n6382 , n6381 );
xor ( n6383 , n3341 , n3401 );
not ( n6384 , n3145 );
not ( n6385 , n3371 );
not ( n6386 , n6385 );
and ( n6387 , n6384 , n6386 );
not ( n6388 , n3124 );
nor ( n6389 , n6388 , n4671 );
nor ( n6390 , n6387 , n6389 );
buf ( n6391 , n6390 );
not ( n6392 , n3788 );
not ( n6393 , n4728 );
or ( n6394 , n6392 , n6393 );
nand ( n6395 , n42 , n3350 );
nand ( n6396 , n6394 , n6395 );
not ( n6397 , n6396 );
not ( n6398 , n4549 );
not ( n6399 , n6398 );
and ( n6400 , n6399 , n36 );
not ( n6401 , n6400 );
and ( n6402 , n6397 , n6401 );
not ( n6403 , n6397 );
and ( n6404 , n6403 , n6400 );
nor ( n6405 , n6402 , n6404 );
not ( n6406 , n6405 );
or ( n6407 , n6391 , n6406 );
or ( n6408 , n6401 , n6397 );
nand ( n6409 , n6407 , n6408 );
not ( n6410 , n6409 );
not ( n6411 , n6410 );
not ( n6412 , n3385 );
not ( n6413 , n3392 );
not ( n6414 , n6413 );
or ( n6415 , n6412 , n6414 );
not ( n6416 , n3385 );
nand ( n6417 , n6416 , n3392 );
nand ( n6418 , n6415 , n6417 );
not ( n6419 , n6418 );
not ( n6420 , n6419 );
and ( n6421 , n6411 , n6420 );
not ( n6422 , n3092 );
buf ( n6423 , n3507 );
and ( n6424 , n6423 , n3096 );
not ( n6425 , n6423 );
and ( n6426 , n6425 , n38 );
nor ( n6427 , n6424 , n6426 );
not ( n6428 , n6427 );
or ( n6429 , n6422 , n6428 );
or ( n6430 , n3114 , n3289 );
nand ( n6431 , n6429 , n6430 );
buf ( n6432 , n4670 );
not ( n6433 , n6432 );
xor ( n6434 , n6431 , n6433 );
not ( n6435 , n4685 );
not ( n6436 , n3225 );
or ( n6437 , n6435 , n6436 );
nand ( n6438 , n3317 , n3380 );
nand ( n6439 , n6437 , n6438 );
buf ( n6440 , n6439 );
and ( n6441 , n6434 , n6440 );
not ( n6442 , n6434 );
not ( n6443 , n6440 );
and ( n6444 , n6442 , n6443 );
nor ( n6445 , n6441 , n6444 );
and ( n6446 , n6418 , n6409 );
not ( n6447 , n6418 );
and ( n6448 , n6447 , n6410 );
or ( n6449 , n6446 , n6448 );
not ( n6450 , n6449 );
and ( n6451 , n6445 , n6450 );
nor ( n6452 , n6421 , n6451 );
not ( n6453 , n3346 );
and ( n6454 , n3398 , n6453 );
not ( n6455 , n3398 );
and ( n6456 , n6455 , n3346 );
nor ( n6457 , n6454 , n6456 );
and ( n6458 , n6440 , n6434 );
not ( n6459 , n6432 );
and ( n6460 , n6459 , n6431 );
nor ( n6461 , n6458 , n6460 );
xnor ( n6462 , n6457 , n6461 );
or ( n6463 , n6452 , n6462 );
or ( n6464 , n6461 , n6457 );
nand ( n6465 , n6463 , n6464 );
or ( n6466 , n6383 , n6465 );
not ( n6467 , n4676 );
not ( n6468 , n6467 );
not ( n6469 , n4690 );
or ( n6470 , n6468 , n6469 );
nand ( n6471 , n4679 , n4689 );
nand ( n6472 , n6470 , n6471 );
not ( n6473 , n4416 );
not ( n6474 , n6427 );
or ( n6475 , n6473 , n6474 );
not ( n6476 , n4743 );
or ( n6477 , n3093 , n6476 );
nand ( n6478 , n6475 , n6477 );
not ( n6479 , n6439 );
and ( n6480 , n6478 , n6479 );
not ( n6481 , n6478 );
and ( n6482 , n6481 , n6439 );
nor ( n6483 , n6480 , n6482 );
xor ( n6484 , n6472 , n6483 );
not ( n6485 , n6484 );
not ( n6486 , n4730 );
not ( n6487 , n4747 );
or ( n6488 , n6486 , n6487 );
nand ( n6489 , n4737 , n4746 );
nand ( n6490 , n6488 , n6489 );
not ( n6491 , n6490 );
not ( n6492 , n6391 );
not ( n6493 , n6405 );
or ( n6494 , n6492 , n6493 );
or ( n6495 , n6391 , n6405 );
nand ( n6496 , n6494 , n6495 );
xor ( n6497 , n6491 , n6496 );
or ( n6498 , n6485 , n6497 );
not ( n6499 , n6496 );
or ( n6500 , n6491 , n6499 );
nand ( n6501 , n6498 , n6500 );
and ( n6502 , n6483 , n6472 );
and ( n6503 , n6443 , n6478 );
nor ( n6504 , n6502 , n6503 );
not ( n6505 , n6504 );
not ( n6506 , n6445 );
not ( n6507 , n6449 );
or ( n6508 , n6506 , n6507 );
or ( n6509 , n6445 , n6449 );
nand ( n6510 , n6508 , n6509 );
not ( n6511 , n6510 );
or ( n6512 , n6505 , n6511 );
or ( n6513 , n6504 , n6510 );
nand ( n6514 , n6512 , n6513 );
and ( n6515 , n6501 , n6514 );
not ( n6516 , n6504 );
and ( n6517 , n6516 , n6510 );
nor ( n6518 , n6515 , n6517 );
xnor ( n6519 , n6452 , n6462 );
nand ( n6520 , n6518 , n6519 );
not ( n6521 , n4694 );
not ( n6522 , n4707 );
or ( n6523 , n6521 , n6522 );
nand ( n6524 , n4608 , n4703 );
nand ( n6525 , n6523 , n6524 );
not ( n6526 , n6525 );
not ( n6527 , n6484 );
not ( n6528 , n6497 );
and ( n6529 , n6527 , n6528 );
and ( n6530 , n6484 , n6497 );
nor ( n6531 , n6529 , n6530 );
or ( n6532 , n6526 , n6531 );
not ( n6533 , n4752 );
or ( n6534 , n6533 , n4712 );
not ( n6535 , n4718 );
or ( n6536 , n6535 , n4748 );
nand ( n6537 , n6534 , n6536 );
not ( n6538 , n6525 );
not ( n6539 , n6531 );
or ( n6540 , n6538 , n6539 );
or ( n6541 , n6525 , n6531 );
nand ( n6542 , n6540 , n6541 );
nand ( n6543 , n6537 , n6542 );
nand ( n6544 , n6532 , n6543 );
not ( n6545 , n6544 );
xnor ( n6546 , n6501 , n6514 );
nand ( n6547 , n6545 , n6546 );
xor ( n6548 , n6537 , n6542 );
not ( n6549 , n6548 );
not ( n6550 , n4656 );
not ( n6551 , n4760 );
or ( n6552 , n6550 , n6551 );
not ( n6553 , n4756 );
nand ( n6554 , n4662 , n6553 );
nand ( n6555 , n6552 , n6554 );
not ( n6556 , n6555 );
nand ( n6557 , n6549 , n6556 );
and ( n6558 , n6547 , n6557 );
and ( n6559 , n6520 , n6558 );
nand ( n6560 , n6380 , n6382 , n6466 , n6559 );
not ( n6561 , n6466 );
not ( n6562 , n6520 );
not ( n6563 , n6546 );
nand ( n6564 , n6544 , n6563 );
and ( n6565 , n6548 , n6555 );
nand ( n6566 , n6547 , n6565 );
nand ( n6567 , n6564 , n6566 );
not ( n6568 , n6567 );
or ( n6569 , n6562 , n6568 );
not ( n6570 , n6519 );
not ( n6571 , n6518 );
nand ( n6572 , n6570 , n6571 );
nand ( n6573 , n6569 , n6572 );
not ( n6574 , n6573 );
or ( n6575 , n6561 , n6574 );
nand ( n6576 , n6383 , n6465 );
nand ( n6577 , n6575 , n6576 );
nand ( n6578 , n6577 , n6382 );
nand ( n6579 , n3406 , n6560 , n6578 );
not ( n6580 , n6579 );
or ( n6581 , n3337 , n6580 );
nand ( n6582 , n6581 , n2 );
not ( n6583 , n3337 );
nor ( n6584 , n6583 , n6579 );
or ( n6585 , n6582 , n6584 );
or ( n6586 , n36 , n55 );
nand ( n6587 , n36 , n55 );
nand ( n6588 , n6586 , n6587 );
not ( n6589 , n36 );
not ( n6590 , n4223 );
or ( n6591 , n6589 , n6590 );
not ( n6592 , n36 );
nand ( n6593 , n6592 , n38 , n37 );
nand ( n6594 , n6591 , n6593 );
not ( n6595 , n6594 );
not ( n6596 , n6595 );
not ( n6597 , n6596 );
not ( n6598 , n6597 );
not ( n6599 , n6598 );
or ( n6600 , n6588 , n6599 );
not ( n6601 , n3144 );
or ( n6602 , n36 , n54 );
nand ( n6603 , n36 , n54 );
nand ( n6604 , n6602 , n6603 );
or ( n6605 , n6601 , n6604 );
nand ( n6606 , n6600 , n6605 );
not ( n6607 , n3229 );
not ( n6608 , n3318 );
and ( n6609 , n6607 , n6608 );
not ( n6610 , n42 );
nand ( n6611 , n6610 , n41 );
not ( n6612 , n41 );
nand ( n6613 , n6612 , n42 );
and ( n6614 , n6611 , n6613 , n3218 );
buf ( n6615 , n6614 );
buf ( n6616 , n6615 );
not ( n6617 , n6616 );
not ( n6618 , n6617 );
and ( n6619 , n40 , n52 );
not ( n6620 , n40 );
not ( n6621 , n52 );
and ( n6622 , n6620 , n6621 );
nor ( n6623 , n6619 , n6622 );
and ( n6624 , n6618 , n6623 );
nor ( n6625 , n6609 , n6624 );
not ( n6626 , n6625 );
and ( n6627 , n6606 , n6626 );
not ( n6628 , n6606 );
and ( n6629 , n6628 , n6625 );
nor ( n6630 , n6627 , n6629 );
not ( n6631 , n38 );
not ( n6632 , n54 );
and ( n6633 , n6631 , n6632 );
and ( n6634 , n38 , n54 );
nor ( n6635 , n6633 , n6634 );
xnor ( n6636 , n38 , n39 );
nor ( n6637 , n6636 , n3087 );
buf ( n6638 , n6637 );
buf ( n6639 , n6638 );
not ( n6640 , n6639 );
not ( n6641 , n6640 );
and ( n6642 , n6635 , n6641 );
not ( n6643 , n53 );
and ( n6644 , n3096 , n6643 );
and ( n6645 , n38 , n53 );
nor ( n6646 , n6644 , n6645 );
and ( n6647 , n4525 , n6646 );
nor ( n6648 , n6642 , n6647 );
nand ( n6649 , n36 , n57 );
xor ( n6650 , n36 , n56 );
not ( n6651 , n6650 );
not ( n6652 , n6598 );
or ( n6653 , n6651 , n6652 );
not ( n6654 , n6588 );
nand ( n6655 , n6654 , n3142 );
nand ( n6656 , n6653 , n6655 );
xor ( n6657 , n6649 , n6656 );
or ( n6658 , n6648 , n6657 );
not ( n6659 , n6656 );
or ( n6660 , n6649 , n6659 );
nand ( n6661 , n6658 , n6660 );
and ( n6662 , n6630 , n6661 );
and ( n6663 , n6626 , n6606 );
nor ( n6664 , n6662 , n6663 );
or ( n6665 , n6604 , n6599 );
or ( n6666 , n36 , n53 );
nand ( n6667 , n36 , n53 );
nand ( n6668 , n6666 , n6667 );
or ( n6669 , n3147 , n6668 );
nand ( n6670 , n6665 , n6669 );
not ( n6671 , n6587 );
xor ( n6672 , n6670 , n6671 );
not ( n6673 , n38 );
not ( n6674 , n52 );
and ( n6675 , n6673 , n6674 );
and ( n6676 , n38 , n52 );
nor ( n6677 , n6675 , n6676 );
and ( n6678 , n6677 , n6641 );
not ( n6679 , n3116 );
nor ( n6680 , n6678 , n6679 );
xnor ( n6681 , n6672 , n6680 );
not ( n6682 , n3318 );
not ( n6683 , n6618 );
not ( n6684 , n6683 );
or ( n6685 , n6682 , n6684 );
nand ( n6686 , n6685 , n40 );
and ( n6687 , n36 , n56 );
not ( n6688 , n6646 );
not ( n6689 , n6641 );
or ( n6690 , n6688 , n6689 );
not ( n6691 , n3114 );
nand ( n6692 , n6691 , n6677 );
nand ( n6693 , n6690 , n6692 );
xor ( n6694 , n6687 , n6693 );
and ( n6695 , n6686 , n6694 );
and ( n6696 , n6687 , n6693 );
nor ( n6697 , n6695 , n6696 );
xnor ( n6698 , n6681 , n6697 );
xnor ( n6699 , n6664 , n6698 );
not ( n6700 , n3350 );
not ( n6701 , n43 );
nand ( n6702 , n6701 , n44 );
not ( n6703 , n44 );
nand ( n6704 , n6703 , n43 );
and ( n6705 , n6702 , n6704 , n3353 );
buf ( n6706 , n6705 );
not ( n6707 , n6706 );
nand ( n6708 , n6700 , n6707 );
nand ( n6709 , n42 , n6708 );
not ( n6710 , n6709 );
and ( n6711 , n36 , n57 );
not ( n6712 , n36 );
not ( n6713 , n57 );
and ( n6714 , n6712 , n6713 );
nor ( n6715 , n6711 , n6714 );
not ( n6716 , n6715 );
not ( n6717 , n6598 );
or ( n6718 , n6716 , n6717 );
nand ( n6719 , n3583 , n6650 );
nand ( n6720 , n6718 , n6719 );
not ( n6721 , n6720 );
not ( n6722 , n6721 );
and ( n6723 , n6710 , n6722 );
and ( n6724 , n6709 , n6721 );
nor ( n6725 , n6723 , n6724 );
not ( n6726 , n6725 );
and ( n6727 , n40 , n53 );
nor ( n6728 , n40 , n53 );
nor ( n6729 , n6727 , n6728 );
and ( n6730 , n6618 , n6729 );
and ( n6731 , n3238 , n6623 );
nor ( n6732 , n6730 , n6731 );
not ( n6733 , n6732 );
and ( n6734 , n6726 , n6733 );
and ( n6735 , n6709 , n6720 );
nor ( n6736 , n6734 , n6735 );
not ( n6737 , n6648 );
and ( n6738 , n6657 , n6737 );
not ( n6739 , n6657 );
and ( n6740 , n6739 , n6648 );
nor ( n6741 , n6738 , n6740 );
and ( n6742 , n6741 , n6625 );
not ( n6743 , n6741 );
and ( n6744 , n6743 , n6626 );
nor ( n6745 , n6742 , n6744 );
or ( n6746 , n6736 , n6745 );
or ( n6747 , n6626 , n6741 );
nand ( n6748 , n6746 , n6747 );
xor ( n6749 , n6661 , n6630 );
xor ( n6750 , n6686 , n6694 );
xor ( n6751 , n6749 , n6750 );
and ( n6752 , n6748 , n6751 );
and ( n6753 , n6750 , n6749 );
nor ( n6754 , n6752 , n6753 );
nand ( n6755 , n6699 , n6754 );
xnor ( n6756 , n6748 , n6751 );
xor ( n6757 , n6732 , n6725 );
not ( n6758 , n6757 );
nand ( n6759 , n36 , n59 );
not ( n6760 , n6759 );
not ( n6761 , n6760 );
xnor ( n6762 , n36 , n58 );
not ( n6763 , n6762 );
not ( n6764 , n6763 );
not ( n6765 , n6598 );
or ( n6766 , n6764 , n6765 );
nand ( n6767 , n3583 , n6715 );
nand ( n6768 , n6766 , n6767 );
not ( n6769 , n6768 );
or ( n6770 , n6761 , n6769 );
and ( n6771 , n42 , n52 );
nor ( n6772 , n42 , n52 );
nor ( n6773 , n6771 , n6772 );
not ( n6774 , n6707 );
and ( n6775 , n6773 , n6774 );
and ( n6776 , n4601 , n42 );
nor ( n6777 , n6775 , n6776 );
not ( n6778 , n6777 );
not ( n6779 , n6759 );
not ( n6780 , n6768 );
or ( n6781 , n6779 , n6780 );
or ( n6782 , n6759 , n6768 );
nand ( n6783 , n6781 , n6782 );
nand ( n6784 , n6778 , n6783 );
nand ( n6785 , n6770 , n6784 );
xnor ( n6786 , n40 , n54 );
not ( n6787 , n6786 );
not ( n6788 , n6617 );
and ( n6789 , n6787 , n6788 );
not ( n6790 , n3237 );
and ( n6791 , n6790 , n6729 );
nor ( n6792 , n6789 , n6791 );
nand ( n6793 , n36 , n58 );
not ( n6794 , n6793 );
and ( n6795 , n38 , n55 );
not ( n6796 , n38 );
not ( n6797 , n55 );
and ( n6798 , n6796 , n6797 );
nor ( n6799 , n6795 , n6798 );
not ( n6800 , n6799 );
not ( n6801 , n6639 );
or ( n6802 , n6800 , n6801 );
nand ( n6803 , n5132 , n6635 );
nand ( n6804 , n6802 , n6803 );
not ( n6805 , n6804 );
or ( n6806 , n6794 , n6805 );
or ( n6807 , n6793 , n6804 );
nand ( n6808 , n6806 , n6807 );
xor ( n6809 , n6792 , n6808 );
xor ( n6810 , n6785 , n6809 );
or ( n6811 , n6758 , n6810 );
not ( n6812 , n6785 );
or ( n6813 , n6812 , n6809 );
nand ( n6814 , n6811 , n6813 );
and ( n6815 , n6745 , n6736 );
not ( n6816 , n6745 );
not ( n6817 , n6736 );
and ( n6818 , n6816 , n6817 );
nor ( n6819 , n6815 , n6818 );
not ( n6820 , n6792 );
not ( n6821 , n6820 );
not ( n6822 , n6808 );
or ( n6823 , n6821 , n6822 );
not ( n6824 , n6804 );
or ( n6825 , n6793 , n6824 );
nand ( n6826 , n6823 , n6825 );
xor ( n6827 , n6819 , n6826 );
and ( n6828 , n6814 , n6827 );
and ( n6829 , n6826 , n6819 );
nor ( n6830 , n6828 , n6829 );
nand ( n6831 , n6756 , n6830 );
not ( n6832 , n6831 );
not ( n6833 , n6814 );
and ( n6834 , n6827 , n6833 );
not ( n6835 , n6827 );
and ( n6836 , n6835 , n6814 );
nor ( n6837 , n6834 , n6836 );
xnor ( n6838 , n36 , n59 );
not ( n6839 , n6597 );
not ( n6840 , n6839 );
or ( n6841 , n6838 , n6840 );
or ( n6842 , n3143 , n6762 );
nand ( n6843 , n6841 , n6842 );
not ( n6844 , n6843 );
nand ( n6845 , n36 , n60 );
not ( n6846 , n6845 );
and ( n6847 , n40 , n55 );
not ( n6848 , n40 );
and ( n6849 , n6848 , n6797 );
nor ( n6850 , n6847 , n6849 );
not ( n6851 , n6850 );
not ( n6852 , n6616 );
or ( n6853 , n6851 , n6852 );
not ( n6854 , n6786 );
nand ( n6855 , n6854 , n3235 );
nand ( n6856 , n6853 , n6855 );
not ( n6857 , n6856 );
or ( n6858 , n6846 , n6857 );
or ( n6859 , n6845 , n6856 );
nand ( n6860 , n6858 , n6859 );
not ( n6861 , n6860 );
or ( n6862 , n6844 , n6861 );
not ( n6863 , n6845 );
nand ( n6864 , n6863 , n6856 );
nand ( n6865 , n6862 , n6864 );
not ( n6866 , n6865 );
not ( n6867 , n4415 );
not ( n6868 , n6799 );
not ( n6869 , n6868 );
and ( n6870 , n6867 , n6869 );
not ( n6871 , n38 );
not ( n6872 , n56 );
and ( n6873 , n6871 , n6872 );
and ( n6874 , n38 , n56 );
nor ( n6875 , n6873 , n6874 );
not ( n6876 , n6640 );
and ( n6877 , n6875 , n6876 );
nor ( n6878 , n6870 , n6877 );
and ( n6879 , n6878 , n6792 );
not ( n6880 , n6878 );
and ( n6881 , n6880 , n6820 );
nor ( n6882 , n6879 , n6881 );
or ( n6883 , n6866 , n6882 );
or ( n6884 , n6820 , n6878 );
nand ( n6885 , n6883 , n6884 );
buf ( n6886 , n6885 );
not ( n6887 , n6886 );
and ( n6888 , n6810 , n6757 );
not ( n6889 , n6810 );
and ( n6890 , n6889 , n6758 );
nor ( n6891 , n6888 , n6890 );
not ( n6892 , n6891 );
not ( n6893 , n6892 );
or ( n6894 , n6887 , n6893 );
nand ( n6895 , n6885 , n6891 );
not ( n6896 , n6895 );
not ( n6897 , n6892 );
nor ( n6898 , n6897 , n6886 );
nor ( n6899 , n6896 , n6898 );
and ( n6900 , n42 , n6643 );
not ( n6901 , n42 );
and ( n6902 , n6901 , n53 );
nor ( n6903 , n6900 , n6902 );
not ( n6904 , n6903 );
not ( n6905 , n6774 );
not ( n6906 , n6905 );
and ( n6907 , n6904 , n6906 );
and ( n6908 , n4601 , n6773 );
nor ( n6909 , n6907 , n6908 );
not ( n6910 , n6909 );
not ( n6911 , n6910 );
not ( n6912 , n3468 );
xor ( n6913 , n45 , n46 );
nand ( n6914 , n3451 , n6913 );
not ( n6915 , n6914 );
not ( n6916 , n6915 );
not ( n6917 , n6916 );
not ( n6918 , n6917 );
not ( n6919 , n6918 );
not ( n6920 , n6919 );
not ( n6921 , n6920 );
or ( n6922 , n6912 , n6921 );
nand ( n6923 , n6922 , n44 );
xor ( n6924 , n38 , n57 );
not ( n6925 , n6924 );
not ( n6926 , n6639 );
or ( n6927 , n6925 , n6926 );
nand ( n6928 , n4321 , n6875 );
nand ( n6929 , n6927 , n6928 );
xor ( n6930 , n6923 , n6929 );
not ( n6931 , n6930 );
or ( n6932 , n6911 , n6931 );
nand ( n6933 , n6923 , n6929 );
nand ( n6934 , n6932 , n6933 );
not ( n6935 , n6934 );
not ( n6936 , n6777 );
not ( n6937 , n6783 );
or ( n6938 , n6936 , n6937 );
not ( n6939 , n6777 );
not ( n6940 , n6783 );
nand ( n6941 , n6939 , n6940 );
nand ( n6942 , n6938 , n6941 );
and ( n6943 , n6935 , n6942 );
not ( n6944 , n6935 );
not ( n6945 , n6942 );
and ( n6946 , n6944 , n6945 );
nor ( n6947 , n6943 , n6946 );
not ( n6948 , n6947 );
not ( n6949 , n6882 );
not ( n6950 , n6949 );
not ( n6951 , n6866 );
or ( n6952 , n6950 , n6951 );
nand ( n6953 , n6865 , n6882 );
nand ( n6954 , n6952 , n6953 );
and ( n6955 , n6948 , n6954 );
and ( n6956 , n6942 , n6934 );
nor ( n6957 , n6955 , n6956 );
buf ( n6958 , n6957 );
or ( n6959 , n6899 , n6958 );
nand ( n6960 , n6894 , n6959 );
not ( n6961 , n6960 );
nand ( n6962 , n6837 , n6961 );
not ( n6963 , n6962 );
not ( n6964 , n6954 );
not ( n6965 , n6947 );
and ( n6966 , n6964 , n6965 );
and ( n6967 , n6954 , n6947 );
nor ( n6968 , n6966 , n6967 );
xor ( n6969 , n6843 , n6860 );
not ( n6970 , n6969 );
not ( n6971 , n6970 );
not ( n6972 , n44 );
not ( n6973 , n4732 );
or ( n6974 , n6972 , n6973 );
and ( n6975 , n44 , n52 );
not ( n6976 , n44 );
and ( n6977 , n6976 , n6621 );
nor ( n6978 , n6975 , n6977 );
nand ( n6979 , n6978 , n6919 );
nand ( n6980 , n6974 , n6979 );
not ( n6981 , n6980 );
xor ( n6982 , n36 , n60 );
not ( n6983 , n6982 );
not ( n6984 , n6839 );
or ( n6985 , n6983 , n6984 );
not ( n6986 , n6838 );
nand ( n6987 , n6986 , n3142 );
nand ( n6988 , n6985 , n6987 );
not ( n6989 , n6988 );
or ( n6990 , n6981 , n6989 );
or ( n6991 , n6980 , n6988 );
xor ( n6992 , n38 , n58 );
not ( n6993 , n6992 );
not ( n6994 , n6639 );
or ( n6995 , n6993 , n6994 );
nand ( n6996 , n3422 , n6924 );
nand ( n6997 , n6995 , n6996 );
nand ( n6998 , n6991 , n6997 );
nand ( n6999 , n6990 , n6998 );
not ( n7000 , n6999 );
xnor ( n7001 , n42 , n54 );
not ( n7002 , n7001 );
not ( n7003 , n7002 );
not ( n7004 , n6774 );
or ( n7005 , n7003 , n7004 );
not ( n7006 , n6903 );
nand ( n7007 , n7006 , n3350 );
nand ( n7008 , n7005 , n7007 );
and ( n7009 , n7000 , n7008 );
not ( n7010 , n7000 );
not ( n7011 , n7008 );
and ( n7012 , n7010 , n7011 );
nor ( n7013 , n7009 , n7012 );
not ( n7014 , n7013 );
and ( n7015 , n6971 , n7014 );
and ( n7016 , n7008 , n6999 );
nor ( n7017 , n7015 , n7016 );
not ( n7018 , n7017 );
and ( n7019 , n6968 , n7018 );
not ( n7020 , n6968 );
and ( n7021 , n7020 , n7017 );
nor ( n7022 , n7019 , n7021 );
and ( n7023 , n36 , n61 );
xor ( n7024 , n40 , n56 );
not ( n7025 , n7024 );
not ( n7026 , n6616 );
or ( n7027 , n7025 , n7026 );
not ( n7028 , n3236 );
not ( n7029 , n6850 );
or ( n7030 , n7028 , n7029 );
nand ( n7031 , n7027 , n7030 );
xor ( n7032 , n7023 , n7031 );
and ( n7033 , n7011 , n7032 );
and ( n7034 , n7023 , n7031 );
nor ( n7035 , n7033 , n7034 );
not ( n7036 , n7035 );
not ( n7037 , n6909 );
not ( n7038 , n6930 );
or ( n7039 , n7037 , n7038 );
or ( n7040 , n6909 , n6930 );
nand ( n7041 , n7039 , n7040 );
not ( n7042 , n7041 );
not ( n7043 , n7042 );
and ( n7044 , n7036 , n7043 );
not ( n7045 , n7035 );
not ( n7046 , n7045 );
not ( n7047 , n7042 );
or ( n7048 , n7046 , n7047 );
nand ( n7049 , n7035 , n7041 );
nand ( n7050 , n7048 , n7049 );
not ( n7051 , n7013 );
nand ( n7052 , n6970 , n7051 );
nand ( n7053 , n6969 , n7013 );
nand ( n7054 , n7052 , n7053 );
and ( n7055 , n7050 , n7054 );
nor ( n7056 , n7044 , n7055 );
xor ( n7057 , n7022 , n7056 );
and ( n7058 , n7032 , n7008 );
not ( n7059 , n7032 );
and ( n7060 , n7059 , n7011 );
nor ( n7061 , n7058 , n7060 );
not ( n7062 , n7061 );
and ( n7063 , n36 , n62 );
not ( n7064 , n7063 );
and ( n7065 , n46 , n52 );
not ( n7066 , n46 );
and ( n7067 , n7066 , n6621 );
nor ( n7068 , n7065 , n7067 );
not ( n7069 , n7068 );
nor ( n7070 , n46 , n47 );
not ( n7071 , n7070 );
nand ( n7072 , n46 , n47 );
nand ( n7073 , n7071 , n3608 , n7072 );
not ( n7074 , n7073 );
buf ( n7075 , n7074 );
not ( n7076 , n7075 );
not ( n7077 , n7076 );
not ( n7078 , n7077 );
or ( n7079 , n7069 , n7078 );
buf ( n7080 , n3609 );
buf ( n7081 , n7080 );
nand ( n7082 , n46 , n7081 );
nand ( n7083 , n7079 , n7082 );
not ( n7084 , n7083 );
or ( n7085 , n7064 , n7084 );
not ( n7086 , n7063 );
not ( n7087 , n7083 );
nand ( n7088 , n7086 , n7087 );
xor ( n7089 , n40 , n58 );
not ( n7090 , n7089 );
not ( n7091 , n6616 );
or ( n7092 , n7090 , n7091 );
and ( n7093 , n40 , n57 );
not ( n7094 , n40 );
and ( n7095 , n7094 , n6713 );
nor ( n7096 , n7093 , n7095 );
nand ( n7097 , n3235 , n7096 );
nand ( n7098 , n7092 , n7097 );
not ( n7099 , n7098 );
xor ( n7100 , n44 , n53 );
not ( n7101 , n7100 );
not ( n7102 , n4248 );
or ( n7103 , n7101 , n7102 );
xor ( n7104 , n44 , n54 );
not ( n7105 , n6916 );
nand ( n7106 , n7104 , n7105 );
nand ( n7107 , n7103 , n7106 );
xor ( n7108 , n38 , n60 );
not ( n7109 , n7108 );
not ( n7110 , n6638 );
or ( n7111 , n7109 , n7110 );
xor ( n7112 , n38 , n59 );
nand ( n7113 , n3112 , n7112 );
nand ( n7114 , n7111 , n7113 );
xor ( n7115 , n7107 , n7114 );
not ( n7116 , n7115 );
or ( n7117 , n7099 , n7116 );
nand ( n7118 , n7107 , n7114 );
nand ( n7119 , n7117 , n7118 );
nand ( n7120 , n7088 , n7119 );
nand ( n7121 , n7085 , n7120 );
not ( n7122 , n7121 );
or ( n7123 , n7062 , n7122 );
buf ( n7124 , n7061 );
or ( n7125 , n7124 , n7121 );
nand ( n7126 , n7123 , n7125 );
not ( n7127 , n7126 );
not ( n7128 , n7112 );
not ( n7129 , n6639 );
or ( n7130 , n7128 , n7129 );
nand ( n7131 , n3422 , n6992 );
nand ( n7132 , n7130 , n7131 );
xor ( n7133 , n36 , n61 );
not ( n7134 , n7133 );
not ( n7135 , n6598 );
or ( n7136 , n7134 , n7135 );
nand ( n7137 , n3583 , n6982 );
nand ( n7138 , n7136 , n7137 );
and ( n7139 , n7132 , n7138 );
not ( n7140 , n7132 );
not ( n7141 , n7138 );
and ( n7142 , n7140 , n7141 );
nor ( n7143 , n7139 , n7142 );
and ( n7144 , n42 , n55 );
not ( n7145 , n42 );
and ( n7146 , n7145 , n6797 );
nor ( n7147 , n7144 , n7146 );
not ( n7148 , n7147 );
not ( n7149 , n6774 );
or ( n7150 , n7148 , n7149 );
not ( n7151 , n3350 );
or ( n7152 , n7151 , n7001 );
nand ( n7153 , n7150 , n7152 );
xor ( n7154 , n7143 , n7153 );
not ( n7155 , n7154 );
xor ( n7156 , n42 , n56 );
not ( n7157 , n7156 );
not ( n7158 , n6774 );
or ( n7159 , n7157 , n7158 );
nand ( n7160 , n3350 , n7147 );
nand ( n7161 , n7159 , n7160 );
not ( n7162 , n7161 );
not ( n7163 , n7162 );
xor ( n7164 , n36 , n62 );
not ( n7165 , n7164 );
not ( n7166 , n6839 );
or ( n7167 , n7165 , n7166 );
nand ( n7168 , n3521 , n7133 );
nand ( n7169 , n7167 , n7168 );
not ( n7170 , n7169 );
nand ( n7171 , n36 , n63 );
not ( n7172 , n7171 );
and ( n7173 , n7170 , n7172 );
and ( n7174 , n7171 , n7169 );
nor ( n7175 , n7173 , n7174 );
not ( n7176 , n7175 );
and ( n7177 , n7163 , n7176 );
not ( n7178 , n7169 );
nor ( n7179 , n7178 , n7171 );
nor ( n7180 , n7177 , n7179 );
not ( n7181 , n6978 );
not ( n7182 , n3467 );
or ( n7183 , n7181 , n7182 );
nand ( n7184 , n6919 , n7100 );
nand ( n7185 , n7183 , n7184 );
not ( n7186 , n7185 );
not ( n7187 , n7080 );
not ( n7188 , n7187 );
not ( n7189 , n7075 );
nand ( n7190 , n7188 , n7189 );
nand ( n7191 , n46 , n7190 );
not ( n7192 , n7191 );
not ( n7193 , n7192 );
and ( n7194 , n7186 , n7193 );
and ( n7195 , n7192 , n7185 );
nor ( n7196 , n7194 , n7195 );
not ( n7197 , n7096 );
not ( n7198 , n6616 );
or ( n7199 , n7197 , n7198 );
nand ( n7200 , n3236 , n7024 );
nand ( n7201 , n7199 , n7200 );
and ( n7202 , n7196 , n7201 );
not ( n7203 , n7196 );
not ( n7204 , n7201 );
and ( n7205 , n7203 , n7204 );
nor ( n7206 , n7202 , n7205 );
not ( n7207 , n7206 );
and ( n7208 , n7180 , n7207 );
not ( n7209 , n7180 );
and ( n7210 , n7209 , n7206 );
nor ( n7211 , n7208 , n7210 );
not ( n7212 , n7211 );
not ( n7213 , n7212 );
or ( n7214 , n7155 , n7213 );
not ( n7215 , n7180 );
nand ( n7216 , n7215 , n7207 );
nand ( n7217 , n7214 , n7216 );
not ( n7218 , n7217 );
or ( n7219 , n7127 , n7218 );
not ( n7220 , n7121 );
or ( n7221 , n7124 , n7220 );
nand ( n7222 , n7219 , n7221 );
not ( n7223 , n7222 );
not ( n7224 , n7054 );
and ( n7225 , n7050 , n7224 );
not ( n7226 , n7050 );
and ( n7227 , n7226 , n7054 );
nor ( n7228 , n7225 , n7227 );
not ( n7229 , n7228 );
not ( n7230 , n7201 );
not ( n7231 , n7196 );
not ( n7232 , n7231 );
or ( n7233 , n7230 , n7232 );
nand ( n7234 , n7191 , n7185 );
nand ( n7235 , n7233 , n7234 );
not ( n7236 , n7235 );
not ( n7237 , n7236 );
xor ( n7238 , n6980 , n6997 );
not ( n7239 , n6988 );
and ( n7240 , n7238 , n7239 );
not ( n7241 , n7238 );
and ( n7242 , n7241 , n6988 );
nor ( n7243 , n7240 , n7242 );
not ( n7244 , n7243 );
not ( n7245 , n7244 );
or ( n7246 , n7237 , n7245 );
nand ( n7247 , n7235 , n7243 );
nand ( n7248 , n7246 , n7247 );
not ( n7249 , n7248 );
nand ( n7250 , n7138 , n7132 );
nand ( n7251 , n7153 , n7143 );
and ( n7252 , n7250 , n7251 );
or ( n7253 , n7249 , n7252 );
nand ( n7254 , n7235 , n7244 );
nand ( n7255 , n7253 , n7254 );
not ( n7256 , n7255 );
and ( n7257 , n7229 , n7256 );
and ( n7258 , n7255 , n7228 );
nor ( n7259 , n7257 , n7258 );
not ( n7260 , n7259 );
not ( n7261 , n7260 );
or ( n7262 , n7223 , n7261 );
not ( n7263 , n7228 );
nand ( n7264 , n7263 , n7255 );
nand ( n7265 , n7262 , n7264 );
nand ( n7266 , n7057 , n7265 );
not ( n7267 , n6957 );
not ( n7268 , n7267 );
not ( n7269 , n6899 );
or ( n7270 , n7268 , n7269 );
not ( n7271 , n6958 );
or ( n7272 , n7271 , n6899 );
nand ( n7273 , n7270 , n7272 );
or ( n7274 , n7056 , n7022 );
or ( n7275 , n7017 , n6968 );
nand ( n7276 , n7274 , n7275 );
nor ( n7277 , n7273 , n7276 );
or ( n7278 , n7266 , n7277 );
nand ( n7279 , n7273 , n7276 );
nand ( n7280 , n7278 , n7279 );
not ( n7281 , n7280 );
or ( n7282 , n6963 , n7281 );
not ( n7283 , n6837 );
nand ( n7284 , n7283 , n6960 );
nand ( n7285 , n7282 , n7284 );
not ( n7286 , n7285 );
or ( n7287 , n6832 , n7286 );
not ( n7288 , n6756 );
not ( n7289 , n6830 );
nand ( n7290 , n7288 , n7289 );
buf ( n7291 , n7290 );
nand ( n7292 , n7287 , n7291 );
nand ( n7293 , n6755 , n7292 );
or ( n7294 , n6699 , n6754 );
not ( n7295 , n7126 );
not ( n7296 , n7217 );
not ( n7297 , n7296 );
or ( n7298 , n7295 , n7297 );
not ( n7299 , n7126 );
nand ( n7300 , n7299 , n7217 );
nand ( n7301 , n7298 , n7300 );
not ( n7302 , n7161 );
not ( n7303 , n7175 );
or ( n7304 , n7302 , n7303 );
or ( n7305 , n7175 , n7161 );
nand ( n7306 , n7304 , n7305 );
not ( n7307 , n7306 );
xor ( n7308 , n48 , n52 );
not ( n7309 , n7308 );
xor ( n7310 , n49 , n50 );
not ( n7311 , n7310 );
and ( n7312 , n3561 , n7311 );
not ( n7313 , n7312 );
not ( n7314 , n7313 );
not ( n7315 , n7314 );
or ( n7316 , n7309 , n7315 );
buf ( n7317 , n7310 );
buf ( n7318 , n7317 );
buf ( n7319 , n7318 );
nand ( n7320 , n48 , n7319 );
nand ( n7321 , n7316 , n7320 );
buf ( n7322 , n7321 );
not ( n7323 , n7322 );
xor ( n7324 , n36 , n63 );
not ( n7325 , n7324 );
not ( n7326 , n6839 );
or ( n7327 , n7325 , n7326 );
nand ( n7328 , n3142 , n7164 );
nand ( n7329 , n7327 , n7328 );
not ( n7330 , n7329 );
or ( n7331 , n7323 , n7330 );
not ( n7332 , n7321 );
not ( n7333 , n7332 );
not ( n7334 , n7329 );
not ( n7335 , n7334 );
or ( n7336 , n7333 , n7335 );
xor ( n7337 , n38 , n61 );
not ( n7338 , n7337 );
not ( n7339 , n6639 );
or ( n7340 , n7338 , n7339 );
nand ( n7341 , n3112 , n7108 );
nand ( n7342 , n7340 , n7341 );
nand ( n7343 , n7336 , n7342 );
nand ( n7344 , n7331 , n7343 );
not ( n7345 , n7344 );
not ( n7346 , n7098 );
not ( n7347 , n7346 );
not ( n7348 , n7115 );
and ( n7349 , n7347 , n7348 );
and ( n7350 , n7346 , n7115 );
nor ( n7351 , n7349 , n7350 );
not ( n7352 , n7351 );
or ( n7353 , n7345 , n7352 );
or ( n7354 , n7344 , n7351 );
nand ( n7355 , n7353 , n7354 );
not ( n7356 , n7355 );
or ( n7357 , n7307 , n7356 );
not ( n7358 , n7351 );
nand ( n7359 , n7344 , n7358 );
nand ( n7360 , n7357 , n7359 );
not ( n7361 , n7360 );
xor ( n7362 , n46 , n53 );
not ( n7363 , n7362 );
not ( n7364 , n7077 );
or ( n7365 , n7363 , n7364 );
nand ( n7366 , n7068 , n7081 );
nand ( n7367 , n7365 , n7366 );
not ( n7368 , n7367 );
not ( n7369 , n7318 );
not ( n7370 , n7369 );
not ( n7371 , n7313 );
or ( n7372 , n7370 , n7371 );
nand ( n7373 , n7372 , n48 );
not ( n7374 , n7373 );
xor ( n7375 , n42 , n57 );
not ( n7376 , n7375 );
not ( n7377 , n6705 );
or ( n7378 , n7376 , n7377 );
nand ( n7379 , n3348 , n7156 );
nand ( n7380 , n7378 , n7379 );
not ( n7381 , n7380 );
not ( n7382 , n7381 );
or ( n7383 , n7374 , n7382 );
not ( n7384 , n7380 );
or ( n7385 , n7373 , n7384 );
nand ( n7386 , n7383 , n7385 );
not ( n7387 , n7386 );
or ( n7388 , n7368 , n7387 );
not ( n7389 , n7384 );
nand ( n7390 , n7373 , n7389 );
nand ( n7391 , n7388 , n7390 );
not ( n7392 , n7391 );
not ( n7393 , n7087 );
xor ( n7394 , n40 , n59 );
not ( n7395 , n7394 );
not ( n7396 , n6615 );
or ( n7397 , n7395 , n7396 );
nand ( n7398 , n3736 , n7089 );
nand ( n7399 , n7397 , n7398 );
not ( n7400 , n7399 );
and ( n7401 , n36 , n64 );
not ( n7402 , n7104 );
not ( n7403 , n4247 );
or ( n7404 , n7402 , n7403 );
not ( n7405 , n6914 );
and ( n7406 , n44 , n55 );
not ( n7407 , n44 );
and ( n7408 , n7407 , n6797 );
nor ( n7409 , n7406 , n7408 );
nand ( n7410 , n7405 , n7409 );
nand ( n7411 , n7404 , n7410 );
and ( n7412 , n7401 , n7411 );
not ( n7413 , n7401 );
not ( n7414 , n7411 );
and ( n7415 , n7413 , n7414 );
nor ( n7416 , n7412 , n7415 );
not ( n7417 , n7416 );
or ( n7418 , n7400 , n7417 );
not ( n7419 , n7414 );
nand ( n7420 , n7401 , n7419 );
nand ( n7421 , n7418 , n7420 );
not ( n7422 , n7421 );
not ( n7423 , n7422 );
or ( n7424 , n7393 , n7423 );
not ( n7425 , n7421 );
or ( n7426 , n7087 , n7425 );
nand ( n7427 , n7424 , n7426 );
not ( n7428 , n7427 );
or ( n7429 , n7392 , n7428 );
not ( n7430 , n7425 );
nand ( n7431 , n7087 , n7430 );
nand ( n7432 , n7429 , n7431 );
not ( n7433 , n7119 );
not ( n7434 , n7063 );
not ( n7435 , n7087 );
and ( n7436 , n7434 , n7435 );
and ( n7437 , n7063 , n7087 );
nor ( n7438 , n7436 , n7437 );
not ( n7439 , n7438 );
and ( n7440 , n7433 , n7439 );
not ( n7441 , n7433 );
and ( n7442 , n7441 , n7438 );
nor ( n7443 , n7440 , n7442 );
and ( n7444 , n7432 , n7443 );
not ( n7445 , n7432 );
not ( n7446 , n7443 );
and ( n7447 , n7445 , n7446 );
nor ( n7448 , n7444 , n7447 );
not ( n7449 , n7448 );
not ( n7450 , n7449 );
or ( n7451 , n7361 , n7450 );
nand ( n7452 , n7446 , n7432 );
nand ( n7453 , n7451 , n7452 );
not ( n7454 , n7252 );
not ( n7455 , n7248 );
or ( n7456 , n7454 , n7455 );
or ( n7457 , n7252 , n7248 );
nand ( n7458 , n7456 , n7457 );
xor ( n7459 , n7453 , n7458 );
not ( n7460 , n7459 );
and ( n7461 , n7301 , n7460 );
not ( n7462 , n7301 );
and ( n7463 , n7462 , n7459 );
nor ( n7464 , n7461 , n7463 );
and ( n7465 , n7355 , n7306 );
not ( n7466 , n7355 );
not ( n7467 , n7306 );
and ( n7468 , n7466 , n7467 );
nor ( n7469 , n7465 , n7468 );
not ( n7470 , n7469 );
not ( n7471 , n7391 );
and ( n7472 , n7427 , n7471 );
not ( n7473 , n7427 );
and ( n7474 , n7473 , n7391 );
nor ( n7475 , n7472 , n7474 );
not ( n7476 , n7475 );
not ( n7477 , n7367 );
not ( n7478 , n7477 );
not ( n7479 , n7386 );
and ( n7480 , n7478 , n7479 );
and ( n7481 , n7477 , n7386 );
nor ( n7482 , n7480 , n7481 );
not ( n7483 , n7482 );
not ( n7484 , n7483 );
xor ( n7485 , n46 , n54 );
not ( n7486 , n7485 );
not ( n7487 , n7075 );
or ( n7488 , n7486 , n7487 );
nand ( n7489 , n7362 , n7080 );
nand ( n7490 , n7488 , n7489 );
not ( n7491 , n7490 );
xor ( n7492 , n42 , n58 );
not ( n7493 , n7492 );
and ( n7494 , n6702 , n6704 , n3353 );
not ( n7495 , n7494 );
or ( n7496 , n7493 , n7495 );
nand ( n7497 , n3355 , n7375 );
nand ( n7498 , n7496 , n7497 );
not ( n7499 , n7498 );
nand ( n7500 , n36 , n65 );
not ( n7501 , n7500 );
and ( n7502 , n7499 , n7501 );
and ( n7503 , n7500 , n7498 );
nor ( n7504 , n7502 , n7503 );
or ( n7505 , n7491 , n7504 );
not ( n7506 , n7500 );
nand ( n7507 , n7506 , n7498 );
nand ( n7508 , n7505 , n7507 );
not ( n7509 , n7508 );
xor ( n7510 , n40 , n60 );
not ( n7511 , n7510 );
not ( n7512 , n6614 );
or ( n7513 , n7511 , n7512 );
nand ( n7514 , n3233 , n7394 );
nand ( n7515 , n7513 , n7514 );
not ( n7516 , n7515 );
not ( n7517 , n7409 );
not ( n7518 , n3464 );
or ( n7519 , n7517 , n7518 );
xor ( n7520 , n44 , n56 );
nand ( n7521 , n7520 , n7405 );
nand ( n7522 , n7519 , n7521 );
not ( n7523 , n7522 );
or ( n7524 , n7516 , n7523 );
not ( n7525 , n7515 );
not ( n7526 , n7525 );
not ( n7527 , n7522 );
not ( n7528 , n7527 );
or ( n7529 , n7526 , n7528 );
xor ( n7530 , n38 , n62 );
not ( n7531 , n7530 );
not ( n7532 , n6638 );
or ( n7533 , n7531 , n7532 );
nand ( n7534 , n3972 , n7337 );
nand ( n7535 , n7533 , n7534 );
nand ( n7536 , n7529 , n7535 );
nand ( n7537 , n7524 , n7536 );
not ( n7538 , n7537 );
not ( n7539 , n7538 );
or ( n7540 , n7509 , n7539 );
or ( n7541 , n7508 , n7538 );
nand ( n7542 , n7540 , n7541 );
not ( n7543 , n7542 );
or ( n7544 , n7484 , n7543 );
nand ( n7545 , n7508 , n7537 );
nand ( n7546 , n7544 , n7545 );
not ( n7547 , n7546 );
or ( n7548 , n7476 , n7547 );
or ( n7549 , n7475 , n7546 );
nand ( n7550 , n7548 , n7549 );
not ( n7551 , n7550 );
or ( n7552 , n7470 , n7551 );
not ( n7553 , n7475 );
nand ( n7554 , n7553 , n7546 );
nand ( n7555 , n7552 , n7554 );
not ( n7556 , n7555 );
not ( n7557 , n7154 );
not ( n7558 , n7557 );
not ( n7559 , n7212 );
or ( n7560 , n7558 , n7559 );
nand ( n7561 , n7154 , n7211 );
nand ( n7562 , n7560 , n7561 );
not ( n7563 , n7360 );
not ( n7564 , n7563 );
not ( n7565 , n7449 );
or ( n7566 , n7564 , n7565 );
nand ( n7567 , n7360 , n7448 );
nand ( n7568 , n7566 , n7567 );
and ( n7569 , n7562 , n7568 );
not ( n7570 , n7562 );
not ( n7571 , n7568 );
and ( n7572 , n7570 , n7571 );
nor ( n7573 , n7569 , n7572 );
not ( n7574 , n7573 );
or ( n7575 , n7556 , n7574 );
not ( n7576 , n7571 );
nand ( n7577 , n7562 , n7576 );
nand ( n7578 , n7575 , n7577 );
not ( n7579 , n7578 );
nand ( n7580 , n7464 , n7579 );
not ( n7581 , n7580 );
not ( n7582 , n7581 );
xor ( n7583 , n42 , n61 );
not ( n7584 , n7583 );
not ( n7585 , n6706 );
or ( n7586 , n7584 , n7585 );
xor ( n7587 , n42 , n60 );
nand ( n7588 , n3350 , n7587 );
nand ( n7589 , n7586 , n7588 );
not ( n7590 , n7589 );
xor ( n7591 , n40 , n63 );
not ( n7592 , n7591 );
not ( n7593 , n6615 );
or ( n7594 , n7592 , n7593 );
xor ( n7595 , n40 , n62 );
nand ( n7596 , n3234 , n7595 );
nand ( n7597 , n7594 , n7596 );
xor ( n7598 , n46 , n57 );
not ( n7599 , n7598 );
not ( n7600 , n7075 );
or ( n7601 , n7599 , n7600 );
xor ( n7602 , n46 , n56 );
nand ( n7603 , n7602 , n7080 );
nand ( n7604 , n7601 , n7603 );
and ( n7605 , n7597 , n7604 );
not ( n7606 , n7597 );
not ( n7607 , n7604 );
and ( n7608 , n7606 , n7607 );
nor ( n7609 , n7605 , n7608 );
not ( n7610 , n7609 );
or ( n7611 , n7590 , n7610 );
not ( n7612 , n7607 );
nand ( n7613 , n7597 , n7612 );
nand ( n7614 , n7611 , n7613 );
not ( n7615 , n7614 );
not ( n7616 , n4224 );
not ( n7617 , n67 );
nand ( n7618 , n7617 , n4230 );
not ( n7619 , n7618 );
or ( n7620 , n7616 , n7619 );
nand ( n7621 , n7620 , n36 );
not ( n7622 , n7621 );
not ( n7623 , n5655 );
xor ( n7624 , n50 , n53 );
not ( n7625 , n7624 );
or ( n7626 , n7623 , n7625 );
xor ( n7627 , n50 , n52 );
nand ( n7628 , n51 , n7627 );
nand ( n7629 , n7626 , n7628 );
nand ( n7630 , n7622 , n7629 );
not ( n7631 , n7630 );
not ( n7632 , n3121 );
xor ( n7633 , n36 , n66 );
not ( n7634 , n7633 );
or ( n7635 , n7632 , n7634 );
nor ( n7636 , n36 , n67 );
not ( n7637 , n7636 );
nand ( n7638 , n36 , n67 );
nand ( n7639 , n7637 , n7638 , n6594 );
nand ( n7640 , n7635 , n7639 );
not ( n7641 , n7640 );
not ( n7642 , n7641 );
not ( n7643 , n7642 );
xor ( n7644 , n48 , n55 );
not ( n7645 , n7644 );
not ( n7646 , n7312 );
or ( n7647 , n7645 , n7646 );
xor ( n7648 , n48 , n54 );
nand ( n7649 , n7318 , n7648 );
nand ( n7650 , n7647 , n7649 );
not ( n7651 , n7650 );
not ( n7652 , n7651 );
not ( n7653 , n7652 );
or ( n7654 , n7643 , n7653 );
not ( n7655 , n7641 );
not ( n7656 , n7651 );
or ( n7657 , n7655 , n7656 );
xor ( n7658 , n44 , n58 );
not ( n7659 , n7658 );
not ( n7660 , n4248 );
or ( n7661 , n7659 , n7660 );
xor ( n7662 , n44 , n59 );
nand ( n7663 , n6917 , n7662 );
nand ( n7664 , n7661 , n7663 );
nand ( n7665 , n7657 , n7664 );
nand ( n7666 , n7654 , n7665 );
not ( n7667 , n7666 );
or ( n7668 , n7631 , n7667 );
or ( n7669 , n7630 , n7666 );
nand ( n7670 , n7668 , n7669 );
not ( n7671 , n7670 );
or ( n7672 , n7615 , n7671 );
not ( n7673 , n7630 );
nand ( n7674 , n7673 , n7666 );
nand ( n7675 , n7672 , n7674 );
not ( n7676 , n7675 );
xor ( n7677 , n36 , n65 );
not ( n7678 , n7677 );
not ( n7679 , n6596 );
or ( n7680 , n7678 , n7679 );
xor ( n7681 , n36 , n64 );
nand ( n7682 , n3141 , n7681 );
nand ( n7683 , n7680 , n7682 );
nand ( n7684 , n36 , n66 );
xor ( n7685 , n7684 , n50 );
xnor ( n7686 , n7683 , n7685 );
not ( n7687 , n7686 );
xor ( n7688 , n42 , n59 );
not ( n7689 , n7688 );
not ( n7690 , n6705 );
or ( n7691 , n7689 , n7690 );
nand ( n7692 , n3348 , n7492 );
nand ( n7693 , n7691 , n7692 );
xor ( n7694 , n46 , n55 );
not ( n7695 , n7694 );
not ( n7696 , n7075 );
or ( n7697 , n7695 , n7696 );
nand ( n7698 , n7485 , n7080 );
nand ( n7699 , n7697 , n7698 );
xor ( n7700 , n7693 , n7699 );
xor ( n7701 , n48 , n53 );
not ( n7702 , n7701 );
not ( n7703 , n7312 );
or ( n7704 , n7702 , n7703 );
nand ( n7705 , n7318 , n7308 );
nand ( n7706 , n7704 , n7705 );
not ( n7707 , n7706 );
not ( n7708 , n7707 );
xnor ( n7709 , n7700 , n7708 );
not ( n7710 , n7709 );
not ( n7711 , n7710 );
or ( n7712 , n7687 , n7711 );
not ( n7713 , n7686 );
nand ( n7714 , n7713 , n7709 );
nand ( n7715 , n7712 , n7714 );
not ( n7716 , n7715 );
or ( n7717 , n7676 , n7716 );
not ( n7718 , n7686 );
nand ( n7719 , n7718 , n7710 );
nand ( n7720 , n7717 , n7719 );
xor ( n7721 , n7515 , n7527 );
xnor ( n7722 , n7721 , n7535 );
not ( n7723 , n7685 );
not ( n7724 , n7683 );
or ( n7725 , n7723 , n7724 );
or ( n7726 , n50 , n7684 );
nand ( n7727 , n7725 , n7726 );
not ( n7728 , n7727 );
nand ( n7729 , n7708 , n7693 );
not ( n7730 , n7707 );
not ( n7731 , n7693 );
not ( n7732 , n7731 );
or ( n7733 , n7730 , n7732 );
nand ( n7734 , n7733 , n7699 );
nand ( n7735 , n7729 , n7734 );
not ( n7736 , n7735 );
not ( n7737 , n7736 );
or ( n7738 , n7728 , n7737 );
not ( n7739 , n7729 );
not ( n7740 , n7734 );
or ( n7741 , n7739 , n7740 );
not ( n7742 , n7727 );
nand ( n7743 , n7741 , n7742 );
nand ( n7744 , n7738 , n7743 );
xor ( n7745 , n7722 , n7744 );
xor ( n7746 , n40 , n61 );
not ( n7747 , n7746 );
not ( n7748 , n6616 );
or ( n7749 , n7747 , n7748 );
nand ( n7750 , n3236 , n7510 );
nand ( n7751 , n7749 , n7750 );
not ( n7752 , n7751 );
xor ( n7753 , n38 , n63 );
not ( n7754 , n7753 );
not ( n7755 , n6638 );
or ( n7756 , n7754 , n7755 );
nand ( n7757 , n4321 , n7530 );
nand ( n7758 , n7756 , n7757 );
not ( n7759 , n7520 );
not ( n7760 , n4248 );
or ( n7761 , n7759 , n7760 );
and ( n7762 , n44 , n57 );
not ( n7763 , n44 );
and ( n7764 , n7763 , n6713 );
nor ( n7765 , n7762 , n7764 );
nand ( n7766 , n6917 , n7765 );
nand ( n7767 , n7761 , n7766 );
not ( n7768 , n7767 );
and ( n7769 , n7758 , n7768 );
not ( n7770 , n7758 );
not ( n7771 , n7768 );
and ( n7772 , n7770 , n7771 );
nor ( n7773 , n7769 , n7772 );
not ( n7774 , n7773 );
or ( n7775 , n7752 , n7774 );
not ( n7776 , n7771 );
nand ( n7777 , n7758 , n7776 );
nand ( n7778 , n7775 , n7777 );
not ( n7779 , n7778 );
xnor ( n7780 , n7745 , n7779 );
xor ( n7781 , n7720 , n7780 );
not ( n7782 , n7781 );
not ( n7783 , n7694 );
not ( n7784 , n7081 );
not ( n7785 , n7784 );
or ( n7786 , n7783 , n7785 );
nand ( n7787 , n7602 , n7077 );
nand ( n7788 , n7786 , n7787 );
not ( n7789 , n7788 );
xor ( n7790 , n38 , n64 );
not ( n7791 , n7790 );
not ( n7792 , n6638 );
or ( n7793 , n7791 , n7792 );
nand ( n7794 , n3112 , n7753 );
nand ( n7795 , n7793 , n7794 );
not ( n7796 , n7795 );
not ( n7797 , n7595 );
not ( n7798 , n6615 );
or ( n7799 , n7797 , n7798 );
nand ( n7800 , n3234 , n7746 );
nand ( n7801 , n7799 , n7800 );
not ( n7802 , n7801 );
not ( n7803 , n7802 );
or ( n7804 , n7796 , n7803 );
not ( n7805 , n7801 );
or ( n7806 , n7805 , n7795 );
nand ( n7807 , n7804 , n7806 );
not ( n7808 , n7807 );
or ( n7809 , n7789 , n7808 );
not ( n7810 , n7805 );
nand ( n7811 , n7810 , n7795 );
nand ( n7812 , n7809 , n7811 );
not ( n7813 , n7812 );
not ( n7814 , n7587 );
not ( n7815 , n6706 );
or ( n7816 , n7814 , n7815 );
nand ( n7817 , n3634 , n7688 );
nand ( n7818 , n7816 , n7817 );
not ( n7819 , n7818 );
not ( n7820 , n7658 );
not ( n7821 , n7405 );
or ( n7822 , n7820 , n7821 );
nand ( n7823 , n7765 , n3464 );
nand ( n7824 , n7822 , n7823 );
not ( n7825 , n7633 );
not ( n7826 , n6595 );
not ( n7827 , n7826 );
or ( n7828 , n7825 , n7827 );
nand ( n7829 , n3121 , n7677 );
nand ( n7830 , n7828 , n7829 );
and ( n7831 , n7824 , n7830 );
not ( n7832 , n7824 );
not ( n7833 , n7830 );
and ( n7834 , n7832 , n7833 );
nor ( n7835 , n7831 , n7834 );
not ( n7836 , n7835 );
or ( n7837 , n7819 , n7836 );
not ( n7838 , n7833 );
nand ( n7839 , n7838 , n7824 );
nand ( n7840 , n7837 , n7839 );
not ( n7841 , n7638 );
not ( n7842 , n5655 );
not ( n7843 , n7627 );
or ( n7844 , n7842 , n7843 );
nand ( n7845 , n7844 , n4042 );
xor ( n7846 , n7841 , n7845 );
not ( n7847 , n7846 );
not ( n7848 , n7648 );
not ( n7849 , n7314 );
or ( n7850 , n7848 , n7849 );
nand ( n7851 , n7319 , n7701 );
nand ( n7852 , n7850 , n7851 );
not ( n7853 , n7852 );
or ( n7854 , n7847 , n7853 );
nand ( n7855 , n7841 , n7845 );
nand ( n7856 , n7854 , n7855 );
and ( n7857 , n7840 , n7856 );
not ( n7858 , n7840 );
not ( n7859 , n7856 );
and ( n7860 , n7858 , n7859 );
nor ( n7861 , n7857 , n7860 );
not ( n7862 , n7861 );
or ( n7863 , n7813 , n7862 );
not ( n7864 , n7859 );
nand ( n7865 , n7864 , n7840 );
nand ( n7866 , n7863 , n7865 );
not ( n7867 , n7490 );
not ( n7868 , n7867 );
and ( n7869 , n7504 , n7868 );
not ( n7870 , n7504 );
and ( n7871 , n7870 , n7867 );
nor ( n7872 , n7869 , n7871 );
not ( n7873 , n7872 );
not ( n7874 , n7322 );
not ( n7875 , n7874 );
not ( n7876 , n7681 );
not ( n7877 , n6596 );
or ( n7878 , n7876 , n7877 );
nand ( n7879 , n3521 , n7324 );
nand ( n7880 , n7878 , n7879 );
and ( n7881 , n7880 , n7767 );
not ( n7882 , n7880 );
and ( n7883 , n7882 , n7768 );
nor ( n7884 , n7881 , n7883 );
not ( n7885 , n7884 );
not ( n7886 , n7885 );
or ( n7887 , n7875 , n7886 );
nand ( n7888 , n7322 , n7884 );
nand ( n7889 , n7887 , n7888 );
not ( n7890 , n7889 );
or ( n7891 , n7873 , n7890 );
or ( n7892 , n7872 , n7889 );
nand ( n7893 , n7891 , n7892 );
not ( n7894 , n7893 );
and ( n7895 , n7866 , n7894 );
not ( n7896 , n7866 );
and ( n7897 , n7896 , n7893 );
nor ( n7898 , n7895 , n7897 );
not ( n7899 , n7898 );
and ( n7900 , n7861 , n7812 );
not ( n7901 , n7861 );
not ( n7902 , n7812 );
and ( n7903 , n7901 , n7902 );
nor ( n7904 , n7900 , n7903 );
not ( n7905 , n7904 );
xor ( n7906 , n7767 , n7758 );
xor ( n7907 , n7906 , n7751 );
xnor ( n7908 , n7788 , n7807 );
xnor ( n7909 , n7846 , n7852 );
not ( n7910 , n7909 );
not ( n7911 , n7818 );
not ( n7912 , n7835 );
not ( n7913 , n7912 );
or ( n7914 , n7911 , n7913 );
not ( n7915 , n7818 );
nand ( n7916 , n7915 , n7835 );
nand ( n7917 , n7914 , n7916 );
nor ( n7918 , n7910 , n7917 );
or ( n7919 , n7908 , n7918 );
not ( n7920 , n7909 );
nand ( n7921 , n7920 , n7917 );
nand ( n7922 , n7919 , n7921 );
not ( n7923 , n7922 );
and ( n7924 , n7907 , n7923 );
not ( n7925 , n7907 );
not ( n7926 , n7923 );
and ( n7927 , n7925 , n7926 );
nor ( n7928 , n7924 , n7927 );
not ( n7929 , n7928 );
or ( n7930 , n7905 , n7929 );
not ( n7931 , n7907 );
nand ( n7932 , n7931 , n7926 );
nand ( n7933 , n7930 , n7932 );
not ( n7934 , n7933 );
or ( n7935 , n7899 , n7934 );
or ( n7936 , n7898 , n7933 );
nand ( n7937 , n7935 , n7936 );
not ( n7938 , n7937 );
or ( n7939 , n7782 , n7938 );
not ( n7940 , n7898 );
nand ( n7941 , n7940 , n7933 );
nand ( n7942 , n7939 , n7941 );
not ( n7943 , n7942 );
not ( n7944 , n7866 );
not ( n7945 , n7893 );
or ( n7946 , n7944 , n7945 );
not ( n7947 , n7872 );
nand ( n7948 , n7947 , n7889 );
nand ( n7949 , n7946 , n7948 );
not ( n7950 , n7722 );
not ( n7951 , n7744 );
or ( n7952 , n7950 , n7951 );
not ( n7953 , n7742 );
nand ( n7954 , n7953 , n7735 );
nand ( n7955 , n7952 , n7954 );
not ( n7956 , n7542 );
not ( n7957 , n7482 );
and ( n7958 , n7956 , n7957 );
and ( n7959 , n7482 , n7542 );
nor ( n7960 , n7958 , n7959 );
xnor ( n7961 , n7955 , n7960 );
xor ( n7962 , n7949 , n7961 );
not ( n7963 , n7962 );
and ( n7964 , n7342 , n7334 );
not ( n7965 , n7342 );
and ( n7966 , n7965 , n7329 );
nor ( n7967 , n7964 , n7966 );
not ( n7968 , n7322 );
xor ( n7969 , n7967 , n7968 );
not ( n7970 , n7968 );
not ( n7971 , n7884 );
or ( n7972 , n7970 , n7971 );
nand ( n7973 , n7880 , n7771 );
nand ( n7974 , n7972 , n7973 );
not ( n7975 , n7974 );
xnor ( n7976 , n7416 , n7399 );
not ( n7977 , n7976 );
and ( n7978 , n7975 , n7977 );
not ( n7979 , n7975 );
and ( n7980 , n7979 , n7976 );
nor ( n7981 , n7978 , n7980 );
xor ( n7982 , n7969 , n7981 );
not ( n7983 , n7982 );
not ( n7984 , n7720 );
not ( n7985 , n7780 );
or ( n7986 , n7984 , n7985 );
not ( n7987 , n7779 );
xor ( n7988 , n7722 , n7744 );
nand ( n7989 , n7987 , n7988 );
nand ( n7990 , n7986 , n7989 );
not ( n7991 , n7990 );
or ( n7992 , n7983 , n7991 );
or ( n7993 , n7982 , n7990 );
nand ( n7994 , n7992 , n7993 );
nand ( n7995 , n7963 , n7994 );
not ( n7996 , n7995 );
not ( n7997 , n7962 );
nor ( n7998 , n7997 , n7994 );
nor ( n7999 , n7996 , n7998 );
nand ( n8000 , n7943 , n7999 );
not ( n8001 , n7259 );
not ( n8002 , n7222 );
and ( n8003 , n8001 , n8002 );
and ( n8004 , n7222 , n7259 );
nor ( n8005 , n8003 , n8004 );
not ( n8006 , n7301 );
not ( n8007 , n7459 );
or ( n8008 , n8006 , n8007 );
nand ( n8009 , n7458 , n7453 );
nand ( n8010 , n8008 , n8009 );
not ( n8011 , n8010 );
nand ( n8012 , n8005 , n8011 );
buf ( n8013 , n8012 );
nand ( n8014 , n7582 , n8000 , n8013 );
nor ( n8015 , n7943 , n7999 );
xnor ( n8016 , n7589 , n7609 );
not ( n8017 , n8016 );
not ( n8018 , n8017 );
xor ( n8019 , n7640 , n7650 );
not ( n8020 , n7664 );
xor ( n8021 , n8019 , n8020 );
not ( n8022 , n8021 );
not ( n8023 , n7662 );
not ( n8024 , n5588 );
or ( n8025 , n8023 , n8024 );
not ( n8026 , n6916 );
xor ( n8027 , n44 , n60 );
nand ( n8028 , n8026 , n8027 );
nand ( n8029 , n8025 , n8028 );
not ( n8030 , n8029 );
not ( n8031 , n8030 );
xor ( n8032 , n42 , n62 );
not ( n8033 , n8032 );
not ( n8034 , n6705 );
or ( n8035 , n8033 , n8034 );
nand ( n8036 , n3348 , n7583 );
nand ( n8037 , n8035 , n8036 );
nor ( n8038 , n8031 , n8037 );
xor ( n8039 , n46 , n58 );
not ( n8040 , n8039 );
not ( n8041 , n7076 );
not ( n8042 , n8041 );
or ( n8043 , n8040 , n8042 );
nand ( n8044 , n7598 , n7187 );
nand ( n8045 , n8043 , n8044 );
not ( n8046 , n8045 );
or ( n8047 , n8038 , n8046 );
nand ( n8048 , n8037 , n8031 );
nand ( n8049 , n8047 , n8048 );
not ( n8050 , n8049 );
or ( n8051 , n8022 , n8050 );
or ( n8052 , n8049 , n8021 );
nand ( n8053 , n8051 , n8052 );
not ( n8054 , n8053 );
or ( n8055 , n8018 , n8054 );
not ( n8056 , n8021 );
nand ( n8057 , n8049 , n8056 );
nand ( n8058 , n8055 , n8057 );
not ( n8059 , n8058 );
xor ( n8060 , n38 , n65 );
not ( n8061 , n8060 );
not ( n8062 , n6638 );
or ( n8063 , n8061 , n8062 );
nand ( n8064 , n3112 , n7790 );
nand ( n8065 , n8063 , n8064 );
not ( n8066 , n8065 );
and ( n8067 , n7629 , n7622 );
not ( n8068 , n7629 );
and ( n8069 , n8068 , n7621 );
or ( n8070 , n8067 , n8069 );
not ( n8071 , n8070 );
or ( n8072 , n8066 , n8071 );
or ( n8073 , n8065 , n8070 );
nand ( n8074 , n8072 , n8073 );
not ( n8075 , n8074 );
xor ( n8076 , n48 , n56 );
not ( n8077 , n8076 );
not ( n8078 , n7313 );
not ( n8079 , n8078 );
or ( n8080 , n8077 , n8079 );
nand ( n8081 , n7318 , n7644 );
nand ( n8082 , n8080 , n8081 );
not ( n8083 , n8082 );
not ( n8084 , n5655 );
xor ( n8085 , n50 , n54 );
not ( n8086 , n8085 );
or ( n8087 , n8084 , n8086 );
nand ( n8088 , n51 , n7624 );
nand ( n8089 , n8087 , n8088 );
nand ( n8090 , n67 , n3121 );
not ( n8091 , n8090 );
and ( n8092 , n8089 , n8091 );
not ( n8093 , n8089 );
not ( n8094 , n8091 );
and ( n8095 , n8093 , n8094 );
nor ( n8096 , n8092 , n8095 );
not ( n8097 , n8096 );
or ( n8098 , n8083 , n8097 );
not ( n8099 , n8094 );
nand ( n8100 , n8099 , n8089 );
nand ( n8101 , n8098 , n8100 );
not ( n8102 , n8101 );
not ( n8103 , n8102 );
not ( n8104 , n8103 );
or ( n8105 , n8075 , n8104 );
not ( n8106 , n8070 );
nand ( n8107 , n8065 , n8106 );
nand ( n8108 , n8105 , n8107 );
not ( n8109 , n8108 );
not ( n8110 , n8109 );
xor ( n8111 , n7614 , n7670 );
not ( n8112 , n8111 );
or ( n8113 , n8110 , n8112 );
or ( n8114 , n8109 , n8111 );
nand ( n8115 , n8113 , n8114 );
not ( n8116 , n8115 );
or ( n8117 , n8059 , n8116 );
not ( n8118 , n8109 );
nand ( n8119 , n8118 , n8111 );
nand ( n8120 , n8117 , n8119 );
not ( n8121 , n8120 );
not ( n8122 , n7715 );
and ( n8123 , n7675 , n8122 );
not ( n8124 , n7675 );
and ( n8125 , n8124 , n7715 );
nor ( n8126 , n8123 , n8125 );
xor ( n8127 , n7907 , n7923 );
xnor ( n8128 , n8127 , n7904 );
and ( n8129 , n8126 , n8128 );
not ( n8130 , n8126 );
not ( n8131 , n8128 );
and ( n8132 , n8130 , n8131 );
nor ( n8133 , n8129 , n8132 );
not ( n8134 , n8133 );
or ( n8135 , n8121 , n8134 );
not ( n8136 , n8126 );
nand ( n8137 , n8136 , n8131 );
nand ( n8138 , n8135 , n8137 );
not ( n8139 , n8138 );
not ( n8140 , n7781 );
nand ( n8141 , n8140 , n7937 );
not ( n8142 , n8141 );
not ( n8143 , n7781 );
nor ( n8144 , n8143 , n7937 );
nor ( n8145 , n8142 , n8144 );
nor ( n8146 , n8139 , n8145 );
nor ( n8147 , n8015 , n8146 );
not ( n8148 , n8147 );
nand ( n8149 , n8139 , n8145 );
not ( n8150 , n8027 );
not ( n8151 , n3727 );
not ( n8152 , n8151 );
or ( n8153 , n8150 , n8152 );
xor ( n8154 , n44 , n61 );
nand ( n8155 , n8154 , n7105 );
nand ( n8156 , n8153 , n8155 );
not ( n8157 , n8156 );
xor ( n8158 , n42 , n63 );
not ( n8159 , n8158 );
not ( n8160 , n6705 );
or ( n8161 , n8159 , n8160 );
nand ( n8162 , n3348 , n8032 );
nand ( n8163 , n8161 , n8162 );
xor ( n8164 , n48 , n57 );
not ( n8165 , n8164 );
not ( n8166 , n7312 );
or ( n8167 , n8165 , n8166 );
buf ( n8168 , n7317 );
nand ( n8169 , n8168 , n8076 );
nand ( n8170 , n8167 , n8169 );
xor ( n8171 , n8163 , n8170 );
not ( n8172 , n8171 );
or ( n8173 , n8157 , n8172 );
nand ( n8174 , n8170 , n8163 );
nand ( n8175 , n8173 , n8174 );
not ( n8176 , n8175 );
xor ( n8177 , n8091 , n8089 );
xnor ( n8178 , n8177 , n8082 );
not ( n8179 , n8178 );
xnor ( n8180 , n59 , n46 );
or ( n8181 , n8180 , n7189 );
nand ( n8182 , n8039 , n7187 );
nand ( n8183 , n8181 , n8182 );
not ( n8184 , n8183 );
xor ( n8185 , n38 , n67 );
not ( n8186 , n8185 );
not ( n8187 , n6637 );
or ( n8188 , n8186 , n8187 );
xor ( n8189 , n38 , n66 );
nand ( n8190 , n3111 , n8189 );
nand ( n8191 , n8188 , n8190 );
xor ( n8192 , n40 , n65 );
not ( n8193 , n8192 );
not ( n8194 , n6614 );
or ( n8195 , n8193 , n8194 );
xor ( n8196 , n40 , n64 );
nand ( n8197 , n3220 , n8196 );
nand ( n8198 , n8195 , n8197 );
and ( n8199 , n8191 , n8198 );
not ( n8200 , n8191 );
not ( n8201 , n8198 );
and ( n8202 , n8200 , n8201 );
nor ( n8203 , n8199 , n8202 );
not ( n8204 , n8203 );
or ( n8205 , n8184 , n8204 );
not ( n8206 , n8201 );
nand ( n8207 , n8206 , n8191 );
nand ( n8208 , n8205 , n8207 );
not ( n8209 , n8208 );
or ( n8210 , n8179 , n8209 );
or ( n8211 , n8178 , n8208 );
nand ( n8212 , n8210 , n8211 );
not ( n8213 , n8212 );
or ( n8214 , n8176 , n8213 );
not ( n8215 , n8178 );
nand ( n8216 , n8215 , n8208 );
nand ( n8217 , n8214 , n8216 );
and ( n8218 , n8074 , n8101 );
not ( n8219 , n8074 );
and ( n8220 , n8219 , n8102 );
nor ( n8221 , n8218 , n8220 );
not ( n8222 , n8221 );
not ( n8223 , n8189 );
not ( n8224 , n6639 );
or ( n8225 , n8223 , n8224 );
nand ( n8226 , n3112 , n8060 );
nand ( n8227 , n8225 , n8226 );
not ( n8228 , n8227 );
not ( n8229 , n8196 );
not ( n8230 , n6614 );
or ( n8231 , n8229 , n8230 );
nand ( n8232 , n3234 , n7591 );
nand ( n8233 , n8231 , n8232 );
not ( n8234 , n5110 );
not ( n8235 , n67 );
nand ( n8236 , n8235 , n5105 );
not ( n8237 , n8236 );
or ( n8238 , n8234 , n8237 );
nand ( n8239 , n8238 , n38 );
not ( n8240 , n8239 );
not ( n8241 , n6264 );
xor ( n8242 , n50 , n55 );
not ( n8243 , n8242 );
or ( n8244 , n8241 , n8243 );
nand ( n8245 , n51 , n8085 );
nand ( n8246 , n8244 , n8245 );
nand ( n8247 , n8240 , n8246 );
xor ( n8248 , n8233 , n8247 );
not ( n8249 , n8248 );
not ( n8250 , n8249 );
or ( n8251 , n8228 , n8250 );
not ( n8252 , n8247 );
nand ( n8253 , n8252 , n8233 );
nand ( n8254 , n8251 , n8253 );
not ( n8255 , n8254 );
not ( n8256 , n8255 );
or ( n8257 , n8222 , n8256 );
not ( n8258 , n8254 );
or ( n8259 , n8258 , n8221 );
nand ( n8260 , n8257 , n8259 );
and ( n8261 , n8217 , n8260 );
not ( n8262 , n8217 );
not ( n8263 , n8260 );
and ( n8264 , n8262 , n8263 );
nor ( n8265 , n8261 , n8264 );
not ( n8266 , n8265 );
not ( n8267 , n8266 );
not ( n8268 , n8267 );
xor ( n8269 , n40 , n66 );
not ( n8270 , n8269 );
not ( n8271 , n6615 );
or ( n8272 , n8270 , n8271 );
nand ( n8273 , n3235 , n8192 );
nand ( n8274 , n8272 , n8273 );
not ( n8275 , n8274 );
xor ( n8276 , n42 , n64 );
not ( n8277 , n8276 );
not ( n8278 , n6705 );
or ( n8279 , n8277 , n8278 );
nand ( n8280 , n3348 , n8158 );
nand ( n8281 , n8279 , n8280 );
not ( n8282 , n6264 );
xor ( n8283 , n50 , n56 );
not ( n8284 , n8283 );
or ( n8285 , n8282 , n8284 );
nand ( n8286 , n51 , n8242 );
nand ( n8287 , n8285 , n8286 );
xor ( n8288 , n8281 , n8287 );
not ( n8289 , n8288 );
or ( n8290 , n8275 , n8289 );
nand ( n8291 , n8287 , n8281 );
nand ( n8292 , n8290 , n8291 );
not ( n8293 , n8292 );
xnor ( n8294 , n8246 , n8240 );
xor ( n8295 , n48 , n58 );
not ( n8296 , n8295 );
not ( n8297 , n7312 );
or ( n8298 , n8296 , n8297 );
nand ( n8299 , n7318 , n8164 );
nand ( n8300 , n8298 , n8299 );
not ( n8301 , n8300 );
and ( n8302 , n67 , n3087 );
not ( n8303 , n8302 );
not ( n8304 , n8303 );
xor ( n8305 , n44 , n62 );
not ( n8306 , n8305 );
nand ( n8307 , n3451 , n6913 );
not ( n8308 , n8307 );
not ( n8309 , n8308 );
or ( n8310 , n8306 , n8309 );
nand ( n8311 , n8154 , n3463 );
nand ( n8312 , n8310 , n8311 );
not ( n8313 , n8312 );
or ( n8314 , n8304 , n8313 );
or ( n8315 , n8303 , n8312 );
nand ( n8316 , n8314 , n8315 );
not ( n8317 , n8316 );
or ( n8318 , n8301 , n8317 );
not ( n8319 , n8303 );
nand ( n8320 , n8319 , n8312 );
nand ( n8321 , n8318 , n8320 );
xnor ( n8322 , n8294 , n8321 );
not ( n8323 , n8322 );
or ( n8324 , n8293 , n8323 );
not ( n8325 , n8294 );
nand ( n8326 , n8325 , n8321 );
nand ( n8327 , n8324 , n8326 );
not ( n8328 , n8327 );
not ( n8329 , n8227 );
and ( n8330 , n8248 , n8329 );
not ( n8331 , n8248 );
and ( n8332 , n8331 , n8227 );
nor ( n8333 , n8330 , n8332 );
not ( n8334 , n8333 );
not ( n8335 , n8334 );
not ( n8336 , n8037 );
not ( n8337 , n8030 );
or ( n8338 , n8336 , n8337 );
or ( n8339 , n8030 , n8037 );
nand ( n8340 , n8338 , n8339 );
and ( n8341 , n8340 , n8046 );
not ( n8342 , n8340 );
and ( n8343 , n8342 , n8045 );
nor ( n8344 , n8341 , n8343 );
not ( n8345 , n8344 );
not ( n8346 , n8345 );
or ( n8347 , n8335 , n8346 );
nand ( n8348 , n8333 , n8344 );
nand ( n8349 , n8347 , n8348 );
not ( n8350 , n8349 );
or ( n8351 , n8328 , n8350 );
nand ( n8352 , n8333 , n8345 );
nand ( n8353 , n8351 , n8352 );
not ( n8354 , n8353 );
not ( n8355 , n8053 );
not ( n8356 , n8016 );
and ( n8357 , n8355 , n8356 );
and ( n8358 , n8016 , n8053 );
nor ( n8359 , n8357 , n8358 );
not ( n8360 , n8359 );
or ( n8361 , n8354 , n8360 );
or ( n8362 , n8359 , n8353 );
nand ( n8363 , n8361 , n8362 );
not ( n8364 , n8363 );
or ( n8365 , n8268 , n8364 );
not ( n8366 , n8359 );
nand ( n8367 , n8366 , n8353 );
nand ( n8368 , n8365 , n8367 );
not ( n8369 , n8115 );
not ( n8370 , n8058 );
not ( n8371 , n8370 );
or ( n8372 , n8369 , n8371 );
or ( n8373 , n8370 , n8115 );
nand ( n8374 , n8372 , n8373 );
not ( n8375 , n8374 );
not ( n8376 , n7921 );
not ( n8377 , n8376 );
buf ( n8378 , n7908 );
not ( n8379 , n8378 );
not ( n8380 , n8379 );
or ( n8381 , n8377 , n8380 );
not ( n8382 , n7910 );
buf ( n8383 , n7917 );
not ( n8384 , n8383 );
nand ( n8385 , n8379 , n8382 , n8384 );
nand ( n8386 , n8381 , n8385 );
not ( n8387 , n8378 );
xor ( n8388 , n8382 , n8383 );
nor ( n8389 , n8387 , n8388 );
nor ( n8390 , n8386 , n8389 );
not ( n8391 , n8390 );
not ( n8392 , n8217 );
not ( n8393 , n8260 );
or ( n8394 , n8392 , n8393 );
not ( n8395 , n8258 );
nand ( n8396 , n8395 , n8221 );
nand ( n8397 , n8394 , n8396 );
not ( n8398 , n8397 );
and ( n8399 , n8391 , n8398 );
and ( n8400 , n8390 , n8397 );
nor ( n8401 , n8399 , n8400 );
not ( n8402 , n8401 );
or ( n8403 , n8375 , n8402 );
or ( n8404 , n8374 , n8401 );
nand ( n8405 , n8403 , n8404 );
nand ( n8406 , n8368 , n8405 );
not ( n8407 , n8406 );
not ( n8408 , n8374 );
not ( n8409 , n8401 );
not ( n8410 , n8409 );
or ( n8411 , n8408 , n8410 );
not ( n8412 , n8390 );
nand ( n8413 , n8412 , n8397 );
nand ( n8414 , n8411 , n8413 );
not ( n8415 , n8414 );
xor ( n8416 , n8126 , n8128 );
xnor ( n8417 , n8416 , n8120 );
nand ( n8418 , n8415 , n8417 );
nand ( n8419 , n8407 , n8418 );
not ( n8420 , n8415 );
not ( n8421 , n8417 );
nand ( n8422 , n8420 , n8421 );
nand ( n8423 , n8419 , n8422 );
nand ( n8424 , n8149 , n8423 );
not ( n8425 , n8424 );
or ( n8426 , n8148 , n8425 );
xor ( n8427 , n7562 , n7568 );
xnor ( n8428 , n8427 , n7555 );
xor ( n8429 , n7469 , n7550 );
not ( n8430 , n8429 );
not ( n8431 , n7969 );
not ( n8432 , n7981 );
not ( n8433 , n8432 );
or ( n8434 , n8431 , n8433 );
or ( n8435 , n7976 , n7975 );
nand ( n8436 , n8434 , n8435 );
not ( n8437 , n8436 );
not ( n8438 , n7949 );
not ( n8439 , n7961 );
or ( n8440 , n8438 , n8439 );
not ( n8441 , n7960 );
nand ( n8442 , n7955 , n8441 );
nand ( n8443 , n8440 , n8442 );
not ( n8444 , n8443 );
not ( n8445 , n8444 );
or ( n8446 , n8437 , n8445 );
not ( n8447 , n8436 );
nand ( n8448 , n8447 , n8443 );
nand ( n8449 , n8446 , n8448 );
not ( n8450 , n8449 );
or ( n8451 , n8430 , n8450 );
nand ( n8452 , n8436 , n8443 );
nand ( n8453 , n8451 , n8452 );
not ( n8454 , n8453 );
nand ( n8455 , n8428 , n8454 );
not ( n8456 , n7962 );
not ( n8457 , n7994 );
or ( n8458 , n8456 , n8457 );
not ( n8459 , n7982 );
nand ( n8460 , n8459 , n7990 );
nand ( n8461 , n8458 , n8460 );
not ( n8462 , n8461 );
not ( n8463 , n8449 );
and ( n8464 , n8429 , n8463 );
not ( n8465 , n8429 );
and ( n8466 , n8465 , n8449 );
nor ( n8467 , n8464 , n8466 );
nand ( n8468 , n8462 , n8467 );
and ( n8469 , n8455 , n8468 );
nand ( n8470 , n8426 , n8469 );
nor ( n8471 , n8014 , n8470 );
not ( n8472 , n8471 );
nor ( n8473 , n8428 , n8454 );
not ( n8474 , n8473 );
not ( n8475 , n8454 );
not ( n8476 , n8428 );
or ( n8477 , n8475 , n8476 );
nor ( n8478 , n8467 , n8462 );
nand ( n8479 , n8477 , n8478 );
nand ( n8480 , n8474 , n8479 );
not ( n8481 , n7464 );
and ( n8482 , n8481 , n7578 );
or ( n8483 , n8480 , n8482 );
and ( n8484 , n8012 , n7580 );
nand ( n8485 , n8483 , n8484 );
not ( n8486 , n8011 );
not ( n8487 , n8005 );
nand ( n8488 , n8486 , n8487 );
nand ( n8489 , n8485 , n8488 );
not ( n8490 , n8489 );
nand ( n8491 , n8000 , n8149 );
not ( n8492 , n8368 );
not ( n8493 , n8405 );
nand ( n8494 , n8492 , n8493 );
and ( n8495 , n8494 , n8418 );
not ( n8496 , n8495 );
nor ( n8497 , n8491 , n8496 );
xor ( n8498 , n8327 , n8349 );
not ( n8499 , n8498 );
not ( n8500 , n8175 );
not ( n8501 , n8500 );
not ( n8502 , n8212 );
and ( n8503 , n8501 , n8502 );
and ( n8504 , n8500 , n8212 );
nor ( n8505 , n8503 , n8504 );
not ( n8506 , n8505 );
not ( n8507 , n8506 );
xor ( n8508 , n46 , n60 );
not ( n8509 , n8508 );
not ( n8510 , n7075 );
or ( n8511 , n8509 , n8510 );
or ( n8512 , n8180 , n7081 );
nand ( n8513 , n8511 , n8512 );
not ( n8514 , n8513 );
not ( n8515 , n8514 );
nand ( n8516 , n41 , n42 );
nand ( n8517 , n40 , n8516 );
not ( n8518 , n8517 );
or ( n8519 , n41 , n42 );
nand ( n8520 , n8519 , n67 );
nand ( n8521 , n8518 , n8520 );
not ( n8522 , n8521 );
xor ( n8523 , n48 , n59 );
not ( n8524 , n8523 );
not ( n8525 , n7310 );
and ( n8526 , n3561 , n8525 );
not ( n8527 , n8526 );
or ( n8528 , n8524 , n8527 );
nand ( n8529 , n7317 , n8295 );
nand ( n8530 , n8528 , n8529 );
and ( n8531 , n8522 , n8530 );
not ( n8532 , n8531 );
or ( n8533 , n8515 , n8532 );
not ( n8534 , n8522 );
not ( n8535 , n8530 );
or ( n8536 , n8534 , n8535 );
nand ( n8537 , n8536 , n8513 );
nand ( n8538 , n8533 , n8537 );
not ( n8539 , n8538 );
not ( n8540 , n8305 );
not ( n8541 , n8151 );
or ( n8542 , n8540 , n8541 );
xor ( n8543 , n44 , n63 );
nand ( n8544 , n8543 , n7105 );
nand ( n8545 , n8542 , n8544 );
not ( n8546 , n8545 );
not ( n8547 , n4888 );
xor ( n8548 , n50 , n57 );
not ( n8549 , n8548 );
or ( n8550 , n8547 , n8549 );
nand ( n8551 , n51 , n8283 );
nand ( n8552 , n8550 , n8551 );
not ( n8553 , n8552 );
not ( n8554 , n8553 );
xor ( n8555 , n42 , n65 );
not ( n8556 , n8555 );
not ( n8557 , n6705 );
or ( n8558 , n8556 , n8557 );
nand ( n8559 , n3348 , n8276 );
nand ( n8560 , n8558 , n8559 );
not ( n8561 , n8560 );
or ( n8562 , n8554 , n8561 );
or ( n8563 , n8553 , n8560 );
nand ( n8564 , n8562 , n8563 );
not ( n8565 , n8564 );
or ( n8566 , n8546 , n8565 );
not ( n8567 , n8553 );
nand ( n8568 , n8567 , n8560 );
nand ( n8569 , n8566 , n8568 );
not ( n8570 , n8569 );
or ( n8571 , n8539 , n8570 );
not ( n8572 , n8514 );
nand ( n8573 , n8572 , n8531 );
nand ( n8574 , n8571 , n8573 );
not ( n8575 , n8574 );
xor ( n8576 , n8156 , n8171 );
not ( n8577 , n8576 );
not ( n8578 , n8577 );
xnor ( n8579 , n8183 , n8203 );
not ( n8580 , n8579 );
not ( n8581 , n8580 );
or ( n8582 , n8578 , n8581 );
nand ( n8583 , n8576 , n8579 );
nand ( n8584 , n8582 , n8583 );
not ( n8585 , n8584 );
or ( n8586 , n8575 , n8585 );
not ( n8587 , n8579 );
nand ( n8588 , n8576 , n8587 );
nand ( n8589 , n8586 , n8588 );
not ( n8590 , n8589 );
not ( n8591 , n8590 );
or ( n8592 , n8507 , n8591 );
nand ( n8593 , n8505 , n8589 );
nand ( n8594 , n8592 , n8593 );
nand ( n8595 , n8499 , n8594 );
not ( n8596 , n8595 );
not ( n8597 , n8498 );
nor ( n8598 , n8594 , n8597 );
nor ( n8599 , n8596 , n8598 );
and ( n8600 , n8584 , n8574 );
not ( n8601 , n8584 );
not ( n8602 , n8574 );
and ( n8603 , n8601 , n8602 );
nor ( n8604 , n8600 , n8603 );
not ( n8605 , n8604 );
not ( n8606 , n8605 );
not ( n8607 , n8606 );
xor ( n8608 , n8292 , n8322 );
not ( n8609 , n8608 );
not ( n8610 , n8281 );
xor ( n8611 , n8287 , n8610 );
xnor ( n8612 , n8611 , n8274 );
not ( n8613 , n8612 );
not ( n8614 , n8312 );
xor ( n8615 , n8302 , n8614 );
xnor ( n8616 , n8615 , n8300 );
not ( n8617 , n8616 );
not ( n8618 , n3220 );
not ( n8619 , n8269 );
or ( n8620 , n8618 , n8619 );
and ( n8621 , n6611 , n6613 , n3218 );
nor ( n8622 , n40 , n67 );
not ( n8623 , n8622 );
nand ( n8624 , n40 , n67 );
nand ( n8625 , n8621 , n8623 , n8624 );
nand ( n8626 , n8620 , n8625 );
xor ( n8627 , n46 , n61 );
not ( n8628 , n8627 );
not ( n8629 , n7073 );
not ( n8630 , n8629 );
or ( n8631 , n8628 , n8630 );
not ( n8632 , n8508 );
or ( n8633 , n8632 , n3609 );
nand ( n8634 , n8631 , n8633 );
not ( n8635 , n8634 );
not ( n8636 , n8635 );
nand ( n8637 , n8626 , n8636 );
not ( n8638 , n8637 );
xor ( n8639 , n8522 , n8530 );
not ( n8640 , n8634 );
nor ( n8641 , n8626 , n8640 );
not ( n8642 , n8641 );
nand ( n8643 , n8626 , n8635 );
nand ( n8644 , n8642 , n8643 );
nand ( n8645 , n8639 , n8644 );
not ( n8646 , n8645 );
nor ( n8647 , n8638 , n8646 );
not ( n8648 , n8647 );
or ( n8649 , n8617 , n8648 );
not ( n8650 , n8637 );
not ( n8651 , n8645 );
or ( n8652 , n8650 , n8651 );
not ( n8653 , n8616 );
nand ( n8654 , n8652 , n8653 );
nand ( n8655 , n8649 , n8654 );
not ( n8656 , n8655 );
or ( n8657 , n8613 , n8656 );
not ( n8658 , n8637 );
not ( n8659 , n8645 );
or ( n8660 , n8658 , n8659 );
nand ( n8661 , n8660 , n8616 );
nand ( n8662 , n8657 , n8661 );
not ( n8663 , n8662 );
not ( n8664 , n8663 );
or ( n8665 , n8609 , n8664 );
not ( n8666 , n8662 );
or ( n8667 , n8608 , n8666 );
nand ( n8668 , n8665 , n8667 );
not ( n8669 , n8668 );
or ( n8670 , n8607 , n8669 );
not ( n8671 , n8666 );
nand ( n8672 , n8608 , n8671 );
nand ( n8673 , n8670 , n8672 );
not ( n8674 , n8673 );
nand ( n8675 , n8599 , n8674 );
not ( n8676 , n8675 );
xor ( n8677 , n8569 , n8538 );
not ( n8678 , n8560 );
xor ( n8679 , n8552 , n8678 );
not ( n8680 , n8545 );
xnor ( n8681 , n8679 , n8680 );
not ( n8682 , n8681 );
not ( n8683 , n8682 );
not ( n8684 , n8627 );
not ( n8685 , n7187 );
or ( n8686 , n8684 , n8685 );
xor ( n8687 , n46 , n62 );
nand ( n8688 , n8687 , n7075 );
nand ( n8689 , n8686 , n8688 );
not ( n8690 , n8689 );
not ( n8691 , n6196 );
xor ( n8692 , n50 , n58 );
not ( n8693 , n8692 );
or ( n8694 , n8691 , n8693 );
nand ( n8695 , n51 , n8548 );
nand ( n8696 , n8694 , n8695 );
not ( n8697 , n8696 );
xor ( n8698 , n42 , n66 );
not ( n8699 , n8698 );
not ( n8700 , n7494 );
or ( n8701 , n8699 , n8700 );
nand ( n8702 , n3355 , n8555 );
nand ( n8703 , n8701 , n8702 );
not ( n8704 , n8703 );
not ( n8705 , n8704 );
or ( n8706 , n8697 , n8705 );
not ( n8707 , n8703 );
or ( n8708 , n8696 , n8707 );
nand ( n8709 , n8706 , n8708 );
not ( n8710 , n8709 );
or ( n8711 , n8690 , n8710 );
not ( n8712 , n8707 );
nand ( n8713 , n8696 , n8712 );
nand ( n8714 , n8711 , n8713 );
nand ( n8715 , n67 , n3220 );
not ( n8716 , n8715 );
not ( n8717 , n8716 );
xor ( n8718 , n48 , n60 );
not ( n8719 , n8718 );
not ( n8720 , n8526 );
or ( n8721 , n8719 , n8720 );
nand ( n8722 , n7317 , n8523 );
nand ( n8723 , n8721 , n8722 );
not ( n8724 , n8723 );
or ( n8725 , n8717 , n8724 );
or ( n8726 , n8716 , n8723 );
not ( n8727 , n8543 );
not ( n8728 , n3726 );
or ( n8729 , n8727 , n8728 );
xor ( n8730 , n44 , n64 );
nand ( n8731 , n8730 , n7405 );
nand ( n8732 , n8729 , n8731 );
nand ( n8733 , n8726 , n8732 );
nand ( n8734 , n8725 , n8733 );
xor ( n8735 , n8714 , n8734 );
not ( n8736 , n8735 );
or ( n8737 , n8683 , n8736 );
not ( n8738 , n8714 );
not ( n8739 , n8738 );
nand ( n8740 , n8734 , n8739 );
nand ( n8741 , n8737 , n8740 );
not ( n8742 , n8741 );
xor ( n8743 , n8677 , n8742 );
xnor ( n8744 , n8655 , n8612 );
xor ( n8745 , n8743 , n8744 );
not ( n8746 , n67 );
not ( n8747 , n8746 );
not ( n8748 , n6706 );
or ( n8749 , n8747 , n8748 );
nand ( n8750 , n3349 , n8698 );
nand ( n8751 , n8749 , n8750 );
not ( n8752 , n8751 );
not ( n8753 , n6264 );
xor ( n8754 , n50 , n59 );
not ( n8755 , n8754 );
or ( n8756 , n8753 , n8755 );
nand ( n8757 , n51 , n8692 );
nand ( n8758 , n8756 , n8757 );
not ( n8759 , n8758 );
not ( n8760 , n8730 );
not ( n8761 , n3464 );
or ( n8762 , n8760 , n8761 );
xor ( n8763 , n44 , n65 );
nand ( n8764 , n6915 , n8763 );
nand ( n8765 , n8762 , n8764 );
not ( n8766 , n8765 );
not ( n8767 , n8766 );
or ( n8768 , n8759 , n8767 );
not ( n8769 , n8765 );
or ( n8770 , n8758 , n8769 );
nand ( n8771 , n8768 , n8770 );
not ( n8772 , n8771 );
or ( n8773 , n8752 , n8772 );
not ( n8774 , n8769 );
nand ( n8775 , n8758 , n8774 );
nand ( n8776 , n8773 , n8775 );
not ( n8777 , n8776 );
not ( n8778 , n8777 );
not ( n8779 , n8778 );
not ( n8780 , n67 );
nand ( n8781 , n8780 , n5688 );
not ( n8782 , n8781 );
not ( n8783 , n5693 );
or ( n8784 , n8782 , n8783 );
nand ( n8785 , n8784 , n42 );
not ( n8786 , n8785 );
xor ( n8787 , n48 , n61 );
not ( n8788 , n8787 );
not ( n8789 , n8526 );
or ( n8790 , n8788 , n8789 );
nand ( n8791 , n7317 , n8718 );
nand ( n8792 , n8790 , n8791 );
nand ( n8793 , n8786 , n8792 );
not ( n8794 , n8793 );
xor ( n8795 , n8715 , n8723 );
xnor ( n8796 , n8795 , n8732 );
not ( n8797 , n8796 );
or ( n8798 , n8794 , n8797 );
or ( n8799 , n8793 , n8796 );
nand ( n8800 , n8798 , n8799 );
not ( n8801 , n8800 );
or ( n8802 , n8779 , n8801 );
not ( n8803 , n8793 );
nand ( n8804 , n8803 , n8796 );
nand ( n8805 , n8802 , n8804 );
not ( n8806 , n8805 );
xor ( n8807 , n8734 , n8738 );
xnor ( n8808 , n8807 , n8681 );
not ( n8809 , n8639 );
not ( n8810 , n8644 );
not ( n8811 , n8810 );
or ( n8812 , n8809 , n8811 );
not ( n8813 , n8639 );
not ( n8814 , n8810 );
nand ( n8815 , n8813 , n8814 );
nand ( n8816 , n8812 , n8815 );
not ( n8817 , n8816 );
and ( n8818 , n8808 , n8817 );
not ( n8819 , n8808 );
and ( n8820 , n8819 , n8816 );
nor ( n8821 , n8818 , n8820 );
not ( n8822 , n8821 );
or ( n8823 , n8806 , n8822 );
not ( n8824 , n8808 );
nand ( n8825 , n8816 , n8824 );
nand ( n8826 , n8823 , n8825 );
nand ( n8827 , n8745 , n8826 );
not ( n8828 , n8677 );
not ( n8829 , n8828 );
not ( n8830 , n8741 );
and ( n8831 , n8829 , n8830 );
and ( n8832 , n8828 , n8741 );
nor ( n8833 , n8831 , n8832 );
or ( n8834 , n8744 , n8833 );
not ( n8835 , n8828 );
nand ( n8836 , n8835 , n8741 );
nand ( n8837 , n8834 , n8836 );
not ( n8838 , n8604 );
not ( n8839 , n8838 );
not ( n8840 , n8668 );
or ( n8841 , n8839 , n8840 );
or ( n8842 , n8605 , n8668 );
nand ( n8843 , n8841 , n8842 );
nor ( n8844 , n8837 , n8843 );
or ( n8845 , n8827 , n8844 );
nand ( n8846 , n8837 , n8843 );
nand ( n8847 , n8845 , n8846 );
not ( n8848 , n8847 );
or ( n8849 , n8676 , n8848 );
not ( n8850 , n8674 );
not ( n8851 , n8599 );
nand ( n8852 , n8850 , n8851 );
nand ( n8853 , n8849 , n8852 );
not ( n8854 , n8265 );
nand ( n8855 , n8854 , n8363 );
not ( n8856 , n8855 );
nor ( n8857 , n8266 , n8363 );
nor ( n8858 , n8856 , n8857 );
not ( n8859 , n8597 );
not ( n8860 , n8859 );
not ( n8861 , n8594 );
or ( n8862 , n8860 , n8861 );
nand ( n8863 , n8506 , n8589 );
nand ( n8864 , n8862 , n8863 );
not ( n8865 , n8864 );
nand ( n8866 , n8858 , n8865 );
nand ( n8867 , n8853 , n8866 );
not ( n8868 , n8675 );
not ( n8869 , n8745 );
not ( n8870 , n8826 );
nand ( n8871 , n8869 , n8870 );
not ( n8872 , n8844 );
nand ( n8873 , n8871 , n8872 );
nor ( n8874 , n8868 , n8873 );
not ( n8875 , n8800 );
not ( n8876 , n8777 );
and ( n8877 , n8875 , n8876 );
and ( n8878 , n8800 , n8777 );
nor ( n8879 , n8877 , n8878 );
not ( n8880 , n8879 );
not ( n8881 , n8880 );
not ( n8882 , n8689 );
xor ( n8883 , n8882 , n8709 );
not ( n8884 , n8883 );
not ( n8885 , n8763 );
not ( n8886 , n4248 );
or ( n8887 , n8885 , n8886 );
xor ( n8888 , n44 , n66 );
nand ( n8889 , n8888 , n7105 );
nand ( n8890 , n8887 , n8889 );
not ( n8891 , n8890 );
nand ( n8892 , n67 , n3348 );
not ( n8893 , n8892 );
not ( n8894 , n8893 );
not ( n8895 , n6196 );
xor ( n8896 , n50 , n60 );
not ( n8897 , n8896 );
or ( n8898 , n8895 , n8897 );
nand ( n8899 , n51 , n8754 );
nand ( n8900 , n8898 , n8899 );
not ( n8901 , n8900 );
not ( n8902 , n8901 );
or ( n8903 , n8894 , n8902 );
not ( n8904 , n8892 );
not ( n8905 , n8900 );
or ( n8906 , n8904 , n8905 );
nand ( n8907 , n8903 , n8906 );
not ( n8908 , n8907 );
or ( n8909 , n8891 , n8908 );
not ( n8910 , n8901 );
nand ( n8911 , n8904 , n8910 );
nand ( n8912 , n8909 , n8911 );
not ( n8913 , n8912 );
xnor ( n8914 , n46 , n63 );
or ( n8915 , n8914 , n7189 );
nand ( n8916 , n8687 , n7187 );
nand ( n8917 , n8915 , n8916 );
not ( n8918 , n8917 );
not ( n8919 , n8785 );
not ( n8920 , n8792 );
and ( n8921 , n8919 , n8920 );
and ( n8922 , n8785 , n8792 );
nor ( n8923 , n8921 , n8922 );
not ( n8924 , n8923 );
or ( n8925 , n8918 , n8924 );
or ( n8926 , n8917 , n8923 );
nand ( n8927 , n8925 , n8926 );
not ( n8928 , n8927 );
or ( n8929 , n8913 , n8928 );
not ( n8930 , n8923 );
nand ( n8931 , n8917 , n8930 );
nand ( n8932 , n8929 , n8931 );
not ( n8933 , n8932 );
or ( n8934 , n8884 , n8933 );
or ( n8935 , n8883 , n8932 );
nand ( n8936 , n8934 , n8935 );
not ( n8937 , n8936 );
or ( n8938 , n8881 , n8937 );
not ( n8939 , n8883 );
nand ( n8940 , n8939 , n8932 );
nand ( n8941 , n8938 , n8940 );
not ( n8942 , n8941 );
xor ( n8943 , n8816 , n8808 );
xnor ( n8944 , n8943 , n8805 );
not ( n8945 , n8944 );
nand ( n8946 , n8942 , n8945 );
not ( n8947 , n8946 );
not ( n8948 , n6196 );
xor ( n8949 , n50 , n61 );
not ( n8950 , n8949 );
or ( n8951 , n8948 , n8950 );
nand ( n8952 , n51 , n8896 );
nand ( n8953 , n8951 , n8952 );
not ( n8954 , n44 );
not ( n8955 , n8954 );
nand ( n8956 , n45 , n46 );
or ( n8957 , n45 , n46 );
nand ( n8958 , n8957 , n67 );
nand ( n8959 , n8955 , n8956 , n8958 );
not ( n8960 , n8959 );
nand ( n8961 , n8953 , n8960 );
not ( n8962 , n8961 );
xor ( n8963 , n48 , n62 );
not ( n8964 , n8963 );
not ( n8965 , n7312 );
or ( n8966 , n8964 , n8965 );
nand ( n8967 , n8168 , n8787 );
nand ( n8968 , n8966 , n8967 );
not ( n8969 , n8968 );
or ( n8970 , n8962 , n8969 );
or ( n8971 , n8961 , n8968 );
nand ( n8972 , n8970 , n8971 );
not ( n8973 , n46 );
not ( n8974 , n64 );
and ( n8975 , n8973 , n8974 );
and ( n8976 , n46 , n64 );
nor ( n8977 , n8975 , n8976 );
not ( n8978 , n8977 );
not ( n8979 , n7075 );
or ( n8980 , n8978 , n8979 );
or ( n8981 , n8914 , n7081 );
nand ( n8982 , n8980 , n8981 );
and ( n8983 , n8972 , n8982 );
not ( n8984 , n8972 );
not ( n8985 , n8982 );
and ( n8986 , n8984 , n8985 );
nor ( n8987 , n8983 , n8986 );
not ( n8988 , n8987 );
xor ( n8989 , n48 , n63 );
not ( n8990 , n8989 );
not ( n8991 , n8526 );
or ( n8992 , n8990 , n8991 );
nand ( n8993 , n8168 , n8963 );
nand ( n8994 , n8992 , n8993 );
not ( n8995 , n8994 );
xor ( n8996 , n46 , n65 );
not ( n8997 , n8996 );
not ( n8998 , n7074 );
or ( n8999 , n8997 , n8998 );
not ( n9000 , n8977 );
or ( n9001 , n7080 , n9000 );
nand ( n9002 , n8999 , n9001 );
not ( n9003 , n9002 );
or ( n9004 , n8995 , n9003 );
not ( n9005 , n8888 );
not ( n9006 , n3467 );
or ( n9007 , n9005 , n9006 );
not ( n9008 , n6918 );
or ( n9009 , n44 , n67 );
nand ( n9010 , n44 , n67 );
nand ( n9011 , n9008 , n9009 , n9010 );
nand ( n9012 , n9007 , n9011 );
not ( n9013 , n8994 );
not ( n9014 , n9002 );
and ( n9015 , n9013 , n9014 );
not ( n9016 , n9013 );
and ( n9017 , n9016 , n9002 );
nor ( n9018 , n9015 , n9017 );
nand ( n9019 , n9012 , n9018 );
nand ( n9020 , n9004 , n9019 );
not ( n9021 , n8890 );
and ( n9022 , n8907 , n9021 );
not ( n9023 , n8907 );
and ( n9024 , n9023 , n8890 );
nor ( n9025 , n9022 , n9024 );
not ( n9026 , n9025 );
and ( n9027 , n9020 , n9026 );
not ( n9028 , n9020 );
and ( n9029 , n9028 , n9025 );
nor ( n9030 , n9027 , n9029 );
not ( n9031 , n9030 );
or ( n9032 , n8988 , n9031 );
not ( n9033 , n9020 );
not ( n9034 , n9033 );
nand ( n9035 , n9026 , n9034 );
nand ( n9036 , n9032 , n9035 );
not ( n9037 , n9036 );
and ( n9038 , n8927 , n8912 );
not ( n9039 , n8927 );
not ( n9040 , n8912 );
and ( n9041 , n9039 , n9040 );
nor ( n9042 , n9038 , n9041 );
not ( n9043 , n8982 );
not ( n9044 , n8972 );
or ( n9045 , n9043 , n9044 );
not ( n9046 , n8961 );
nand ( n9047 , n9046 , n8968 );
nand ( n9048 , n9045 , n9047 );
not ( n9049 , n9048 );
not ( n9050 , n9049 );
not ( n9051 , n8771 );
and ( n9052 , n8751 , n9051 );
not ( n9053 , n8751 );
and ( n9054 , n9053 , n8771 );
nor ( n9055 , n9052 , n9054 );
not ( n9056 , n9055 );
not ( n9057 , n9056 );
or ( n9058 , n9050 , n9057 );
nand ( n9059 , n9048 , n9055 );
nand ( n9060 , n9058 , n9059 );
xnor ( n9061 , n9042 , n9060 );
nor ( n9062 , n9037 , n9061 );
xor ( n9063 , n9012 , n9018 );
not ( n9064 , n9063 );
and ( n9065 , n8953 , n8959 );
not ( n9066 , n8953 );
and ( n9067 , n9066 , n8960 );
nor ( n9068 , n9065 , n9067 );
not ( n9069 , n9068 );
xor ( n9070 , n48 , n64 );
not ( n9071 , n9070 );
not ( n9072 , n7314 );
or ( n9073 , n9071 , n9072 );
nand ( n9074 , n7319 , n8989 );
nand ( n9075 , n9073 , n9074 );
not ( n9076 , n9075 );
and ( n9077 , n67 , n4247 );
not ( n9078 , n4031 );
not ( n9079 , n9078 );
xor ( n9080 , n50 , n62 );
not ( n9081 , n9080 );
or ( n9082 , n9079 , n9081 );
nand ( n9083 , n51 , n8949 );
nand ( n9084 , n9082 , n9083 );
and ( n9085 , n9077 , n9084 );
not ( n9086 , n9077 );
not ( n9087 , n9084 );
and ( n9088 , n9086 , n9087 );
nor ( n9089 , n9085 , n9088 );
not ( n9090 , n9089 );
or ( n9091 , n9076 , n9090 );
not ( n9092 , n9087 );
nand ( n9093 , n9077 , n9092 );
nand ( n9094 , n9091 , n9093 );
not ( n9095 , n9094 );
or ( n9096 , n9069 , n9095 );
or ( n9097 , n9068 , n9094 );
nand ( n9098 , n9096 , n9097 );
not ( n9099 , n9098 );
or ( n9100 , n9064 , n9099 );
not ( n9101 , n9068 );
nand ( n9102 , n9101 , n9094 );
nand ( n9103 , n9100 , n9102 );
not ( n9104 , n9103 );
xor ( n9105 , n9025 , n9033 );
xnor ( n9106 , n9105 , n8987 );
nor ( n9107 , n9104 , n9106 );
or ( n9108 , n9062 , n9107 );
nand ( n9109 , n9037 , n9061 );
nand ( n9110 , n9108 , n9109 );
not ( n9111 , n9110 );
not ( n9112 , n8879 );
not ( n9113 , n8936 );
and ( n9114 , n9112 , n9113 );
and ( n9115 , n8879 , n8936 );
nor ( n9116 , n9114 , n9115 );
not ( n9117 , n9042 );
not ( n9118 , n9060 );
or ( n9119 , n9117 , n9118 );
nand ( n9120 , n9048 , n9056 );
nand ( n9121 , n9119 , n9120 );
not ( n9122 , n9121 );
nand ( n9123 , n9116 , n9122 );
nand ( n9124 , n9111 , n9123 );
not ( n9125 , n9122 );
not ( n9126 , n9116 );
nand ( n9127 , n9125 , n9126 );
not ( n9128 , n8942 );
nand ( n9129 , n9128 , n8944 );
nand ( n9130 , n9124 , n9127 , n9129 );
not ( n9131 , n9130 );
or ( n9132 , n8947 , n9131 );
nand ( n9133 , n47 , n48 );
or ( n9134 , n47 , n48 );
nand ( n9135 , n9134 , n67 );
nand ( n9136 , n9133 , n46 , n9135 );
not ( n9137 , n9136 );
not ( n9138 , n6264 );
xor ( n9139 , n50 , n63 );
not ( n9140 , n9139 );
or ( n9141 , n9138 , n9140 );
nand ( n9142 , n51 , n9080 );
nand ( n9143 , n9141 , n9142 );
nand ( n9144 , n9137 , n9143 );
not ( n9145 , n8996 );
not ( n9146 , n7784 );
or ( n9147 , n9145 , n9146 );
xor ( n9148 , n46 , n66 );
nand ( n9149 , n9148 , n7077 );
nand ( n9150 , n9147 , n9149 );
and ( n9151 , n9144 , n9150 );
and ( n9152 , n9089 , n9075 );
not ( n9153 , n9089 );
not ( n9154 , n9075 );
and ( n9155 , n9153 , n9154 );
nor ( n9156 , n9152 , n9155 );
xor ( n9157 , n9144 , n9150 );
and ( n9158 , n9156 , n9157 );
nor ( n9159 , n9151 , n9158 );
not ( n9160 , n9063 );
and ( n9161 , n9098 , n9160 );
not ( n9162 , n9098 );
and ( n9163 , n9162 , n9063 );
nor ( n9164 , n9161 , n9163 );
nand ( n9165 , n9159 , n9164 );
not ( n9166 , n9165 );
not ( n9167 , n9136 );
not ( n9168 , n9143 );
or ( n9169 , n9167 , n9168 );
or ( n9170 , n9136 , n9143 );
nand ( n9171 , n9169 , n9170 );
not ( n9172 , n9171 );
not ( n9173 , n9148 );
not ( n9174 , n7080 );
not ( n9175 , n9174 );
or ( n9176 , n9173 , n9175 );
xor ( n9177 , n46 , n67 );
nand ( n9178 , n9177 , n7074 );
nand ( n9179 , n9176 , n9178 );
xor ( n9180 , n48 , n65 );
not ( n9181 , n9180 );
not ( n9182 , n8526 );
or ( n9183 , n9181 , n9182 );
nand ( n9184 , n8168 , n9070 );
nand ( n9185 , n9183 , n9184 );
and ( n9186 , n9179 , n9185 );
not ( n9187 , n9179 );
not ( n9188 , n9185 );
and ( n9189 , n9187 , n9188 );
nor ( n9190 , n9186 , n9189 );
not ( n9191 , n9190 );
or ( n9192 , n9172 , n9191 );
not ( n9193 , n9188 );
nand ( n9194 , n9193 , n9179 );
nand ( n9195 , n9192 , n9194 );
not ( n9196 , n9195 );
xor ( n9197 , n9156 , n9157 );
nand ( n9198 , n9196 , n9197 );
not ( n9199 , n9198 );
not ( n9200 , n6236 );
nand ( n9201 , n8746 , n6231 );
not ( n9202 , n9201 );
or ( n9203 , n9200 , n9202 );
nand ( n9204 , n9203 , n48 );
not ( n9205 , n9204 );
not ( n9206 , n4031 );
not ( n9207 , n9206 );
xor ( n9208 , n50 , n65 );
not ( n9209 , n9208 );
or ( n9210 , n9207 , n9209 );
xor ( n9211 , n50 , n64 );
nand ( n9212 , n51 , n9211 );
nand ( n9213 , n9210 , n9212 );
and ( n9214 , n9205 , n9213 );
xor ( n9215 , n48 , n66 );
not ( n9216 , n9215 );
not ( n9217 , n7314 );
or ( n9218 , n9216 , n9217 );
nand ( n9219 , n7319 , n9180 );
nand ( n9220 , n9218 , n9219 );
not ( n9221 , n9220 );
not ( n9222 , n9221 );
nand ( n9223 , n67 , n9174 );
not ( n9224 , n9223 );
not ( n9225 , n5655 );
not ( n9226 , n9211 );
or ( n9227 , n9225 , n9226 );
nand ( n9228 , n51 , n9139 );
nand ( n9229 , n9227 , n9228 );
not ( n9230 , n9229 );
and ( n9231 , n9224 , n9230 );
and ( n9232 , n9223 , n9229 );
nor ( n9233 , n9231 , n9232 );
not ( n9234 , n9233 );
not ( n9235 , n9234 );
or ( n9236 , n9222 , n9235 );
nand ( n9237 , n9220 , n9233 );
nand ( n9238 , n9236 , n9237 );
nor ( n9239 , n9214 , n9238 );
nand ( n9240 , n50 , n67 );
and ( n9241 , n67 , n7318 );
not ( n9242 , n4888 );
xor ( n9243 , n50 , n66 );
not ( n9244 , n9243 );
or ( n9245 , n9242 , n9244 );
nand ( n9246 , n51 , n9208 );
nand ( n9247 , n9245 , n9246 );
or ( n9248 , n9241 , n9247 );
not ( n9249 , n9243 );
nand ( n9250 , n6277 , n9249 );
nand ( n9251 , n9248 , n9250 );
or ( n9252 , n9240 , n9251 );
nand ( n9253 , n9241 , n9247 );
nand ( n9254 , n9252 , n9253 );
not ( n9255 , n9254 );
xor ( n9256 , n9205 , n9213 );
not ( n9257 , n8746 );
not ( n9258 , n7314 );
or ( n9259 , n9257 , n9258 );
nand ( n9260 , n7319 , n9215 );
nand ( n9261 , n9259 , n9260 );
nor ( n9262 , n9256 , n9261 );
or ( n9263 , n9255 , n9262 );
nand ( n9264 , n9261 , n9256 );
nand ( n9265 , n9263 , n9264 );
not ( n9266 , n9265 );
or ( n9267 , n9239 , n9266 );
nand ( n9268 , n9214 , n9238 );
nand ( n9269 , n9267 , n9268 );
not ( n9270 , n9269 );
not ( n9271 , n9220 );
not ( n9272 , n9234 );
or ( n9273 , n9271 , n9272 );
not ( n9274 , n9223 );
nand ( n9275 , n9274 , n9229 );
nand ( n9276 , n9273 , n9275 );
not ( n9277 , n9276 );
not ( n9278 , n9277 );
not ( n9279 , n9171 );
not ( n9280 , n9190 );
not ( n9281 , n9280 );
or ( n9282 , n9279 , n9281 );
not ( n9283 , n9171 );
nand ( n9284 , n9283 , n9190 );
nand ( n9285 , n9282 , n9284 );
not ( n9286 , n9285 );
or ( n9287 , n9278 , n9286 );
or ( n9288 , n9277 , n9285 );
nand ( n9289 , n9287 , n9288 );
not ( n9290 , n9289 );
or ( n9291 , n9270 , n9290 );
not ( n9292 , n9277 );
nand ( n9293 , n9292 , n9285 );
nand ( n9294 , n9291 , n9293 );
not ( n9295 , n9294 );
or ( n9296 , n9199 , n9295 );
not ( n9297 , n9196 );
not ( n9298 , n9197 );
nand ( n9299 , n9297 , n9298 );
nand ( n9300 , n9296 , n9299 );
not ( n9301 , n9300 );
or ( n9302 , n9166 , n9301 );
not ( n9303 , n9159 );
not ( n9304 , n9164 );
nand ( n9305 , n9303 , n9304 );
nand ( n9306 , n9302 , n9305 );
nand ( n9307 , n9306 , n9123 );
not ( n9308 , n9307 );
nand ( n9309 , n9104 , n9106 );
and ( n9310 , n9309 , n9109 );
nand ( n9311 , n9308 , n9310 , n8946 );
nand ( n9312 , n9132 , n9311 );
nand ( n9313 , n8874 , n8866 , n9312 );
not ( n9314 , n8858 );
not ( n9315 , n8865 );
nand ( n9316 , n9314 , n9315 );
nand ( n9317 , n8867 , n9313 , n9316 );
not ( n9318 , n9317 );
not ( n9319 , n9318 );
and ( n9320 , n8455 , n7580 , n8468 );
nand ( n9321 , n8497 , n8013 , n9319 , n9320 );
nand ( n9322 , n8472 , n8490 , n9321 );
nor ( n9323 , n7057 , n7265 );
nor ( n9324 , n7277 , n9323 );
and ( n9325 , n6962 , n9324 );
nand ( n9326 , n9322 , n9325 );
not ( n9327 , n9326 );
nand ( n9328 , n9327 , n6755 , n6831 );
nand ( n9329 , n7293 , n7294 , n9328 );
and ( n9330 , n6680 , n6672 );
and ( n9331 , n6671 , n6670 );
nor ( n9332 , n9330 , n9331 );
xnor ( n9333 , n6680 , n9332 );
or ( n9334 , n6668 , n6599 );
or ( n9335 , n36 , n52 );
nand ( n9336 , n36 , n52 );
nand ( n9337 , n9335 , n9336 );
or ( n9338 , n3149 , n9337 );
nand ( n9339 , n9334 , n9338 );
or ( n9340 , n3210 , n6641 );
nand ( n9341 , n9340 , n38 );
not ( n9342 , n6603 );
xor ( n9343 , n9341 , n9342 );
xnor ( n9344 , n9339 , n9343 );
xor ( n9345 , n9333 , n9344 );
or ( n9346 , n6664 , n6698 );
or ( n9347 , n6697 , n6681 );
nand ( n9348 , n9346 , n9347 );
nand ( n9349 , n9345 , n9348 );
not ( n9350 , n9345 );
not ( n9351 , n9348 );
nand ( n9352 , n9350 , n9351 );
and ( n9353 , n9349 , n9352 );
xnor ( n9354 , n9329 , n9353 );
or ( n9355 , n9354 , n2 );
nand ( n9356 , n6585 , n9355 );
not ( n9357 , n9356 );
or ( n9358 , n3203 , n3215 );
or ( n9359 , n3208 , n3214 );
nand ( n9360 , n9358 , n9359 );
not ( n9361 , n3188 );
not ( n9362 , n3201 );
or ( n9363 , n9361 , n9362 );
nand ( n9364 , n36 , n3191 );
nand ( n9365 , n9363 , n9364 );
and ( n9366 , n9365 , n3162 );
not ( n9367 , n9365 );
not ( n9368 , n3162 );
and ( n9369 , n9367 , n9368 );
nor ( n9370 , n9366 , n9369 );
xor ( n9371 , n9360 , n9370 );
or ( n9372 , n3216 , n3187 );
or ( n9373 , n3182 , n3184 );
nand ( n9374 , n9372 , n9373 );
nand ( n9375 , n9371 , n9374 );
not ( n9376 , n9371 );
not ( n9377 , n9374 );
nand ( n9378 , n9376 , n9377 );
and ( n9379 , n9375 , n9378 );
not ( n9380 , n9379 );
not ( n9381 , n3336 );
not ( n9382 , n6579 );
or ( n9383 , n9381 , n9382 );
nand ( n9384 , n9383 , n3333 );
not ( n9385 , n9384 );
or ( n9386 , n9380 , n9385 );
nand ( n9387 , n9386 , n2 );
nor ( n9388 , n9379 , n9384 );
or ( n9389 , n9387 , n9388 );
or ( n9390 , n9337 , n6599 );
nand ( n9391 , n9390 , n9364 );
xor ( n9392 , n9391 , n6667 );
not ( n9393 , n9392 );
and ( n9394 , n9339 , n9343 );
and ( n9395 , n9342 , n9341 );
nor ( n9396 , n9394 , n9395 );
not ( n9397 , n9396 );
or ( n9398 , n9393 , n9397 );
or ( n9399 , n9392 , n9396 );
nand ( n9400 , n9398 , n9399 );
or ( n9401 , n9344 , n9333 );
or ( n9402 , n6680 , n9332 );
nand ( n9403 , n9401 , n9402 );
nand ( n9404 , n9400 , n9403 );
not ( n9405 , n9400 );
not ( n9406 , n9403 );
nand ( n9407 , n9405 , n9406 );
and ( n9408 , n9404 , n9407 );
not ( n9409 , n9352 );
not ( n9410 , n9329 );
or ( n9411 , n9409 , n9410 );
nand ( n9412 , n9411 , n9349 );
xor ( n9413 , n9408 , n9412 );
not ( n9414 , n2 );
nand ( n9415 , n9413 , n9414 );
nand ( n9416 , n9389 , n9415 );
nand ( n9417 , n9357 , n9416 );
not ( n9418 , n9417 );
not ( n9419 , n2 );
not ( n9420 , n6466 );
nand ( n9421 , n4817 , n5356 , n5360 );
not ( n9422 , n5364 );
nand ( n9423 , n4766 , n6377 , n9421 , n9422 );
nand ( n9424 , n6559 , n9423 );
not ( n9425 , n9424 );
not ( n9426 , n9425 );
or ( n9427 , n9420 , n9426 );
not ( n9428 , n6577 );
nand ( n9429 , n9427 , n9428 );
not ( n9430 , n3405 );
nand ( n9431 , n9430 , n6381 );
not ( n9432 , n9431 );
and ( n9433 , n9429 , n9432 );
not ( n9434 , n9429 );
and ( n9435 , n9434 , n9431 );
nor ( n9436 , n9433 , n9435 );
not ( n9437 , n9436 );
or ( n9438 , n9419 , n9437 );
and ( n9439 , n7294 , n6755 );
not ( n9440 , n9439 );
not ( n9441 , n9326 );
nand ( n9442 , n9441 , n6831 );
not ( n9443 , n7292 );
nand ( n9444 , n9440 , n9442 , n9443 );
not ( n9445 , n9439 );
nand ( n9446 , n9442 , n9443 );
not ( n9447 , n9446 );
or ( n9448 , n9445 , n9447 );
nand ( n9449 , n9448 , n9414 );
not ( n9450 , n9449 );
nand ( n9451 , n9444 , n9450 );
nand ( n9452 , n9438 , n9451 );
not ( n9453 , n9452 );
nand ( n9454 , n9453 , n9356 );
not ( n9455 , n9454 );
nor ( n9456 , n9418 , n9455 );
not ( n9457 , n9456 );
not ( n9458 , n9457 );
buf ( n9459 , n9416 );
not ( n9460 , n9459 );
not ( n9461 , n9378 );
not ( n9462 , n9384 );
or ( n9463 , n9461 , n9462 );
nand ( n9464 , n9463 , n9375 );
not ( n9465 , n9464 );
not ( n9466 , n3191 );
not ( n9467 , n3188 );
and ( n9468 , n9466 , n9467 );
nor ( n9469 , n9468 , n3126 );
not ( n9470 , n9469 );
not ( n9471 , n3200 );
and ( n9472 , n9471 , n9368 );
and ( n9473 , n3162 , n3200 );
nor ( n9474 , n9472 , n9473 );
not ( n9475 , n9474 );
and ( n9476 , n9470 , n9475 );
and ( n9477 , n9469 , n9474 );
nor ( n9478 , n9476 , n9477 );
not ( n9479 , n9478 );
and ( n9480 , n9370 , n9360 );
and ( n9481 , n3162 , n9365 );
nor ( n9482 , n9480 , n9481 );
not ( n9483 , n9482 );
or ( n9484 , n9479 , n9483 );
or ( n9485 , n9478 , n9482 );
nand ( n9486 , n9484 , n9485 );
nand ( n9487 , n9465 , n2 , n9486 );
not ( n9488 , n9486 );
nand ( n9489 , n2 , n9488 , n9464 );
not ( n9490 , n6667 );
not ( n9491 , n9336 );
not ( n9492 , n6599 );
or ( n9493 , n3191 , n9492 );
nand ( n9494 , n9493 , n36 );
not ( n9495 , n9494 );
or ( n9496 , n9491 , n9495 );
or ( n9497 , n9336 , n9494 );
nand ( n9498 , n9496 , n9497 );
not ( n9499 , n9498 );
or ( n9500 , n9490 , n9499 );
or ( n9501 , n6667 , n9498 );
nand ( n9502 , n9500 , n9501 );
not ( n9503 , n9502 );
not ( n9504 , n9396 );
and ( n9505 , n9392 , n9504 );
and ( n9506 , n6667 , n9391 );
nor ( n9507 , n9505 , n9506 );
not ( n9508 , n9507 );
or ( n9509 , n9503 , n9508 );
or ( n9510 , n9502 , n9507 );
nand ( n9511 , n9509 , n9510 );
not ( n9512 , n9407 );
not ( n9513 , n9412 );
or ( n9514 , n9512 , n9513 );
nand ( n9515 , n9514 , n9404 );
nor ( n9516 , n9511 , n9515 );
not ( n9517 , n9516 );
nand ( n9518 , n9511 , n9515 );
nand ( n9519 , n9517 , n9518 , n9414 );
nand ( n9520 , n9487 , n9489 , n9519 );
nand ( n9521 , n9460 , n9520 );
not ( n9522 , n6565 );
nand ( n9523 , n6378 , n6557 );
nand ( n9524 , n9522 , n9523 );
not ( n9525 , n9524 );
and ( n9526 , n6564 , n6547 );
nor ( n9527 , n9414 , n9526 );
not ( n9528 , n9527 );
or ( n9529 , n9525 , n9528 );
not ( n9530 , n9323 );
not ( n9531 , n9530 );
not ( n9532 , n8471 );
nand ( n9533 , n9532 , n8490 , n9321 );
not ( n9534 , n9533 );
or ( n9535 , n9531 , n9534 );
nand ( n9536 , n9535 , n7266 );
not ( n9537 , n7279 );
nor ( n9538 , n9537 , n7277 );
nor ( n9539 , n2 , n9538 );
nand ( n9540 , n9536 , n9539 );
nand ( n9541 , n9529 , n9540 );
not ( n9542 , n9541 );
not ( n9543 , n9523 );
not ( n9544 , n9543 );
nand ( n9545 , n2 , n9526 , n9522 , n9544 );
not ( n9546 , n9536 );
nand ( n9547 , n9546 , n9414 , n9538 );
nand ( n9548 , n9542 , n9545 , n9547 );
not ( n9549 , n9548 );
not ( n9550 , n9414 );
nand ( n9551 , n7266 , n9530 );
not ( n9552 , n9551 );
and ( n9553 , n9533 , n9552 );
not ( n9554 , n9533 );
and ( n9555 , n9554 , n9551 );
nor ( n9556 , n9553 , n9555 );
not ( n9557 , n9556 );
or ( n9558 , n9550 , n9557 );
nand ( n9559 , n9522 , n6557 );
not ( n9560 , n9559 );
nand ( n9561 , n9560 , n9423 );
not ( n9562 , n9423 );
nand ( n9563 , n9559 , n9562 );
nand ( n9564 , n9561 , n2 , n9563 );
nand ( n9565 , n9558 , n9564 );
nor ( n9566 , n9549 , n9565 );
not ( n9567 , n9566 );
not ( n9568 , n9542 );
not ( n9569 , n9543 );
nand ( n9570 , n9569 , n2 , n9526 , n9522 );
nand ( n9571 , n9570 , n9547 );
nor ( n9572 , n9568 , n9571 );
and ( n9573 , n7284 , n6962 );
not ( n9574 , n9573 );
buf ( n9575 , n9324 );
nand ( n9576 , n9322 , n9575 );
not ( n9577 , n7280 );
nand ( n9578 , n9574 , n9576 , n9577 );
not ( n9579 , n9573 );
nand ( n9580 , n9576 , n9577 );
not ( n9581 , n9580 );
or ( n9582 , n9579 , n9581 );
nand ( n9583 , n9582 , n9414 );
not ( n9584 , n9583 );
nand ( n9585 , n9578 , n9584 );
nand ( n9586 , n6572 , n6520 );
nand ( n9587 , n9423 , n6558 );
not ( n9588 , n6567 );
nand ( n9589 , n9587 , n9588 );
nand ( n9590 , n2 , n9586 , n9589 );
not ( n9591 , n9586 );
nand ( n9592 , n9591 , n2 , n9587 , n9588 );
nand ( n9593 , n9585 , n9590 , n9592 );
nand ( n9594 , n9572 , n9593 );
nand ( n9595 , n9567 , n9594 );
not ( n9596 , n9595 );
not ( n9597 , n85 );
not ( n9598 , n8494 );
not ( n9599 , n9318 );
not ( n9600 , n9599 );
or ( n9601 , n9598 , n9600 );
nand ( n9602 , n9601 , n8406 );
not ( n9603 , n8418 );
not ( n9604 , n8422 );
nor ( n9605 , n9603 , n9604 );
buf ( n9606 , n9605 );
nor ( n9607 , n9602 , n9606 );
not ( n9608 , n9607 );
nand ( n9609 , n9606 , n9602 );
nand ( n9610 , n9608 , n9609 , n9414 );
not ( n9611 , n9610 );
not ( n9612 , n9611 );
not ( n9613 , n9414 );
not ( n9614 , n6369 );
not ( n9615 , n9614 );
not ( n9616 , n6367 );
or ( n9617 , n9615 , n9616 );
buf ( n9618 , n5342 );
nand ( n9619 , n9617 , n9618 );
nand ( n9620 , n5345 , n6371 );
nand ( n9621 , n9613 , n9619 , n9620 );
nor ( n9622 , n9619 , n9620 );
nand ( n9623 , n2 , n9622 );
nand ( n9624 , n9597 , n9612 , n9621 , n9623 );
not ( n9625 , n4981 );
not ( n9626 , n5351 );
nor ( n9627 , n9625 , n9626 );
not ( n9628 , n9627 );
not ( n9629 , n9628 );
nand ( n9630 , n5766 , n6333 , n6348 );
nand ( n9631 , n9630 , n6363 , n6366 );
not ( n9632 , n9631 );
not ( n9633 , n6372 );
not ( n9634 , n9633 );
or ( n9635 , n9632 , n9634 );
not ( n9636 , n5346 );
nand ( n9637 , n9635 , n9636 );
not ( n9638 , n9637 );
not ( n9639 , n9638 );
or ( n9640 , n9629 , n9639 );
not ( n9641 , n9627 );
not ( n9642 , n9637 );
or ( n9643 , n9641 , n9642 );
nand ( n9644 , n9643 , n2 );
not ( n9645 , n9644 );
nand ( n9646 , n9640 , n9645 );
not ( n9647 , n8146 );
nand ( n9648 , n9647 , n8149 );
not ( n9649 , n9648 );
not ( n9650 , n9317 );
not ( n9651 , n8495 );
or ( n9652 , n9650 , n9651 );
not ( n9653 , n8423 );
nand ( n9654 , n9652 , n9653 );
not ( n9655 , n9654 );
or ( n9656 , n9649 , n9655 );
or ( n9657 , n9648 , n9654 );
nand ( n9658 , n9656 , n9657 );
nand ( n9659 , n9658 , n9414 );
nand ( n9660 , n9646 , n9659 );
and ( n9661 , n84 , n9660 );
not ( n9662 , n9661 );
nand ( n9663 , n248 , n9659 , n9646 );
nand ( n9664 , n9662 , n9663 );
and ( n9665 , n9624 , n9664 );
nand ( n9666 , n9610 , n9623 , n9621 );
nand ( n9667 , n85 , n9666 );
and ( n9668 , n2 , n9619 , n9620 );
nor ( n9669 , n9611 , n9668 );
and ( n9670 , n2 , n9622 );
nor ( n9671 , n9670 , n85 );
nand ( n9672 , n9669 , n9671 );
and ( n9673 , n9667 , n9672 );
not ( n9674 , n6369 );
nand ( n9675 , n9674 , n5342 );
not ( n9676 , n9675 );
not ( n9677 , n9631 );
not ( n9678 , n9677 );
or ( n9679 , n9676 , n9678 );
nand ( n9680 , n9679 , n2 );
not ( n9681 , n6367 );
nor ( n9682 , n9681 , n9675 );
or ( n9683 , n9680 , n9682 );
not ( n9684 , n8494 );
not ( n9685 , n9684 );
and ( n9686 , n8406 , n9685 );
and ( n9687 , n9686 , n9317 );
not ( n9688 , n9687 );
not ( n9689 , n9686 );
nand ( n9690 , n9689 , n9318 );
nand ( n9691 , n9688 , n9414 , n9690 );
nand ( n9692 , n9683 , n9691 );
nor ( n9693 , n86 , n9692 );
nor ( n9694 , n9673 , n9693 );
nor ( n9695 , n9665 , n9694 );
not ( n9696 , n9695 );
nand ( n9697 , n9672 , n9667 , n9693 );
not ( n9698 , n87 );
not ( n9699 , n5542 );
not ( n9700 , n9699 );
not ( n9701 , n9700 );
not ( n9702 , n5747 );
not ( n9703 , n5765 );
nor ( n9704 , n9702 , n9703 );
not ( n9705 , n9704 );
not ( n9706 , n6333 );
or ( n9707 , n9705 , n9706 );
not ( n9708 , n6359 );
nand ( n9709 , n9707 , n9708 );
not ( n9710 , n9709 );
or ( n9711 , n9701 , n9710 );
nand ( n9712 , n9711 , n6352 );
nand ( n9713 , n6366 , n6348 );
nor ( n9714 , n9712 , n9713 );
and ( n9715 , n2 , n9714 );
not ( n9716 , n8873 );
not ( n9717 , n9716 );
not ( n9718 , n9312 );
or ( n9719 , n9717 , n9718 );
not ( n9720 , n8847 );
nand ( n9721 , n9719 , n9720 );
not ( n9722 , n9721 );
not ( n9723 , n8868 );
not ( n9724 , n9723 );
or ( n9725 , n9722 , n9724 );
not ( n9726 , n8852 );
not ( n9727 , n9726 );
nand ( n9728 , n9725 , n9727 );
nand ( n9729 , n9316 , n8866 );
and ( n9730 , n9414 , n9728 , n9729 );
nor ( n9731 , n9715 , n9730 );
not ( n9732 , n9728 );
not ( n9733 , n9729 );
and ( n9734 , n9414 , n9732 , n9733 );
not ( n9735 , n9734 );
not ( n9736 , n9414 );
buf ( n9737 , n9713 );
nand ( n9738 , n9736 , n9712 , n9737 );
nand ( n9739 , n9698 , n9731 , n9735 , n9738 );
buf ( n9740 , n9739 );
nor ( n9741 , n9692 , n86 );
not ( n9742 , n9741 );
nand ( n9743 , n86 , n9692 );
nand ( n9744 , n9742 , n9743 );
nand ( n9745 , n9740 , n9744 );
nand ( n9746 , n9712 , n2 , n9713 );
not ( n9747 , n9746 );
nor ( n9748 , n9747 , n9734 );
and ( n9749 , n9748 , n9731 );
not ( n9750 , n87 );
nor ( n9751 , n9749 , n9750 );
not ( n9752 , n9751 );
nand ( n9753 , n9752 , n9739 );
not ( n9754 , n88 );
not ( n9755 , n9699 );
nand ( n9756 , n9755 , n6352 );
not ( n9757 , n9756 );
not ( n9758 , n9709 );
or ( n9759 , n9757 , n9758 );
nand ( n9760 , n9759 , n2 );
not ( n9761 , n9721 );
not ( n9762 , n9726 );
nand ( n9763 , n9762 , n9723 );
not ( n9764 , n9763 );
or ( n9765 , n9761 , n9764 );
nand ( n9766 , n9765 , n9414 );
nand ( n9767 , n9760 , n9766 );
not ( n9768 , n9756 );
not ( n9769 , n9768 );
not ( n9770 , n9709 );
not ( n9771 , n9770 );
or ( n9772 , n9769 , n9771 );
nand ( n9773 , n9772 , n2 );
or ( n9774 , n9721 , n9763 );
nand ( n9775 , n9774 , n9414 );
nand ( n9776 , n9773 , n9775 );
nand ( n9777 , n9754 , n9767 , n9776 );
nand ( n9778 , n9753 , n9777 );
nand ( n9779 , n9745 , n9778 );
not ( n9780 , n9744 );
not ( n9781 , n9740 );
nand ( n9782 , n9780 , n9781 );
nand ( n9783 , n9697 , n9779 , n9782 );
not ( n9784 , n9783 );
or ( n9785 , n9696 , n9784 );
not ( n9786 , n9624 );
not ( n9787 , n9664 );
nand ( n9788 , n9786 , n9787 );
nand ( n9789 , n9785 , n9788 );
and ( n9790 , n9754 , n9767 , n9776 );
not ( n9791 , n9790 );
not ( n9792 , n9414 );
not ( n9793 , n8871 );
not ( n9794 , n9312 );
or ( n9795 , n9793 , n9794 );
nand ( n9796 , n9795 , n8827 );
not ( n9797 , n9796 );
not ( n9798 , n8846 );
not ( n9799 , n8872 );
nor ( n9800 , n9798 , n9799 );
nor ( n9801 , n9797 , n9800 );
not ( n9802 , n9801 );
or ( n9803 , n9792 , n9802 );
not ( n9804 , n9703 );
nand ( n9805 , n9804 , n6358 );
not ( n9806 , n5747 );
not ( n9807 , n9806 );
not ( n9808 , n9807 );
not ( n9809 , n6333 );
or ( n9810 , n9808 , n9809 );
nand ( n9811 , n9810 , n6354 );
nand ( n9812 , n9805 , n2 , n9811 );
nand ( n9813 , n9803 , n9812 );
not ( n9814 , n9813 );
nor ( n9815 , n9811 , n9805 );
and ( n9816 , n2 , n9815 );
not ( n9817 , n2 );
not ( n9818 , n9800 );
nor ( n9819 , n9796 , n9818 );
and ( n9820 , n9817 , n9819 );
nor ( n9821 , n9816 , n9820 );
not ( n9822 , n89 );
nand ( n9823 , n9814 , n9821 , n9822 );
not ( n9824 , n9823 );
not ( n9825 , n9767 );
not ( n9826 , n9776 );
or ( n9827 , n9825 , n9826 );
nand ( n9828 , n9827 , n88 );
nand ( n9829 , n9791 , n9824 , n9828 );
not ( n9830 , n91 );
not ( n9831 , n9123 );
not ( n9832 , n9831 );
not ( n9833 , n9832 );
buf ( n9834 , n9110 );
nand ( n9835 , n9306 , n9310 );
nand ( n9836 , n9834 , n9835 );
not ( n9837 , n9836 );
or ( n9838 , n9833 , n9837 );
nand ( n9839 , n9838 , n9127 );
not ( n9840 , n9129 );
not ( n9841 , n9840 );
nand ( n9842 , n9841 , n8946 );
nand ( n9843 , n9839 , n9842 , n9414 );
not ( n9844 , n9843 );
not ( n9845 , n9844 );
not ( n9846 , n5854 );
not ( n9847 , n9846 );
buf ( n9848 , n5935 );
nand ( n9849 , n9847 , n9848 );
not ( n9850 , n6080 );
nand ( n9851 , n6072 , n6070 );
nand ( n9852 , n9851 , n6330 );
not ( n9853 , n9852 );
or ( n9854 , n9850 , n9853 );
nand ( n9855 , n9854 , n5934 );
nand ( n9856 , n2 , n9849 , n9855 );
not ( n9857 , n9839 );
not ( n9858 , n9842 );
nand ( n9859 , n9857 , n9858 , n9414 );
not ( n9860 , n9855 );
not ( n9861 , n9849 );
nand ( n9862 , n9860 , n2 , n9861 );
nand ( n9863 , n9845 , n9856 , n9859 , n9862 );
not ( n9864 , n9863 );
or ( n9865 , n9830 , n9864 );
nand ( n9866 , n9856 , n9859 );
not ( n9867 , n9866 );
not ( n9868 , n91 );
nor ( n9869 , n9414 , n9849 , n9855 );
nor ( n9870 , n9869 , n9844 );
nand ( n9871 , n9867 , n9868 , n9870 );
nand ( n9872 , n9865 , n9871 );
not ( n9873 , n6079 );
nand ( n9874 , n9873 , n5934 );
not ( n9875 , n9874 );
not ( n9876 , n9852 );
and ( n9877 , n9875 , n9876 );
and ( n9878 , n9874 , n9852 );
nor ( n9879 , n9877 , n9878 );
nor ( n9880 , n9879 , n9414 );
not ( n9881 , n9127 );
nor ( n9882 , n9881 , n9831 );
not ( n9883 , n9882 );
not ( n9884 , n9836 );
or ( n9885 , n9883 , n9884 );
nand ( n9886 , n9885 , n9414 );
nor ( n9887 , n9836 , n9882 );
nor ( n9888 , n9886 , n9887 );
nor ( n9889 , n9880 , n9888 );
not ( n9890 , n92 );
nand ( n9891 , n9889 , n9890 );
nand ( n9892 , n9872 , n9891 );
not ( n9893 , n9414 );
and ( n9894 , n8871 , n8827 );
xor ( n9895 , n9894 , n9312 );
not ( n9896 , n9895 );
or ( n9897 , n9893 , n9896 );
not ( n9898 , n6354 );
nor ( n9899 , n9898 , n9806 );
nor ( n9900 , n6333 , n9899 );
not ( n9901 , n9900 );
nand ( n9902 , n6333 , n9899 );
nand ( n9903 , n9901 , n2 , n9902 );
nand ( n9904 , n9897 , n9903 );
not ( n9905 , n9904 );
not ( n9906 , n90 );
nand ( n9907 , n9905 , n9906 );
not ( n9908 , n9907 );
buf ( n9909 , n9871 );
nand ( n9910 , n90 , n9904 );
not ( n9911 , n9910 );
nor ( n9912 , n9908 , n9909 , n9911 );
or ( n9913 , n9892 , n9912 );
nor ( n9914 , n90 , n9904 );
not ( n9915 , n9914 );
nand ( n9916 , n9915 , n9910 );
nand ( n9917 , n9909 , n9916 );
nand ( n9918 , n9913 , n9917 );
not ( n9919 , n9813 );
and ( n9920 , n9821 , n9919 );
nor ( n9921 , n9920 , n9822 );
not ( n9922 , n9921 );
not ( n9923 , n9907 );
nand ( n9924 , n9922 , n9923 , n9823 );
nand ( n9925 , n9829 , n9918 , n9924 );
not ( n9926 , n9921 );
nand ( n9927 , n9926 , n9823 );
and ( n9928 , n9927 , n9907 );
nand ( n9929 , n9824 , n9828 , n9777 );
nand ( n9930 , n9928 , n9929 );
not ( n9931 , n9828 );
not ( n9932 , n9777 );
or ( n9933 , n9931 , n9932 );
not ( n9934 , n9824 );
nand ( n9935 , n9933 , n9934 );
nand ( n9936 , n9925 , n9930 , n9935 );
not ( n9937 , n9936 );
not ( n9938 , n2 );
not ( n9939 , n6068 );
not ( n9940 , n6328 );
nand ( n9941 , n9939 , n9940 );
not ( n9942 , n9941 );
not ( n9943 , n6326 );
or ( n9944 , n9942 , n9943 );
or ( n9945 , n9941 , n6326 );
nand ( n9946 , n9944 , n9945 );
not ( n9947 , n9946 );
or ( n9948 , n9938 , n9947 );
not ( n9949 , n9309 );
nor ( n9950 , n9104 , n9106 );
nor ( n9951 , n9949 , n9950 );
not ( n9952 , n9951 );
not ( n9953 , n9952 );
not ( n9954 , n9306 );
not ( n9955 , n9954 );
or ( n9956 , n9953 , n9955 );
not ( n9957 , n9951 );
not ( n9958 , n9306 );
or ( n9959 , n9957 , n9958 );
nand ( n9960 , n9959 , n9414 );
not ( n9961 , n9960 );
nand ( n9962 , n9956 , n9961 );
nand ( n9963 , n9948 , n9962 );
nor ( n9964 , n94 , n9963 );
not ( n9965 , n9964 );
nand ( n9966 , n94 , n9963 );
nand ( n9967 , n9965 , n9966 );
not ( n9968 , n9414 );
nand ( n9969 , n9305 , n9165 );
not ( n9970 , n9969 );
not ( n9971 , n9300 );
or ( n9972 , n9970 , n9971 );
or ( n9973 , n9969 , n9300 );
nand ( n9974 , n9972 , n9973 );
not ( n9975 , n9974 );
or ( n9976 , n9968 , n9975 );
not ( n9977 , n6320 );
not ( n9978 , n6325 );
not ( n9979 , n9978 );
nand ( n9980 , n9979 , n6135 );
nor ( n9981 , n9977 , n9980 );
not ( n9982 , n9981 );
nand ( n9983 , n9977 , n9980 );
nand ( n9984 , n9982 , n9983 , n2 );
nand ( n9985 , n9976 , n9984 );
and ( n9986 , n9967 , n9985 );
not ( n9987 , n95 );
nor ( n9988 , n9985 , n9987 );
nand ( n9989 , n9967 , n9988 );
not ( n9990 , n9989 );
nor ( n9991 , n9986 , n9990 );
not ( n9992 , n9991 );
not ( n9993 , n93 );
not ( n9994 , n6072 );
not ( n9995 , n6000 );
not ( n9996 , n5994 );
nor ( n9997 , n9995 , n9996 );
nor ( n9998 , n9994 , n9997 );
not ( n9999 , n9940 );
not ( n10000 , n6326 );
or ( n10001 , n9999 , n10000 );
nand ( n10002 , n10001 , n6069 );
nor ( n10003 , n9998 , n10002 );
not ( n10004 , n9998 );
not ( n10005 , n10002 );
or ( n10006 , n10004 , n10005 );
nand ( n10007 , n10006 , n2 );
or ( n10008 , n10003 , n10007 );
not ( n10009 , n9062 );
and ( n10010 , n10009 , n9109 );
not ( n10011 , n9309 );
not ( n10012 , n9306 );
or ( n10013 , n10011 , n10012 );
not ( n10014 , n9950 );
nand ( n10015 , n10013 , n10014 );
xor ( n10016 , n10010 , n10015 );
nand ( n10017 , n10016 , n9414 );
nand ( n10018 , n10008 , n10017 );
not ( n10019 , n10018 );
and ( n10020 , n9993 , n10019 );
not ( n10021 , n9880 );
not ( n10022 , n9888 );
and ( n10023 , n10021 , n10022 );
nor ( n10024 , n10023 , n9890 );
not ( n10025 , n10024 );
nand ( n10026 , n10025 , n9891 );
not ( n10027 , n10026 );
nand ( n10028 , n10020 , n10027 );
xor ( n10029 , n9993 , n10019 );
not ( n10030 , n9964 );
not ( n10031 , n10030 );
nand ( n10032 , n10029 , n10031 );
nand ( n10033 , n9992 , n10028 , n10032 );
not ( n10034 , n96 );
not ( n10035 , n9414 );
nand ( n10036 , n9299 , n9198 );
not ( n10037 , n10036 );
not ( n10038 , n9294 );
or ( n10039 , n10037 , n10038 );
or ( n10040 , n10036 , n9294 );
nand ( n10041 , n10039 , n10040 );
not ( n10042 , n10041 );
or ( n10043 , n10035 , n10042 );
not ( n10044 , n6314 );
nand ( n10045 , n6319 , n6183 );
nor ( n10046 , n10044 , n10045 );
not ( n10047 , n10046 );
not ( n10048 , n6314 );
nand ( n10049 , n10048 , n10045 );
nand ( n10050 , n10047 , n10049 , n2 );
nand ( n10051 , n10043 , n10050 );
not ( n10052 , n10051 );
nand ( n10053 , n10034 , n10052 );
not ( n10054 , n10053 );
not ( n10055 , n97 );
not ( n10056 , n6223 );
not ( n10057 , n6312 );
or ( n10058 , n10056 , n10057 );
or ( n10059 , n6223 , n6312 );
nand ( n10060 , n10058 , n10059 );
and ( n10061 , n6308 , n10060 );
or ( n10062 , n6308 , n10060 );
nand ( n10063 , n10062 , n2 );
or ( n10064 , n10061 , n10063 );
xnor ( n10065 , n9289 , n9269 );
or ( n10066 , n2 , n10065 );
nand ( n10067 , n10064 , n10066 );
not ( n10068 , n10067 );
nand ( n10069 , n10055 , n10068 );
not ( n10070 , n10069 );
not ( n10071 , n98 );
not ( n10072 , n9414 );
not ( n10073 , n9239 );
nand ( n10074 , n9268 , n10073 );
and ( n10075 , n10074 , n9266 );
not ( n10076 , n10074 );
and ( n10077 , n10076 , n9265 );
nor ( n10078 , n10075 , n10077 );
not ( n10079 , n10078 );
or ( n10080 , n10072 , n10079 );
not ( n10081 , n6260 );
not ( n10082 , n6261 );
nor ( n10083 , n10081 , n10082 );
nor ( n10084 , n6306 , n10083 );
not ( n10085 , n10084 );
nand ( n10086 , n6306 , n10083 );
nand ( n10087 , n10085 , n2 , n10086 );
nand ( n10088 , n10080 , n10087 );
not ( n10089 , n10088 );
or ( n10090 , n10071 , n10089 );
not ( n10091 , n9414 );
not ( n10092 , n9255 );
not ( n10093 , n9264 );
nor ( n10094 , n10093 , n9262 );
not ( n10095 , n10094 );
or ( n10096 , n10092 , n10095 );
or ( n10097 , n9255 , n10094 );
nand ( n10098 , n10096 , n10097 );
not ( n10099 , n10098 );
or ( n10100 , n10091 , n10099 );
not ( n10101 , n6284 );
nand ( n10102 , n6305 , n6302 );
nor ( n10103 , n10101 , n10102 );
not ( n10104 , n10103 );
nand ( n10105 , n10101 , n10102 );
nand ( n10106 , n10104 , n10105 , n2 );
nand ( n10107 , n10100 , n10106 );
and ( n10108 , n99 , n10107 );
not ( n10109 , n98 );
not ( n10110 , n10109 );
not ( n10111 , n10088 );
or ( n10112 , n10110 , n10111 );
or ( n10113 , n10109 , n10088 );
nand ( n10114 , n10112 , n10113 );
nand ( n10115 , n10108 , n10114 );
nand ( n10116 , n10090 , n10115 );
not ( n10117 , n10116 );
or ( n10118 , n10070 , n10117 );
nand ( n10119 , n97 , n10067 );
nand ( n10120 , n10118 , n10119 );
not ( n10121 , n10120 );
or ( n10122 , n10054 , n10121 );
nand ( n10123 , n96 , n10051 );
nand ( n10124 , n10122 , n10123 );
nand ( n10125 , n9987 , n9985 );
and ( n10126 , n10124 , n10125 );
nor ( n10127 , n9967 , n9985 );
not ( n10128 , n10127 );
nand ( n10129 , n10126 , n10128 );
not ( n10130 , n10129 );
nand ( n10131 , n10028 , n10130 , n10032 );
not ( n10132 , n10020 );
not ( n10133 , n10027 );
or ( n10134 , n10132 , n10133 );
not ( n10135 , n10029 );
nand ( n10136 , n10135 , n10030 );
not ( n10137 , n10136 );
nand ( n10138 , n10134 , n10137 );
not ( n10139 , n10020 );
nand ( n10140 , n10139 , n10026 );
nand ( n10141 , n10033 , n10131 , n10138 , n10140 );
nor ( n10142 , n9872 , n9891 );
nor ( n10143 , n9916 , n9909 );
nor ( n10144 , n10142 , n10143 );
nand ( n10145 , n10141 , n10144 , n9829 , n9924 );
nand ( n10146 , n9937 , n10145 );
not ( n10147 , n9753 );
nand ( n10148 , n10147 , n9790 );
nand ( n10149 , n10148 , n9782 );
not ( n10150 , n10149 );
nand ( n10151 , n9788 , n10146 , n10150 , n9697 );
nand ( n10152 , n9789 , n10151 );
buf ( n10153 , n10152 );
not ( n10154 , n4816 );
nand ( n10155 , n10154 , n4981 , n5346 );
not ( n10156 , n6374 );
not ( n10157 , n5351 );
not ( n10158 , n4816 );
nand ( n10159 , n10157 , n10158 );
nand ( n10160 , n10155 , n5353 , n10156 , n10159 );
not ( n10161 , n10160 );
not ( n10162 , n5358 );
not ( n10163 , n10162 );
or ( n10164 , n10161 , n10163 );
not ( n10165 , n4361 );
nand ( n10166 , n10164 , n10165 );
not ( n10167 , n4519 );
nor ( n10168 , n10167 , n5359 );
nor ( n10169 , n10166 , n10168 );
not ( n10170 , n10169 );
nand ( n10171 , n10166 , n10168 );
nand ( n10172 , n10170 , n10171 , n2 );
not ( n10173 , n8473 );
nand ( n10174 , n10173 , n8455 );
not ( n10175 , n10174 );
not ( n10176 , n8468 );
not ( n10177 , n8146 );
not ( n10178 , n10177 );
not ( n10179 , n8424 );
or ( n10180 , n10178 , n10179 );
buf ( n10181 , n8000 );
nand ( n10182 , n10180 , n10181 );
not ( n10183 , n8015 );
nand ( n10184 , n9319 , n8497 );
nand ( n10185 , n10182 , n10183 , n10184 );
not ( n10186 , n10185 );
or ( n10187 , n10176 , n10186 );
not ( n10188 , n8478 );
buf ( n10189 , n10188 );
nand ( n10190 , n10187 , n10189 );
not ( n10191 , n10190 );
or ( n10192 , n10175 , n10191 );
or ( n10193 , n10174 , n10190 );
nand ( n10194 , n10192 , n10193 );
nand ( n10195 , n10194 , n9414 );
nand ( n10196 , n10172 , n10195 );
not ( n10197 , n10196 );
not ( n10198 , n10160 );
nand ( n10199 , n10165 , n10162 );
nor ( n10200 , n10198 , n10199 );
not ( n10201 , n10200 );
nand ( n10202 , n10198 , n10199 );
nand ( n10203 , n10201 , n10202 , n2 );
and ( n10204 , n10188 , n8468 );
not ( n10205 , n10204 );
and ( n10206 , n10182 , n10183 , n10184 );
not ( n10207 , n10206 );
or ( n10208 , n10205 , n10207 );
or ( n10209 , n10204 , n10206 );
nand ( n10210 , n10208 , n10209 );
nand ( n10211 , n9414 , n10210 );
nand ( n10212 , n10203 , n10211 );
not ( n10213 , n10212 );
not ( n10214 , n10213 );
nor ( n10215 , n10197 , n10214 );
not ( n10216 , n10215 );
not ( n10217 , n2 );
not ( n10218 , n6375 );
not ( n10219 , n10218 );
nand ( n10220 , n4646 , n10219 );
not ( n10221 , n10220 );
not ( n10222 , n5360 );
not ( n10223 , n10160 );
or ( n10224 , n10222 , n10223 );
buf ( n10225 , n4521 );
buf ( n10226 , n10225 );
nand ( n10227 , n10224 , n10226 );
not ( n10228 , n10227 );
or ( n10229 , n10221 , n10228 );
or ( n10230 , n10220 , n10227 );
nand ( n10231 , n10229 , n10230 );
not ( n10232 , n10231 );
or ( n10233 , n10217 , n10232 );
not ( n10234 , n8469 );
not ( n10235 , n10185 );
or ( n10236 , n10234 , n10235 );
buf ( n10237 , n8480 );
not ( n10238 , n10237 );
nand ( n10239 , n10236 , n10238 );
buf ( n10240 , n8482 );
not ( n10241 , n7581 );
not ( n10242 , n10241 );
nor ( n10243 , n10240 , n10242 );
nor ( n10244 , n10239 , n10243 );
not ( n10245 , n10244 );
nand ( n10246 , n10239 , n10243 );
nand ( n10247 , n10245 , n9414 , n10246 );
nand ( n10248 , n10233 , n10247 );
not ( n10249 , n10196 );
nand ( n10250 , n10248 , n10249 );
not ( n10251 , n9638 );
buf ( n10252 , n4981 );
nand ( n10253 , n10251 , n10252 );
not ( n10254 , n10253 );
not ( n10255 , n10157 );
not ( n10256 , n10255 );
or ( n10257 , n10254 , n10256 );
and ( n10258 , n5353 , n10158 );
nor ( n10259 , n10258 , n9414 );
nand ( n10260 , n10257 , n10259 );
not ( n10261 , n10177 );
nand ( n10262 , n8149 , n9654 );
not ( n10263 , n10262 );
or ( n10264 , n10261 , n10263 );
and ( n10265 , n10183 , n10181 );
nor ( n10266 , n10265 , n2 );
nand ( n10267 , n10264 , n10266 );
nand ( n10268 , n10260 , n10267 );
not ( n10269 , n9414 );
not ( n10270 , n5355 );
not ( n10271 , n10158 );
nor ( n10272 , n10270 , n10271 );
nand ( n10273 , n10269 , n10272 , n10253 );
and ( n10274 , n9414 , n8147 );
nand ( n10275 , n10274 , n10181 , n10262 );
nand ( n10276 , n10273 , n10275 );
nor ( n10277 , n10268 , n10276 );
not ( n10278 , n10277 );
not ( n10279 , n9663 );
nand ( n10280 , n10278 , n10279 );
not ( n10281 , n10280 );
and ( n10282 , n10260 , n10267 , n10273 , n10275 );
not ( n10283 , n10282 );
nor ( n10284 , n10283 , n10213 );
nor ( n10285 , n10281 , n10284 );
nand ( n10286 , n10216 , n10250 , n10285 );
not ( n10287 , n10286 );
not ( n10288 , n9565 );
not ( n10289 , n2 );
nor ( n10290 , n10225 , n10218 );
not ( n10291 , n10290 );
nand ( n10292 , n10160 , n6376 );
nand ( n10293 , n10291 , n10292 , n4646 );
nand ( n10294 , n9422 , n4763 );
not ( n10295 , n10294 );
and ( n10296 , n10293 , n10295 );
not ( n10297 , n10293 );
and ( n10298 , n10297 , n10294 );
nor ( n10299 , n10296 , n10298 );
not ( n10300 , n10299 );
or ( n10301 , n10289 , n10300 );
and ( n10302 , n8488 , n8013 );
not ( n10303 , n10302 );
nand ( n10304 , n10185 , n9320 );
and ( n10305 , n10237 , n10241 );
nor ( n10306 , n10305 , n10240 );
nand ( n10307 , n10303 , n10304 , n10306 );
not ( n10308 , n10302 );
nand ( n10309 , n10304 , n10306 );
not ( n10310 , n10309 );
or ( n10311 , n10308 , n10310 );
nand ( n10312 , n10311 , n9414 );
not ( n10313 , n10312 );
nand ( n10314 , n10307 , n10313 );
nand ( n10315 , n10301 , n10314 );
or ( n10316 , n10288 , n10315 );
not ( n10317 , n10248 );
nand ( n10318 , n10317 , n10315 );
nand ( n10319 , n10316 , n10318 );
not ( n10320 , n10319 );
nand ( n10321 , n9596 , n10153 , n10287 , n10320 );
not ( n10322 , n10321 );
buf ( n10323 , n10322 );
not ( n10324 , n2 );
not ( n10325 , n6573 );
nand ( n10326 , n9424 , n10325 );
nand ( n10327 , n6576 , n6466 );
not ( n10328 , n10327 );
and ( n10329 , n10326 , n10328 );
not ( n10330 , n10326 );
and ( n10331 , n10330 , n10327 );
nor ( n10332 , n10329 , n10331 );
not ( n10333 , n10332 );
or ( n10334 , n10324 , n10333 );
not ( n10335 , n9326 );
not ( n10336 , n7285 );
and ( n10337 , n7290 , n6831 );
nand ( n10338 , n10336 , n10337 );
not ( n10339 , n10338 );
not ( n10340 , n10339 );
or ( n10341 , n10335 , n10340 );
nand ( n10342 , n10341 , n10337 );
nand ( n10343 , n10336 , n9326 , n10338 );
nand ( n10344 , n10342 , n9414 , n10343 );
nand ( n10345 , n10334 , n10344 );
not ( n10346 , n10345 );
and ( n10347 , n9452 , n10346 );
not ( n10348 , n9593 );
and ( n10349 , n10348 , n10345 );
nor ( n10350 , n10347 , n10349 );
not ( n10351 , n10350 );
not ( n10352 , n10351 );
nand ( n10353 , n9458 , n9521 , n10323 , n10352 );
not ( n10354 , n10353 );
not ( n10355 , n10354 );
not ( n10356 , n9520 );
not ( n10357 , n10356 );
not ( n10358 , n9460 );
nor ( n10359 , n10357 , n10358 );
buf ( n10360 , n9357 );
nor ( n10361 , n10360 , n9459 );
not ( n10362 , n10361 );
not ( n10363 , n10345 );
nand ( n10364 , n9593 , n10363 );
not ( n10365 , n10364 );
nand ( n10366 , n9452 , n10346 );
nand ( n10367 , n10365 , n10366 );
not ( n10368 , n10346 );
nand ( n10369 , n9453 , n10368 );
nand ( n10370 , n10367 , n10369 );
nand ( n10371 , n9456 , n10370 );
nand ( n10372 , n9452 , n9357 );
not ( n10373 , n10372 );
nand ( n10374 , n10360 , n9459 );
nand ( n10375 , n10373 , n10374 );
nand ( n10376 , n10362 , n10371 , n10375 );
not ( n10377 , n10248 );
not ( n10378 , n10377 );
not ( n10379 , n10315 );
not ( n10380 , n10379 );
or ( n10381 , n10378 , n10380 );
nand ( n10382 , n10381 , n10288 );
or ( n10383 , n10382 , n9595 );
not ( n10384 , n9568 );
nand ( n10385 , n10384 , n9565 , n9570 , n9547 );
not ( n10386 , n10385 );
nand ( n10387 , n10386 , n9594 );
nand ( n10388 , n10383 , n10387 );
not ( n10389 , n10388 );
not ( n10390 , n9595 );
not ( n10391 , n10249 );
not ( n10392 , n10212 );
nand ( n10393 , n10392 , n10277 );
not ( n10394 , n10279 );
nor ( n10395 , n10393 , n10394 );
not ( n10396 , n10395 );
or ( n10397 , n10391 , n10396 );
nand ( n10398 , n10397 , n10377 );
not ( n10399 , n10398 );
nand ( n10400 , n10390 , n10399 , n10320 );
or ( n10401 , n9593 , n9572 );
nand ( n10402 , n10389 , n10400 , n10401 );
buf ( n10403 , n10402 );
nor ( n10404 , n10376 , n10403 );
nand ( n10405 , n10355 , n1 , n10359 , n10404 );
nand ( n10406 , n3086 , n10405 );
not ( n10407 , n10349 );
buf ( n10408 , n10364 );
nand ( n10409 , n10407 , n10408 );
not ( n10410 , n10409 );
nor ( n10411 , n10410 , n237 );
not ( n10412 , n10411 );
nand ( n10413 , n10389 , n10400 , n10401 );
nor ( n10414 , n10322 , n10413 );
not ( n10415 , n10414 );
not ( n10416 , n10415 );
or ( n10417 , n10412 , n10416 );
nor ( n10418 , n10409 , n237 );
not ( n10419 , n10418 );
not ( n10420 , n10414 );
or ( n10421 , n10419 , n10420 );
and ( n10422 , n3061 , n2994 );
nor ( n10423 , n2947 , n10422 );
not ( n10424 , n10423 );
nand ( n10425 , n2947 , n10422 );
nand ( n10426 , n10424 , n237 , n10425 );
nand ( n10427 , n10421 , n10426 );
not ( n10428 , n10427 );
nand ( n10429 , n10417 , n10428 );
buf ( n10430 , n10429 );
nand ( n10431 , n10406 , n10430 );
not ( n10432 , n10431 );
buf ( n10433 , n10148 );
not ( n10434 , n10433 );
not ( n10435 , n10434 );
not ( n10436 , n9778 );
not ( n10437 , n10436 );
nand ( n10438 , n10435 , n10437 );
not ( n10439 , n10438 );
buf ( n10440 , n10146 );
buf ( n10441 , n10440 );
not ( n10442 , n10441 );
nand ( n10443 , n1 , n10439 , n10442 );
nand ( n10444 , n1 , n10438 , n10441 );
and ( n10445 , n2909 , n2363 );
xnor ( n10446 , n2904 , n10445 );
or ( n10447 , n1 , n10446 );
nand ( n10448 , n10443 , n10444 , n10447 );
not ( n10449 , n10141 );
not ( n10450 , n10449 );
not ( n10451 , n9892 );
nor ( n10452 , n10451 , n10142 );
nor ( n10453 , n10450 , n10452 );
not ( n10454 , n10452 );
not ( n10455 , n10141 );
or ( n10456 , n10454 , n10455 );
nand ( n10457 , n10456 , n1 );
or ( n10458 , n10453 , n10457 );
and ( n10459 , n2887 , n2656 );
or ( n10460 , n10459 , n2884 );
nand ( n10461 , n10459 , n2884 );
nand ( n10462 , n10460 , n10461 , n237 );
nand ( n10463 , n10458 , n10462 );
nand ( n10464 , n16 , n10463 );
or ( n10465 , n16 , n10463 );
not ( n10466 , n10028 );
not ( n10467 , n10140 );
nor ( n10468 , n10466 , n10467 );
not ( n10469 , n10468 );
nand ( n10470 , n9991 , n10129 );
not ( n10471 , n10470 );
not ( n10472 , n10032 );
or ( n10473 , n10471 , n10472 );
nand ( n10474 , n10473 , n10136 );
not ( n10475 , n10474 );
nor ( n10476 , n10469 , n10475 );
or ( n10477 , n10468 , n10474 );
nand ( n10478 , n10477 , n1 );
or ( n10479 , n10476 , n10478 );
buf ( n10480 , n2880 );
and ( n10481 , n2883 , n2711 );
or ( n10482 , n10480 , n10481 );
and ( n10483 , n10480 , n10481 );
nor ( n10484 , n10483 , n1 );
nand ( n10485 , n10482 , n10484 );
nand ( n10486 , n10479 , n10485 );
not ( n10487 , n10486 );
nand ( n10488 , n10487 , n2801 );
not ( n10489 , n237 );
not ( n10490 , n2799 );
nor ( n10491 , n10490 , n2797 );
xor ( n10492 , n2876 , n10491 );
not ( n10493 , n10492 );
or ( n10494 , n10489 , n10493 );
nor ( n10495 , n10126 , n9988 );
not ( n10496 , n10127 );
not ( n10497 , n9986 );
nand ( n10498 , n10496 , n10497 );
nor ( n10499 , n10495 , n10498 );
not ( n10500 , n10499 );
nand ( n10501 , n10498 , n10495 );
nand ( n10502 , n10500 , n10501 , n1 );
nand ( n10503 , n10494 , n10502 );
nand ( n10504 , n19 , n10503 );
not ( n10505 , n10504 );
nand ( n10506 , n18 , n10505 );
not ( n10507 , n2878 );
nand ( n10508 , n2761 , n2763 );
and ( n10509 , n10507 , n10508 );
nor ( n10510 , n10507 , n10508 );
nor ( n10511 , n10509 , n1 , n10510 );
not ( n10512 , n10511 );
not ( n10513 , n10470 );
not ( n10514 , n10032 );
not ( n10515 , n10514 );
nand ( n10516 , n10515 , n10136 );
not ( n10517 , n10516 );
nand ( n10518 , n1 , n10513 , n10517 );
nand ( n10519 , n1 , n10470 , n10516 );
nand ( n10520 , n10512 , n10518 , n10519 );
not ( n10521 , n18 );
nand ( n10522 , n10521 , n10504 );
nand ( n10523 , n10520 , n10522 );
nand ( n10524 , n10506 , n10523 );
nand ( n10525 , n10488 , n10524 );
nand ( n10526 , n17 , n10486 );
nand ( n10527 , n10525 , n10526 );
nand ( n10528 , n10465 , n10527 );
nand ( n10529 , n10464 , n10528 );
not ( n10530 , n10142 );
not ( n10531 , n10530 );
not ( n10532 , n10141 );
or ( n10533 , n10531 , n10532 );
buf ( n10534 , n9892 );
nand ( n10535 , n10533 , n10534 );
not ( n10536 , n10535 );
not ( n10537 , n9917 );
nor ( n10538 , n10537 , n10143 );
not ( n10539 , n10538 );
nor ( n10540 , n10536 , n10539 );
or ( n10541 , n10535 , n10538 );
nand ( n10542 , n10541 , n1 );
or ( n10543 , n10540 , n10542 );
nand ( n10544 , n2892 , n2609 );
not ( n10545 , n10544 );
not ( n10546 , n2888 );
or ( n10547 , n10545 , n10546 );
or ( n10548 , n10544 , n2888 );
nand ( n10549 , n10547 , n10548 );
nand ( n10550 , n237 , n10549 );
nand ( n10551 , n10543 , n10550 );
not ( n10552 , n10551 );
not ( n10553 , n15 );
nand ( n10554 , n10552 , n10553 );
not ( n10555 , n237 );
and ( n10556 , n2898 , n2542 );
xor ( n10557 , n10556 , n2893 );
not ( n10558 , n10557 );
or ( n10559 , n10555 , n10558 );
not ( n10560 , n10144 );
not ( n10561 , n10141 );
or ( n10562 , n10560 , n10561 );
not ( n10563 , n9918 );
nand ( n10564 , n10562 , n10563 );
not ( n10565 , n10564 );
not ( n10566 , n9924 );
nor ( n10567 , n10566 , n9928 );
not ( n10568 , n10567 );
nand ( n10569 , n10565 , n10568 );
not ( n10570 , n10567 );
not ( n10571 , n10564 );
or ( n10572 , n10570 , n10571 );
nand ( n10573 , n10572 , n1 );
not ( n10574 , n10573 );
nand ( n10575 , n10569 , n10574 );
nand ( n10576 , n10559 , n10575 );
nand ( n10577 , n10529 , n10554 , n10576 );
and ( n10578 , n15 , n10551 );
nand ( n10579 , n10578 , n10576 );
and ( n10580 , n10577 , n10579 );
not ( n10581 , n9935 );
not ( n10582 , n9929 );
nor ( n10583 , n10581 , n10582 );
not ( n10584 , n10583 );
not ( n10585 , n10564 );
not ( n10586 , n9924 );
or ( n10587 , n10585 , n10586 );
not ( n10588 , n9928 );
nand ( n10589 , n10587 , n10588 );
and ( n10590 , n1 , n10584 , n10589 );
not ( n10591 , n237 );
and ( n10592 , n2903 , n2461 );
xor ( n10593 , n10592 , n2899 );
not ( n10594 , n10593 );
or ( n10595 , n10591 , n10594 );
not ( n10596 , n10589 );
nand ( n10597 , n1 , n10583 , n10596 );
nand ( n10598 , n10595 , n10597 );
nor ( n10599 , n10590 , n10598 );
nor ( n10600 , n10580 , n10599 );
nand ( n10601 , n10448 , n10600 );
not ( n10602 , n10601 );
not ( n10603 , n237 );
nor ( n10604 , n2157 , n2928 );
buf ( n10605 , n2201 );
not ( n10606 , n2189 );
nand ( n10607 , n10605 , n10606 );
xor ( n10608 , n10604 , n10607 );
not ( n10609 , n10608 );
or ( n10610 , n10603 , n10609 );
not ( n10611 , n10280 );
not ( n10612 , n10282 );
not ( n10613 , n10394 );
nor ( n10614 , n10612 , n10613 );
nor ( n10615 , n10611 , n10614 );
nor ( n10616 , n10152 , n10615 );
not ( n10617 , n10616 );
nand ( n10618 , n10152 , n10615 );
nand ( n10619 , n10617 , n10618 , n1 );
nand ( n10620 , n10610 , n10619 );
buf ( n10621 , n9782 );
not ( n10622 , n10621 );
not ( n10623 , n10622 );
nand ( n10624 , n10623 , n9745 );
not ( n10625 , n10624 );
not ( n10626 , n10145 );
and ( n10627 , n10433 , n10626 );
not ( n10628 , n10148 );
not ( n10629 , n9936 );
or ( n10630 , n10628 , n10629 );
nand ( n10631 , n10630 , n10437 );
nor ( n10632 , n10627 , n10631 );
not ( n10633 , n10632 );
or ( n10634 , n10625 , n10633 );
nand ( n10635 , n10634 , n1 );
not ( n10636 , n10631 );
not ( n10637 , n10627 );
and ( n10638 , n10636 , n10637 );
nor ( n10639 , n10638 , n10624 );
or ( n10640 , n10635 , n10639 );
xor ( n10641 , n2921 , n2910 );
nand ( n10642 , n237 , n10641 );
nand ( n10643 , n10640 , n10642 );
not ( n10644 , n9694 );
not ( n10645 , n10644 );
not ( n10646 , n9697 );
nor ( n10647 , n10645 , n10646 );
not ( n10648 , n10647 );
nand ( n10649 , n10150 , n10626 );
not ( n10650 , n9745 );
not ( n10651 , n10436 );
not ( n10652 , n10651 );
or ( n10653 , n10650 , n10652 );
nand ( n10654 , n10653 , n10621 );
nand ( n10655 , n10150 , n9936 );
nand ( n10656 , n10649 , n10654 , n10655 );
not ( n10657 , n10656 );
or ( n10658 , n10648 , n10657 );
nand ( n10659 , n10658 , n1 );
nor ( n10660 , n10656 , n10647 );
or ( n10661 , n10659 , n10660 );
buf ( n10662 , n2113 );
nand ( n10663 , n10662 , n2217 );
not ( n10664 , n10663 );
not ( n10665 , n2926 );
or ( n10666 , n10664 , n10665 );
or ( n10667 , n10663 , n2926 );
nand ( n10668 , n10666 , n10667 );
nand ( n10669 , n237 , n10668 );
nand ( n10670 , n10661 , n10669 );
and ( n10671 , n10643 , n10670 );
not ( n10672 , n237 );
not ( n10673 , n2154 );
nand ( n10674 , n10673 , n2156 );
not ( n10675 , n10674 );
nand ( n10676 , n10662 , n2927 );
not ( n10677 , n10676 );
or ( n10678 , n10675 , n10677 );
or ( n10679 , n10674 , n10676 );
nand ( n10680 , n10678 , n10679 );
not ( n10681 , n10680 );
or ( n10682 , n10672 , n10681 );
nand ( n10683 , n9783 , n10644 );
not ( n10684 , n10683 );
not ( n10685 , n10646 );
nand ( n10686 , n10440 , n10150 , n10685 );
and ( n10687 , n10684 , n10686 );
not ( n10688 , n9624 );
nor ( n10689 , n10688 , n9787 );
not ( n10690 , n10689 );
nand ( n10691 , n10690 , n9788 );
nor ( n10692 , n10687 , n10691 );
not ( n10693 , n10692 );
nand ( n10694 , n10691 , n10684 , n10686 );
nand ( n10695 , n10693 , n1 , n10694 );
nand ( n10696 , n10682 , n10695 );
and ( n10697 , n10620 , n10671 , n10696 );
not ( n10698 , n10213 );
xnor ( n10699 , n10282 , n10698 );
not ( n10700 , n10699 );
nand ( n10701 , n10152 , n10280 );
not ( n10702 , n10614 );
nand ( n10703 , n1 , n10700 , n10701 , n10702 );
not ( n10704 , n2203 );
nor ( n10705 , n10704 , n2198 );
not ( n10706 , n10606 );
not ( n10707 , n10604 );
not ( n10708 , n10707 );
or ( n10709 , n10706 , n10708 );
nand ( n10710 , n10709 , n10605 );
nor ( n10711 , n10705 , n10710 );
not ( n10712 , n10711 );
nand ( n10713 , n10705 , n10710 );
nand ( n10714 , n10712 , n237 , n10713 );
nand ( n10715 , n10701 , n10702 );
nand ( n10716 , n1 , n10699 , n10715 );
nand ( n10717 , n10703 , n10714 , n10716 );
nand ( n10718 , n10602 , n10697 , n10717 );
not ( n10719 , n10718 );
not ( n10720 , n10152 );
not ( n10721 , n10286 );
not ( n10722 , n10721 );
or ( n10723 , n10720 , n10722 );
nand ( n10724 , n10723 , n10398 );
buf ( n10725 , n10724 );
not ( n10726 , n10318 );
buf ( n10727 , n10315 );
not ( n10728 , n10727 );
not ( n10729 , n10377 );
nand ( n10730 , n10728 , n10729 );
not ( n10731 , n10730 );
nor ( n10732 , n10726 , n10731 );
nand ( n10733 , n10725 , n10732 );
not ( n10734 , n10733 );
or ( n10735 , n10725 , n10732 );
nand ( n10736 , n10735 , n1 );
or ( n10737 , n10734 , n10736 );
nand ( n10738 , n2934 , n1297 );
not ( n10739 , n10738 );
not ( n10740 , n2930 );
or ( n10741 , n10739 , n10740 );
or ( n10742 , n10738 , n2930 );
nand ( n10743 , n10741 , n10742 );
nand ( n10744 , n237 , n10743 );
nand ( n10745 , n10737 , n10744 );
not ( n10746 , n10698 );
not ( n10747 , n10249 );
nor ( n10748 , n10746 , n10747 );
not ( n10749 , n10748 );
not ( n10750 , n10152 );
not ( n10751 , n10285 );
or ( n10752 , n10750 , n10751 );
nor ( n10753 , n10698 , n10282 );
nor ( n10754 , n10393 , n10613 );
nor ( n10755 , n10753 , n10754 );
nand ( n10756 , n10752 , n10755 );
not ( n10757 , n10215 );
buf ( n10758 , n10757 );
nand ( n10759 , n10756 , n10758 );
and ( n10760 , n10749 , n10759 );
xor ( n10761 , n10747 , n10729 );
nor ( n10762 , n10760 , n10761 );
not ( n10763 , n10761 );
nand ( n10764 , n10749 , n10759 );
or ( n10765 , n10763 , n10764 );
nand ( n10766 , n10765 , n1 );
or ( n10767 , n10762 , n10766 );
and ( n10768 , n2212 , n1405 );
not ( n10769 , n2208 );
or ( n10770 , n10768 , n10769 );
not ( n10771 , n2199 );
not ( n10772 , n10707 );
or ( n10773 , n10771 , n10772 );
not ( n10774 , n2204 );
nand ( n10775 , n10773 , n10774 );
or ( n10776 , n10770 , n10775 );
nand ( n10777 , n10775 , n10768 , n1712 );
and ( n10778 , n10768 , n10769 );
nor ( n10779 , n1712 , n10768 , n10769 );
nor ( n10780 , n10778 , n10779 , n1 );
nand ( n10781 , n10776 , n10777 , n10780 );
nand ( n10782 , n10767 , n10781 );
not ( n10783 , n10757 );
nor ( n10784 , n10783 , n10748 );
nor ( n10785 , n10756 , n10784 );
not ( n10786 , n10785 );
nand ( n10787 , n10756 , n10784 );
nand ( n10788 , n10786 , n10787 , n1 );
nand ( n10789 , n2208 , n1712 );
not ( n10790 , n10789 );
not ( n10791 , n10775 );
or ( n10792 , n10790 , n10791 );
or ( n10793 , n10789 , n10775 );
nand ( n10794 , n10792 , n10793 );
nand ( n10795 , n237 , n10794 );
nand ( n10796 , n10788 , n10795 );
nand ( n10797 , n10719 , n10745 , n10782 , n10796 );
not ( n10798 , n10797 );
not ( n10799 , n10319 );
and ( n10800 , n10153 , n10799 , n10287 );
not ( n10801 , n10399 );
not ( n10802 , n10799 );
or ( n10803 , n10801 , n10802 );
nand ( n10804 , n10803 , n10382 );
nor ( n10805 , n10800 , n10804 );
not ( n10806 , n10805 );
not ( n10807 , n10385 );
not ( n10808 , n10807 );
not ( n10809 , n10808 );
not ( n10810 , n9566 );
buf ( n10811 , n10810 );
not ( n10812 , n10811 );
nor ( n10813 , n10809 , n10812 );
nor ( n10814 , n10813 , n237 );
nand ( n10815 , n10806 , n10814 );
nand ( n10816 , n2941 , n843 );
not ( n10817 , n10816 );
nand ( n10818 , n1304 , n2930 );
not ( n10819 , n2937 );
nand ( n10820 , n10818 , n10819 );
not ( n10821 , n10820 );
not ( n10822 , n10821 );
or ( n10823 , n10817 , n10822 );
not ( n10824 , n10816 );
not ( n10825 , n10824 );
not ( n10826 , n10820 );
or ( n10827 , n10825 , n10826 );
nand ( n10828 , n10827 , n237 );
not ( n10829 , n10828 );
nand ( n10830 , n10823 , n10829 );
nand ( n10831 , n1 , n10805 , n10813 );
nand ( n10832 , n10815 , n10830 , n10831 );
not ( n10833 , n10832 );
not ( n10834 , n10833 );
buf ( n10835 , n10727 );
and ( n10836 , n10835 , n9565 );
not ( n10837 , n10835 );
and ( n10838 , n10837 , n10288 );
or ( n10839 , n10836 , n10838 );
not ( n10840 , n10839 );
not ( n10841 , n10318 );
not ( n10842 , n10724 );
or ( n10843 , n10841 , n10842 );
nand ( n10844 , n10843 , n10730 );
not ( n10845 , n10844 );
nor ( n10846 , n10840 , n10845 );
or ( n10847 , n10839 , n10844 );
nand ( n10848 , n10847 , n1 );
or ( n10849 , n10846 , n10848 );
not ( n10850 , n1297 );
not ( n10851 , n2930 );
or ( n10852 , n10850 , n10851 );
nand ( n10853 , n10852 , n2934 );
not ( n10854 , n10853 );
not ( n10855 , n1303 );
nand ( n10856 , n10855 , n2936 );
not ( n10857 , n10856 );
or ( n10858 , n10854 , n10857 );
or ( n10859 , n10853 , n10856 );
nand ( n10860 , n10858 , n10859 );
nand ( n10861 , n237 , n10860 );
nand ( n10862 , n10849 , n10861 );
not ( n10863 , n10862 );
not ( n10864 , n10863 );
nand ( n10865 , n10834 , n10864 );
nand ( n10866 , n10153 , n10287 , n10799 , n10811 );
and ( n10867 , n10399 , n10799 , n10811 );
not ( n10868 , n10810 );
nor ( n10869 , n10868 , n10382 );
nor ( n10870 , n10867 , n10869 );
not ( n10871 , n10807 );
and ( n10872 , n10866 , n10870 , n10871 );
nand ( n10873 , n10401 , n9594 );
nor ( n10874 , n10872 , n10873 );
not ( n10875 , n10874 );
nand ( n10876 , n10873 , n10870 , n10866 , n10871 );
nand ( n10877 , n10875 , n10876 , n1 );
not ( n10878 , n2944 );
nand ( n10879 , n10878 , n667 );
not ( n10880 , n10879 );
not ( n10881 , n2942 );
not ( n10882 , n2931 );
nand ( n10883 , n10881 , n10882 );
not ( n10884 , n10883 );
or ( n10885 , n10880 , n10884 );
or ( n10886 , n10879 , n10883 );
nand ( n10887 , n10885 , n10886 );
nand ( n10888 , n237 , n10887 );
nand ( n10889 , n10877 , n10888 );
not ( n10890 , n10889 );
nor ( n10891 , n10865 , n10890 );
nand ( n10892 , n10798 , n10891 );
not ( n10893 , n10892 );
nor ( n10894 , n3057 , n281 );
not ( n10895 , n10894 );
not ( n10896 , n319 );
nor ( n10897 , n3049 , n3039 );
and ( n10898 , n10897 , n2994 );
nand ( n10899 , n10896 , n10898 );
or ( n10900 , n2932 , n10899 );
nand ( n10901 , n10900 , n3053 );
not ( n10902 , n3061 );
and ( n10903 , n10897 , n10902 );
or ( n10904 , n3049 , n3066 );
nand ( n10905 , n10904 , n3059 );
nor ( n10906 , n10903 , n10905 );
not ( n10907 , n2945 );
nand ( n10908 , n10898 , n10907 );
and ( n10909 , n10906 , n10908 );
nor ( n10910 , n10909 , n319 );
nor ( n10911 , n10901 , n10910 );
nand ( n10912 , n10895 , n10911 );
not ( n10913 , n10912 );
not ( n10914 , n10911 );
and ( n10915 , n10894 , n10914 );
nor ( n10916 , n10915 , n1 );
not ( n10917 , n10916 );
or ( n10918 , n10913 , n10917 );
nor ( n10919 , n10351 , n9457 );
nand ( n10920 , n10357 , n9521 , n10323 , n10919 );
not ( n10921 , n10920 );
not ( n10922 , n10376 );
not ( n10923 , n10403 );
nand ( n10924 , n10359 , n10353 , n10922 , n10923 );
not ( n10925 , n10924 );
or ( n10926 , n10921 , n10925 );
nand ( n10927 , n10926 , n1 );
nand ( n10928 , n10918 , n10927 );
and ( n10929 , n10893 , n10928 );
not ( n10930 , n3065 );
nand ( n10931 , n10930 , n3033 );
not ( n10932 , n3038 );
not ( n10933 , n2994 );
not ( n10934 , n2946 );
or ( n10935 , n10933 , n10934 );
nand ( n10936 , n10935 , n3061 );
not ( n10937 , n10936 );
or ( n10938 , n10932 , n10937 );
not ( n10939 , n3063 );
nand ( n10940 , n10938 , n10939 );
not ( n10941 , n10940 );
and ( n10942 , n10931 , n10941 );
not ( n10943 , n10931 );
not ( n10944 , n10943 );
not ( n10945 , n10940 );
or ( n10946 , n10944 , n10945 );
nand ( n10947 , n10946 , n237 );
nor ( n10948 , n10942 , n10947 );
not ( n10949 , n10948 );
not ( n10950 , n10350 );
not ( n10951 , n10402 );
or ( n10952 , n10950 , n10951 );
not ( n10953 , n10370 );
nand ( n10954 , n10952 , n10953 );
not ( n10955 , n10954 );
not ( n10956 , n9455 );
not ( n10957 , n10956 );
not ( n10958 , n10372 );
nor ( n10959 , n10957 , n10958 );
not ( n10960 , n10321 );
not ( n10961 , n10351 );
nand ( n10962 , n10960 , n10961 );
nand ( n10963 , n10955 , n1 , n10959 , n10962 );
not ( n10964 , n10962 );
or ( n10965 , n10964 , n10954 );
nor ( n10966 , n237 , n10959 );
nand ( n10967 , n10965 , n10966 );
nand ( n10968 , n10949 , n10963 , n10967 );
not ( n10969 , n10968 );
not ( n10970 , n10408 );
nand ( n10971 , n10960 , n10407 );
not ( n10972 , n10971 );
or ( n10973 , n10970 , n10972 );
not ( n10974 , n10369 );
not ( n10975 , n10974 );
nand ( n10976 , n10975 , n10366 );
not ( n10977 , n10976 );
nand ( n10978 , n10973 , n10977 );
nand ( n10979 , n10978 , n1 );
not ( n10980 , n10322 );
not ( n10981 , n10407 );
or ( n10982 , n10980 , n10981 );
nand ( n10983 , n10982 , n10408 );
not ( n10984 , n10407 );
not ( n10985 , n10402 );
or ( n10986 , n10984 , n10985 );
nand ( n10987 , n10986 , n10976 );
nor ( n10988 , n10983 , n10987 );
nor ( n10989 , n10979 , n10988 );
and ( n10990 , n10407 , n10403 );
nand ( n10991 , n10990 , n10977 );
and ( n10992 , n10989 , n10991 );
nand ( n10993 , n10939 , n3038 );
not ( n10994 , n10936 );
not ( n10995 , n10994 );
and ( n10996 , n10993 , n10995 );
not ( n10997 , n10993 );
and ( n10998 , n10997 , n10994 );
nor ( n10999 , n10996 , n10998 );
nor ( n11000 , n10999 , n1 );
nor ( n11001 , n10992 , n11000 );
nor ( n11002 , n10969 , n11001 );
nand ( n11003 , n10415 , n10919 );
nand ( n11004 , n10922 , n11003 );
nand ( n11005 , n10358 , n10356 );
nand ( n11006 , n9521 , n11005 );
not ( n11007 , n11006 );
or ( n11008 , n11004 , n11007 );
nand ( n11009 , n11008 , n1 );
and ( n11010 , n10922 , n11003 );
nor ( n11011 , n11010 , n11006 );
or ( n11012 , n11009 , n11011 );
not ( n11013 , n3053 );
nor ( n11014 , n11013 , n319 );
not ( n11015 , n2947 );
not ( n11016 , n10898 );
or ( n11017 , n11015 , n11016 );
nand ( n11018 , n11017 , n10906 );
nor ( n11019 , n11014 , n11018 );
not ( n11020 , n11019 );
nand ( n11021 , n11014 , n11018 );
nand ( n11022 , n11020 , n11021 , n237 );
nand ( n11023 , n11012 , n11022 );
not ( n11024 , n10956 );
not ( n11025 , n10370 );
or ( n11026 , n11024 , n11025 );
not ( n11027 , n10958 );
nand ( n11028 , n11026 , n11027 );
not ( n11029 , n11028 );
not ( n11030 , n10414 );
nand ( n11031 , n11030 , n10956 , n10961 );
nand ( n11032 , n11029 , n11031 );
not ( n11033 , n10361 );
nand ( n11034 , n11033 , n10374 );
nand ( n11035 , n11032 , n1 , n11034 );
not ( n11036 , n11034 );
nand ( n11037 , n1 , n11036 , n11029 , n11031 );
and ( n11038 , n3059 , n3050 );
not ( n11039 , n3067 );
nand ( n11040 , n3041 , n11039 );
nor ( n11041 , n11038 , n11040 );
not ( n11042 , n11041 );
nand ( n11043 , n11038 , n11040 );
nand ( n11044 , n11042 , n237 , n11043 );
nand ( n11045 , n11035 , n11037 , n11044 );
nand ( n11046 , n11002 , n11023 , n11045 );
not ( n11047 , n11046 );
nand ( n11048 , n10432 , n10929 , n11047 );
not ( n11049 , n3 );
and ( n11050 , n237 , n11049 );
and ( n11051 , n1 , n3 );
nor ( n11052 , n11050 , n11051 );
and ( n11053 , n11052 , n9414 );
not ( n11054 , n11052 );
and ( n11055 , n11054 , n2 );
or ( n11056 , n11053 , n11055 );
buf ( n11057 , n11056 );
buf ( n11058 , n11057 );
not ( n11059 , n237 );
not ( n11060 , n3058 );
nand ( n11061 , n320 , n10905 );
not ( n11062 , n11061 );
or ( n11063 , n11060 , n11062 );
nand ( n11064 , n11063 , n3078 );
and ( n11065 , n3078 , n320 );
nand ( n11066 , n11065 , n10995 , n10897 );
nand ( n11067 , n11064 , n3077 , n11066 );
not ( n11068 , n11067 );
or ( n11069 , n11059 , n11068 );
nand ( n11070 , n11069 , n10405 );
nand ( n11071 , n11048 , n11058 , n11070 );
not ( n11072 , n3198 );
not ( n11073 , n11072 );
not ( n11074 , n11073 );
nand ( n11075 , n40 , n11074 );
not ( n11076 , n3906 );
nand ( n11077 , n4530 , n11076 );
not ( n11078 , n11077 );
not ( n11079 , n11078 );
not ( n11080 , n4530 );
not ( n11081 , n3482 );
nand ( n11082 , n11080 , n11081 );
nand ( n11083 , n11079 , n11082 );
buf ( n11084 , n11083 );
not ( n11085 , n11084 );
buf ( n11086 , n11085 );
not ( n11087 , n11086 );
not ( n11088 , n11087 );
buf ( n11089 , n11088 );
buf ( n11090 , n11089 );
not ( n11091 , n11090 );
and ( n11092 , n3258 , n3271 );
not ( n11093 , n11092 );
nand ( n11094 , n3259 , n3275 );
nand ( n11095 , n11093 , n11083 , n11094 );
not ( n11096 , n11095 );
not ( n11097 , n11096 );
not ( n11098 , n11097 );
not ( n11099 , n11098 );
not ( n11100 , n11099 );
not ( n11101 , n11100 );
and ( n11102 , n11091 , n11101 );
not ( n11103 , n3315 );
not ( n11104 , n11103 );
not ( n11105 , n11104 );
not ( n11106 , n11105 );
not ( n11107 , n11106 );
nor ( n11108 , n11102 , n11107 );
and ( n11109 , n37 , n3207 );
not ( n11110 , n37 );
and ( n11111 , n11110 , n3206 );
nor ( n11112 , n11109 , n11111 );
not ( n11113 , n3271 );
nand ( n11114 , n11113 , n4617 );
not ( n11115 , n11114 );
nor ( n11116 , n6423 , n4739 );
nor ( n11117 , n11115 , n11116 );
not ( n11118 , n11117 );
not ( n11119 , n3286 );
nand ( n11120 , n11119 , n6423 );
not ( n11121 , n6423 );
nand ( n11122 , n3134 , n11121 );
nand ( n11123 , n11118 , n11120 , n11122 );
not ( n11124 , n11123 );
not ( n11125 , n11124 );
not ( n11126 , n11125 );
not ( n11127 , n11126 );
not ( n11128 , n11127 );
and ( n11129 , n11112 , n11128 );
not ( n11130 , n3207 );
and ( n11131 , n3126 , n11130 );
not ( n11132 , n3208 );
nor ( n11133 , n11131 , n11132 );
not ( n11134 , n11117 );
not ( n11135 , n11134 );
not ( n11136 , n11135 );
not ( n11137 , n11136 );
not ( n11138 , n11137 );
not ( n11139 , n11138 );
not ( n11140 , n11139 );
not ( n11141 , n11140 );
and ( n11142 , n11133 , n11141 );
nor ( n11143 , n11129 , n11142 );
xnor ( n11144 , n11108 , n11143 );
or ( n11145 , n11075 , n11144 );
or ( n11146 , n11108 , n11143 );
nand ( n11147 , n11145 , n11146 );
not ( n11148 , n3198 );
nand ( n11149 , n39 , n11148 );
nand ( n11150 , n3192 , n3292 );
nand ( n11151 , n3106 , n3157 );
xnor ( n11152 , n4024 , n3132 );
and ( n11153 , n11150 , n11151 , n11152 );
not ( n11154 , n11153 );
not ( n11155 , n11154 );
not ( n11156 , n11155 );
not ( n11157 , n11156 );
not ( n11158 , n11157 );
not ( n11159 , n11158 );
and ( n11160 , n3108 , n11159 );
and ( n11161 , n11110 , n11073 );
nand ( n11162 , n37 , n11072 );
not ( n11163 , n11162 );
nor ( n11164 , n11161 , n11163 );
not ( n11165 , n11152 );
and ( n11166 , n11164 , n11165 );
nor ( n11167 , n11160 , n11166 );
xnor ( n11168 , n11149 , n11167 );
not ( n11169 , n11128 );
not ( n11170 , n11169 );
and ( n11171 , n11133 , n11170 );
not ( n11172 , n11130 );
not ( n11173 , n11141 );
not ( n11174 , n11173 );
and ( n11175 , n11172 , n11174 );
nor ( n11176 , n11171 , n11175 );
not ( n11177 , n11176 );
and ( n11178 , n11168 , n11177 );
not ( n11179 , n11168 );
and ( n11180 , n11179 , n11176 );
nor ( n11181 , n11178 , n11180 );
xor ( n11182 , n11147 , n11181 );
and ( n11183 , n3126 , n11105 );
nor ( n11184 , n11183 , n3316 );
and ( n11185 , n11184 , n11100 );
and ( n11186 , n11106 , n11090 );
nor ( n11187 , n11185 , n11186 );
not ( n11188 , n39 );
and ( n11189 , n11188 , n11073 );
not ( n11190 , n11149 );
nor ( n11191 , n11189 , n11190 );
and ( n11192 , n11191 , n11159 );
and ( n11193 , n3108 , n11165 );
nor ( n11194 , n11192 , n11193 );
xnor ( n11195 , n11187 , n11194 );
not ( n11196 , n11191 );
not ( n11197 , n11165 );
or ( n11198 , n11196 , n11197 );
or ( n11199 , n3229 , n3197 );
nand ( n11200 , n11199 , n3230 );
not ( n11201 , n11200 );
or ( n11202 , n11201 , n11158 );
nand ( n11203 , n11198 , n11202 );
buf ( n11204 , n3290 );
or ( n11205 , n11204 , n11127 );
not ( n11206 , n11112 );
or ( n11207 , n11206 , n11140 );
nand ( n11208 , n11205 , n11207 );
and ( n11209 , n41 , n3193 );
xor ( n11210 , n11208 , n11209 );
and ( n11211 , n11203 , n11210 );
and ( n11212 , n11209 , n11208 );
nor ( n11213 , n11211 , n11212 );
or ( n11214 , n11195 , n11213 );
or ( n11215 , n11187 , n11194 );
nand ( n11216 , n11214 , n11215 );
xnor ( n11217 , n11182 , n11216 );
not ( n11218 , n11217 );
xor ( n11219 , n11210 , n11203 );
not ( n11220 , n41 );
and ( n11221 , n11220 , n3194 );
nor ( n11222 , n11221 , n11209 );
and ( n11223 , n11222 , n11157 );
and ( n11224 , n11200 , n11165 );
nor ( n11225 , n11223 , n11224 );
and ( n11226 , n37 , n11104 );
and ( n11227 , n11110 , n11103 );
nor ( n11228 , n11226 , n11227 );
not ( n11229 , n11099 );
and ( n11230 , n11228 , n11229 );
and ( n11231 , n11184 , n11089 );
nor ( n11232 , n11230 , n11231 );
not ( n11233 , n4545 );
not ( n11234 , n3415 );
or ( n11235 , n11233 , n11234 );
nand ( n11236 , n3433 , n3414 );
nand ( n11237 , n11235 , n11236 );
buf ( n11238 , n11237 );
not ( n11239 , n11238 );
not ( n11240 , n11239 );
not ( n11241 , n11240 );
not ( n11242 , n11241 );
not ( n11243 , n4420 );
and ( n11244 , n3433 , n11243 );
not ( n11245 , n11244 );
nand ( n11246 , n6398 , n4666 );
nand ( n11247 , n11245 , n11246 , n11237 );
not ( n11248 , n11247 );
not ( n11249 , n11248 );
not ( n11250 , n11249 );
not ( n11251 , n11250 );
not ( n11252 , n11251 );
not ( n11253 , n11252 );
and ( n11254 , n11242 , n11253 );
buf ( n11255 , n4420 );
not ( n11256 , n11255 );
buf ( n11257 , n11256 );
buf ( n11258 , n11257 );
not ( n11259 , n11258 );
nor ( n11260 , n11254 , n11259 );
xnor ( n11261 , n11232 , n11260 );
or ( n11262 , n11225 , n11261 );
or ( n11263 , n11260 , n11232 );
nand ( n11264 , n11262 , n11263 );
xor ( n11265 , n11264 , n11187 );
and ( n11266 , n11219 , n11265 );
and ( n11267 , n11187 , n11264 );
nor ( n11268 , n11266 , n11267 );
xnor ( n11269 , n11075 , n11144 );
xnor ( n11270 , n11195 , n11213 );
xnor ( n11271 , n11269 , n11270 );
or ( n11272 , n11268 , n11271 );
or ( n11273 , n11269 , n11270 );
nand ( n11274 , n11272 , n11273 );
nand ( n11275 , n11218 , n11274 );
not ( n11276 , n11274 );
nand ( n11277 , n11217 , n11276 );
nand ( n11278 , n11275 , n11277 );
xor ( n11279 , n11271 , n11268 );
and ( n11280 , n39 , n3205 );
and ( n11281 , n11188 , n3204 );
nor ( n11282 , n11280 , n11281 );
not ( n11283 , n11282 );
not ( n11284 , n11128 );
or ( n11285 , n11283 , n11284 );
or ( n11286 , n11204 , n11140 );
nand ( n11287 , n11285 , n11286 );
nor ( n11288 , n3502 , n11073 );
xor ( n11289 , n11287 , n11288 );
not ( n11290 , n6476 );
not ( n11291 , n11099 );
and ( n11292 , n11290 , n11291 );
not ( n11293 , n11087 );
and ( n11294 , n11228 , n11293 );
nor ( n11295 , n11292 , n11294 );
not ( n11296 , n11295 );
and ( n11297 , n11289 , n11296 );
not ( n11298 , n11289 );
and ( n11299 , n11298 , n11295 );
nor ( n11300 , n11297 , n11299 );
xor ( n11301 , n11261 , n11225 );
not ( n11302 , n11259 );
not ( n11303 , n11242 );
and ( n11304 , n11302 , n11303 );
not ( n11305 , n11253 );
and ( n11306 , n11305 , n4672 );
nor ( n11307 , n11304 , n11306 );
nand ( n11308 , n43 , n3106 );
not ( n11309 , n3104 );
or ( n11310 , n3502 , n11309 );
nand ( n11311 , n11310 , n4727 );
and ( n11312 , n11311 , n11155 );
and ( n11313 , n11222 , n11165 );
nor ( n11314 , n11312 , n11313 );
xnor ( n11315 , n11308 , n11314 );
or ( n11316 , n11307 , n11315 );
or ( n11317 , n11308 , n11314 );
nand ( n11318 , n11316 , n11317 );
xor ( n11319 , n11301 , n11318 );
and ( n11320 , n11300 , n11319 );
and ( n11321 , n11318 , n11301 );
nor ( n11322 , n11320 , n11321 );
and ( n11323 , n11296 , n11289 );
and ( n11324 , n11288 , n11287 );
nor ( n11325 , n11323 , n11324 );
xnor ( n11326 , n11219 , n11265 );
xnor ( n11327 , n11325 , n11326 );
or ( n11328 , n11322 , n11327 );
or ( n11329 , n11325 , n11326 );
nand ( n11330 , n11328 , n11329 );
nor ( n11331 , n11279 , n11330 );
xor ( n11332 , n11327 , n11322 );
nand ( n11333 , n44 , n11072 );
not ( n11334 , n6476 );
not ( n11335 , n11087 );
and ( n11336 , n11334 , n11335 );
and ( n11337 , n39 , n3315 );
not ( n11338 , n3314 );
not ( n11339 , n11338 );
and ( n11340 , n11188 , n11339 );
nor ( n11341 , n11337 , n11340 );
and ( n11342 , n11341 , n11098 );
nor ( n11343 , n11336 , n11342 );
not ( n11344 , n43 );
and ( n11345 , n11344 , n3104 );
not ( n11346 , n11308 );
nor ( n11347 , n11345 , n11346 );
and ( n11348 , n11347 , n11155 );
and ( n11349 , n11311 , n11165 );
nor ( n11350 , n11348 , n11349 );
xnor ( n11351 , n11343 , n11350 );
or ( n11352 , n11333 , n11351 );
or ( n11353 , n11343 , n11350 );
nand ( n11354 , n11352 , n11353 );
not ( n11355 , n4685 );
or ( n11356 , n11355 , n11125 );
not ( n11357 , n11282 );
or ( n11358 , n11357 , n11138 );
nand ( n11359 , n11356 , n11358 );
and ( n11360 , n11359 , n11295 );
not ( n11361 , n11359 );
and ( n11362 , n11361 , n11296 );
nor ( n11363 , n11360 , n11362 );
xor ( n11364 , n11354 , n11363 );
and ( n11365 , n41 , n3136 );
and ( n11366 , n11220 , n3135 );
nor ( n11367 , n11365 , n11366 );
and ( n11368 , n11367 , n11126 );
and ( n11369 , n4685 , n11139 );
nor ( n11370 , n11368 , n11369 );
not ( n11371 , n11251 );
and ( n11372 , n37 , n11258 );
not ( n11373 , n11258 );
and ( n11374 , n11110 , n11373 );
nor ( n11375 , n11372 , n11374 );
and ( n11376 , n11371 , n11375 );
and ( n11377 , n4672 , n11241 );
nor ( n11378 , n11376 , n11377 );
not ( n11379 , n3547 );
not ( n11380 , n4593 );
or ( n11381 , n11379 , n11380 );
not ( n11382 , n3544 );
not ( n11383 , n3528 );
nand ( n11384 , n11382 , n11383 );
nand ( n11385 , n11381 , n11384 );
not ( n11386 , n11385 );
not ( n11387 , n11386 );
buf ( n11388 , n11387 );
nor ( n11389 , n4437 , n4594 );
not ( n11390 , n11389 );
nand ( n11391 , n4437 , n4594 );
nand ( n11392 , n11390 , n11391 , n11385 );
not ( n11393 , n11392 );
not ( n11394 , n11393 );
not ( n11395 , n11394 );
not ( n11396 , n11395 );
and ( n11397 , n11388 , n11396 );
not ( n11398 , n4678 );
not ( n11399 , n11398 );
not ( n11400 , n11399 );
nor ( n11401 , n11397 , n11400 );
xnor ( n11402 , n11378 , n11401 );
or ( n11403 , n11370 , n11402 );
or ( n11404 , n11401 , n11378 );
nand ( n11405 , n11403 , n11404 );
xor ( n11406 , n11315 , n11307 );
xor ( n11407 , n11405 , n11406 );
and ( n11408 , n11364 , n11407 );
and ( n11409 , n11406 , n11405 );
nor ( n11410 , n11408 , n11409 );
and ( n11411 , n11363 , n11354 );
and ( n11412 , n11295 , n11359 );
nor ( n11413 , n11411 , n11412 );
xnor ( n11414 , n11300 , n11319 );
xnor ( n11415 , n11413 , n11414 );
or ( n11416 , n11410 , n11415 );
or ( n11417 , n11413 , n11414 );
nand ( n11418 , n11416 , n11417 );
nand ( n11419 , n11332 , n11418 );
or ( n11420 , n11331 , n11419 );
nand ( n11421 , n11279 , n11330 );
nand ( n11422 , n11420 , n11421 );
buf ( n11423 , n11422 );
not ( n11424 , n11423 );
nand ( n11425 , n45 , n3103 );
not ( n11426 , n11097 );
and ( n11427 , n4375 , n11426 );
and ( n11428 , n11341 , n11293 );
nor ( n11429 , n11427 , n11428 );
xnor ( n11430 , n11425 , n11429 );
not ( n11431 , n4424 );
not ( n11432 , n11431 );
and ( n11433 , n11252 , n11432 );
and ( n11434 , n11375 , n11241 );
nor ( n11435 , n11433 , n11434 );
and ( n11436 , n11430 , n11435 );
not ( n11437 , n11430 );
not ( n11438 , n11435 );
and ( n11439 , n11437 , n11438 );
nor ( n11440 , n11436 , n11439 );
not ( n11441 , n46 );
nor ( n11442 , n11441 , n3196 );
buf ( n11443 , n11382 );
not ( n11444 , n11443 );
not ( n11445 , n11444 );
not ( n11446 , n11445 );
nand ( n11447 , n3126 , n11446 );
and ( n11448 , n4462 , n11447 );
not ( n11449 , n11448 );
not ( n11450 , n11449 );
not ( n11451 , n5076 );
nand ( n11452 , n11451 , n3692 );
not ( n11453 , n3852 );
nand ( n11454 , n11453 , n3518 );
not ( n11455 , n3544 );
not ( n11456 , n5076 );
or ( n11457 , n11455 , n11456 );
or ( n11458 , n3518 , n3547 );
nand ( n11459 , n11457 , n11458 );
and ( n11460 , n11452 , n11454 , n11459 );
not ( n11461 , n11460 );
not ( n11462 , n11461 );
not ( n11463 , n11462 );
not ( n11464 , n11463 );
not ( n11465 , n11464 );
not ( n11466 , n11465 );
and ( n11467 , n11450 , n11466 );
not ( n11468 , n11446 );
not ( n11469 , n11454 );
not ( n11470 , n11469 );
nand ( n11471 , n11470 , n11452 );
not ( n11472 , n11471 );
not ( n11473 , n11472 );
and ( n11474 , n11468 , n11473 );
nor ( n11475 , n11467 , n11474 );
not ( n11476 , n11475 );
and ( n11477 , n11442 , n11476 );
not ( n11478 , n11442 );
and ( n11479 , n11478 , n11475 );
nor ( n11480 , n11477 , n11479 );
not ( n11481 , n3287 );
xor ( n11482 , n11481 , n44 );
not ( n11483 , n11125 );
and ( n11484 , n11482 , n11483 );
and ( n11485 , n43 , n3136 );
and ( n11486 , n11344 , n3135 );
nor ( n11487 , n11485 , n11486 );
and ( n11488 , n11487 , n11137 );
nor ( n11489 , n11484 , n11488 );
not ( n11490 , n3419 );
not ( n11491 , n11490 );
not ( n11492 , n11394 );
and ( n11493 , n11491 , n11492 );
and ( n11494 , n37 , n11399 );
buf ( n11495 , n4437 );
not ( n11496 , n11495 );
and ( n11497 , n11110 , n11496 );
nor ( n11498 , n11494 , n11497 );
not ( n11499 , n11387 );
and ( n11500 , n11498 , n11499 );
nor ( n11501 , n11493 , n11500 );
not ( n11502 , n3314 );
and ( n11503 , n11502 , n42 );
not ( n11504 , n11502 );
and ( n11505 , n11504 , n3502 );
nor ( n11506 , n11503 , n11505 );
not ( n11507 , n11506 );
not ( n11508 , n11096 );
or ( n11509 , n11507 , n11508 );
not ( n11510 , n3314 );
and ( n11511 , n41 , n11510 );
not ( n11512 , n3313 );
and ( n11513 , n11220 , n11512 );
nor ( n11514 , n11511 , n11513 );
nand ( n11515 , n11514 , n11086 );
nand ( n11516 , n11509 , n11515 );
and ( n11517 , n11501 , n11516 );
not ( n11518 , n11501 );
not ( n11519 , n11516 );
and ( n11520 , n11518 , n11519 );
nor ( n11521 , n11517 , n11520 );
or ( n11522 , n11489 , n11521 );
or ( n11523 , n11519 , n11501 );
nand ( n11524 , n11522 , n11523 );
and ( n11525 , n11480 , n11524 );
and ( n11526 , n11442 , n11476 );
nor ( n11527 , n11525 , n11526 );
xnor ( n11528 , n11440 , n11527 );
and ( n11529 , n3194 , n44 );
not ( n11530 , n3194 );
not ( n11531 , n44 );
and ( n11532 , n11530 , n11531 );
nor ( n11533 , n11529 , n11532 );
not ( n11534 , n11533 );
not ( n11535 , n11152 );
and ( n11536 , n11534 , n11535 );
or ( n11537 , n45 , n3103 );
nand ( n11538 , n11537 , n11425 );
not ( n11539 , n11538 );
and ( n11540 , n11539 , n11157 );
nor ( n11541 , n11536 , n11540 );
or ( n11542 , n3502 , n11481 );
nand ( n11543 , n11542 , n4408 );
nand ( n11544 , n11543 , n11135 );
nand ( n11545 , n11487 , n11124 );
and ( n11546 , n11544 , n11545 );
not ( n11547 , n11431 );
not ( n11548 , n11240 );
and ( n11549 , n11547 , n11548 );
not ( n11550 , n4665 );
buf ( n11551 , n11550 );
and ( n11552 , n11551 , n11188 );
not ( n11553 , n11551 );
and ( n11554 , n11553 , n39 );
nor ( n11555 , n11552 , n11554 );
and ( n11556 , n11555 , n11250 );
nor ( n11557 , n11549 , n11556 );
xnor ( n11558 , n11546 , n11557 );
xor ( n11559 , n11541 , n11558 );
and ( n11560 , n47 , n3103 );
not ( n11561 , n11560 );
not ( n11562 , n11238 );
nand ( n11563 , n11555 , n11562 );
not ( n11564 , n11550 );
and ( n11565 , n3229 , n11564 );
and ( n11566 , n40 , n11550 );
nor ( n11567 , n11565 , n11566 );
not ( n11568 , n11567 );
nand ( n11569 , n11568 , n11248 );
and ( n11570 , n11563 , n11569 );
not ( n11571 , n11153 );
not ( n11572 , n3623 );
or ( n11573 , n11571 , n11572 );
or ( n11574 , n11538 , n11152 );
nand ( n11575 , n11573 , n11574 );
and ( n11576 , n11570 , n11575 );
not ( n11577 , n11570 );
not ( n11578 , n11575 );
and ( n11579 , n11577 , n11578 );
nor ( n11580 , n11576 , n11579 );
or ( n11581 , n11561 , n11580 );
or ( n11582 , n11570 , n11578 );
nand ( n11583 , n11581 , n11582 );
xor ( n11584 , n11559 , n11583 );
not ( n11585 , n11473 );
not ( n11586 , n11465 );
not ( n11587 , n11586 );
and ( n11588 , n11585 , n11587 );
not ( n11589 , n11468 );
nor ( n11590 , n11588 , n11589 );
not ( n11591 , n11396 );
and ( n11592 , n11591 , n11498 );
and ( n11593 , n3126 , n11400 );
nor ( n11594 , n11593 , n4679 );
not ( n11595 , n11388 );
and ( n11596 , n11594 , n11595 );
nor ( n11597 , n11592 , n11596 );
xnor ( n11598 , n11590 , n11597 );
and ( n11599 , n11514 , n11100 );
and ( n11600 , n4375 , n11090 );
nor ( n11601 , n11599 , n11600 );
xor ( n11602 , n11598 , n11601 );
and ( n11603 , n11584 , n11602 );
and ( n11604 , n11583 , n11559 );
nor ( n11605 , n11603 , n11604 );
or ( n11606 , n11528 , n11605 );
or ( n11607 , n11440 , n11527 );
nand ( n11608 , n11606 , n11607 );
not ( n11609 , n11608 );
or ( n11610 , n11438 , n11430 );
or ( n11611 , n11425 , n11429 );
nand ( n11612 , n11610 , n11611 );
xor ( n11613 , n11402 , n11370 );
xor ( n11614 , n11612 , n11613 );
xor ( n11615 , n11351 , n11333 );
and ( n11616 , n11594 , n11591 );
not ( n11617 , n11400 );
and ( n11618 , n11617 , n11595 );
nor ( n11619 , n11616 , n11618 );
not ( n11620 , n11533 );
not ( n11621 , n11154 );
and ( n11622 , n11620 , n11621 );
and ( n11623 , n11347 , n11165 );
nor ( n11624 , n11622 , n11623 );
not ( n11625 , n11543 );
not ( n11626 , n11124 );
or ( n11627 , n11625 , n11626 );
nand ( n11628 , n11367 , n11135 );
nand ( n11629 , n11627 , n11628 );
and ( n11630 , n11624 , n11629 );
not ( n11631 , n11624 );
not ( n11632 , n11629 );
and ( n11633 , n11631 , n11632 );
nor ( n11634 , n11630 , n11633 );
or ( n11635 , n11619 , n11634 );
or ( n11636 , n11624 , n11632 );
nand ( n11637 , n11635 , n11636 );
and ( n11638 , n11637 , n11438 );
not ( n11639 , n11637 );
and ( n11640 , n11639 , n11435 );
nor ( n11641 , n11638 , n11640 );
xor ( n11642 , n11615 , n11641 );
xnor ( n11643 , n11614 , n11642 );
xor ( n11644 , n11634 , n11619 );
or ( n11645 , n11541 , n11558 );
or ( n11646 , n11557 , n11546 );
nand ( n11647 , n11645 , n11646 );
or ( n11648 , n11601 , n11598 );
or ( n11649 , n11590 , n11597 );
nand ( n11650 , n11648 , n11649 );
xor ( n11651 , n11647 , n11650 );
and ( n11652 , n11644 , n11651 );
and ( n11653 , n11650 , n11647 );
nor ( n11654 , n11652 , n11653 );
xor ( n11655 , n11643 , n11654 );
not ( n11656 , n11655 );
or ( n11657 , n11609 , n11656 );
or ( n11658 , n11654 , n11643 );
nand ( n11659 , n11657 , n11658 );
xnor ( n11660 , n11407 , n11364 );
and ( n11661 , n11615 , n11641 );
and ( n11662 , n11438 , n11637 );
nor ( n11663 , n11661 , n11662 );
xnor ( n11664 , n11660 , n11663 );
and ( n11665 , n11614 , n11642 );
and ( n11666 , n11612 , n11613 );
nor ( n11667 , n11665 , n11666 );
xor ( n11668 , n11664 , n11667 );
nor ( n11669 , n11659 , n11668 );
not ( n11670 , n11669 );
xnor ( n11671 , n11655 , n11608 );
xor ( n11672 , n11561 , n11580 );
and ( n11673 , n45 , n11481 );
not ( n11674 , n45 );
and ( n11675 , n11674 , n11119 );
nor ( n11676 , n11673 , n11675 );
not ( n11677 , n11676 );
not ( n11678 , n11123 );
not ( n11679 , n11678 );
or ( n11680 , n11677 , n11679 );
not ( n11681 , n11134 );
nand ( n11682 , n11482 , n11681 );
nand ( n11683 , n11680 , n11682 );
not ( n11684 , n11683 );
not ( n11685 , n11490 );
not ( n11686 , n11388 );
and ( n11687 , n11685 , n11686 );
and ( n11688 , n11188 , n11496 );
not ( n11689 , n11188 );
and ( n11690 , n11689 , n11495 );
nor ( n11691 , n11688 , n11690 );
and ( n11692 , n11691 , n11395 );
nor ( n11693 , n11687 , n11692 );
xnor ( n11694 , n11684 , n11693 );
not ( n11695 , n47 );
and ( n11696 , n11695 , n3194 );
nor ( n11697 , n11696 , n11560 );
not ( n11698 , n11156 );
and ( n11699 , n11697 , n11698 );
and ( n11700 , n3623 , n11165 );
nor ( n11701 , n11699 , n11700 );
or ( n11702 , n11694 , n11701 );
or ( n11703 , n11693 , n11684 );
nand ( n11704 , n11702 , n11703 );
xor ( n11705 , n11672 , n11704 );
xor ( n11706 , n11521 , n11489 );
and ( n11707 , n11705 , n11706 );
and ( n11708 , n11704 , n11672 );
nor ( n11709 , n11707 , n11708 );
and ( n11710 , n43 , n11338 );
and ( n11711 , n11344 , n3314 );
nor ( n11712 , n11710 , n11711 );
and ( n11713 , n11712 , n11098 );
and ( n11714 , n11506 , n11088 );
nor ( n11715 , n11713 , n11714 );
nand ( n11716 , n48 , n3195 );
not ( n11717 , n11567 );
not ( n11718 , n11238 );
and ( n11719 , n11717 , n11718 );
and ( n11720 , n11550 , n11220 );
not ( n11721 , n11550 );
and ( n11722 , n11721 , n41 );
nor ( n11723 , n11720 , n11722 );
and ( n11724 , n11723 , n11248 );
nor ( n11725 , n11719 , n11724 );
xnor ( n11726 , n11716 , n11725 );
or ( n11727 , n11715 , n11726 );
or ( n11728 , n11716 , n11725 );
nand ( n11729 , n11727 , n11728 );
not ( n11730 , n3774 );
buf ( n11731 , n11730 );
not ( n11732 , n11731 );
not ( n11733 , n11732 );
not ( n11734 , n3774 );
not ( n11735 , n11453 );
nand ( n11736 , n11734 , n11735 );
not ( n11737 , n11736 );
not ( n11738 , n11737 );
not ( n11739 , n11738 );
not ( n11740 , n11739 );
and ( n11741 , n11733 , n11740 );
not ( n11742 , n11735 );
not ( n11743 , n11742 );
not ( n11744 , n11743 );
nor ( n11745 , n11741 , n11744 );
and ( n11746 , n11444 , n11110 );
not ( n11747 , n11444 );
and ( n11748 , n11747 , n37 );
nor ( n11749 , n11746 , n11748 );
and ( n11750 , n11749 , n11464 );
and ( n11751 , n11448 , n11473 );
nor ( n11752 , n11750 , n11751 );
nand ( n11753 , n11745 , n11752 );
and ( n11754 , n11753 , n11475 );
not ( n11755 , n11753 );
and ( n11756 , n11755 , n11476 );
nor ( n11757 , n11754 , n11756 );
and ( n11758 , n11729 , n11757 );
and ( n11759 , n11475 , n11753 );
nor ( n11760 , n11758 , n11759 );
xnor ( n11761 , n11524 , n11480 );
xnor ( n11762 , n11760 , n11761 );
or ( n11763 , n11709 , n11762 );
or ( n11764 , n11760 , n11761 );
nand ( n11765 , n11763 , n11764 );
xor ( n11766 , n11605 , n11528 );
xor ( n11767 , n11651 , n11644 );
xor ( n11768 , n11766 , n11767 );
and ( n11769 , n11765 , n11768 );
and ( n11770 , n11767 , n11766 );
nor ( n11771 , n11769 , n11770 );
or ( n11772 , n11671 , n11771 );
not ( n11773 , n11772 );
and ( n11774 , n11670 , n11773 );
nand ( n11775 , n11668 , n11659 );
not ( n11776 , n11775 );
nor ( n11777 , n11774 , n11776 );
xor ( n11778 , n11415 , n11410 );
or ( n11779 , n11667 , n11664 );
or ( n11780 , n11663 , n11660 );
nand ( n11781 , n11779 , n11780 );
nor ( n11782 , n11778 , n11781 );
or ( n11783 , n11777 , n11782 );
nand ( n11784 , n11778 , n11781 );
nand ( n11785 , n11783 , n11784 );
not ( n11786 , n11785 );
buf ( n11787 , n11669 );
nor ( n11788 , n11787 , n11782 );
xor ( n11789 , n11726 , n11715 );
xor ( n11790 , n11694 , n11701 );
or ( n11791 , n11745 , n11752 );
nand ( n11792 , n11791 , n11753 );
xor ( n11793 , n11790 , n11792 );
and ( n11794 , n11789 , n11793 );
and ( n11795 , n11792 , n11790 );
nor ( n11796 , n11794 , n11795 );
and ( n11797 , n3559 , n11155 );
and ( n11798 , n11697 , n11165 );
nor ( n11799 , n11797 , n11798 );
not ( n11800 , n11394 );
not ( n11801 , n3229 );
not ( n11802 , n4440 );
or ( n11803 , n11801 , n11802 );
or ( n11804 , n3229 , n4440 );
nand ( n11805 , n11803 , n11804 );
not ( n11806 , n11805 );
and ( n11807 , n11800 , n11806 );
not ( n11808 , n11387 );
and ( n11809 , n11808 , n11691 );
nor ( n11810 , n11807 , n11809 );
not ( n11811 , n3777 );
not ( n11812 , n11678 );
or ( n11813 , n11811 , n11812 );
not ( n11814 , n11134 );
nand ( n11815 , n11676 , n11814 );
nand ( n11816 , n11813 , n11815 );
xor ( n11817 , n11810 , n11816 );
or ( n11818 , n11799 , n11817 );
not ( n11819 , n11816 );
or ( n11820 , n11810 , n11819 );
nand ( n11821 , n11818 , n11820 );
not ( n11822 , n11737 );
not ( n11823 , n3854 );
or ( n11824 , n11822 , n11823 );
not ( n11825 , n3774 );
not ( n11826 , n11825 );
not ( n11827 , n11826 );
or ( n11828 , n11744 , n11827 );
nand ( n11829 , n11824 , n11828 );
not ( n11830 , n11829 );
not ( n11831 , n11749 );
not ( n11832 , n11831 );
not ( n11833 , n11472 );
and ( n11834 , n11832 , n11833 );
not ( n11835 , n11443 );
and ( n11836 , n11835 , n3096 );
not ( n11837 , n11835 );
and ( n11838 , n11837 , n38 );
nor ( n11839 , n11836 , n11838 );
not ( n11840 , n11463 );
and ( n11841 , n11839 , n11840 );
nor ( n11842 , n11834 , n11841 );
nor ( n11843 , n11830 , n11842 );
not ( n11844 , n11843 );
and ( n11845 , n4373 , n44 );
not ( n11846 , n4373 );
not ( n11847 , n44 );
and ( n11848 , n11846 , n11847 );
nor ( n11849 , n11845 , n11848 );
not ( n11850 , n11849 );
not ( n11851 , n11097 );
and ( n11852 , n11850 , n11851 );
not ( n11853 , n11087 );
and ( n11854 , n11712 , n11853 );
nor ( n11855 , n11852 , n11854 );
and ( n11856 , n11550 , n42 );
not ( n11857 , n11550 );
and ( n11858 , n11857 , n3502 );
nor ( n11859 , n11856 , n11858 );
not ( n11860 , n11859 );
not ( n11861 , n11860 );
not ( n11862 , n11248 );
or ( n11863 , n11861 , n11862 );
not ( n11864 , n11237 );
nand ( n11865 , n11723 , n11864 );
nand ( n11866 , n11863 , n11865 );
nand ( n11867 , n49 , n3106 );
xor ( n11868 , n11866 , n11867 );
or ( n11869 , n11855 , n11868 );
not ( n11870 , n11866 );
or ( n11871 , n11867 , n11870 );
nand ( n11872 , n11869 , n11871 );
not ( n11873 , n11872 );
not ( n11874 , n11873 );
or ( n11875 , n11844 , n11874 );
not ( n11876 , n11843 );
nand ( n11877 , n11876 , n11872 );
nand ( n11878 , n11875 , n11877 );
and ( n11879 , n11821 , n11878 );
not ( n11880 , n11873 );
and ( n11881 , n11843 , n11880 );
nor ( n11882 , n11879 , n11881 );
xnor ( n11883 , n11757 , n11729 );
xnor ( n11884 , n11882 , n11883 );
or ( n11885 , n11796 , n11884 );
or ( n11886 , n11883 , n11882 );
nand ( n11887 , n11885 , n11886 );
xor ( n11888 , n11709 , n11762 );
xor ( n11889 , n11584 , n11602 );
xor ( n11890 , n11888 , n11889 );
and ( n11891 , n11887 , n11890 );
and ( n11892 , n11889 , n11888 );
nor ( n11893 , n11891 , n11892 );
xnor ( n11894 , n11768 , n11765 );
nand ( n11895 , n11893 , n11894 );
xor ( n11896 , n11868 , n11855 );
not ( n11897 , n3777 );
not ( n11898 , n11897 );
not ( n11899 , n11136 );
and ( n11900 , n11898 , n11899 );
and ( n11901 , n47 , n11481 );
and ( n11902 , n11695 , n3287 );
nor ( n11903 , n11901 , n11902 );
and ( n11904 , n11903 , n11124 );
nor ( n11905 , n11900 , n11904 );
not ( n11906 , n11905 );
not ( n11907 , n11906 );
and ( n11908 , n45 , n3313 );
and ( n11909 , n11674 , n4373 );
nor ( n11910 , n11908 , n11909 );
not ( n11911 , n11910 );
not ( n11912 , n11096 );
or ( n11913 , n11911 , n11912 );
not ( n11914 , n11849 );
nand ( n11915 , n11914 , n11085 );
nand ( n11916 , n11913 , n11915 );
not ( n11917 , n11916 );
not ( n11918 , n11917 );
and ( n11919 , n11496 , n11220 );
not ( n11920 , n11496 );
and ( n11921 , n11920 , n41 );
nor ( n11922 , n11919 , n11921 );
not ( n11923 , n11392 );
buf ( n11924 , n11923 );
and ( n11925 , n11922 , n11924 );
not ( n11926 , n11386 );
nor ( n11927 , n11805 , n11926 );
nor ( n11928 , n11925 , n11927 );
not ( n11929 , n11928 );
not ( n11930 , n11929 );
or ( n11931 , n11918 , n11930 );
not ( n11932 , n11916 );
or ( n11933 , n11932 , n11929 );
nand ( n11934 , n11931 , n11933 );
not ( n11935 , n11934 );
or ( n11936 , n11907 , n11935 );
or ( n11937 , n11932 , n11928 );
nand ( n11938 , n11936 , n11937 );
xor ( n11939 , n11817 , n11799 );
xor ( n11940 , n11938 , n11939 );
and ( n11941 , n11896 , n11940 );
and ( n11942 , n11938 , n11939 );
nor ( n11943 , n11941 , n11942 );
not ( n11944 , n11829 );
not ( n11945 , n11842 );
and ( n11946 , n11944 , n11945 );
and ( n11947 , n11842 , n11829 );
nor ( n11948 , n11946 , n11947 );
not ( n11949 , n11948 );
and ( n11950 , n11551 , n11344 );
not ( n11951 , n11551 );
and ( n11952 , n11951 , n43 );
nor ( n11953 , n11950 , n11952 );
not ( n11954 , n11953 );
not ( n11955 , n11248 );
or ( n11956 , n11954 , n11955 );
or ( n11957 , n11859 , n11238 );
nand ( n11958 , n11956 , n11957 );
not ( n11959 , n11958 );
nand ( n11960 , n50 , n11309 );
not ( n11961 , n11960 );
and ( n11962 , n11188 , n11835 );
and ( n11963 , n39 , n4461 );
nor ( n11964 , n11962 , n11963 );
not ( n11965 , n11964 );
not ( n11966 , n11461 );
not ( n11967 , n11966 );
or ( n11968 , n11965 , n11967 );
nand ( n11969 , n11839 , n11471 );
nand ( n11970 , n11968 , n11969 );
not ( n11971 , n11970 );
or ( n11972 , n11961 , n11971 );
or ( n11973 , n11960 , n11970 );
nand ( n11974 , n11972 , n11973 );
not ( n11975 , n11974 );
or ( n11976 , n11959 , n11975 );
not ( n11977 , n11960 );
nand ( n11978 , n11977 , n11970 );
nand ( n11979 , n11976 , n11978 );
nand ( n11980 , n11949 , n11979 );
not ( n11981 , n11878 );
and ( n11982 , n11821 , n11981 );
not ( n11983 , n11821 );
and ( n11984 , n11983 , n11878 );
nor ( n11985 , n11982 , n11984 );
not ( n11986 , n11985 );
and ( n11987 , n11980 , n11986 );
not ( n11988 , n11980 );
and ( n11989 , n11988 , n11985 );
nor ( n11990 , n11987 , n11989 );
or ( n11991 , n11943 , n11990 );
or ( n11992 , n11980 , n11985 );
nand ( n11993 , n11991 , n11992 );
xor ( n11994 , n11705 , n11706 );
xor ( n11995 , n11993 , n11994 );
xor ( n11996 , n11796 , n11884 );
xnor ( n11997 , n11995 , n11996 );
xor ( n11998 , n11793 , n11789 );
not ( n11999 , n11735 );
and ( n12000 , n11999 , n11110 );
not ( n12001 , n11999 );
and ( n12002 , n12001 , n37 );
nor ( n12003 , n12000 , n12002 );
and ( n12004 , n11739 , n12003 );
and ( n12005 , n11732 , n3854 );
nor ( n12006 , n12004 , n12005 );
not ( n12007 , n12006 );
or ( n12008 , n49 , n3103 );
nand ( n12009 , n12008 , n11867 );
not ( n12010 , n12009 );
not ( n12011 , n11154 );
and ( n12012 , n12010 , n12011 );
and ( n12013 , n3559 , n11165 );
nor ( n12014 , n12012 , n12013 );
not ( n12015 , n12014 );
and ( n12016 , n12007 , n12015 );
or ( n12017 , n3229 , n11443 );
nand ( n12018 , n12017 , n3948 );
and ( n12019 , n12018 , n11464 );
and ( n12020 , n11964 , n11473 );
nor ( n12021 , n12019 , n12020 );
nand ( n12022 , n11826 , n12003 );
and ( n12023 , n3096 , n11999 );
not ( n12024 , n3096 );
not ( n12025 , n11742 );
and ( n12026 , n12024 , n12025 );
nor ( n12027 , n12023 , n12026 );
nand ( n12028 , n11737 , n12027 );
and ( n12029 , n12022 , n12028 );
nand ( n12030 , n51 , n3193 );
xnor ( n12031 , n12029 , n12030 );
or ( n12032 , n12021 , n12031 );
or ( n12033 , n12030 , n12029 );
nand ( n12034 , n12032 , n12033 );
xor ( n12035 , n12014 , n12006 );
and ( n12036 , n12034 , n12035 );
nor ( n12037 , n12016 , n12036 );
xor ( n12038 , n11948 , n11979 );
xnor ( n12039 , n12037 , n12038 );
xnor ( n12040 , n11974 , n11958 );
not ( n12041 , n12040 );
and ( n12042 , n11496 , n42 );
not ( n12043 , n11496 );
and ( n12044 , n12043 , n3502 );
nor ( n12045 , n12042 , n12044 );
not ( n12046 , n12045 );
and ( n12047 , n12046 , n11395 );
and ( n12048 , n11922 , n11499 );
nor ( n12049 , n12047 , n12048 );
not ( n12050 , n12049 );
not ( n12051 , n12050 );
not ( n12052 , n4173 );
not ( n12053 , n11096 );
or ( n12054 , n12052 , n12053 );
not ( n12055 , n11084 );
nand ( n12056 , n11910 , n12055 );
nand ( n12057 , n12054 , n12056 );
not ( n12058 , n3911 );
not ( n12059 , n11248 );
or ( n12060 , n12058 , n12059 );
not ( n12061 , n11238 );
nand ( n12062 , n11953 , n12061 );
nand ( n12063 , n12060 , n12062 );
xor ( n12064 , n12057 , n12063 );
not ( n12065 , n12064 );
or ( n12066 , n12051 , n12065 );
nand ( n12067 , n12057 , n12063 );
nand ( n12068 , n12066 , n12067 );
not ( n12069 , n11906 );
not ( n12070 , n11934 );
not ( n12071 , n12070 );
or ( n12072 , n12069 , n12071 );
nand ( n12073 , n11905 , n11934 );
nand ( n12074 , n12072 , n12073 );
not ( n12075 , n12074 );
and ( n12076 , n12068 , n12075 );
not ( n12077 , n12068 );
and ( n12078 , n12077 , n12074 );
nor ( n12079 , n12076 , n12078 );
not ( n12080 , n12079 );
and ( n12081 , n12041 , n12080 );
and ( n12082 , n12068 , n12074 );
nor ( n12083 , n12081 , n12082 );
or ( n12084 , n12039 , n12083 );
or ( n12085 , n12037 , n12038 );
nand ( n12086 , n12084 , n12085 );
xor ( n12087 , n11998 , n12086 );
xor ( n12088 , n11943 , n11990 );
and ( n12089 , n12087 , n12088 );
and ( n12090 , n11998 , n12086 );
nor ( n12091 , n12089 , n12090 );
nand ( n12092 , n11997 , n12091 );
xnor ( n12093 , n12087 , n12088 );
xnor ( n12094 , n12034 , n12035 );
not ( n12095 , n12009 );
not ( n12096 , n11152 );
and ( n12097 , n12095 , n12096 );
and ( n12098 , n4039 , n11153 );
nor ( n12099 , n12097 , n12098 );
not ( n12100 , n12099 );
not ( n12101 , n12100 );
not ( n12102 , n12101 );
not ( n12103 , n4019 );
not ( n12104 , n11678 );
or ( n12105 , n12103 , n12104 );
nand ( n12106 , n11903 , n11681 );
nand ( n12107 , n12105 , n12106 );
not ( n12108 , n12107 );
not ( n12109 , n12108 );
and ( n12110 , n12102 , n12109 );
not ( n12111 , n51 );
nand ( n12112 , n12111 , n3287 );
and ( n12113 , n3160 , n12112 );
not ( n12114 , n51 );
nor ( n12115 , n12114 , n11119 );
nor ( n12116 , n12113 , n12115 , n3104 );
not ( n12117 , n11738 );
not ( n12118 , n12117 );
and ( n12119 , n11999 , n11188 );
not ( n12120 , n11999 );
and ( n12121 , n12120 , n39 );
nor ( n12122 , n12119 , n12121 );
not ( n12123 , n12122 );
or ( n12124 , n12118 , n12123 );
nand ( n12125 , n11732 , n12027 );
nand ( n12126 , n12124 , n12125 );
and ( n12127 , n12116 , n12126 );
not ( n12128 , n12100 );
not ( n12129 , n12108 );
or ( n12130 , n12128 , n12129 );
nand ( n12131 , n12107 , n12101 );
nand ( n12132 , n12130 , n12131 );
and ( n12133 , n12127 , n12132 );
nor ( n12134 , n12110 , n12133 );
xnor ( n12135 , n12094 , n12134 );
xor ( n12136 , n12031 , n12021 );
and ( n12137 , n4039 , n11165 );
not ( n12138 , n51 );
and ( n12139 , n12138 , n3194 );
not ( n12140 , n12030 );
nor ( n12141 , n12139 , n12140 , n11154 );
nor ( n12142 , n12137 , n12141 );
not ( n12143 , n12045 );
not ( n12144 , n11387 );
and ( n12145 , n12143 , n12144 );
and ( n12146 , n43 , n11495 );
and ( n12147 , n11344 , n11398 );
nor ( n12148 , n12146 , n12147 );
and ( n12149 , n12148 , n11924 );
nor ( n12150 , n12145 , n12149 );
and ( n12151 , n49 , n11481 );
not ( n12152 , n49 );
and ( n12153 , n12152 , n11119 );
nor ( n12154 , n12151 , n12153 );
not ( n12155 , n12154 );
not ( n12156 , n11678 );
or ( n12157 , n12155 , n12156 );
not ( n12158 , n4019 );
not ( n12159 , n11681 );
or ( n12160 , n12158 , n12159 );
nand ( n12161 , n12157 , n12160 );
and ( n12162 , n12150 , n12161 );
not ( n12163 , n12150 );
not ( n12164 , n12161 );
and ( n12165 , n12163 , n12164 );
nor ( n12166 , n12162 , n12165 );
or ( n12167 , n12142 , n12166 );
or ( n12168 , n12150 , n12164 );
nand ( n12169 , n12167 , n12168 );
not ( n12170 , n4173 );
not ( n12171 , n12170 );
not ( n12172 , n11087 );
and ( n12173 , n12171 , n12172 );
and ( n12174 , n4373 , n11695 );
not ( n12175 , n4373 );
and ( n12176 , n12175 , n47 );
nor ( n12177 , n12174 , n12176 );
and ( n12178 , n12177 , n11098 );
nor ( n12179 , n12173 , n12178 );
nand ( n12180 , n12018 , n11471 );
and ( n12181 , n11444 , n11220 );
not ( n12182 , n11444 );
and ( n12183 , n12182 , n41 );
nor ( n12184 , n12181 , n12183 );
nand ( n12185 , n12184 , n11966 );
and ( n12186 , n12180 , n12185 );
and ( n12187 , n11551 , n11674 );
not ( n12188 , n11551 );
and ( n12189 , n12188 , n45 );
nor ( n12190 , n12187 , n12189 );
not ( n12191 , n12190 );
not ( n12192 , n11248 );
or ( n12193 , n12191 , n12192 );
not ( n12194 , n3911 );
or ( n12195 , n12194 , n11238 );
nand ( n12196 , n12193 , n12195 );
and ( n12197 , n12186 , n12196 );
not ( n12198 , n12186 );
not ( n12199 , n12196 );
and ( n12200 , n12198 , n12199 );
nor ( n12201 , n12197 , n12200 );
or ( n12202 , n12179 , n12201 );
or ( n12203 , n12186 , n12199 );
nand ( n12204 , n12202 , n12203 );
xor ( n12205 , n12169 , n12204 );
and ( n12206 , n12136 , n12205 );
and ( n12207 , n12204 , n12169 );
nor ( n12208 , n12206 , n12207 );
or ( n12209 , n12135 , n12208 );
or ( n12210 , n12134 , n12094 );
nand ( n12211 , n12209 , n12210 );
xor ( n12212 , n12039 , n12083 );
xor ( n12213 , n11940 , n11896 );
xor ( n12214 , n12212 , n12213 );
and ( n12215 , n12211 , n12214 );
and ( n12216 , n12213 , n12212 );
nor ( n12217 , n12215 , n12216 );
nor ( n12218 , n12093 , n12217 );
and ( n12219 , n12092 , n12218 );
nor ( n12220 , n11997 , n12091 );
nor ( n12221 , n12219 , n12220 );
not ( n12222 , n12221 );
and ( n12223 , n11996 , n11995 );
and ( n12224 , n11994 , n11993 );
nor ( n12225 , n12223 , n12224 );
xnor ( n12226 , n11890 , n11887 );
nand ( n12227 , n12225 , n12226 );
nand ( n12228 , n12222 , n12227 );
nor ( n12229 , n12225 , n12226 );
not ( n12230 , n12229 );
nand ( n12231 , n12228 , n12230 );
and ( n12232 , n11895 , n12231 );
xor ( n12233 , n12214 , n12211 );
xor ( n12234 , n12135 , n12208 );
not ( n12235 , n11249 );
buf ( n12236 , n4856 );
buf ( n12237 , n12236 );
and ( n12238 , n12235 , n12237 );
and ( n12239 , n12190 , n11239 );
nor ( n12240 , n12238 , n12239 );
not ( n12241 , n12240 );
not ( n12242 , n12241 );
and ( n12243 , n51 , n11165 );
not ( n12244 , n42 );
not ( n12245 , n11835 );
or ( n12246 , n12244 , n12245 );
nand ( n12247 , n12246 , n4833 );
not ( n12248 , n12247 );
not ( n12249 , n11966 );
or ( n12250 , n12248 , n12249 );
nand ( n12251 , n12184 , n11471 );
nand ( n12252 , n12250 , n12251 );
xor ( n12253 , n12243 , n12252 );
not ( n12254 , n12253 );
or ( n12255 , n12242 , n12254 );
nand ( n12256 , n12243 , n12252 );
nand ( n12257 , n12255 , n12256 );
xor ( n12258 , n12116 , n12126 );
xor ( n12259 , n12257 , n12258 );
not ( n12260 , n11678 );
not ( n12261 , n12260 );
xor ( n12262 , n11119 , n50 );
not ( n12263 , n12262 );
and ( n12264 , n12261 , n12263 );
and ( n12265 , n12154 , n11135 );
nor ( n12266 , n12264 , n12265 );
not ( n12267 , n12266 );
not ( n12268 , n12267 );
not ( n12269 , n11738 );
not ( n12270 , n5013 );
not ( n12271 , n12270 );
and ( n12272 , n12269 , n12271 );
and ( n12273 , n11732 , n12122 );
nor ( n12274 , n12272 , n12273 );
not ( n12275 , n12274 );
xor ( n12276 , n3272 , n48 );
not ( n12277 , n12276 );
not ( n12278 , n11096 );
or ( n12279 , n12277 , n12278 );
not ( n12280 , n11084 );
nand ( n12281 , n12177 , n12280 );
nand ( n12282 , n12279 , n12281 );
not ( n12283 , n12282 );
and ( n12284 , n12275 , n12283 );
and ( n12285 , n12274 , n12282 );
nor ( n12286 , n12284 , n12285 );
or ( n12287 , n12268 , n12286 );
not ( n12288 , n12282 );
or ( n12289 , n12274 , n12288 );
nand ( n12290 , n12287 , n12289 );
and ( n12291 , n12259 , n12290 );
and ( n12292 , n12258 , n12257 );
nor ( n12293 , n12291 , n12292 );
and ( n12294 , n12064 , n12049 );
not ( n12295 , n12064 );
and ( n12296 , n12295 , n12050 );
nor ( n12297 , n12294 , n12296 );
not ( n12298 , n12127 );
and ( n12299 , n12132 , n12298 );
not ( n12300 , n12132 );
and ( n12301 , n12300 , n12127 );
nor ( n12302 , n12299 , n12301 );
xnor ( n12303 , n12297 , n12302 );
or ( n12304 , n12293 , n12303 );
or ( n12305 , n12302 , n12297 );
nand ( n12306 , n12304 , n12305 );
xor ( n12307 , n12079 , n12040 );
xor ( n12308 , n12306 , n12307 );
and ( n12309 , n12234 , n12308 );
and ( n12310 , n12307 , n12306 );
nor ( n12311 , n12309 , n12310 );
not ( n12312 , n12311 );
and ( n12313 , n12233 , n12312 );
not ( n12314 , n12313 );
nand ( n12315 , n51 , n11114 );
not ( n12316 , n11116 );
and ( n12317 , n12315 , n3136 , n12316 );
and ( n12318 , n11444 , n11344 );
not ( n12319 , n11444 );
and ( n12320 , n12319 , n43 );
nor ( n12321 , n12318 , n12320 );
not ( n12322 , n12321 );
not ( n12323 , n11966 );
or ( n12324 , n12322 , n12323 );
nand ( n12325 , n12247 , n11471 );
nand ( n12326 , n12324 , n12325 );
and ( n12327 , n12317 , n12326 );
not ( n12328 , n12148 );
not ( n12329 , n11499 );
or ( n12330 , n12328 , n12329 );
xor ( n12331 , n11398 , n44 );
or ( n12332 , n12331 , n11394 );
nand ( n12333 , n12330 , n12332 );
xor ( n12334 , n12327 , n12333 );
not ( n12335 , n11739 );
and ( n12336 , n41 , n11743 );
not ( n12337 , n3693 );
and ( n12338 , n11220 , n12337 );
nor ( n12339 , n12336 , n12338 );
not ( n12340 , n12339 );
or ( n12341 , n12335 , n12340 );
or ( n12342 , n11733 , n12270 );
nand ( n12343 , n12341 , n12342 );
not ( n12344 , n12343 );
and ( n12345 , n3272 , n49 );
not ( n12346 , n3272 );
and ( n12347 , n12346 , n12152 );
nor ( n12348 , n12345 , n12347 );
not ( n12349 , n12348 );
not ( n12350 , n11096 );
or ( n12351 , n12349 , n12350 );
nand ( n12352 , n12276 , n12055 );
nand ( n12353 , n12351 , n12352 );
not ( n12354 , n12353 );
and ( n12355 , n47 , n11256 );
and ( n12356 , n11695 , n11255 );
nor ( n12357 , n12355 , n12356 );
not ( n12358 , n12357 );
not ( n12359 , n11244 );
nand ( n12360 , n12359 , n11246 , n11237 );
not ( n12361 , n12360 );
not ( n12362 , n12361 );
or ( n12363 , n12358 , n12362 );
nand ( n12364 , n12236 , n11864 );
nand ( n12365 , n12363 , n12364 );
not ( n12366 , n12365 );
not ( n12367 , n12366 );
or ( n12368 , n12354 , n12367 );
or ( n12369 , n12353 , n12366 );
nand ( n12370 , n12368 , n12369 );
not ( n12371 , n12370 );
or ( n12372 , n12344 , n12371 );
not ( n12373 , n12353 );
or ( n12374 , n12373 , n12366 );
nand ( n12375 , n12372 , n12374 );
and ( n12376 , n12334 , n12375 );
and ( n12377 , n12333 , n12327 );
nor ( n12378 , n12376 , n12377 );
xnor ( n12379 , n12179 , n12201 );
xnor ( n12380 , n12142 , n12166 );
xnor ( n12381 , n12379 , n12380 );
or ( n12382 , n12378 , n12381 );
or ( n12383 , n12379 , n12380 );
nand ( n12384 , n12382 , n12383 );
xor ( n12385 , n12293 , n12303 );
xor ( n12386 , n12136 , n12205 );
xor ( n12387 , n12385 , n12386 );
xor ( n12388 , n12384 , n12387 );
not ( n12389 , n12388 );
xor ( n12390 , n12381 , n12378 );
xor ( n12391 , n12259 , n12290 );
and ( n12392 , n45 , n11399 );
and ( n12393 , n11496 , n11674 );
nor ( n12394 , n12392 , n12393 );
and ( n12395 , n12394 , n11923 );
not ( n12396 , n12331 );
and ( n12397 , n12396 , n11808 );
nor ( n12398 , n12395 , n12397 );
not ( n12399 , n12398 );
not ( n12400 , n12115 );
and ( n12401 , n12112 , n12400 , n11124 );
nor ( n12402 , n12262 , n11134 );
nor ( n12403 , n12401 , n12402 );
not ( n12404 , n12403 );
and ( n12405 , n12399 , n12404 );
not ( n12406 , n12317 );
not ( n12407 , n12326 );
not ( n12408 , n12407 );
or ( n12409 , n12406 , n12408 );
or ( n12410 , n12317 , n12407 );
nand ( n12411 , n12409 , n12410 );
xor ( n12412 , n12398 , n12403 );
and ( n12413 , n12411 , n12412 );
nor ( n12414 , n12405 , n12413 );
and ( n12415 , n12253 , n12240 );
not ( n12416 , n12253 );
and ( n12417 , n12416 , n12241 );
nor ( n12418 , n12415 , n12417 );
and ( n12419 , n12286 , n12267 );
not ( n12420 , n12286 );
and ( n12421 , n12420 , n12266 );
nor ( n12422 , n12419 , n12421 );
xnor ( n12423 , n12418 , n12422 );
or ( n12424 , n12414 , n12423 );
or ( n12425 , n12418 , n12422 );
nand ( n12426 , n12424 , n12425 );
xor ( n12427 , n12391 , n12426 );
and ( n12428 , n12390 , n12427 );
and ( n12429 , n12391 , n12426 );
nor ( n12430 , n12428 , n12429 );
nand ( n12431 , n12389 , n12430 );
not ( n12432 , n12431 );
not ( n12433 , n5406 );
not ( n12434 , n12433 );
not ( n12435 , n11388 );
and ( n12436 , n12434 , n12435 );
and ( n12437 , n4678 , n47 );
not ( n12438 , n4678 );
and ( n12439 , n12438 , n11695 );
nor ( n12440 , n12437 , n12439 );
and ( n12441 , n11395 , n12440 );
nor ( n12442 , n12436 , n12441 );
nand ( n12443 , n51 , n11082 );
and ( n12444 , n12443 , n3315 , n11077 );
not ( n12445 , n12444 );
and ( n12446 , n45 , n11445 );
not ( n12447 , n45 );
and ( n12448 , n12447 , n11835 );
nor ( n12449 , n12446 , n12448 );
not ( n12450 , n12449 );
not ( n12451 , n11462 );
or ( n12452 , n12450 , n12451 );
xor ( n12453 , n11443 , n44 );
nand ( n12454 , n12453 , n11471 );
nand ( n12455 , n12452 , n12454 );
not ( n12456 , n12455 );
not ( n12457 , n12456 );
and ( n12458 , n12445 , n12457 );
and ( n12459 , n12444 , n12456 );
nor ( n12460 , n12458 , n12459 );
not ( n12461 , n12460 );
and ( n12462 , n12442 , n12461 );
not ( n12463 , n12442 );
and ( n12464 , n12463 , n12460 );
nor ( n12465 , n12462 , n12464 );
nand ( n12466 , n51 , n12055 );
not ( n12467 , n12466 );
not ( n12468 , n11826 );
not ( n12469 , n43 );
not ( n12470 , n3693 );
not ( n12471 , n12470 );
or ( n12472 , n12469 , n12471 );
or ( n12473 , n43 , n12337 );
nand ( n12474 , n12472 , n12473 );
not ( n12475 , n12474 );
or ( n12476 , n12468 , n12475 );
nand ( n12477 , n11737 , n5585 );
nand ( n12478 , n12476 , n12477 );
not ( n12479 , n12478 );
and ( n12480 , n12467 , n12479 );
and ( n12481 , n12466 , n12478 );
nor ( n12482 , n12480 , n12481 );
not ( n12483 , n12482 );
not ( n12484 , n4666 );
and ( n12485 , n12484 , n12152 );
and ( n12486 , n11255 , n49 );
nor ( n12487 , n12485 , n12486 );
not ( n12488 , n12487 );
not ( n12489 , n11238 );
and ( n12490 , n12488 , n12489 );
and ( n12491 , n12361 , n5564 );
nor ( n12492 , n12490 , n12491 );
not ( n12493 , n12492 );
and ( n12494 , n12483 , n12493 );
not ( n12495 , n12466 );
and ( n12496 , n12495 , n12478 );
nor ( n12497 , n12494 , n12496 );
not ( n12498 , n12497 );
and ( n12499 , n12465 , n12498 );
not ( n12500 , n12465 );
and ( n12501 , n12500 , n12497 );
nor ( n12502 , n12499 , n12501 );
not ( n12503 , n12502 );
not ( n12504 , n12474 );
or ( n12505 , n11740 , n12504 );
not ( n12506 , n5209 );
or ( n12507 , n11733 , n12506 );
nand ( n12508 , n12505 , n12507 );
not ( n12509 , n12487 );
not ( n12510 , n12360 );
and ( n12511 , n12509 , n12510 );
and ( n12512 , n5239 , n11864 );
nor ( n12513 , n12511 , n12512 );
not ( n12514 , n12513 );
not ( n12515 , n5197 );
not ( n12516 , n11086 );
or ( n12517 , n12515 , n12516 );
not ( n12518 , n51 );
nand ( n12519 , n12518 , n3314 );
nand ( n12520 , n51 , n11338 );
nand ( n12521 , n12519 , n12520 , n11096 );
nand ( n12522 , n12517 , n12521 );
not ( n12523 , n12522 );
or ( n12524 , n12514 , n12523 );
or ( n12525 , n12513 , n12522 );
nand ( n12526 , n12524 , n12525 );
not ( n12527 , n12526 );
and ( n12528 , n12508 , n12527 );
not ( n12529 , n12508 );
and ( n12530 , n12529 , n12526 );
or ( n12531 , n12528 , n12530 );
not ( n12532 , n4440 );
nand ( n12533 , n51 , n12532 );
not ( n12534 , n51 );
nand ( n12535 , n12534 , n4440 );
nand ( n12536 , n6399 , n12535 );
and ( n12537 , n12533 , n11257 , n12536 );
not ( n12538 , n3692 );
and ( n12539 , n11674 , n12538 );
not ( n12540 , n11674 );
and ( n12541 , n12540 , n3693 );
nor ( n12542 , n12539 , n12541 );
not ( n12543 , n12542 );
or ( n12544 , n11738 , n12543 );
not ( n12545 , n5585 );
or ( n12546 , n11731 , n12545 );
nand ( n12547 , n12544 , n12546 );
nand ( n12548 , n12537 , n12547 );
not ( n12549 , n12548 );
xor ( n12550 , n11443 , n46 );
not ( n12551 , n12550 );
not ( n12552 , n11966 );
or ( n12553 , n12551 , n12552 );
nand ( n12554 , n12449 , n11471 );
nand ( n12555 , n12553 , n12554 );
not ( n12556 , n5704 );
not ( n12557 , n11923 );
or ( n12558 , n12556 , n12557 );
nand ( n12559 , n12440 , n11386 );
nand ( n12560 , n12558 , n12559 );
not ( n12561 , n12560 );
and ( n12562 , n12555 , n12561 );
not ( n12563 , n12555 );
and ( n12564 , n12563 , n12560 );
nor ( n12565 , n12562 , n12564 );
not ( n12566 , n12565 );
and ( n12567 , n12549 , n12566 );
and ( n12568 , n12555 , n12560 );
nor ( n12569 , n12567 , n12568 );
and ( n12570 , n12531 , n12569 );
not ( n12571 , n12531 );
not ( n12572 , n12569 );
and ( n12573 , n12571 , n12572 );
nor ( n12574 , n12570 , n12573 );
not ( n12575 , n12574 );
and ( n12576 , n12503 , n12575 );
and ( n12577 , n12572 , n12531 );
nor ( n12578 , n12576 , n12577 );
not ( n12579 , n12513 );
nand ( n12580 , n12579 , n12522 );
nand ( n12581 , n12508 , n12526 );
and ( n12582 , n12580 , n12581 );
nand ( n12583 , n12444 , n12455 );
not ( n12584 , n12583 );
and ( n12585 , n12582 , n12584 );
not ( n12586 , n12582 );
and ( n12587 , n12586 , n12583 );
nor ( n12588 , n12585 , n12587 );
not ( n12589 , n12453 );
not ( n12590 , n11462 );
or ( n12591 , n12589 , n12590 );
nand ( n12592 , n12321 , n11471 );
nand ( n12593 , n12591 , n12592 );
and ( n12594 , n51 , n11117 );
and ( n12595 , n12593 , n12594 );
not ( n12596 , n12593 );
not ( n12597 , n12594 );
and ( n12598 , n12596 , n12597 );
nor ( n12599 , n12595 , n12598 );
not ( n12600 , n5239 );
not ( n12601 , n12361 );
or ( n12602 , n12600 , n12601 );
nand ( n12603 , n12357 , n11864 );
nand ( n12604 , n12602 , n12603 );
xnor ( n12605 , n12599 , n12604 );
and ( n12606 , n12588 , n12605 );
not ( n12607 , n12588 );
not ( n12608 , n12605 );
and ( n12609 , n12607 , n12608 );
or ( n12610 , n12606 , n12609 );
or ( n12611 , n12497 , n12465 );
not ( n12612 , n12461 );
or ( n12613 , n12442 , n12612 );
nand ( n12614 , n12611 , n12613 );
not ( n12615 , n11738 );
not ( n12616 , n12506 );
and ( n12617 , n12615 , n12616 );
not ( n12618 , n11731 );
and ( n12619 , n12618 , n12339 );
nor ( n12620 , n12617 , n12619 );
not ( n12621 , n12620 );
not ( n12622 , n5197 );
not ( n12623 , n11096 );
or ( n12624 , n12622 , n12623 );
nand ( n12625 , n12348 , n12280 );
nand ( n12626 , n12624 , n12625 );
not ( n12627 , n12626 );
or ( n12628 , n12621 , n12627 );
or ( n12629 , n12620 , n12626 );
nand ( n12630 , n12628 , n12629 );
not ( n12631 , n5406 );
not ( n12632 , n11924 );
or ( n12633 , n12631 , n12632 );
nand ( n12634 , n12394 , n11499 );
nand ( n12635 , n12633 , n12634 );
buf ( n12636 , n12635 );
xor ( n12637 , n12630 , n12636 );
not ( n12638 , n12637 );
and ( n12639 , n12614 , n12638 );
not ( n12640 , n12614 );
and ( n12641 , n12640 , n12637 );
nor ( n12642 , n12639 , n12641 );
not ( n12643 , n12642 );
and ( n12644 , n12610 , n12643 );
not ( n12645 , n12610 );
and ( n12646 , n12645 , n12642 );
nor ( n12647 , n12644 , n12646 );
or ( n12648 , n12578 , n12647 );
xor ( n12649 , n12578 , n12647 );
not ( n12650 , n11388 );
not ( n12651 , n5704 );
not ( n12652 , n12651 );
and ( n12653 , n12650 , n12652 );
and ( n12654 , n49 , n11495 );
not ( n12655 , n49 );
and ( n12656 , n12655 , n11398 );
nor ( n12657 , n12654 , n12656 );
and ( n12658 , n12657 , n11924 );
nor ( n12659 , n12653 , n12658 );
not ( n12660 , n12659 );
not ( n12661 , n12660 );
not ( n12662 , n4460 );
and ( n12663 , n47 , n12662 );
not ( n12664 , n47 );
and ( n12665 , n12664 , n4461 );
nor ( n12666 , n12663 , n12665 );
not ( n12667 , n12666 );
not ( n12668 , n12667 );
not ( n12669 , n11460 );
or ( n12670 , n12668 , n12669 );
nand ( n12671 , n11454 , n11452 );
nand ( n12672 , n12550 , n12671 );
nand ( n12673 , n12670 , n12672 );
not ( n12674 , n5564 );
not ( n12675 , n11864 );
or ( n12676 , n12674 , n12675 );
not ( n12677 , n51 );
nand ( n12678 , n12677 , n11551 );
nand ( n12679 , n51 , n11564 );
not ( n12680 , n12360 );
nand ( n12681 , n12678 , n12679 , n12680 );
nand ( n12682 , n12676 , n12681 );
xor ( n12683 , n12673 , n12682 );
not ( n12684 , n12683 );
or ( n12685 , n12661 , n12684 );
nand ( n12686 , n12673 , n12682 );
nand ( n12687 , n12685 , n12686 );
not ( n12688 , n12687 );
not ( n12689 , n12492 );
and ( n12690 , n12482 , n12689 );
not ( n12691 , n12482 );
and ( n12692 , n12691 , n12492 );
nor ( n12693 , n12690 , n12692 );
not ( n12694 , n12693 );
and ( n12695 , n12688 , n12694 );
and ( n12696 , n12693 , n12687 );
nor ( n12697 , n12695 , n12696 );
not ( n12698 , n12697 );
xnor ( n12699 , n12548 , n12565 );
not ( n12700 , n12699 );
and ( n12701 , n12698 , n12700 );
not ( n12702 , n12693 );
and ( n12703 , n12702 , n12687 );
nor ( n12704 , n12701 , n12703 );
xnor ( n12705 , n12502 , n12574 );
xor ( n12706 , n12704 , n12705 );
not ( n12707 , n12706 );
not ( n12708 , n48 );
and ( n12709 , n12708 , n11835 );
not ( n12710 , n12708 );
and ( n12711 , n12710 , n4461 );
nor ( n12712 , n12709 , n12711 );
not ( n12713 , n12712 );
not ( n12714 , n11966 );
or ( n12715 , n12713 , n12714 );
or ( n12716 , n11472 , n12666 );
nand ( n12717 , n12715 , n12716 );
not ( n12718 , n12717 );
not ( n12719 , n11737 );
buf ( n12720 , n5898 );
not ( n12721 , n12720 );
or ( n12722 , n12719 , n12721 );
nand ( n12723 , n11826 , n12542 );
nand ( n12724 , n12722 , n12723 );
not ( n12725 , n11237 );
and ( n12726 , n12725 , n51 );
xor ( n12727 , n12724 , n12726 );
not ( n12728 , n12727 );
or ( n12729 , n12718 , n12728 );
nand ( n12730 , n12726 , n12724 );
nand ( n12731 , n12729 , n12730 );
not ( n12732 , n12537 );
and ( n12733 , n12547 , n12732 );
not ( n12734 , n12547 );
and ( n12735 , n12734 , n12537 );
nor ( n12736 , n12733 , n12735 );
not ( n12737 , n12736 );
and ( n12738 , n12731 , n12737 );
not ( n12739 , n12731 );
and ( n12740 , n12739 , n12736 );
nor ( n12741 , n12738 , n12740 );
not ( n12742 , n12741 );
not ( n12743 , n12659 );
not ( n12744 , n12683 );
and ( n12745 , n12743 , n12744 );
and ( n12746 , n12659 , n12683 );
nor ( n12747 , n12745 , n12746 );
or ( n12748 , n12742 , n12747 );
not ( n12749 , n12731 );
or ( n12750 , n12736 , n12749 );
nand ( n12751 , n12748 , n12750 );
not ( n12752 , n12751 );
xnor ( n12753 , n12697 , n12699 );
nand ( n12754 , n12752 , n12753 );
not ( n12755 , n12754 );
nand ( n12756 , n51 , n11443 );
not ( n12757 , n51 );
nand ( n12758 , n12757 , n12662 );
nand ( n12759 , n4594 , n12758 );
and ( n12760 , n12756 , n11399 , n12759 );
not ( n12761 , n11826 );
not ( n12762 , n12720 );
or ( n12763 , n12761 , n12762 );
and ( n12764 , n11695 , n12538 );
not ( n12765 , n11695 );
and ( n12766 , n12765 , n3693 );
nor ( n12767 , n12764 , n12766 );
nand ( n12768 , n11737 , n12767 );
nand ( n12769 , n12763 , n12768 );
nand ( n12770 , n12760 , n12769 );
and ( n12771 , n4678 , n50 );
not ( n12772 , n4678 );
not ( n12773 , n50 );
and ( n12774 , n12772 , n12773 );
nor ( n12775 , n12771 , n12774 );
and ( n12776 , n12775 , n11923 );
and ( n12777 , n12657 , n11386 );
nor ( n12778 , n12776 , n12777 );
not ( n12779 , n12778 );
and ( n12780 , n12770 , n12779 );
not ( n12781 , n12770 );
and ( n12782 , n12781 , n12778 );
nor ( n12783 , n12780 , n12782 );
xor ( n12784 , n12727 , n12717 );
not ( n12785 , n12784 );
or ( n12786 , n12783 , n12785 );
or ( n12787 , n12770 , n12778 );
nand ( n12788 , n12786 , n12787 );
not ( n12789 , n12788 );
and ( n12790 , n12747 , n12741 );
not ( n12791 , n12747 );
and ( n12792 , n12791 , n12742 );
nor ( n12793 , n12790 , n12792 );
nand ( n12794 , n12789 , n12793 );
not ( n12795 , n12794 );
xnor ( n12796 , n12760 , n12769 );
not ( n12797 , n12796 );
and ( n12798 , n11443 , n49 );
not ( n12799 , n11443 );
and ( n12800 , n12799 , n12152 );
nor ( n12801 , n12798 , n12800 );
not ( n12802 , n12801 );
not ( n12803 , n11462 );
or ( n12804 , n12802 , n12803 );
nand ( n12805 , n12712 , n12671 );
nand ( n12806 , n12804 , n12805 );
not ( n12807 , n12806 );
not ( n12808 , n12775 );
not ( n12809 , n11386 );
or ( n12810 , n12808 , n12809 );
nand ( n12811 , n12535 , n12533 , n11393 );
nand ( n12812 , n12810 , n12811 );
not ( n12813 , n12812 );
not ( n12814 , n12813 );
or ( n12815 , n12807 , n12814 );
or ( n12816 , n12806 , n12813 );
nand ( n12817 , n12815 , n12816 );
and ( n12818 , n12797 , n12817 );
and ( n12819 , n12806 , n12812 );
nor ( n12820 , n12818 , n12819 );
and ( n12821 , n12783 , n12784 );
not ( n12822 , n12783 );
and ( n12823 , n12822 , n12785 );
nor ( n12824 , n12821 , n12823 );
nand ( n12825 , n12820 , n12824 );
not ( n12826 , n12825 );
not ( n12827 , n11731 );
not ( n12828 , n12767 );
not ( n12829 , n12828 );
and ( n12830 , n12827 , n12829 );
not ( n12831 , n11738 );
and ( n12832 , n12831 , n6014 );
nor ( n12833 , n12830 , n12832 );
not ( n12834 , n12833 );
not ( n12835 , n51 );
nor ( n12836 , n12835 , n11385 );
not ( n12837 , n12836 );
xor ( n12838 , n11443 , n50 );
not ( n12839 , n12838 );
not ( n12840 , n11460 );
or ( n12841 , n12839 , n12840 );
nand ( n12842 , n12801 , n12671 );
nand ( n12843 , n12841 , n12842 );
not ( n12844 , n12843 );
not ( n12845 , n12844 );
or ( n12846 , n12837 , n12845 );
not ( n12847 , n12836 );
nand ( n12848 , n12847 , n12843 );
nand ( n12849 , n12846 , n12848 );
and ( n12850 , n12834 , n12849 );
and ( n12851 , n12836 , n12843 );
nor ( n12852 , n12850 , n12851 );
not ( n12853 , n12817 );
not ( n12854 , n12796 );
and ( n12855 , n12853 , n12854 );
and ( n12856 , n12796 , n12817 );
nor ( n12857 , n12855 , n12856 );
nand ( n12858 , n12852 , n12857 );
not ( n12859 , n12858 );
nand ( n12860 , n51 , n3693 );
not ( n12861 , n51 );
not ( n12862 , n12861 );
not ( n12863 , n12538 );
or ( n12864 , n12862 , n12863 );
not ( n12865 , n11451 );
nand ( n12866 , n12864 , n12865 );
and ( n12867 , n12860 , n11445 , n12866 );
not ( n12868 , n11737 );
and ( n12869 , n49 , n11735 );
not ( n12870 , n49 );
and ( n12871 , n12870 , n12538 );
nor ( n12872 , n12869 , n12871 );
not ( n12873 , n12872 );
or ( n12874 , n12868 , n12873 );
not ( n12875 , n11825 );
nand ( n12876 , n12875 , n6014 );
nand ( n12877 , n12874 , n12876 );
nand ( n12878 , n12867 , n12877 );
not ( n12879 , n12878 );
not ( n12880 , n12833 );
not ( n12881 , n12849 );
or ( n12882 , n12880 , n12881 );
or ( n12883 , n12833 , n12849 );
nand ( n12884 , n12882 , n12883 );
nor ( n12885 , n12879 , n12884 );
nand ( n12886 , n51 , n3774 );
and ( n12887 , n11743 , n12886 );
not ( n12888 , n51 );
not ( n12889 , n12888 );
not ( n12890 , n11737 );
or ( n12891 , n12889 , n12890 );
nand ( n12892 , n12875 , n6210 );
nand ( n12893 , n12891 , n12892 );
nand ( n12894 , n12887 , n12893 );
and ( n12895 , n51 , n12671 );
not ( n12896 , n11730 );
not ( n12897 , n12896 );
not ( n12898 , n12872 );
or ( n12899 , n12897 , n12898 );
nand ( n12900 , n11737 , n6210 );
nand ( n12901 , n12899 , n12900 );
nor ( n12902 , n12895 , n12901 );
or ( n12903 , n12894 , n12902 );
nand ( n12904 , n12895 , n12901 );
nand ( n12905 , n12903 , n12904 );
not ( n12906 , n12758 );
nor ( n12907 , n12906 , n11461 );
and ( n12908 , n12756 , n12907 );
and ( n12909 , n12838 , n11471 );
nor ( n12910 , n12908 , n12909 );
nor ( n12911 , n12867 , n12877 );
not ( n12912 , n12911 );
nand ( n12913 , n12912 , n12878 );
nand ( n12914 , n12910 , n12913 );
and ( n12915 , n12905 , n12914 );
nor ( n12916 , n12913 , n12910 );
nor ( n12917 , n12915 , n12916 );
or ( n12918 , n12885 , n12917 );
nand ( n12919 , n12879 , n12884 );
nand ( n12920 , n12918 , n12919 );
not ( n12921 , n12920 );
or ( n12922 , n12859 , n12921 );
not ( n12923 , n12852 );
not ( n12924 , n12857 );
nand ( n12925 , n12923 , n12924 );
nand ( n12926 , n12922 , n12925 );
not ( n12927 , n12926 );
or ( n12928 , n12826 , n12927 );
not ( n12929 , n12820 );
not ( n12930 , n12824 );
nand ( n12931 , n12929 , n12930 );
nand ( n12932 , n12928 , n12931 );
not ( n12933 , n12932 );
or ( n12934 , n12795 , n12933 );
not ( n12935 , n12793 );
nand ( n12936 , n12788 , n12935 );
nand ( n12937 , n12934 , n12936 );
not ( n12938 , n12937 );
or ( n12939 , n12755 , n12938 );
not ( n12940 , n12753 );
nand ( n12941 , n12751 , n12940 );
nand ( n12942 , n12939 , n12941 );
not ( n12943 , n12942 );
or ( n12944 , n12707 , n12943 );
or ( n12945 , n12704 , n12705 );
nand ( n12946 , n12944 , n12945 );
nand ( n12947 , n12649 , n12946 );
nand ( n12948 , n12648 , n12947 );
not ( n12949 , n12948 );
xor ( n12950 , n12412 , n12411 );
xnor ( n12951 , n12370 , n12343 );
not ( n12952 , n12635 );
not ( n12953 , n12630 );
or ( n12954 , n12952 , n12953 );
not ( n12955 , n12620 );
nand ( n12956 , n12955 , n12626 );
nand ( n12957 , n12954 , n12956 );
not ( n12958 , n12604 );
not ( n12959 , n12599 );
or ( n12960 , n12958 , n12959 );
nand ( n12961 , n12594 , n12593 );
nand ( n12962 , n12960 , n12961 );
not ( n12963 , n12962 );
and ( n12964 , n12957 , n12963 );
not ( n12965 , n12957 );
and ( n12966 , n12965 , n12962 );
nor ( n12967 , n12964 , n12966 );
xor ( n12968 , n12951 , n12967 );
xor ( n12969 , n12950 , n12968 );
or ( n12970 , n12605 , n12588 );
or ( n12971 , n12583 , n12582 );
nand ( n12972 , n12970 , n12971 );
not ( n12973 , n12972 );
and ( n12974 , n12969 , n12973 );
not ( n12975 , n12969 );
and ( n12976 , n12975 , n12972 );
nor ( n12977 , n12974 , n12976 );
not ( n12978 , n12642 );
not ( n12979 , n12610 );
and ( n12980 , n12978 , n12979 );
and ( n12981 , n12637 , n12614 );
nor ( n12982 , n12980 , n12981 );
not ( n12983 , n12982 );
and ( n12984 , n12977 , n12983 );
not ( n12985 , n12977 );
and ( n12986 , n12985 , n12982 );
nor ( n12987 , n12984 , n12986 );
or ( n12988 , n12949 , n12987 );
or ( n12989 , n12982 , n12977 );
nand ( n12990 , n12988 , n12989 );
not ( n12991 , n12990 );
and ( n12992 , n12969 , n12972 );
and ( n12993 , n12950 , n12968 );
nor ( n12994 , n12992 , n12993 );
xnor ( n12995 , n12414 , n12423 );
not ( n12996 , n12951 );
not ( n12997 , n12967 );
and ( n12998 , n12996 , n12997 );
and ( n12999 , n12962 , n12957 );
nor ( n13000 , n12998 , n12999 );
xnor ( n13001 , n12375 , n12334 );
xnor ( n13002 , n13000 , n13001 );
xnor ( n13003 , n12995 , n13002 );
xor ( n13004 , n12994 , n13003 );
not ( n13005 , n13004 );
or ( n13006 , n12991 , n13005 );
or ( n13007 , n12994 , n13003 );
nand ( n13008 , n13006 , n13007 );
not ( n13009 , n13008 );
or ( n13010 , n12995 , n13002 );
or ( n13011 , n13001 , n13000 );
nand ( n13012 , n13010 , n13011 );
not ( n13013 , n13012 );
xnor ( n13014 , n12390 , n12427 );
not ( n13015 , n13014 );
or ( n13016 , n13013 , n13015 );
or ( n13017 , n13012 , n13014 );
nand ( n13018 , n13016 , n13017 );
not ( n13019 , n13018 );
or ( n13020 , n13009 , n13019 );
not ( n13021 , n13014 );
nand ( n13022 , n13021 , n13012 );
nand ( n13023 , n13020 , n13022 );
not ( n13024 , n13023 );
or ( n13025 , n12432 , n13024 );
not ( n13026 , n12430 );
nand ( n13027 , n13026 , n12388 );
nand ( n13028 , n13025 , n13027 );
xnor ( n13029 , n12308 , n12234 );
and ( n13030 , n12384 , n12387 );
and ( n13031 , n12386 , n12385 );
nor ( n13032 , n13030 , n13031 );
nor ( n13033 , n13029 , n13032 );
or ( n13034 , n13028 , n13033 );
nand ( n13035 , n13029 , n13032 );
nand ( n13036 , n13034 , n13035 );
nand ( n13037 , n12314 , n13036 );
not ( n13038 , n12233 );
nand ( n13039 , n13038 , n12311 );
or ( n13040 , n12313 , n13039 );
nand ( n13041 , n13037 , n11895 , n13040 );
nand ( n13042 , n12093 , n12217 );
nand ( n13043 , n13042 , n12092 );
not ( n13044 , n13043 );
nand ( n13045 , n13044 , n12227 );
or ( n13046 , n13041 , n13045 );
or ( n13047 , n11893 , n11894 );
nand ( n13048 , n13046 , n13047 );
nor ( n13049 , n12232 , n13048 );
and ( n13050 , n11671 , n11771 );
nor ( n13051 , n13049 , n13050 );
nand ( n13052 , n11788 , n13051 );
nand ( n13053 , n11786 , n13052 );
nor ( n13054 , n11332 , n11418 );
nor ( n13055 , n11331 , n13054 );
nand ( n13056 , n13053 , n13055 );
nand ( n13057 , n11424 , n13056 );
not ( n13058 , n13057 );
nand ( n13059 , n11278 , n13058 );
not ( n13060 , n11058 );
not ( n13061 , n11278 );
nand ( n13062 , n13061 , n13057 );
nand ( n13063 , n13059 , n13060 , n13062 );
not ( n13064 , n11058 );
nor ( n13065 , n13064 , n11070 );
not ( n13066 , n10431 );
nand ( n13067 , n13065 , n11047 , n10929 , n13066 );
nand ( n13068 , n11071 , n13063 , n13067 );
not ( n13069 , n13054 );
nand ( n13070 , n13069 , n11419 );
not ( n13071 , n13053 );
buf ( n13072 , n13071 );
and ( n13073 , n13070 , n13072 );
or ( n13074 , n13070 , n13072 );
not ( n13075 , n11058 );
nand ( n13076 , n13074 , n13075 );
nor ( n13077 , n13073 , n13076 );
not ( n13078 , n13077 );
not ( n13079 , n10928 );
not ( n13080 , n13079 );
and ( n13081 , n10429 , n10889 , n10832 , n10862 );
not ( n13082 , n10797 );
nand ( n13083 , n13081 , n13082 );
not ( n13084 , n13083 );
not ( n13085 , n11046 );
nand ( n13086 , n13084 , n13085 );
nand ( n13087 , n13080 , n11058 , n13086 );
not ( n13088 , n11046 );
nand ( n13089 , n11058 , n13079 , n13084 , n13088 );
nand ( n13090 , n13078 , n13087 , n13089 );
not ( n13091 , n11784 );
nor ( n13092 , n13091 , n11782 );
not ( n13093 , n13051 );
and ( n13094 , n13093 , n11772 );
and ( n13095 , n13092 , n11775 , n13094 );
buf ( n13096 , n11787 );
nor ( n13097 , n13094 , n13096 , n13092 );
nor ( n13098 , n13095 , n13097 );
or ( n13099 , n11776 , n13092 );
not ( n13100 , n11775 );
not ( n13101 , n13096 );
or ( n13102 , n13100 , n13101 );
nand ( n13103 , n13102 , n13092 );
nand ( n13104 , n13099 , n13103 );
and ( n13105 , n13098 , n13104 );
nor ( n13106 , n13105 , n11058 );
not ( n13107 , n13106 );
not ( n13108 , n13081 );
not ( n13109 , n13108 );
not ( n13110 , n237 );
not ( n13111 , n10999 );
not ( n13112 , n13111 );
or ( n13113 , n13110 , n13112 );
nand ( n13114 , n10989 , n10991 );
nand ( n13115 , n13113 , n13114 );
and ( n13116 , n13082 , n10968 , n13115 );
nand ( n13117 , n13109 , n13116 );
not ( n13118 , n13117 );
buf ( n13119 , n11045 );
buf ( n13120 , n13119 );
nand ( n13121 , n13118 , n13120 );
not ( n13122 , n11023 );
buf ( n13123 , n13122 );
not ( n13124 , n13123 );
nand ( n13125 , n13121 , n11058 , n13124 );
not ( n13126 , n13117 );
nand ( n13127 , n13126 , n13123 , n13120 , n11058 );
nand ( n13128 , n13107 , n13125 , n13127 );
or ( n13129 , n13071 , n13054 );
nand ( n13130 , n13129 , n11419 );
not ( n13131 , n11331 );
nand ( n13132 , n13131 , n11421 );
not ( n13133 , n13132 );
nor ( n13134 , n13130 , n13133 );
not ( n13135 , n13130 );
nor ( n13136 , n13135 , n13132 );
or ( n13137 , n13134 , n11058 , n13136 );
nor ( n13138 , n13122 , n13108 );
nand ( n13139 , n13138 , n10928 , n13119 );
and ( n13140 , n11058 , n10406 );
and ( n13141 , n13139 , n13140 );
not ( n13142 , n13139 );
not ( n13143 , n11058 );
not ( n13144 , n10406 );
not ( n13145 , n13144 );
or ( n13146 , n13143 , n13145 );
nand ( n13147 , n13146 , n13116 );
and ( n13148 , n13142 , n13147 );
nor ( n13149 , n13141 , n13148 );
and ( n13150 , n11058 , n10406 );
nor ( n13151 , n13150 , n13116 );
or ( n13152 , n13149 , n13151 );
nand ( n13153 , n13137 , n13152 );
buf ( n13154 , n10969 );
not ( n13155 , n13154 );
not ( n13156 , n13155 );
buf ( n13157 , n13115 );
nand ( n13158 , n13084 , n13157 );
not ( n13159 , n13158 );
not ( n13160 , n13159 );
or ( n13161 , n13156 , n13160 );
not ( n13162 , n13154 );
not ( n13163 , n13158 );
or ( n13164 , n13162 , n13163 );
nand ( n13165 , n13164 , n11058 );
not ( n13166 , n13165 );
nand ( n13167 , n13161 , n13166 );
not ( n13168 , n11058 );
buf ( n13169 , n13049 );
not ( n13170 , n13169 );
not ( n13171 , n11772 );
nor ( n13172 , n13171 , n13050 );
not ( n13173 , n13172 );
or ( n13174 , n13170 , n13173 );
or ( n13175 , n13169 , n13172 );
nand ( n13176 , n13174 , n13175 );
nand ( n13177 , n13168 , n13176 );
nand ( n13178 , n13167 , n13177 );
buf ( n13179 , n10798 );
nor ( n13180 , n13144 , n13108 );
and ( n13181 , n10928 , n11070 );
and ( n13182 , n13179 , n13088 , n13180 , n13181 );
not ( n13183 , n10405 );
and ( n13184 , n11058 , n13183 );
not ( n13185 , n13184 );
or ( n13186 , n13182 , n13185 );
not ( n13187 , n11277 );
not ( n13188 , n13057 );
or ( n13189 , n13187 , n13188 );
nand ( n13190 , n13189 , n11275 );
and ( n13191 , n11164 , n11159 );
and ( n13192 , n3201 , n11165 );
nor ( n13193 , n13191 , n13192 );
and ( n13194 , n11173 , n11169 );
nor ( n13195 , n13194 , n11130 );
xnor ( n13196 , n13193 , n13195 );
xor ( n13197 , n13196 , n3107 );
or ( n13198 , n11176 , n13197 );
nand ( n13199 , n11176 , n13197 );
nand ( n13200 , n13198 , n13199 );
or ( n13201 , n11177 , n11168 );
or ( n13202 , n11149 , n11167 );
nand ( n13203 , n13201 , n13202 );
xnor ( n13204 , n13200 , n13203 );
and ( n13205 , n11216 , n11182 );
and ( n13206 , n11147 , n11181 );
nor ( n13207 , n13205 , n13206 );
nor ( n13208 , n13204 , n13207 );
and ( n13209 , n13204 , n13207 );
nor ( n13210 , n13208 , n13209 );
xnor ( n13211 , n13190 , n13210 );
or ( n13212 , n13211 , n11058 );
nand ( n13213 , n13186 , n13212 );
not ( n13214 , n13036 );
and ( n13215 , n13039 , n13214 );
nor ( n13216 , n13215 , n12313 );
or ( n13217 , n13216 , n13043 );
nand ( n13218 , n13217 , n12221 );
buf ( n13219 , n12230 );
buf ( n13220 , n13219 );
not ( n13221 , n13220 );
and ( n13222 , n13047 , n11895 );
or ( n13223 , n13218 , n13221 , n13222 );
and ( n13224 , n13218 , n12227 , n13222 );
not ( n13225 , n13220 );
or ( n13226 , n12227 , n13225 , n13222 );
not ( n13227 , n13219 );
and ( n13228 , n13227 , n13222 );
nor ( n13229 , n13228 , n11057 );
nand ( n13230 , n13226 , n13229 );
nor ( n13231 , n13224 , n13230 );
nand ( n13232 , n13223 , n13231 );
nor ( n13233 , n13084 , n13157 );
not ( n13234 , n13233 );
not ( n13235 , n13159 );
nand ( n13236 , n13234 , n11058 , n13235 );
nand ( n13237 , n13232 , n13236 );
not ( n13238 , n11162 );
not ( n13239 , n9471 );
or ( n13240 , n11165 , n11159 );
nand ( n13241 , n13240 , n11074 );
not ( n13242 , n13241 );
or ( n13243 , n13239 , n13242 );
or ( n13244 , n9471 , n13241 );
nand ( n13245 , n13243 , n13244 );
not ( n13246 , n13245 );
or ( n13247 , n13238 , n13246 );
or ( n13248 , n11162 , n13245 );
nand ( n13249 , n13247 , n13248 );
not ( n13250 , n13249 );
and ( n13251 , n3201 , n11159 );
and ( n13252 , n11074 , n11165 );
nor ( n13253 , n13251 , n13252 );
not ( n13254 , n13253 );
and ( n13255 , n11162 , n13254 );
not ( n13256 , n11162 );
and ( n13257 , n13256 , n13253 );
nor ( n13258 , n13255 , n13257 );
or ( n13259 , n3107 , n13196 );
or ( n13260 , n13195 , n13193 );
nand ( n13261 , n13259 , n13260 );
and ( n13262 , n13258 , n13261 );
and ( n13263 , n11162 , n13254 );
nor ( n13264 , n13262 , n13263 );
not ( n13265 , n13264 );
and ( n13266 , n13250 , n13265 );
and ( n13267 , n13249 , n13264 );
nor ( n13268 , n13266 , n13267 );
not ( n13269 , n13268 );
xor ( n13270 , n13261 , n13258 );
not ( n13271 , n13270 );
and ( n13272 , n13203 , n13200 );
and ( n13273 , n11177 , n13197 );
nor ( n13274 , n13272 , n13273 );
nand ( n13275 , n13271 , n13274 );
not ( n13276 , n11277 );
nor ( n13277 , n13276 , n13209 );
not ( n13278 , n13277 );
not ( n13279 , n11422 );
or ( n13280 , n13278 , n13279 );
not ( n13281 , n13209 );
not ( n13282 , n11275 );
and ( n13283 , n13281 , n13282 );
nor ( n13284 , n13283 , n13208 );
nand ( n13285 , n13280 , n13284 );
and ( n13286 , n13275 , n13285 );
not ( n13287 , n13286 );
not ( n13288 , n13274 );
nand ( n13289 , n13270 , n13288 );
not ( n13290 , n13056 );
buf ( n13291 , n13277 );
buf ( n13292 , n13291 );
nand ( n13293 , n13290 , n13275 , n13292 );
nand ( n13294 , n13287 , n13289 , n13293 );
nand ( n13295 , n13269 , n13294 );
not ( n13296 , n13295 );
not ( n13297 , n13294 );
and ( n13298 , n13268 , n13297 );
nor ( n13299 , n13298 , n11058 );
not ( n13300 , n13299 );
or ( n13301 , n13296 , n13300 );
not ( n13302 , n13084 );
not ( n13303 , n11046 );
not ( n13304 , n13303 );
or ( n13305 , n13302 , n13304 );
nand ( n13306 , n13305 , n13184 );
nand ( n13307 , n13301 , n13306 );
not ( n13308 , n11058 );
not ( n13309 , n13308 );
nand ( n13310 , n13289 , n13275 );
and ( n13311 , n13310 , n13291 );
and ( n13312 , n11423 , n13311 );
not ( n13313 , n13284 );
and ( n13314 , n13310 , n13313 );
nor ( n13315 , n13312 , n13314 );
and ( n13316 , n13311 , n13055 );
not ( n13317 , n13052 );
nand ( n13318 , n13316 , n13317 );
not ( n13319 , n13292 );
not ( n13320 , n13057 );
or ( n13321 , n13319 , n13320 );
nor ( n13322 , n13310 , n13313 );
nand ( n13323 , n13321 , n13322 );
nand ( n13324 , n13316 , n11785 );
nand ( n13325 , n13315 , n13318 , n13323 , n13324 );
not ( n13326 , n13325 );
or ( n13327 , n13309 , n13326 );
nand ( n13328 , n13327 , n13306 );
not ( n13329 , n13120 );
nand ( n13330 , n11058 , n13329 , n13126 );
nand ( n13331 , n13120 , n11058 , n13117 );
not ( n13332 , n13096 );
nand ( n13333 , n13332 , n11775 );
or ( n13334 , n13094 , n13333 );
nand ( n13335 , n13094 , n13333 );
not ( n13336 , n11058 );
nand ( n13337 , n13334 , n13335 , n13336 );
nand ( n13338 , n13330 , n13331 , n13337 );
not ( n13339 , n12220 );
nand ( n13340 , n13339 , n12092 );
not ( n13341 , n13340 );
not ( n13342 , n13042 );
or ( n13343 , n13342 , n13216 );
not ( n13344 , n12218 );
nand ( n13345 , n13343 , n13344 );
not ( n13346 , n13345 );
and ( n13347 , n13341 , n13346 );
and ( n13348 , n13340 , n13345 );
nor ( n13349 , n13347 , n13348 );
or ( n13350 , n11058 , n13349 );
not ( n13351 , n10890 );
not ( n13352 , n13351 );
not ( n13353 , n13352 );
buf ( n13354 , n10718 );
not ( n13355 , n13354 );
nor ( n13356 , n13353 , n13355 );
not ( n13357 , n13356 );
not ( n13358 , n13352 );
not ( n13359 , n10833 );
not ( n13360 , n10863 );
and ( n13361 , n10796 , n13359 , n13360 );
not ( n13362 , n10745 );
not ( n13363 , n10782 );
nor ( n13364 , n13362 , n13363 );
nand ( n13365 , n13361 , n13364 );
not ( n13366 , n13365 );
or ( n13367 , n13358 , n13366 );
nand ( n13368 , n13367 , n11058 );
not ( n13369 , n13368 );
not ( n13370 , n13354 );
nand ( n13371 , n13353 , n13370 , n13361 , n13364 );
nand ( n13372 , n13357 , n13369 , n13371 );
nand ( n13373 , n13350 , n13372 );
not ( n13374 , n13306 );
not ( n13375 , n13362 );
not ( n13376 , n13363 );
nand ( n13377 , n13375 , n13376 );
not ( n13378 , n10717 );
not ( n13379 , n13378 );
not ( n13380 , n10697 );
not ( n13381 , n13380 );
not ( n13382 , n10601 );
nand ( n13383 , n13379 , n13381 , n13382 );
nand ( n13384 , n11057 , n10796 );
nor ( n13385 , n13377 , n13383 , n13384 );
nand ( n13386 , n13385 , n13109 );
buf ( n13387 , n13183 );
not ( n13388 , n13387 );
not ( n13389 , n11047 );
nor ( n13390 , n13386 , n13388 , n13389 );
buf ( n13391 , n10430 );
not ( n13392 , n13391 );
nand ( n13393 , n13392 , n11058 , n13179 , n10891 );
not ( n13394 , n11058 );
not ( n13395 , n13391 );
nor ( n13396 , n13394 , n13395 );
nand ( n13397 , n10892 , n13396 );
and ( n13398 , n13220 , n12227 );
or ( n13399 , n13398 , n13218 );
nand ( n13400 , n13398 , n13218 );
not ( n13401 , n11058 );
nand ( n13402 , n13399 , n13400 , n13401 );
nand ( n13403 , n13393 , n13397 , n13402 );
not ( n13404 , n13359 );
not ( n13405 , n13179 );
buf ( n13406 , n13360 );
not ( n13407 , n13406 );
or ( n13408 , n13405 , n13407 );
nand ( n13409 , n13408 , n11057 );
or ( n13410 , n13404 , n13409 );
nor ( n13411 , n12218 , n13342 );
and ( n13412 , n13411 , n13216 );
nor ( n13413 , n13411 , n13216 );
nor ( n13414 , n13412 , n13413 );
or ( n13415 , n11058 , n13414 );
nand ( n13416 , n13404 , n11058 , n13179 , n13406 );
nand ( n13417 , n13410 , n13415 , n13416 );
and ( n13418 , n13405 , n13406 );
not ( n13419 , n13405 );
not ( n13420 , n13406 );
and ( n13421 , n13419 , n13420 );
nor ( n13422 , n13418 , n13421 );
not ( n13423 , n13375 );
not ( n13424 , n13380 );
not ( n13425 , n13378 );
and ( n13426 , n13424 , n10796 , n13382 , n13425 );
nand ( n13427 , n13423 , n11057 , n13426 , n13376 );
not ( n13428 , n13426 );
not ( n13429 , n13376 );
or ( n13430 , n13428 , n13429 );
not ( n13431 , n13362 );
and ( n13432 , n11057 , n13431 );
nand ( n13433 , n13430 , n13432 );
not ( n13434 , n11057 );
buf ( n13435 , n13028 );
not ( n13436 , n13435 );
not ( n13437 , n13033 );
nand ( n13438 , n13437 , n13035 );
not ( n13439 , n13438 );
or ( n13440 , n13436 , n13439 );
or ( n13441 , n13435 , n13438 );
nand ( n13442 , n13440 , n13441 );
nand ( n13443 , n13434 , n13442 );
nand ( n13444 , n13427 , n13433 , n13443 );
not ( n13445 , n11057 );
and ( n13446 , n12430 , n12388 );
not ( n13447 , n13023 );
and ( n13448 , n13446 , n13447 );
and ( n13449 , n13027 , n12431 );
nor ( n13450 , n13449 , n13447 );
nor ( n13451 , n13023 , n12430 , n12388 );
nor ( n13452 , n13448 , n13450 , n13451 );
and ( n13453 , n13445 , n13452 );
not ( n13454 , n13445 );
not ( n13455 , n13426 );
not ( n13456 , n13363 );
and ( n13457 , n13455 , n13456 );
and ( n13458 , n13426 , n13363 );
nor ( n13459 , n13457 , n13458 );
and ( n13460 , n13454 , n13459 );
nor ( n13461 , n13453 , n13460 );
not ( n13462 , n11057 );
not ( n13463 , n13462 );
xor ( n13464 , n13008 , n13018 );
not ( n13465 , n13464 );
or ( n13466 , n13463 , n13465 );
not ( n13467 , n10796 );
xor ( n13468 , n13354 , n13467 );
nand ( n13469 , n13468 , n11057 );
nand ( n13470 , n13466 , n13469 );
not ( n13471 , n11057 );
not ( n13472 , n13471 );
xor ( n13473 , n12990 , n13004 );
not ( n13474 , n13473 );
or ( n13475 , n13472 , n13474 );
nand ( n13476 , n13381 , n13382 );
not ( n13477 , n13379 );
nand ( n13478 , n13476 , n13477 );
nand ( n13479 , n13478 , n11057 , n13383 );
nand ( n13480 , n13475 , n13479 );
not ( n13481 , n10620 );
not ( n13482 , n13481 );
not ( n13483 , n10696 );
nand ( n13484 , n10671 , n13382 );
nor ( n13485 , n13483 , n13484 );
not ( n13486 , n13485 );
nand ( n13487 , n13482 , n13486 );
nand ( n13488 , n13481 , n13485 );
and ( n13489 , n13487 , n11057 , n13488 );
not ( n13490 , n12949 );
buf ( n13491 , n12987 );
and ( n13492 , n13490 , n13491 );
nor ( n13493 , n13490 , n13491 );
nor ( n13494 , n13492 , n11057 , n13493 );
nor ( n13495 , n13489 , n13494 );
or ( n13496 , n12649 , n12946 );
not ( n13497 , n11057 );
nand ( n13498 , n13496 , n13497 , n12947 );
nand ( n13499 , n13484 , n11057 , n10696 );
not ( n13500 , n13484 );
nand ( n13501 , n13483 , n11057 , n13500 );
nand ( n13502 , n13498 , n13499 , n13501 );
and ( n13503 , n10643 , n13382 );
buf ( n13504 , n10670 );
nor ( n13505 , n13503 , n13504 );
not ( n13506 , n13503 );
not ( n13507 , n13504 );
or ( n13508 , n13506 , n13507 );
nand ( n13509 , n13508 , n11057 );
or ( n13510 , n13505 , n13509 );
xnor ( n13511 , n12942 , n12706 );
or ( n13512 , n11057 , n13511 );
nand ( n13513 , n13510 , n13512 );
not ( n13514 , n11057 );
not ( n13515 , n13514 );
nand ( n13516 , n12941 , n12754 );
not ( n13517 , n13516 );
not ( n13518 , n12937 );
or ( n13519 , n13517 , n13518 );
or ( n13520 , n13516 , n12937 );
nand ( n13521 , n13519 , n13520 );
not ( n13522 , n13521 );
or ( n13523 , n13515 , n13522 );
nor ( n13524 , n10643 , n13382 );
not ( n13525 , n13524 );
not ( n13526 , n13503 );
nand ( n13527 , n13525 , n11057 , n13526 );
nand ( n13528 , n13523 , n13527 );
not ( n13529 , n11057 );
not ( n13530 , n13529 );
and ( n13531 , n12936 , n12794 );
xor ( n13532 , n13531 , n12932 );
not ( n13533 , n13532 );
or ( n13534 , n13530 , n13533 );
not ( n13535 , n13382 );
not ( n13536 , n10448 );
not ( n13537 , n10600 );
nand ( n13538 , n13536 , n13537 );
nand ( n13539 , n13535 , n13538 , n11057 );
nand ( n13540 , n13534 , n13539 );
not ( n13541 , n10599 );
nand ( n13542 , n10577 , n10579 );
nor ( n13543 , n13541 , n13542 );
nand ( n13544 , n11057 , n13537 );
or ( n13545 , n13543 , n13544 );
nand ( n13546 , n12931 , n12825 );
not ( n13547 , n13546 );
not ( n13548 , n12926 );
and ( n13549 , n13547 , n13548 );
and ( n13550 , n13546 , n12926 );
nor ( n13551 , n13549 , n13550 );
or ( n13552 , n11057 , n13551 );
nand ( n13553 , n13545 , n13552 );
not ( n13554 , n10554 );
not ( n13555 , n13554 );
nand ( n13556 , n13555 , n10529 );
not ( n13557 , n10578 );
nand ( n13558 , n13556 , n13557 );
and ( n13559 , n10576 , n13558 );
or ( n13560 , n10576 , n13558 );
nand ( n13561 , n13560 , n11057 );
or ( n13562 , n13559 , n13561 );
and ( n13563 , n12925 , n12858 );
xnor ( n13564 , n12920 , n13563 );
or ( n13565 , n11057 , n13564 );
nand ( n13566 , n13562 , n13565 );
not ( n13567 , n13554 );
nand ( n13568 , n13567 , n13557 );
not ( n13569 , n13568 );
not ( n13570 , n10529 );
not ( n13571 , n13570 );
nor ( n13572 , n13569 , n13571 );
or ( n13573 , n13568 , n13570 );
nand ( n13574 , n13573 , n11056 );
or ( n13575 , n13572 , n13574 );
not ( n13576 , n12917 );
not ( n13577 , n12919 );
nor ( n13578 , n13577 , n12885 );
not ( n13579 , n13578 );
and ( n13580 , n13576 , n13579 );
and ( n13581 , n12917 , n13578 );
nor ( n13582 , n13580 , n13581 );
or ( n13583 , n11057 , n13582 );
nand ( n13584 , n13575 , n13583 );
not ( n13585 , n10464 );
not ( n13586 , n10465 );
nor ( n13587 , n13585 , n13586 );
nor ( n13588 , n10527 , n13587 );
not ( n13589 , n10527 );
not ( n13590 , n13587 );
or ( n13591 , n13589 , n13590 );
nand ( n13592 , n13591 , n11056 );
or ( n13593 , n13588 , n13592 );
not ( n13594 , n12905 );
not ( n13595 , n12916 );
nand ( n13596 , n13595 , n12914 );
not ( n13597 , n13596 );
and ( n13598 , n13594 , n13597 );
and ( n13599 , n12905 , n13596 );
nor ( n13600 , n13598 , n13599 );
or ( n13601 , n11056 , n13600 );
nand ( n13602 , n13593 , n13601 );
or ( n13603 , n12887 , n12893 );
not ( n13604 , n11056 );
nand ( n13605 , n13603 , n13604 , n12894 );
not ( n13606 , n10520 );
not ( n13607 , n13606 );
not ( n13608 , n10522 );
nand ( n13609 , n13607 , n13608 );
not ( n13610 , n10505 );
nand ( n13611 , n18 , n13606 , n13610 );
not ( n13612 , n13606 );
not ( n13613 , n13612 );
not ( n13614 , n10506 );
or ( n13615 , n13613 , n13614 );
or ( n13616 , n18 , n13610 );
nand ( n13617 , n13616 , n13606 );
nand ( n13618 , n13615 , n13617 );
nand ( n13619 , n13609 , n13611 , n13618 );
nand ( n13620 , n11056 , n13619 );
nand ( n13621 , n13605 , n13620 );
not ( n13622 , n13214 );
buf ( n13623 , n12233 );
and ( n13624 , n13622 , n13623 , n12311 );
or ( n13625 , n13214 , n13623 , n12311 );
not ( n13626 , n13039 );
or ( n13627 , n12313 , n13626 );
nand ( n13628 , n13627 , n13214 );
nand ( n13629 , n13625 , n13628 );
nor ( n13630 , n13624 , n13629 );
not ( n13631 , n10488 );
not ( n13632 , n13631 );
buf ( n13633 , n10526 );
nand ( n13634 , n13632 , n13633 );
not ( n13635 , n13634 );
not ( n13636 , n10524 );
not ( n13637 , n13636 );
nor ( n13638 , n13635 , n13637 );
or ( n13639 , n13634 , n13636 );
nand ( n13640 , n13639 , n11056 );
or ( n13641 , n13638 , n13640 );
not ( n13642 , n12894 );
not ( n13643 , n12904 );
nor ( n13644 , n13643 , n12902 );
not ( n13645 , n13644 );
and ( n13646 , n13642 , n13645 );
and ( n13647 , n12894 , n13644 );
nor ( n13648 , n13646 , n13647 );
or ( n13649 , n11056 , n13648 );
nand ( n13650 , n13641 , n13649 );
or ( n13651 , n12886 , n11056 );
or ( n13652 , n19 , n10503 );
nand ( n13653 , n13652 , n11056 , n13610 );
nand ( n13654 , n13651 , n13653 );
nand ( n13655 , n2819 , n2820 );
and ( n13656 , n2874 , n13655 );
nor ( n13657 , n2874 , n13655 );
nor ( n13658 , n13656 , n1 , n13657 );
not ( n13659 , n10125 );
nor ( n13660 , n13659 , n9988 );
nor ( n13661 , n237 , n10124 , n13660 );
not ( n13662 , n10124 );
not ( n13663 , n13660 );
nor ( n13664 , n237 , n13662 , n13663 );
nor ( n13665 , n13658 , n13661 , n13664 );
not ( n13666 , n2870 );
nand ( n13667 , n2873 , n2840 );
not ( n13668 , n13667 );
and ( n13669 , n13666 , n13668 );
and ( n13670 , n2870 , n13667 );
nor ( n13671 , n13669 , n13670 );
or ( n13672 , n1 , n13671 );
and ( n13673 , n10123 , n10053 );
or ( n13674 , n10120 , n13673 );
nand ( n13675 , n10120 , n13673 );
nand ( n13676 , n13674 , n13675 , n1 );
nand ( n13677 , n13672 , n13676 );
xnor ( n13678 , n2866 , n2842 );
or ( n13679 , n1 , n13678 );
and ( n13680 , n10119 , n10069 );
or ( n13681 , n10116 , n13680 );
and ( n13682 , n10116 , n13680 );
nor ( n13683 , n13682 , n237 );
nand ( n13684 , n13681 , n13683 );
nand ( n13685 , n13679 , n13684 );
xnor ( n13686 , n2855 , n2845 );
or ( n13687 , n1 , n13686 );
or ( n13688 , n10108 , n10114 );
nand ( n13689 , n13688 , n1 , n10115 );
nand ( n13690 , n13687 , n13689 );
nor ( n13691 , n99 , n10107 );
or ( n13692 , n13691 , n237 , n10108 );
not ( n13693 , n19 );
not ( n13694 , n2847 );
and ( n13695 , n13693 , n13694 );
and ( n13696 , n19 , n2847 );
nor ( n13697 , n13695 , n13696 );
or ( n13698 , n1 , n13697 );
nand ( n13699 , n13692 , n13698 );
and ( n13700 , n11058 , n13422 );
not ( n13701 , n11058 );
and ( n13702 , n13701 , n13630 );
nor ( n13703 , n13700 , n13702 );
buf ( n13704 , n13387 );
buf ( n13705 , n13387 );
not ( n13706 , n13392 );
endmodule
