module top ( g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 );
input g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 ;
output g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 ;

wire n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , 
     n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , 
     n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , 
     n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , 
     n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , 
     n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , 
     n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , 
     n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , 
     n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , 
     n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , 
     n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , 
     n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , 
     n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , 
     n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , 
     n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , 
     n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , 
     n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , 
     n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , 
     n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , 
     n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , 
     n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , 
     n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , 
     n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , 
     n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , 
     n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , 
     n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , 
     n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , 
     n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , 
     n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , 
     n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , 
     n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , 
     n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , 
     n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , 
     n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , 
     n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , 
     n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , 
     n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , 
     n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , 
     n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , 
     n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , 
     n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , 
     n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , 
     n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , 
     n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , 
     n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , 
     n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , 
     n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , 
     n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , 
     n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , 
     n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , 
     n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , 
     n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , 
     n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , 
     n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , 
     n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , 
     n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , 
     n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , 
     n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , 
     n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , 
     n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , 
     n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , 
     n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , 
     n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , 
     n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , 
     n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , 
     n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , 
     n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , 
     n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , 
     n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , 
     n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , 
     n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , 
     n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , 
     n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , 
     n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , 
     n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , 
     n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , 
     n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , 
     n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , 
     n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , 
     n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , 
     n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , 
     n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , 
     n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , 
     n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , 
     n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , 
     n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , 
     n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , 
     n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , 
     n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , 
     n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , 
     n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , 
     n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , 
     n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , 
     n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , 
     n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , 
     n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , 
     n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , 
     n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , 
     n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , 
     n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , 
     n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , 
     n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , 
     n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , 
     n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , 
     n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , 
     n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , 
     n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , 
     n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , 
     n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , 
     n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , 
     n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , 
     n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , 
     n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , 
     n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , 
     n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , 
     n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , 
     n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , 
     n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , 
     n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , 
     n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , 
     n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , 
     n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , 
     n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , 
     n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , 
     n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , 
     n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , 
     n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , 
     n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , 
     n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , 
     n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , 
     n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , 
     n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , 
     n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , 
     n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , 
     n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , 
     n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , 
     n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , 
     n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , 
     n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , 
     n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , 
     n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , 
     n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , 
     n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , 
     n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , 
     n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , 
     n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , 
     n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , 
     n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , 
     n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , 
     n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , 
     n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , 
     n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , 
     n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , 
     n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , 
     n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , 
     n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , 
     n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , 
     n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , 
     n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , 
     n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , 
     n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , 
     n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , 
     n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , 
     n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , 
     n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , 
     n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , 
     n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , 
     n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , 
     n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , 
     n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , 
     n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , 
     n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , 
     n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , 
     n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , 
     n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , 
     n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , 
     n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , 
     n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , 
     n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , 
     n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , 
     n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , 
     n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , 
     n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , 
     n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , 
     n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , 
     n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , 
     n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , 
     n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , 
     n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , 
     n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , 
     n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , 
     n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , 
     n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , 
     n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , 
     n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , 
     n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , 
     n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , 
     n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , 
     n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , 
     n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , 
     n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , 
     n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 ;
wire t_0 , t_1 , t_2 , t_3 , t_4 , t_5 , t_6 , t_7 ;
buf ( n1  , g0 );
buf ( n2  , g1 );
buf ( n3  , g2 );
buf ( n4  , g3 );
buf ( n5  , g4 );
buf ( n6  , g5 );
buf ( n7  , g6 );
buf ( n8  , g7 );
buf ( n9  , g8 );
buf ( n10  , g9 );
buf ( n11  , g10 );
buf ( n12  , g11 );
buf ( n13  , g12 );
buf ( n14  , g13 );
buf ( n15  , g14 );
buf ( n16  , g15 );
buf ( n17  , g16 );
buf ( n18  , g17 );
buf ( n19  , g18 );
buf ( n20  , g19 );
buf ( n21  , g20 );
buf ( n22  , g21 );
buf ( n23  , g22 );
buf ( n24  , g23 );
buf ( n25  , g24 );
buf ( n26  , g25 );
buf ( n27  , g26 );
buf ( n28  , g27 );
buf ( n29  , g28 );
buf ( n30  , g29 );
buf ( n31  , g30 );
buf ( n32  , g31 );
buf ( n33  , g32 );
buf ( n34  , g33 );
buf ( n35  , g34 );
buf ( n36  , g35 );
buf ( n37  , g36 );
buf ( n38  , g37 );
buf ( n39  , g38 );
buf ( n40  , g39 );
buf ( n41  , g40 );
buf ( n42  , g41 );
buf ( n43  , g42 );
buf ( n44  , g43 );
buf ( n45  , g44 );
buf ( n46  , g45 );
buf ( n47  , g46 );
buf ( n48  , g47 );
buf ( g48 , n49  );
buf ( g49 , n50  );
buf ( g50 , n51  );
buf ( g51 , n52  );
buf ( g52 , n53  );
buf ( g53 , n54  );
buf ( g54 , n55  );
buf ( g55 , n56  );
buf ( g56 , n57  );
buf ( g57 , n58  );
buf ( g58 , n59  );
buf ( g59 , n60  );
buf ( g60 , n61  );
buf ( g61 , n62  );
buf ( g62 , n63  );
buf ( g63 , n64  );
buf ( g64 , n65  );
buf ( g65 , n66  );
buf ( g66 , n67  );
buf ( g67 , n68  );
buf ( g68 , n69  );
buf ( g69 , n70  );
buf ( g70 , n71  );
buf ( g71 , n72  );
buf ( g72 , n73  );
buf ( g73 , n74  );
buf ( g74 , n75  );
buf ( g75 , n76  );
buf ( g76 , n77  );
buf ( g77 , n78  );
buf ( g78 , n79  );
buf ( g79 , n80  );
buf ( g80 , n81  );
buf ( g81 , n82  );
buf ( g82 , n83  );
buf ( g83 , n84  );
buf ( g84 , n85  );
buf ( g85 , n86  );
buf ( g86 , n87  );
buf ( g87 , n88  );
buf ( g88 , n89  );
buf ( g89 , n90  );
buf ( g90 , n91  );
buf ( g91 , n92  );
buf ( g92 , n93  );
buf ( g93 , n94  );
buf ( g94 , n95  );
buf ( g95 , n96  );
buf ( g96 , n97  );
buf ( g97 , n98  );
buf ( n49 , 1'b0 );
buf ( n50 , 1'b0 );
buf ( n51 , 1'b0 );
buf ( n52 , 1'b0 );
buf ( n53 , 1'b0 );
buf ( n54 , 1'b0 );
buf ( n55 , 1'b0 );
buf ( n56 , 1'b0 );
buf ( n57 , 1'b0 );
buf ( n58 , 1'b0 );
buf ( n59 , 1'b0 );
buf ( n60 , 1'b0 );
buf ( n61 , 1'b0 );
buf ( n62 , 1'b0 );
buf ( n63 , 1'b0 );
buf ( n64 , 1'b0 );
buf ( n65 , 1'b0 );
buf ( n66 , n1787 );
buf ( n67 , n1605 );
buf ( n68 , n1623 );
buf ( n69 , n1799 );
buf ( n70 , n1827 );
buf ( n71 , n1838 );
buf ( n72 , n1860 );
buf ( n73 , n1876 );
buf ( n74 , n1888 );
buf ( n75 , n1902 );
buf ( n76 , n1931 );
buf ( n77 , n1943 );
buf ( n78 , n1968 );
buf ( n79 , n1993 );
buf ( n80 , n2017 );
buf ( n81 , n2005 );
buf ( n82 , n2013 );
buf ( n83 , n2015 );
buf ( n84 , n1785 );
buf ( n85 , n1808 );
buf ( n86 , n1819 );
buf ( n87 , n1833 );
buf ( n88 , n1844 );
buf ( n89 , n1851 );
buf ( n90 , n1866 );
buf ( n91 , n1891 );
buf ( n92 , n1910 );
buf ( n93 , n1921 );
buf ( n94 , n1949 );
buf ( n95 , n1955 );
buf ( n96 , n1972 );
buf ( n97 , n1980 );
buf ( n98 , n1995 );
nand ( n118 , n4 , n17 );
nand ( n119 , n2 , n19 );
xor ( n120 , n118 , n119 );
nand ( n121 , n3 , n18 );
and ( n122 , n120 , n121 );
and ( n123 , n118 , n119 );
or ( n124 , n122 , n123 );
nand ( n125 , n2 , n18 );
xor ( n126 , n124 , n125 );
nand ( n127 , n3 , n17 );
and ( n128 , n126 , n127 );
and ( n129 , n124 , n125 );
or ( n130 , n128 , n129 );
nand ( n131 , n1 , n18 );
xor ( n132 , n130 , n131 );
nand ( n133 , n2 , n17 );
and ( n134 , n132 , n133 );
and ( n135 , n130 , n131 );
or ( n136 , n134 , n135 );
nand ( n137 , n1 , n17 );
xor ( n138 , n136 , n137 );
nand ( n139 , n2 , n21 );
nand ( n140 , n3 , n20 );
xor ( n141 , n139 , n140 );
nand ( n142 , n4 , n19 );
and ( n143 , n141 , n142 );
and ( n144 , n139 , n140 );
or ( n145 , n143 , n144 );
nand ( n146 , n2 , n20 );
xor ( n147 , n145 , n146 );
nand ( n148 , n3 , n19 );
and ( n149 , n147 , n148 );
and ( n150 , n145 , n146 );
or ( n151 , n149 , n150 );
nand ( n152 , n5 , n17 );
nand ( n153 , n1 , n21 );
xor ( n154 , n152 , n153 );
nand ( n155 , n4 , n18 );
and ( n156 , n154 , n155 );
and ( n157 , n152 , n153 );
or ( n158 , n156 , n157 );
xor ( n159 , n151 , n158 );
xor ( n160 , n118 , n119 );
xor ( n161 , n160 , n121 );
and ( n162 , n159 , n161 );
and ( n163 , n151 , n158 );
or ( n164 , n162 , n163 );
nand ( n165 , n1 , n19 );
xor ( n166 , n164 , n165 );
xor ( n167 , n124 , n125 );
xor ( n168 , n167 , n127 );
and ( n169 , n166 , n168 );
and ( n170 , n164 , n165 );
or ( n171 , n169 , n170 );
xor ( n172 , n130 , n131 );
xor ( n173 , n172 , n133 );
xor ( n174 , n171 , n173 );
not ( n175 , n174 );
xor ( n176 , n164 , n165 );
xor ( n177 , n176 , n168 );
nand ( n178 , n2 , n22 );
nand ( n179 , n3 , n21 );
xor ( n180 , n178 , n179 );
nand ( n181 , n4 , n20 );
and ( n182 , n180 , n181 );
and ( n183 , n178 , n179 );
or ( n184 , n182 , n183 );
xor ( n185 , n139 , n140 );
xor ( n186 , n185 , n142 );
xor ( n187 , n184 , n186 );
nand ( n188 , n5 , n19 );
not ( n189 , n188 );
nand ( n190 , n6 , n18 );
not ( n191 , n190 );
nand ( n192 , n189 , n191 );
and ( n193 , n187 , n192 );
and ( n194 , n184 , n186 );
or ( n195 , n193 , n194 );
xor ( n196 , n152 , n153 );
xor ( n197 , n196 , n155 );
xor ( n198 , n195 , n197 );
xor ( n199 , n145 , n146 );
xor ( n200 , n199 , n148 );
and ( n201 , n198 , n200 );
and ( n202 , n195 , n197 );
or ( n203 , n201 , n202 );
nand ( n204 , n1 , n20 );
xor ( n205 , n203 , n204 );
xor ( n206 , n151 , n158 );
xor ( n207 , n206 , n161 );
and ( n208 , n205 , n207 );
and ( n209 , n203 , n204 );
or ( n210 , n208 , n209 );
xor ( n211 , n177 , n210 );
not ( n212 , n211 );
xor ( n213 , n203 , n204 );
xor ( n214 , n213 , n207 );
xor ( n215 , n195 , n197 );
xor ( n216 , n215 , n200 );
nand ( n217 , n6 , n17 );
nand ( n218 , n1 , n22 );
xor ( n219 , n217 , n218 );
nand ( n220 , n5 , n18 );
and ( n221 , n219 , n220 );
and ( n222 , n217 , n218 );
or ( n223 , n221 , n222 );
xor ( n224 , n216 , n223 );
not ( n225 , n191 );
not ( n226 , n188 );
and ( n227 , n225 , n226 );
and ( n228 , n188 , n191 );
nor ( n229 , n227 , n228 );
not ( n230 , n229 );
nand ( n231 , n4 , n21 );
nand ( n232 , n3 , n22 );
nor ( n233 , n231 , n232 );
not ( n234 , n233 );
not ( n235 , n231 );
not ( n236 , n232 );
or ( n237 , n235 , n236 );
nand ( n238 , n2 , n23 );
not ( n239 , n238 );
nand ( n240 , n237 , n239 );
nand ( n241 , n234 , n240 );
not ( n242 , n241 );
not ( n243 , n242 );
and ( n244 , n230 , n243 );
and ( n245 , n229 , n242 );
xor ( n246 , n178 , n179 );
xor ( n247 , n246 , n181 );
nor ( n248 , n245 , n247 );
nor ( n249 , n244 , n248 );
xor ( n250 , n184 , n186 );
xor ( n251 , n250 , n192 );
xor ( n252 , n249 , n251 );
xor ( n253 , n217 , n218 );
xor ( n254 , n253 , n220 );
and ( n255 , n252 , n254 );
and ( n256 , n249 , n251 );
or ( n257 , n255 , n256 );
and ( n258 , n224 , n257 );
and ( n259 , n216 , n223 );
or ( n260 , n258 , n259 );
xor ( n261 , n214 , n260 );
not ( n262 , n261 );
xor ( n263 , n216 , n223 );
xor ( n264 , n263 , n257 );
xor ( n265 , n249 , n251 );
xor ( n266 , n265 , n254 );
nand ( n267 , n7 , n17 );
not ( n268 , n267 );
nand ( n269 , n1 , n23 );
not ( n270 , n269 );
and ( n271 , n268 , n270 );
and ( n272 , n267 , n269 );
nand ( n273 , n5 , n20 );
nand ( n274 , n6 , n19 );
xor ( n275 , n273 , n274 );
nand ( n276 , n7 , n18 );
and ( n277 , n275 , n276 );
and ( n278 , n273 , n274 );
or ( n279 , n277 , n278 );
nor ( n280 , n272 , n279 );
nor ( n281 , n271 , n280 );
xor ( n282 , n266 , n281 );
not ( n283 , n238 );
xor ( n284 , n232 , n231 );
not ( n285 , n284 );
and ( n286 , n283 , n285 );
and ( n287 , n238 , n284 );
nor ( n288 , n286 , n287 );
not ( n289 , n288 );
nand ( n290 , n4 , n22 );
nand ( n291 , n3 , n23 );
nor ( n292 , n290 , n291 );
not ( n293 , n292 );
not ( n294 , n290 );
not ( n295 , n291 );
or ( n296 , n294 , n295 );
nand ( n297 , n2 , n24 );
not ( n298 , n297 );
nand ( n299 , n296 , n298 );
nand ( n300 , n293 , n299 );
not ( n301 , n300 );
xor ( n302 , n273 , n274 );
xor ( n303 , n302 , n276 );
nand ( n304 , n301 , n303 );
and ( n305 , n289 , n304 );
nor ( n306 , n301 , n303 );
nor ( n307 , n305 , n306 );
xor ( n308 , n267 , n269 );
not ( n309 , n308 );
not ( n310 , n279 );
and ( n311 , n309 , n310 );
and ( n312 , n308 , n279 );
nor ( n313 , n311 , n312 );
xor ( n314 , n307 , n313 );
not ( n315 , n247 );
not ( n316 , n229 );
not ( n317 , n241 );
or ( n318 , n316 , n317 );
or ( n319 , n229 , n241 );
nand ( n320 , n318 , n319 );
not ( n321 , n320 );
and ( n322 , n315 , n321 );
and ( n323 , n247 , n320 );
nor ( n324 , n322 , n323 );
and ( n325 , n314 , n324 );
and ( n326 , n307 , n313 );
or ( n327 , n325 , n326 );
and ( n328 , n282 , n327 );
and ( n329 , n266 , n281 );
or ( n330 , n328 , n329 );
xor ( n331 , n264 , n330 );
not ( n332 , n331 );
xor ( n333 , n266 , n281 );
xor ( n334 , n333 , n327 );
nand ( n335 , n8 , n17 );
nand ( n336 , n1 , n24 );
xor ( n337 , n335 , n336 );
nand ( n338 , n4 , n23 );
nand ( n339 , n3 , n24 );
nor ( n340 , n338 , n339 );
not ( n341 , n340 );
nand ( n342 , n5 , n21 );
nand ( n343 , n341 , n342 );
not ( n344 , n343 );
not ( n345 , n291 );
not ( n346 , n290 );
not ( n347 , n346 );
or ( n348 , n345 , n347 );
or ( n349 , n346 , n291 );
nand ( n350 , n348 , n349 );
and ( n351 , n350 , n298 );
not ( n352 , n350 );
and ( n353 , n352 , n297 );
nor ( n354 , n351 , n353 );
not ( n355 , n354 );
or ( n356 , n344 , n355 );
not ( n357 , n342 );
nand ( n358 , n357 , n340 );
nand ( n359 , n356 , n358 );
and ( n360 , n337 , n359 );
not ( n361 , n337 );
not ( n362 , n359 );
and ( n363 , n361 , n362 );
xor ( n364 , n300 , n303 );
xnor ( n365 , n364 , n288 );
nor ( n366 , n363 , n365 );
nor ( n367 , n360 , n366 );
xor ( n368 , n307 , n313 );
xor ( n369 , n368 , n324 );
xor ( n370 , n367 , n369 );
or ( n371 , n335 , n336 );
and ( n372 , n370 , n371 );
and ( n373 , n367 , n369 );
or ( n374 , n372 , n373 );
xor ( n375 , n334 , n374 );
not ( n376 , n375 );
xor ( n377 , n367 , n369 );
xor ( n378 , n377 , n371 );
nand ( n379 , n6 , n20 );
nand ( n380 , n7 , n19 );
xor ( n381 , n379 , n380 );
nand ( n382 , n8 , n18 );
xor ( n383 , n381 , n382 );
nand ( n384 , n5 , n22 );
not ( n385 , n338 );
not ( n386 , n385 );
not ( n387 , n339 );
and ( n388 , n386 , n387 );
not ( n389 , n338 );
and ( n390 , n339 , n389 );
nor ( n391 , n388 , n390 );
nor ( n392 , n384 , n391 );
not ( n393 , n392 );
not ( n394 , n384 );
not ( n395 , n391 );
or ( n396 , n394 , n395 );
nand ( n397 , n6 , n22 );
not ( n398 , n397 );
not ( n399 , n398 );
nand ( n400 , n5 , n23 );
not ( n401 , n400 );
not ( n402 , n401 );
or ( n403 , n399 , n402 );
not ( n404 , n397 );
not ( n405 , n400 );
or ( n406 , n404 , n405 );
nand ( n407 , n4 , n24 );
not ( n408 , n407 );
nand ( n409 , n406 , n408 );
nand ( n410 , n403 , n409 );
nand ( n411 , n396 , n410 );
nand ( n412 , n393 , n411 );
not ( n413 , n412 );
nand ( n414 , n383 , n413 );
and ( n415 , n340 , n342 );
not ( n416 , n340 );
and ( n417 , n416 , n357 );
nor ( n418 , n415 , n417 );
not ( n419 , n354 );
and ( n420 , n418 , n419 );
not ( n421 , n418 );
and ( n422 , n421 , n354 );
or ( n423 , n420 , n422 );
not ( n424 , n423 );
and ( n425 , n414 , n424 );
not ( n426 , n383 );
and ( n427 , n426 , n412 );
nor ( n428 , n425 , n427 );
xor ( n429 , n379 , n380 );
and ( n430 , n429 , n382 );
and ( n431 , n379 , n380 );
or ( n432 , n430 , n431 );
xor ( n433 , n428 , n432 );
not ( n434 , n359 );
xor ( n435 , n337 , n434 );
xnor ( n436 , n435 , n365 );
and ( n437 , n433 , n436 );
and ( n438 , n428 , n432 );
or ( n439 , n437 , n438 );
and ( n440 , n378 , n439 );
not ( n441 , n378 );
not ( n442 , n439 );
and ( n443 , n441 , n442 );
nor ( n444 , n440 , n443 );
not ( n445 , n444 );
nand ( n446 , n7 , n20 );
nand ( n447 , n6 , n21 );
nor ( n448 , n446 , n447 );
not ( n449 , n448 );
xor ( n450 , n426 , n412 );
and ( n451 , n450 , n424 );
not ( n452 , n450 );
and ( n453 , n452 , n423 );
nor ( n454 , n451 , n453 );
not ( n455 , n454 );
or ( n456 , n449 , n455 );
or ( n457 , n448 , n454 );
and ( n458 , n446 , n447 );
not ( n459 , n446 );
not ( n460 , n447 );
and ( n461 , n459 , n460 );
or ( n462 , n458 , n461 );
not ( n463 , n462 );
not ( n464 , n463 );
xor ( n465 , n384 , n410 );
xnor ( n466 , n465 , n391 );
not ( n467 , n466 );
not ( n468 , n467 );
or ( n469 , n464 , n468 );
not ( n470 , n462 );
not ( n471 , n466 );
or ( n472 , n470 , n471 );
nand ( n473 , n7 , n21 );
not ( n474 , n473 );
not ( n475 , n474 );
nand ( n476 , n7 , n22 );
not ( n477 , n476 );
not ( n478 , n477 );
nand ( n479 , n6 , n23 );
not ( n480 , n479 );
not ( n481 , n480 );
or ( n482 , n478 , n481 );
not ( n483 , n479 );
not ( n484 , n476 );
or ( n485 , n483 , n484 );
nand ( n486 , n5 , n24 );
not ( n487 , n486 );
nand ( n488 , n485 , n487 );
nand ( n489 , n482 , n488 );
not ( n490 , n489 );
or ( n491 , n475 , n490 );
not ( n492 , n473 );
not ( n493 , n489 );
not ( n494 , n493 );
or ( n495 , n492 , n494 );
nand ( n496 , n5 , n23 );
nand ( n497 , n6 , n22 );
xor ( n498 , n496 , n497 );
and ( n499 , n498 , n408 );
not ( n500 , n498 );
not ( n501 , n408 );
and ( n502 , n500 , n501 );
nor ( n503 , n499 , n502 );
nand ( n504 , n495 , n503 );
nand ( n505 , n491 , n504 );
nand ( n506 , n472 , n505 );
nand ( n507 , n469 , n506 );
nand ( n508 , n457 , n507 );
nand ( n509 , n456 , n508 );
xor ( n510 , n428 , n432 );
xor ( n511 , n510 , n436 );
xnor ( n512 , n509 , n511 );
not ( n513 , n512 );
and ( n514 , n8 , n21 );
not ( n515 , n514 );
nand ( n516 , n8 , n22 );
not ( n517 , n516 );
not ( n518 , n517 );
nand ( n519 , n7 , n23 );
not ( n520 , n519 );
not ( n521 , n520 );
or ( n522 , n518 , n521 );
not ( n523 , n516 );
not ( n524 , n519 );
or ( n525 , n523 , n524 );
nand ( n526 , n6 , n24 );
not ( n527 , n526 );
nand ( n528 , n525 , n527 );
nand ( n529 , n522 , n528 );
not ( n530 , n529 );
or ( n531 , n515 , n530 );
or ( n532 , n514 , n529 );
nand ( n533 , n5 , n24 );
nand ( n534 , n6 , n23 );
xor ( n535 , n533 , n534 );
not ( n536 , n476 );
xor ( n537 , n535 , n536 );
nand ( n538 , n532 , n537 );
nand ( n539 , n531 , n538 );
nand ( n540 , n8 , n20 );
not ( n541 , n540 );
and ( n542 , n539 , n541 );
not ( n543 , n539 );
and ( n544 , n543 , n540 );
nor ( n545 , n542 , n544 );
not ( n546 , n473 );
not ( n547 , n489 );
or ( n548 , n546 , n547 );
or ( n549 , n473 , n489 );
nand ( n550 , n548 , n549 );
not ( n551 , n503 );
and ( n552 , n550 , n551 );
not ( n553 , n550 );
and ( n554 , n553 , n503 );
nor ( n555 , n552 , n554 );
not ( n556 , n555 );
not ( n557 , n556 );
and ( n558 , n545 , n557 );
not ( n559 , n545 );
and ( n560 , n559 , n556 );
nor ( n561 , n558 , n560 );
not ( n562 , n561 );
nand ( n563 , n8 , n23 );
not ( n564 , n563 );
nand ( n565 , n7 , n24 );
not ( n566 , n565 );
and ( n567 , n564 , n566 );
not ( n568 , n567 );
not ( n569 , n519 );
not ( n570 , n517 );
or ( n571 , n569 , n570 );
or ( n572 , n517 , n519 );
nand ( n573 , n571 , n572 );
and ( n574 , n573 , n526 );
not ( n575 , n573 );
and ( n576 , n575 , n527 );
nor ( n577 , n574 , n576 );
nor ( n578 , n568 , n577 );
xor ( n579 , n514 , n529 );
not ( n580 , n537 );
xor ( n581 , n579 , n580 );
not ( n582 , n581 );
and ( n583 , n578 , n582 );
and ( n584 , n562 , n583 );
not ( n585 , n584 );
nand ( n586 , n8 , n19 );
not ( n587 , n586 );
xor ( n588 , n462 , n505 );
xnor ( n589 , n588 , n466 );
nand ( n590 , n540 , n555 );
and ( n591 , n590 , n539 );
nor ( n592 , n540 , n555 );
nor ( n593 , n591 , n592 );
xnor ( n594 , n589 , n593 );
not ( n595 , n594 );
not ( n596 , n595 );
or ( n597 , n587 , n596 );
not ( n598 , n586 );
nand ( n599 , n598 , n594 );
nand ( n600 , n597 , n599 );
not ( n601 , n600 );
or ( n602 , n585 , n601 );
not ( n603 , n586 );
nand ( n604 , n603 , n595 );
nand ( n605 , n602 , n604 );
not ( n606 , n605 );
nor ( n607 , n589 , n593 );
not ( n608 , n607 );
not ( n609 , n448 );
xor ( n610 , n609 , n507 );
xnor ( n611 , n610 , n454 );
not ( n612 , n611 );
not ( n613 , n612 );
or ( n614 , n608 , n613 );
not ( n615 , n607 );
nand ( n616 , n615 , n611 );
nand ( n617 , n614 , n616 );
not ( n618 , n617 );
or ( n619 , n606 , n618 );
nand ( n620 , n607 , n611 );
nand ( n621 , n619 , n620 );
not ( n622 , n621 );
or ( n623 , n513 , n622 );
not ( n624 , n509 );
or ( n625 , n624 , n511 );
nand ( n626 , n623 , n625 );
not ( n627 , n626 );
or ( n628 , n445 , n627 );
not ( n629 , n378 );
nand ( n630 , n442 , n629 );
nand ( n631 , n628 , n630 );
not ( n632 , n631 );
or ( n633 , n376 , n632 );
or ( n634 , n374 , n334 );
nand ( n635 , n633 , n634 );
not ( n636 , n635 );
or ( n637 , n332 , n636 );
or ( n638 , n330 , n264 );
nand ( n639 , n637 , n638 );
not ( n640 , n639 );
or ( n641 , n262 , n640 );
or ( n642 , n260 , n214 );
nand ( n643 , n641 , n642 );
not ( n644 , n643 );
or ( n645 , n212 , n644 );
or ( n646 , n177 , n210 );
nand ( n647 , n645 , n646 );
not ( n648 , n647 );
or ( n649 , n175 , n648 );
or ( n650 , n173 , n171 );
nand ( n651 , n649 , n650 );
or ( n652 , n137 , n136 );
nand ( n653 , t_0 , n652 );
nand ( n654 , n12 , n25 );
nand ( n655 , n10 , n27 );
xor ( n656 , n654 , n655 );
nand ( n657 , n11 , n26 );
and ( n658 , n656 , n657 );
and ( n659 , n654 , n655 );
or ( n660 , n658 , n659 );
nand ( n661 , n10 , n26 );
xor ( n662 , n660 , n661 );
nand ( n663 , n11 , n25 );
and ( n664 , n662 , n663 );
and ( n665 , n660 , n661 );
or ( n666 , n664 , n665 );
nand ( n667 , n9 , n26 );
xor ( n668 , n666 , n667 );
nand ( n669 , n10 , n25 );
and ( n670 , n668 , n669 );
and ( n671 , n666 , n667 );
or ( n672 , n670 , n671 );
nand ( n673 , n9 , n25 );
xor ( n674 , n672 , n673 );
not ( n675 , n674 );
nand ( n676 , n10 , n29 );
nand ( n677 , n11 , n28 );
xor ( n678 , n676 , n677 );
nand ( n679 , n12 , n27 );
and ( n680 , n678 , n679 );
and ( n681 , n676 , n677 );
or ( n682 , n680 , n681 );
nand ( n683 , n10 , n28 );
xor ( n684 , n682 , n683 );
nand ( n685 , n11 , n27 );
and ( n686 , n684 , n685 );
and ( n687 , n682 , n683 );
or ( n688 , n686 , n687 );
nand ( n689 , n13 , n25 );
nand ( n690 , n9 , n29 );
xor ( n691 , n689 , n690 );
nand ( n692 , n12 , n26 );
and ( n693 , n691 , n692 );
and ( n694 , n689 , n690 );
or ( n695 , n693 , n694 );
xor ( n696 , n688 , n695 );
xor ( n697 , n654 , n655 );
xor ( n698 , n697 , n657 );
and ( n699 , n696 , n698 );
and ( n700 , n688 , n695 );
or ( n701 , n699 , n700 );
nand ( n702 , n9 , n27 );
xor ( n703 , n701 , n702 );
xor ( n704 , n660 , n661 );
xor ( n705 , n704 , n663 );
and ( n706 , n703 , n705 );
and ( n707 , n701 , n702 );
or ( n708 , n706 , n707 );
xor ( n709 , n666 , n667 );
xor ( n710 , n709 , n669 );
xor ( n711 , n708 , n710 );
xor ( n712 , n701 , n702 );
xor ( n713 , n712 , n705 );
nand ( n714 , n10 , n30 );
not ( n715 , n714 );
nand ( n716 , n12 , n28 );
nand ( n717 , n11 , n29 );
nand ( n718 , n716 , n717 );
and ( n719 , n715 , n718 );
nor ( n720 , n716 , n717 );
nor ( n721 , n719 , n720 );
nand ( n722 , n14 , n26 );
nand ( n723 , n13 , n27 );
or ( n724 , n722 , n723 );
xor ( n725 , n721 , n724 );
xor ( n726 , n676 , n677 );
xor ( n727 , n726 , n679 );
and ( n728 , n725 , n727 );
and ( n729 , n721 , n724 );
or ( n730 , n728 , n729 );
xor ( n731 , n682 , n683 );
xor ( n732 , n731 , n685 );
xor ( n733 , n730 , n732 );
xor ( n734 , n689 , n690 );
xor ( n735 , n734 , n692 );
and ( n736 , n733 , n735 );
and ( n737 , n730 , n732 );
or ( n738 , n736 , n737 );
nand ( n739 , n9 , n28 );
xor ( n740 , n738 , n739 );
xor ( n741 , n688 , n695 );
xor ( n742 , n741 , n698 );
and ( n743 , n740 , n742 );
and ( n744 , n738 , n739 );
or ( n745 , n743 , n744 );
xor ( n746 , n713 , n745 );
not ( n747 , n746 );
xor ( n748 , n730 , n732 );
xor ( n749 , n748 , n735 );
nand ( n750 , n14 , n25 );
nand ( n751 , n9 , n30 );
xor ( n752 , n750 , n751 );
nand ( n753 , n13 , n26 );
and ( n754 , n752 , n753 );
and ( n755 , n750 , n751 );
or ( n756 , n754 , n755 );
xor ( n757 , n749 , n756 );
and ( n758 , n722 , n723 );
not ( n759 , n722 );
not ( n760 , n723 );
and ( n761 , n759 , n760 );
or ( n762 , n758 , n761 );
nand ( n763 , n12 , n29 );
not ( n764 , n763 );
nand ( n765 , n11 , n30 );
not ( n766 , n765 );
nand ( n767 , n764 , n766 );
not ( n768 , n763 );
not ( n769 , n765 );
or ( n770 , n768 , n769 );
nand ( n771 , n10 , n31 );
not ( n772 , n771 );
nand ( n773 , n770 , n772 );
nand ( n774 , n767 , n773 );
not ( n775 , n774 );
nand ( n776 , n762 , n775 );
xor ( n777 , n717 , n716 );
and ( n778 , n777 , n714 );
not ( n779 , n777 );
and ( n780 , n779 , n715 );
nor ( n781 , n778 , n780 );
not ( n782 , n781 );
and ( n783 , n776 , n782 );
nor ( n784 , n762 , n775 );
nor ( n785 , n783 , n784 );
xor ( n786 , n721 , n724 );
xor ( n787 , n786 , n727 );
xor ( n788 , n785 , n787 );
xor ( n789 , n750 , n751 );
xor ( n790 , n789 , n753 );
and ( n791 , n788 , n790 );
and ( n792 , n785 , n787 );
or ( n793 , n791 , n792 );
and ( n794 , n757 , n793 );
and ( n795 , n749 , n756 );
or ( n796 , n794 , n795 );
xor ( n797 , n738 , n739 );
xor ( n798 , n797 , n742 );
xor ( n799 , n796 , n798 );
not ( n800 , n799 );
xor ( n801 , n749 , n756 );
xor ( n802 , n801 , n793 );
xor ( n803 , n785 , n787 );
xor ( n804 , n803 , n790 );
nand ( n805 , n15 , n25 );
not ( n806 , n805 );
nand ( n807 , n9 , n31 );
not ( n808 , n807 );
and ( n809 , n806 , n808 );
and ( n810 , n805 , n807 );
nand ( n811 , n15 , n26 );
not ( n812 , n811 );
nand ( n813 , n14 , n27 );
not ( n814 , n813 );
and ( n815 , n812 , n814 );
nand ( n816 , n13 , n28 );
not ( n817 , n816 );
nand ( n818 , n811 , n813 );
and ( n819 , n817 , n818 );
nor ( n820 , n815 , n819 );
nor ( n821 , n810 , n820 );
nor ( n822 , n809 , n821 );
xor ( n823 , n804 , n822 );
not ( n824 , n771 );
not ( n825 , n765 );
not ( n826 , n764 );
or ( n827 , n825 , n826 );
or ( n828 , n764 , n765 );
nand ( n829 , n827 , n828 );
not ( n830 , n829 );
and ( n831 , n824 , n830 );
and ( n832 , n771 , n829 );
nor ( n833 , n831 , n832 );
not ( n834 , n833 );
nand ( n835 , n12 , n30 );
not ( n836 , n835 );
not ( n837 , n836 );
nand ( n838 , n11 , n31 );
not ( n839 , n838 );
not ( n840 , n839 );
or ( n841 , n837 , n840 );
nand ( n842 , n10 , n32 );
not ( n843 , n842 );
nand ( n844 , n835 , n838 );
nand ( n845 , n843 , n844 );
nand ( n846 , n841 , n845 );
not ( n847 , n846 );
not ( n848 , n816 );
xor ( n849 , n813 , n811 );
not ( n850 , n849 );
or ( n851 , n848 , n850 );
or ( n852 , n816 , n849 );
nand ( n853 , n851 , n852 );
not ( n854 , n853 );
nand ( n855 , n847 , n854 );
and ( n856 , n834 , n855 );
and ( n857 , n846 , n853 );
nor ( n858 , n856 , n857 );
xor ( n859 , n805 , n807 );
not ( n860 , n859 );
not ( n861 , n820 );
and ( n862 , n860 , n861 );
and ( n863 , n859 , n820 );
nor ( n864 , n862 , n863 );
xor ( n865 , n858 , n864 );
not ( n866 , n762 );
not ( n867 , n774 );
or ( n868 , n866 , n867 );
or ( n869 , n762 , n774 );
nand ( n870 , n868 , n869 );
and ( n871 , n870 , n781 );
not ( n872 , n870 );
and ( n873 , n872 , n782 );
nor ( n874 , n871 , n873 );
and ( n875 , n865 , n874 );
and ( n876 , n858 , n864 );
or ( n877 , n875 , n876 );
and ( n878 , n823 , n877 );
and ( n879 , n804 , n822 );
or ( n880 , n878 , n879 );
xor ( n881 , n802 , n880 );
not ( n882 , n881 );
nand ( n883 , n16 , n25 );
nand ( n884 , n9 , n32 );
nor ( n885 , n883 , n884 );
not ( n886 , n885 );
not ( n887 , n886 );
xnor ( n888 , n883 , n884 );
not ( n889 , n888 );
nand ( n890 , n13 , n29 );
nand ( n891 , n12 , n31 );
nand ( n892 , n11 , n32 );
nor ( n893 , n891 , n892 );
not ( n894 , n893 );
nand ( n895 , n890 , n894 );
not ( n896 , n895 );
not ( n897 , n838 );
not ( n898 , n835 );
not ( n899 , n898 );
or ( n900 , n897 , n899 );
or ( n901 , n836 , n838 );
nand ( n902 , n900 , n901 );
and ( n903 , n902 , n843 );
not ( n904 , n902 );
and ( n905 , n904 , n842 );
nor ( n906 , n903 , n905 );
not ( n907 , n906 );
or ( n908 , n896 , n907 );
not ( n909 , n890 );
nand ( n910 , n909 , n893 );
nand ( n911 , n908 , n910 );
nand ( n912 , n889 , n911 );
not ( n913 , n888 );
not ( n914 , n911 );
not ( n915 , n914 );
or ( n916 , n913 , n915 );
xor ( n917 , n846 , n853 );
and ( n918 , n917 , n834 );
not ( n919 , n917 );
and ( n920 , n919 , n833 );
nor ( n921 , n918 , n920 );
nand ( n922 , n916 , n921 );
and ( n923 , n912 , n922 );
not ( n924 , n923 );
and ( n925 , n887 , n924 );
and ( n926 , n886 , n923 );
xor ( n927 , n858 , n864 );
xor ( n928 , n927 , n874 );
nor ( n929 , n926 , n928 );
nor ( n930 , n925 , n929 );
xor ( n931 , n804 , n822 );
xor ( n932 , n931 , n877 );
xor ( n933 , n930 , n932 );
not ( n934 , n933 );
not ( n935 , n885 );
not ( n936 , n923 );
or ( n937 , n935 , n936 );
or ( n938 , n885 , n923 );
nand ( n939 , n937 , n938 );
not ( n940 , n939 );
not ( n941 , n928 );
and ( n942 , n940 , n941 );
and ( n943 , n928 , n939 );
nor ( n944 , n942 , n943 );
nand ( n945 , n14 , n28 );
nand ( n946 , n15 , n27 );
xor ( n947 , n945 , n946 );
nand ( n948 , n16 , n26 );
and ( n949 , n947 , n948 );
and ( n950 , n945 , n946 );
or ( n951 , n949 , n950 );
not ( n952 , n921 );
not ( n953 , n888 );
not ( n954 , n911 );
and ( n955 , n953 , n954 );
and ( n956 , n888 , n911 );
nor ( n957 , n955 , n956 );
xnor ( n958 , n952 , n957 );
nor ( n959 , n951 , n958 );
and ( n960 , n951 , n958 );
xor ( n961 , n945 , n946 );
xor ( n962 , n961 , n948 );
not ( n963 , n909 );
not ( n964 , n894 );
or ( n965 , n963 , n964 );
nand ( n966 , n890 , n893 );
nand ( n967 , n965 , n966 );
not ( n968 , n906 );
and ( n969 , n967 , n968 );
not ( n970 , n967 );
and ( n971 , n970 , n906 );
nor ( n972 , n969 , n971 );
nor ( n973 , n962 , n972 );
not ( n974 , n973 );
not ( n975 , n962 );
not ( n976 , n972 );
or ( n977 , n975 , n976 );
nand ( n978 , n13 , n30 );
not ( n979 , n978 );
not ( n980 , n979 );
not ( n981 , n891 );
not ( n982 , n981 );
nand ( n983 , n11 , n32 );
not ( n984 , n983 );
and ( n985 , n982 , n984 );
and ( n986 , n892 , n981 );
nor ( n987 , n985 , n986 );
not ( n988 , n987 );
not ( n989 , n988 );
or ( n990 , n980 , n989 );
not ( n991 , n978 );
not ( n992 , n987 );
or ( n993 , n991 , n992 );
nand ( n994 , n14 , n30 );
not ( n995 , n994 );
not ( n996 , n995 );
nand ( n997 , n13 , n31 );
not ( n998 , n997 );
not ( n999 , n998 );
or ( n1000 , n996 , n999 );
not ( n1001 , n994 );
not ( n1002 , n997 );
or ( n1003 , n1001 , n1002 );
nand ( n1004 , n12 , n32 );
not ( n1005 , n1004 );
nand ( n1006 , n1003 , n1005 );
nand ( n1007 , n1000 , n1006 );
nand ( n1008 , n993 , n1007 );
nand ( n1009 , n990 , n1008 );
nand ( n1010 , n977 , n1009 );
nand ( n1011 , n974 , n1010 );
not ( n1012 , n1011 );
nor ( n1013 , n960 , n1012 );
nor ( n1014 , n959 , n1013 );
and ( n1015 , n944 , n1014 );
not ( n1016 , n944 );
not ( n1017 , n1014 );
and ( n1018 , n1016 , n1017 );
nor ( n1019 , n1015 , n1018 );
not ( n1020 , n1019 );
nand ( n1021 , n15 , n28 );
nand ( n1022 , n14 , n29 );
or ( n1023 , n1021 , n1022 );
not ( n1024 , n1023 );
not ( n1025 , n962 );
not ( n1026 , n1009 );
and ( n1027 , n1025 , n1026 );
and ( n1028 , n962 , n1009 );
nor ( n1029 , n1027 , n1028 );
not ( n1030 , n972 );
and ( n1031 , n1029 , n1030 );
not ( n1032 , n1029 );
and ( n1033 , n1032 , n972 );
nor ( n1034 , n1031 , n1033 );
not ( n1035 , n1034 );
and ( n1036 , n1024 , n1035 );
and ( n1037 , n1023 , n1034 );
and ( n1038 , n1021 , n1022 );
not ( n1039 , n1021 );
not ( n1040 , n1022 );
and ( n1041 , n1039 , n1040 );
or ( n1042 , n1038 , n1041 );
not ( n1043 , n1042 );
not ( n1044 , n1043 );
xor ( n1045 , n978 , n1007 );
xnor ( n1046 , n1045 , n987 );
not ( n1047 , n1046 );
not ( n1048 , n1047 );
or ( n1049 , n1044 , n1048 );
not ( n1050 , n1042 );
not ( n1051 , n1046 );
or ( n1052 , n1050 , n1051 );
nand ( n1053 , n15 , n29 );
not ( n1054 , n1053 );
not ( n1055 , n1054 );
nand ( n1056 , n15 , n30 );
not ( n1057 , n1056 );
not ( n1058 , n1057 );
nand ( n1059 , n14 , n31 );
not ( n1060 , n1059 );
not ( n1061 , n1060 );
or ( n1062 , n1058 , n1061 );
not ( n1063 , n1056 );
not ( n1064 , n1059 );
or ( n1065 , n1063 , n1064 );
nand ( n1066 , n13 , n32 );
not ( n1067 , n1066 );
nand ( n1068 , n1065 , n1067 );
nand ( n1069 , n1062 , n1068 );
not ( n1070 , n1069 );
or ( n1071 , n1055 , n1070 );
or ( n1072 , n1054 , n1069 );
nand ( n1073 , n14 , n30 );
not ( n1074 , n1073 );
not ( n1075 , n1074 );
nand ( n1076 , n13 , n31 );
not ( n1077 , n1076 );
and ( n1078 , n1075 , n1077 );
and ( n1079 , n1076 , n1074 );
nor ( n1080 , n1078 , n1079 );
nand ( n1081 , n12 , n32 );
and ( n1082 , n1080 , n1081 );
not ( n1083 , n1080 );
not ( n1084 , n1081 );
and ( n1085 , n1083 , n1084 );
nor ( n1086 , n1082 , n1085 );
nand ( n1087 , n1072 , n1086 );
nand ( n1088 , n1071 , n1087 );
nand ( n1089 , n1052 , n1088 );
nand ( n1090 , n1049 , n1089 );
not ( n1091 , n1090 );
nor ( n1092 , n1037 , n1091 );
nor ( n1093 , n1036 , n1092 );
not ( n1094 , n1093 );
not ( n1095 , n1094 );
xor ( n1096 , n951 , n1011 );
xor ( n1097 , n1096 , n958 );
not ( n1098 , n1097 );
not ( n1099 , n1098 );
or ( n1100 , n1095 , n1099 );
nand ( n1101 , n1093 , n1097 );
nand ( n1102 , n1100 , n1101 );
not ( n1103 , n1102 );
nand ( n1104 , n16 , n28 );
not ( n1105 , n1104 );
not ( n1106 , n1105 );
xor ( n1107 , n1054 , n1069 );
xnor ( n1108 , n1107 , n1086 );
not ( n1109 , n1108 );
not ( n1110 , n1109 );
or ( n1111 , n1106 , n1110 );
not ( n1112 , n1104 );
not ( n1113 , n1108 );
or ( n1114 , n1112 , n1113 );
and ( n1115 , n16 , n29 );
not ( n1116 , n1115 );
nand ( n1117 , n14 , n31 );
not ( n1118 , n1117 );
not ( n1119 , n1118 );
nand ( n1120 , n15 , n30 );
not ( n1121 , n1120 );
and ( n1122 , n1119 , n1121 );
not ( n1123 , n1117 );
and ( n1124 , n1120 , n1123 );
nor ( n1125 , n1122 , n1124 );
not ( n1126 , n1067 );
and ( n1127 , n1125 , n1126 );
not ( n1128 , n1125 );
and ( n1129 , n1128 , n1067 );
nor ( n1130 , n1127 , n1129 );
not ( n1131 , n1130 );
or ( n1132 , n1116 , n1131 );
or ( n1133 , n1115 , n1130 );
nand ( n1134 , n16 , n30 );
not ( n1135 , n1134 );
not ( n1136 , n1135 );
nand ( n1137 , n14 , n32 );
not ( n1138 , n1137 );
not ( n1139 , n1138 );
or ( n1140 , n1136 , n1139 );
not ( n1141 , n1134 );
not ( n1142 , n1137 );
or ( n1143 , n1141 , n1142 );
nand ( n1144 , n15 , n31 );
not ( n1145 , n1144 );
nand ( n1146 , n1143 , n1145 );
nand ( n1147 , n1140 , n1146 );
nand ( n1148 , n1133 , n1147 );
nand ( n1149 , n1132 , n1148 );
nand ( n1150 , n1114 , n1149 );
nand ( n1151 , n1111 , n1150 );
not ( n1152 , n1151 );
xor ( n1153 , n1042 , n1088 );
xnor ( n1154 , n1153 , n1046 );
nor ( n1155 , n1152 , n1154 );
buf ( n1156 , n1155 );
not ( n1157 , n1156 );
not ( n1158 , n1090 );
not ( n1159 , n1023 );
and ( n1160 , n1158 , n1159 );
and ( n1161 , n1023 , n1090 );
nor ( n1162 , n1160 , n1161 );
and ( n1163 , n1162 , n1034 );
not ( n1164 , n1162 );
and ( n1165 , n1164 , n1035 );
nor ( n1166 , n1163 , n1165 );
not ( n1167 , n1166 );
not ( n1168 , n1167 );
or ( n1169 , n1157 , n1168 );
not ( n1170 , n1155 );
nand ( n1171 , n1170 , n1166 );
nand ( n1172 , n1169 , n1171 );
not ( n1173 , n1172 );
not ( n1174 , n1134 );
not ( n1175 , n1144 );
not ( n1176 , n1175 );
or ( n1177 , n1174 , n1176 );
or ( n1178 , n1145 , n1134 );
nand ( n1179 , n1177 , n1178 );
and ( n1180 , n1179 , n1137 );
not ( n1181 , n1179 );
and ( n1182 , n1181 , n1138 );
nor ( n1183 , n1180 , n1182 );
not ( n1184 , n1183 );
nand ( n1185 , n16 , n31 );
not ( n1186 , n1185 );
nand ( n1187 , n15 , n32 );
not ( n1188 , n1187 );
and ( n1189 , n1186 , n1188 );
nand ( n1190 , n1184 , n1189 );
xor ( n1191 , n1147 , n1115 );
xnor ( n1192 , n1191 , n1130 );
or ( n1193 , n1190 , n1192 );
and ( n1194 , n1149 , n1105 );
not ( n1195 , n1149 );
and ( n1196 , n1195 , n1104 );
nor ( n1197 , n1194 , n1196 );
and ( n1198 , n1197 , n1108 );
not ( n1199 , n1197 );
and ( n1200 , n1199 , n1109 );
nor ( n1201 , n1198 , n1200 );
nor ( n1202 , n1193 , n1201 );
not ( n1203 , n1202 );
nand ( n1204 , n16 , n27 );
not ( n1205 , n1204 );
not ( n1206 , n1154 );
and ( n1207 , n1152 , n1206 );
not ( n1208 , n1152 );
and ( n1209 , n1208 , n1154 );
nor ( n1210 , n1207 , n1209 );
not ( n1211 , n1210 );
not ( n1212 , n1211 );
or ( n1213 , n1205 , n1212 );
not ( n1214 , n1204 );
nand ( n1215 , n1214 , n1210 );
nand ( n1216 , n1213 , n1215 );
not ( n1217 , n1216 );
or ( n1218 , n1203 , n1217 );
not ( n1219 , n1204 );
nand ( n1220 , n1219 , n1211 );
nand ( n1221 , n1218 , n1220 );
not ( n1222 , n1221 );
or ( n1223 , n1173 , n1222 );
nand ( n1224 , n1156 , n1166 );
nand ( n1225 , n1223 , n1224 );
not ( n1226 , n1225 );
or ( n1227 , n1103 , n1226 );
nand ( n1228 , n1094 , n1097 );
nand ( n1229 , n1227 , n1228 );
not ( n1230 , n1229 );
or ( n1231 , n1020 , n1230 );
not ( n1232 , n944 );
nand ( n1233 , n1017 , n1232 );
nand ( n1234 , n1231 , n1233 );
not ( n1235 , n1234 );
or ( n1236 , n934 , n1235 );
or ( n1237 , n930 , n932 );
nand ( n1238 , n1236 , n1237 );
not ( n1239 , n1238 );
or ( n1240 , n882 , n1239 );
or ( n1241 , n880 , n802 );
nand ( n1242 , n1240 , n1241 );
not ( n1243 , n1242 );
or ( n1244 , n800 , n1243 );
or ( n1245 , n796 , n798 );
nand ( n1246 , n1244 , n1245 );
not ( n1247 , n1246 );
or ( n1248 , n747 , n1247 );
or ( n1249 , n713 , n745 );
nand ( n1250 , n1248 , n1249 );
or ( n1251 , n710 , n708 );
nand ( n1252 , t_2 , n1251 );
not ( n1253 , n1252 );
or ( n1254 , n675 , n1253 );
or ( n1255 , n673 , n672 );
nand ( n1256 , n1254 , n1255 );
not ( n1257 , n1256 );
or ( n1258 , n1257 , n653 );
nand ( n1259 , t_3 , n1258 );
not ( n1260 , n25 );
and ( n1261 , n17 , n1260 );
not ( n1262 , n17 );
and ( n1263 , n25 , n1262 );
nor ( n1264 , n1261 , n1263 );
not ( n1265 , n1264 );
not ( n1266 , n18 );
not ( n1267 , n26 );
or ( n1268 , n1266 , n1267 );
or ( n1269 , n18 , n26 );
not ( n1270 , n19 );
not ( n1271 , n27 );
or ( n1272 , n1270 , n1271 );
or ( n1273 , n19 , n27 );
not ( n1274 , n20 );
not ( n1275 , n28 );
or ( n1276 , n1274 , n1275 );
or ( n1277 , n20 , n28 );
not ( n1278 , n21 );
not ( n1279 , n29 );
or ( n1280 , n1278 , n1279 );
or ( n1281 , n21 , n29 );
not ( n1282 , n22 );
not ( n1283 , n30 );
or ( n1284 , n1282 , n1283 );
not ( n1285 , n22 );
not ( n1286 , n1285 );
not ( n1287 , n30 );
not ( n1288 , n1287 );
or ( n1289 , n1286 , n1288 );
not ( n1290 , n23 );
not ( n1291 , n31 );
or ( n1292 , n1290 , n1291 );
nand ( n1293 , n24 , n32 );
not ( n1294 , n1293 );
nor ( n1295 , n23 , n31 );
not ( n1296 , n1295 );
nand ( n1297 , n1294 , n1296 );
nand ( n1298 , n1292 , n1297 );
nand ( n1299 , n1289 , n1298 );
nand ( n1300 , n1284 , n1299 );
nand ( n1301 , n1281 , n1300 );
nand ( n1302 , n1280 , n1301 );
nand ( n1303 , n1277 , n1302 );
nand ( n1304 , n1276 , n1303 );
nand ( n1305 , n1273 , n1304 );
nand ( n1306 , n1272 , n1305 );
nand ( n1307 , n1269 , n1306 );
nand ( n1308 , n1268 , n1307 );
not ( n1309 , n1308 );
or ( n1310 , n1265 , n1309 );
or ( n1311 , n1264 , n1308 );
nand ( n1312 , n1310 , n1311 );
nand ( n1313 , n8 , n24 );
not ( n1314 , n1313 );
not ( n1315 , n1314 );
nand ( n1316 , n16 , n32 );
not ( n1317 , n1316 );
and ( n1318 , n1315 , n1317 );
and ( n1319 , n1316 , n1314 );
nor ( n1320 , n1318 , n1319 );
not ( n1321 , n1320 );
buf ( n1322 , n1321 );
buf ( n1323 , n1322 );
not ( n1324 , n1323 );
not ( n1325 , n1324 );
not ( n1326 , n1325 );
not ( n1327 , n1326 );
not ( n1328 , n1327 );
and ( n1329 , n1312 , n1328 );
not ( n1330 , n1328 );
not ( n1331 , n9 );
and ( n1332 , n1 , n1331 );
not ( n1333 , n1 );
and ( n1334 , n9 , n1333 );
nor ( n1335 , n1332 , n1334 );
not ( n1336 , n1335 );
not ( n1337 , n2 );
not ( n1338 , n10 );
or ( n1339 , n1337 , n1338 );
or ( n1340 , n2 , n10 );
not ( n1341 , n3 );
not ( n1342 , n11 );
or ( n1343 , n1341 , n1342 );
or ( n1344 , n3 , n11 );
not ( n1345 , n4 );
not ( n1346 , n12 );
or ( n1347 , n1345 , n1346 );
or ( n1348 , n4 , n12 );
not ( n1349 , n5 );
not ( n1350 , n13 );
or ( n1351 , n1349 , n1350 );
or ( n1352 , n5 , n13 );
not ( n1353 , n6 );
not ( n1354 , n14 );
or ( n1355 , n1353 , n1354 );
or ( n1356 , n6 , n14 );
not ( n1357 , n7 );
not ( n1358 , n15 );
or ( n1359 , n1357 , n1358 );
nand ( n1360 , n8 , n16 );
not ( n1361 , n1360 );
nor ( n1362 , n7 , n15 );
not ( n1363 , n1362 );
nand ( n1364 , n1361 , n1363 );
nand ( n1365 , n1359 , n1364 );
nand ( n1366 , n1356 , n1365 );
nand ( n1367 , n1355 , n1366 );
nand ( n1368 , n1352 , n1367 );
nand ( n1369 , n1351 , n1368 );
nand ( n1370 , n1348 , n1369 );
nand ( n1371 , n1347 , n1370 );
nand ( n1372 , n1344 , n1371 );
nand ( n1373 , n1343 , n1372 );
nand ( n1374 , n1340 , n1373 );
nand ( n1375 , n1339 , n1374 );
not ( n1376 , n1375 );
or ( n1377 , n1336 , n1376 );
or ( n1378 , n1335 , n1375 );
nand ( n1379 , n1377 , n1378 );
and ( n1380 , n1330 , n1379 );
nor ( n1381 , n1329 , n1380 );
not ( n1382 , n512 );
not ( n1383 , n621 );
not ( n1384 , n1383 );
or ( n1385 , n1382 , n1384 );
not ( n1386 , n512 );
nand ( n1387 , n1386 , n621 );
nand ( n1388 , n1385 , n1387 );
not ( n1389 , n1388 );
nand ( n1390 , n1381 , n1389 );
xnor ( n1391 , n3 , n11 );
not ( n1392 , n1391 );
not ( n1393 , n1371 );
or ( n1394 , n1392 , n1393 );
or ( n1395 , n1391 , n1371 );
nand ( n1396 , n1394 , n1395 );
and ( n1397 , n1325 , n1396 );
not ( n1398 , n1325 );
xnor ( n1399 , n19 , n27 );
not ( n1400 , n1399 );
not ( n1401 , n1304 );
or ( n1402 , n1400 , n1401 );
or ( n1403 , n1399 , n1304 );
nand ( n1404 , n1402 , n1403 );
and ( n1405 , n1398 , n1404 );
nor ( n1406 , n1397 , n1405 );
not ( n1407 , n1406 );
xnor ( n1408 , n4 , n12 );
not ( n1409 , n1408 );
not ( n1410 , n1369 );
or ( n1411 , n1409 , n1410 );
or ( n1412 , n1408 , n1369 );
nand ( n1413 , n1411 , n1412 );
and ( n1414 , n1323 , n1413 );
not ( n1415 , n1323 );
xnor ( n1416 , n20 , n28 );
not ( n1417 , n1416 );
not ( n1418 , n1302 );
or ( n1419 , n1417 , n1418 );
or ( n1420 , n1416 , n1302 );
nand ( n1421 , n1419 , n1420 );
and ( n1422 , n1415 , n1421 );
nor ( n1423 , n1414 , n1422 );
not ( n1424 , n1423 );
not ( n1425 , n583 );
not ( n1426 , n561 );
and ( n1427 , n1425 , n1426 );
and ( n1428 , n583 , n561 );
nor ( n1429 , n1427 , n1428 );
not ( n1430 , n1429 );
and ( n1431 , n1424 , n1430 );
and ( n1432 , n1423 , n1429 );
xnor ( n1433 , n5 , n13 );
not ( n1434 , n1433 );
not ( n1435 , n1367 );
or ( n1436 , n1434 , n1435 );
or ( n1437 , n1433 , n1367 );
nand ( n1438 , n1436 , n1437 );
and ( n1439 , n1323 , n1438 );
not ( n1440 , n1323 );
xnor ( n1441 , n21 , n29 );
not ( n1442 , n1441 );
not ( n1443 , n1300 );
or ( n1444 , n1442 , n1443 );
or ( n1445 , n1441 , n1300 );
nand ( n1446 , n1444 , n1445 );
and ( n1447 , n1440 , n1446 );
nor ( n1448 , n1439 , n1447 );
not ( n1449 , n1448 );
not ( n1450 , n578 );
and ( n1451 , n581 , n1450 );
not ( n1452 , n581 );
and ( n1453 , n1452 , n578 );
or ( n1454 , n1451 , n1453 );
not ( n1455 , n1454 );
and ( n1456 , n1449 , n1455 );
nand ( n1457 , n1448 , n1454 );
and ( n1458 , n577 , n567 );
not ( n1459 , n577 );
and ( n1460 , n1459 , n568 );
nor ( n1461 , n1458 , n1460 );
xor ( n1462 , n14 , n6 );
xor ( n1463 , n1365 , n1462 );
and ( n1464 , n1322 , n1463 );
not ( n1465 , n1322 );
and ( n1466 , n30 , n1285 );
not ( n1467 , n30 );
and ( n1468 , n1467 , n22 );
nor ( n1469 , n1466 , n1468 );
not ( n1470 , n1469 );
not ( n1471 , n1298 );
or ( n1472 , n1470 , n1471 );
or ( n1473 , n1469 , n1298 );
nand ( n1474 , n1472 , n1473 );
and ( n1475 , n1465 , n1474 );
nor ( n1476 , n1464 , n1475 );
and ( n1477 , n1461 , n1476 );
and ( n1478 , n564 , n565 );
not ( n1479 , n564 );
and ( n1480 , n1479 , n566 );
nor ( n1481 , n1478 , n1480 );
not ( n1482 , n1360 );
xor ( n1483 , n7 , n15 );
not ( n1484 , n1483 );
or ( n1485 , n1482 , n1484 );
or ( n1486 , n1360 , n1483 );
nand ( n1487 , n1485 , n1486 );
and ( n1488 , n1322 , n1487 );
not ( n1489 , n1293 );
xor ( n1490 , n23 , n31 );
not ( n1491 , n1490 );
or ( n1492 , n1489 , n1491 );
or ( n1493 , n1293 , n1490 );
nand ( n1494 , n1492 , n1493 );
and ( n1495 , n1320 , n1494 );
nor ( n1496 , n1488 , n1495 );
nor ( n1497 , n1481 , n1496 );
and ( n1498 , n1481 , n1496 );
not ( n1499 , n1314 );
not ( n1500 , n1499 );
xor ( n1501 , n16 , n8 );
not ( n1502 , n1501 );
not ( n1503 , n1321 );
or ( n1504 , n1502 , n1503 );
xor ( n1505 , n24 , n32 );
nand ( n1506 , n1505 , n1320 );
nand ( n1507 , n1504 , n1506 );
nand ( n1508 , n1500 , n1507 );
nor ( n1509 , n1498 , n1508 );
nor ( n1510 , n1497 , n1509 );
or ( n1511 , n1477 , n1510 );
or ( n1512 , n1461 , n1476 );
nand ( n1513 , n1511 , n1512 );
and ( n1514 , n1457 , n1513 );
nor ( n1515 , n1456 , n1514 );
nor ( n1516 , n1432 , n1515 );
nor ( n1517 , n1431 , n1516 );
not ( n1518 , n1517 );
and ( n1519 , n1407 , n1518 );
and ( n1520 , n1406 , n1517 );
buf ( n1521 , n600 );
and ( n1522 , n1521 , n584 );
not ( n1523 , n1521 );
not ( n1524 , n584 );
and ( n1525 , n1523 , n1524 );
nor ( n1526 , n1522 , n1525 );
not ( n1527 , n1526 );
nor ( n1528 , n1520 , n1527 );
nor ( n1529 , n1519 , n1528 );
not ( n1530 , n1326 );
xnor ( n1531 , n2 , n10 );
not ( n1532 , n1531 );
not ( n1533 , n1373 );
or ( n1534 , n1532 , n1533 );
or ( n1535 , n1531 , n1373 );
nand ( n1536 , n1534 , n1535 );
and ( n1537 , n1530 , n1536 );
not ( n1538 , n1530 );
xnor ( n1539 , n18 , n26 );
not ( n1540 , n1539 );
not ( n1541 , n1306 );
or ( n1542 , n1540 , n1541 );
or ( n1543 , n1539 , n1306 );
nand ( n1544 , n1542 , n1543 );
and ( n1545 , n1538 , n1544 );
nor ( n1546 , n1537 , n1545 );
not ( n1547 , n1546 );
not ( n1548 , n617 );
and ( n1549 , n605 , n1548 );
not ( n1550 , n605 );
and ( n1551 , n1550 , n617 );
or ( n1552 , n1549 , n1551 );
nor ( n1553 , n1547 , n1552 );
or ( n1554 , n1529 , n1553 );
not ( n1555 , n1546 );
nand ( n1556 , n1555 , n1552 );
nand ( n1557 , n1554 , n1556 );
and ( n1558 , n1390 , n1557 );
nor ( n1559 , n1381 , n1389 );
nor ( n1560 , n1558 , n1559 );
and ( n1561 , n1333 , n1331 );
and ( n1562 , n1 , n9 );
nor ( n1563 , n1562 , n1375 );
nor ( n1564 , n1561 , n1328 , n1563 );
and ( n1565 , n1262 , n1260 );
and ( n1566 , n17 , n25 );
nor ( n1567 , n1566 , n1308 );
nor ( n1568 , n1565 , n1327 , n1567 );
or ( n1569 , n1564 , n1568 );
not ( n1570 , n444 );
not ( n1571 , n626 );
not ( n1572 , n1571 );
or ( n1573 , n1570 , n1572 );
not ( n1574 , n444 );
nand ( n1575 , n1574 , n626 );
nand ( n1576 , n1573 , n1575 );
nor ( n1577 , n1569 , n1576 );
or ( n1578 , n1560 , n1577 );
nand ( n1579 , n1576 , n1569 );
nand ( n1580 , n1578 , n1579 );
xor ( n1581 , n375 , n631 );
and ( n1582 , n1580 , n1581 );
xor ( n1583 , n331 , n635 );
nand ( n1584 , n1582 , n1583 );
not ( n1585 , n1584 );
buf ( n1586 , n639 );
xor ( n1587 , n1586 , n261 );
nand ( n1588 , n1585 , n1587 );
not ( n1589 , n1588 );
buf ( n1590 , n643 );
xor ( n1591 , n1590 , n211 );
nand ( n1592 , n1589 , n1591 );
not ( n1593 , n1592 );
xor ( n1594 , n647 , n174 );
nand ( n1595 , n1593 , n1594 );
not ( n1596 , n1595 );
not ( n1597 , n138 );
nand ( n1598 , n1597 , n651 );
nand ( n1599 , t_1 , n1598 );
nand ( n1600 , n1596 , n1599 );
not ( n1601 , n1600 );
and ( n1602 , n1259 , n1601 );
not ( n1603 , n1259 );
and ( n1604 , n1603 , n1600 );
nor ( n1605 , n1602 , n1604 );
not ( n1606 , n1595 );
not ( n1607 , n1599 );
or ( n1608 , n1606 , n1607 );
or ( n1609 , n1595 , n1599 );
nand ( n1610 , n1608 , n1609 );
not ( n1611 , n1252 );
and ( n1612 , n1611 , n674 );
not ( n1613 , n1611 );
not ( n1614 , n674 );
and ( n1615 , n1613 , n1614 );
nor ( n1616 , n1612 , n1615 );
not ( n1617 , n1616 );
not ( n1618 , n1617 );
not ( n1619 , n1618 );
and ( n1620 , n1610 , n1619 );
not ( n1621 , n1610 );
and ( n1622 , n1621 , n1618 );
nor ( n1623 , n1620 , n1622 );
buf ( n1624 , n1234 );
buf ( n1625 , n933 );
xor ( n1626 , n1624 , n1625 );
nor ( n1627 , n1499 , n1316 );
not ( n1628 , n1627 );
xor ( n1629 , n1186 , n1188 );
not ( n1630 , n1629 );
not ( n1631 , n1481 );
or ( n1632 , n1630 , n1631 );
or ( n1633 , n1481 , n1629 );
nand ( n1634 , n1632 , n1633 );
not ( n1635 , n1634 );
not ( n1636 , n1635 );
or ( n1637 , n1628 , n1636 );
not ( n1638 , n1627 );
nand ( n1639 , n1638 , n1634 );
nand ( n1640 , n1637 , n1639 );
not ( n1641 , n1640 );
not ( n1642 , n1641 );
not ( n1643 , n1642 );
not ( n1644 , n1643 );
not ( n1645 , n1644 );
not ( n1646 , n1645 );
not ( n1647 , n1646 );
buf ( n1648 , n1229 );
and ( n1649 , n1648 , n1019 );
not ( n1650 , n1648 );
not ( n1651 , n1019 );
and ( n1652 , n1650 , n1651 );
nor ( n1653 , n1649 , n1652 );
nand ( n1654 , n1647 , n1653 );
nand ( n1655 , t_7 , n1654 );
buf ( n1656 , n1653 );
nor ( n1657 , n1655 , n1656 );
and ( n1658 , n1221 , n1172 );
not ( n1659 , n1221 );
not ( n1660 , n1172 );
and ( n1661 , n1659 , n1660 );
nor ( n1662 , n1658 , n1661 );
not ( n1663 , n1662 );
not ( n1664 , n1663 );
not ( n1665 , n1664 );
not ( n1666 , n1645 );
not ( n1667 , n1666 );
not ( n1668 , n1552 );
or ( n1669 , n1667 , n1668 );
nand ( n1670 , n1645 , n1662 );
nand ( n1671 , n1669 , n1670 );
not ( n1672 , n1671 );
or ( n1673 , n1665 , n1672 );
or ( n1674 , n1664 , n1671 );
and ( n1675 , n1216 , n1202 );
not ( n1676 , n1216 );
not ( n1677 , n1202 );
and ( n1678 , n1676 , n1677 );
nor ( n1679 , n1675 , n1678 );
not ( n1680 , n1679 );
not ( n1681 , n1680 );
not ( n1682 , n1681 );
and ( n1683 , n1644 , n1526 );
not ( n1684 , n1644 );
and ( n1685 , n1684 , n1679 );
nor ( n1686 , n1683 , n1685 );
not ( n1687 , n1686 );
not ( n1688 , n1687 );
or ( n1689 , n1682 , n1688 );
xor ( n1690 , n1201 , n1193 );
not ( n1691 , n1690 );
and ( n1692 , n1643 , n1690 );
not ( n1693 , n1429 );
and ( n1694 , n1642 , n1693 );
nor ( n1695 , n1692 , n1694 );
not ( n1696 , n1695 );
not ( n1697 , n1696 );
or ( n1698 , n1691 , n1697 );
xor ( n1699 , n1190 , n1192 );
not ( n1700 , n1699 );
and ( n1701 , n1641 , n1699 );
not ( n1702 , n1454 );
and ( n1703 , n1640 , n1702 );
nor ( n1704 , n1701 , n1703 );
not ( n1705 , n1704 );
not ( n1706 , n1705 );
or ( n1707 , n1700 , n1706 );
not ( n1708 , n1699 );
nand ( n1709 , n1708 , n1704 );
xor ( n1710 , n1189 , n1183 );
and ( n1711 , n1640 , n1461 );
not ( n1712 , n1640 );
and ( n1713 , n1712 , n1710 );
or ( n1714 , n1711 , n1713 );
and ( n1715 , n1710 , n1714 );
not ( n1716 , n1629 );
not ( n1717 , n1716 );
not ( n1718 , n1481 );
and ( n1719 , n1718 , n1640 );
nor ( n1720 , n1716 , n1640 );
nor ( n1721 , n1719 , n1720 );
not ( n1722 , n1721 );
and ( n1723 , n1717 , n1722 );
not ( n1724 , n1316 );
not ( n1725 , n1724 );
or ( n1726 , n1725 , n1640 );
nand ( n1727 , n1500 , n1640 );
nand ( n1728 , n1726 , n1727 );
not ( n1729 , n1728 );
not ( n1730 , n1724 );
nor ( n1731 , n1729 , n1730 );
nand ( n1732 , n1716 , n1721 );
and ( n1733 , n1731 , n1732 );
nor ( n1734 , n1723 , n1733 );
or ( n1735 , n1715 , n1734 );
or ( n1736 , n1710 , n1714 );
nand ( n1737 , n1735 , n1736 );
nand ( n1738 , n1709 , n1737 );
nand ( n1739 , n1707 , n1738 );
not ( n1740 , n1690 );
nand ( n1741 , n1740 , n1695 );
nand ( n1742 , n1739 , n1741 );
nand ( n1743 , n1698 , n1742 );
nand ( n1744 , n1680 , n1686 );
nand ( n1745 , n1743 , n1744 );
nand ( n1746 , n1689 , n1745 );
nand ( n1747 , n1674 , n1746 );
nand ( n1748 , n1673 , n1747 );
xor ( n1749 , n1225 , n1102 );
not ( n1750 , n1749 );
not ( n1751 , n1646 );
not ( n1752 , n1388 );
or ( n1753 , n1751 , n1752 );
not ( n1754 , n1646 );
nand ( n1755 , n1754 , n1749 );
nand ( n1756 , n1753 , n1755 );
not ( n1757 , n1756 );
nand ( n1758 , n1750 , n1757 );
and ( n1759 , n1748 , n1758 );
and ( n1760 , n1749 , n1756 );
nor ( n1761 , n1759 , n1760 );
or ( n1762 , n1657 , n1761 );
nand ( n1763 , n1655 , n1656 );
nand ( n1764 , n1762 , n1763 );
nand ( n1765 , n1626 , n1764 );
not ( n1766 , n1765 );
and ( n1767 , n1246 , n746 );
not ( n1768 , n1246 );
not ( n1769 , n746 );
and ( n1770 , n1768 , n1769 );
nor ( n1771 , n1767 , n1770 );
xor ( n1772 , n1242 , n799 );
buf ( n1773 , n1238 );
buf ( n1774 , n881 );
xnor ( n1775 , n1773 , n1774 );
not ( n1776 , n1775 );
nand ( n1777 , n1766 , n1771 , n1772 , n1776 );
not ( n1778 , n711 );
and ( n1779 , n1250 , n1778 );
not ( n1780 , n1250 );
and ( n1781 , n1780 , n711 );
nor ( n1782 , n1779 , n1781 );
nor ( n1783 , n1777 , n1782 );
buf ( n1784 , n1599 );
nor ( n1785 , t_4 , n1784 );
not ( n1786 , n653 );
nor ( n1787 , n1600 , n1786 );
buf ( n1788 , n1592 );
not ( n1789 , n1788 );
and ( n1790 , n1594 , n1789 );
not ( n1791 , n1594 );
and ( n1792 , n1791 , n1788 );
nor ( n1793 , n1790 , n1792 );
buf ( n1794 , n1782 );
not ( n1795 , n1794 );
and ( n1796 , n1793 , n1795 );
not ( n1797 , n1793 );
and ( n1798 , n1797 , n1794 );
nor ( n1799 , n1796 , n1798 );
not ( n1800 , n1783 );
nor ( n1801 , n1800 , n1616 );
buf ( n1802 , n1777 );
not ( n1803 , n1794 );
and ( n1804 , n1802 , n1803 );
not ( n1805 , n1802 );
and ( n1806 , n1805 , n1794 );
nor ( n1807 , n1804 , n1806 );
nor ( n1808 , n1807 , n1594 );
buf ( n1809 , n1765 );
nor ( n1810 , n1775 , n1809 );
nand ( n1811 , n1772 , n1810 );
and ( n1812 , n1811 , n1771 );
not ( n1813 , n1811 );
not ( n1814 , n1771 );
and ( n1815 , n1813 , n1814 );
nor ( n1816 , n1812 , n1815 );
buf ( n1817 , n1591 );
buf ( n1818 , n1817 );
nor ( n1819 , n1816 , n1818 );
and ( n1820 , n1817 , n1588 );
not ( n1821 , n1817 );
and ( n1822 , n1821 , n1589 );
nor ( n1823 , n1820 , n1822 );
and ( n1824 , n1823 , n1814 );
not ( n1825 , n1823 );
and ( n1826 , n1825 , n1771 );
nor ( n1827 , n1824 , n1826 );
not ( n1828 , n1772 );
and ( n1829 , n1810 , n1828 );
not ( n1830 , n1810 );
and ( n1831 , n1830 , n1772 );
nor ( n1832 , n1829 , n1831 );
nor ( n1833 , n1832 , n1587 );
xnor ( n1834 , n1584 , n1587 );
and ( n1835 , n1834 , n1772 );
not ( n1836 , n1834 );
and ( n1837 , n1836 , n1828 );
nor ( n1838 , n1835 , n1837 );
buf ( n1839 , n1809 );
and ( n1840 , n1839 , n1776 );
not ( n1841 , n1839 );
and ( n1842 , n1841 , n1775 );
nor ( n1843 , n1840 , n1842 );
nor ( n1844 , n1583 , n1843 );
buf ( n1845 , n1764 );
not ( n1846 , n1626 );
and ( n1847 , n1845 , n1846 );
not ( n1848 , n1845 );
and ( n1849 , n1848 , n1626 );
nor ( n1850 , n1847 , n1849 );
nor ( n1851 , n1581 , n1850 );
and ( n1852 , n1583 , n1776 );
not ( n1853 , n1583 );
and ( n1854 , n1853 , n1775 );
nor ( n1855 , n1852 , n1854 );
and ( n1856 , n1855 , n1582 );
not ( n1857 , n1855 );
not ( n1858 , n1582 );
and ( n1859 , n1857 , n1858 );
nor ( n1860 , n1856 , n1859 );
buf ( n1861 , n1655 );
and ( n1862 , n1861 , n1656 );
nor ( n1863 , n1862 , t_5 );
and ( n1864 , n1761 , n1863 );
nor ( n1865 , n1864 , t_6 );
nor ( n1866 , n1576 , n1865 );
and ( n1867 , n1581 , n1846 );
not ( n1868 , n1581 );
and ( n1869 , n1868 , n1626 );
nor ( n1870 , n1867 , n1869 );
buf ( n1871 , n1580 );
not ( n1872 , n1871 );
and ( n1873 , n1870 , n1872 );
not ( n1874 , n1870 );
and ( n1875 , n1874 , n1871 );
nor ( n1876 , n1873 , n1875 );
not ( n1877 , n1560 );
and ( n1878 , n1877 , n1656 );
not ( n1879 , n1877 );
not ( n1880 , n1656 );
and ( n1881 , n1879 , n1880 );
nor ( n1882 , n1878 , n1881 );
xnor ( n1883 , n1576 , n1569 );
not ( n1884 , n1883 );
and ( n1885 , n1882 , n1884 );
not ( n1886 , n1882 );
and ( n1887 , n1886 , n1883 );
nor ( n1888 , n1885 , n1887 );
xor ( n1889 , n1749 , n1756 );
xnor ( n1890 , n1748 , n1889 );
nor ( n1891 , n1388 , n1890 );
and ( n1892 , n1557 , n1749 );
not ( n1893 , n1557 );
and ( n1894 , n1893 , n1750 );
nor ( n1895 , n1892 , n1894 );
and ( n1896 , n1381 , n1388 );
not ( n1897 , n1381 );
and ( n1898 , n1897 , n1389 );
nor ( n1899 , n1896 , n1898 );
or ( n1900 , n1895 , n1899 );
nand ( n1901 , n1895 , n1899 );
nand ( n1902 , n1900 , n1901 );
not ( n1903 , n1663 );
and ( n1904 , n1671 , n1903 );
not ( n1905 , n1671 );
and ( n1906 , n1905 , n1663 );
nor ( n1907 , n1904 , n1906 );
not ( n1908 , n1746 );
xor ( n1909 , n1907 , n1908 );
nor ( n1910 , n1909 , n1552 );
not ( n1911 , n1527 );
not ( n1912 , n1743 );
not ( n1913 , n1680 );
and ( n1914 , n1687 , n1913 );
not ( n1915 , n1687 );
and ( n1916 , n1915 , n1680 );
nor ( n1917 , n1914 , n1916 );
and ( n1918 , n1912 , n1917 );
nor ( n1919 , n1912 , n1917 );
nor ( n1920 , n1918 , n1919 );
nor ( n1921 , n1911 , n1920 );
xor ( n1922 , n1546 , n1552 );
not ( n1923 , n1922 );
and ( n1924 , n1529 , n1663 );
not ( n1925 , n1529 );
and ( n1926 , n1925 , n1664 );
nor ( n1927 , n1924 , n1926 );
not ( n1928 , n1927 );
or ( n1929 , n1923 , n1928 );
or ( n1930 , n1922 , n1927 );
nand ( n1931 , n1929 , n1930 );
xor ( n1932 , n1406 , n1911 );
not ( n1933 , n1932 );
buf ( n1934 , n1517 );
not ( n1935 , n1934 );
not ( n1936 , n1913 );
or ( n1937 , n1935 , n1936 );
or ( n1938 , n1934 , n1913 );
nand ( n1939 , n1937 , n1938 );
not ( n1940 , n1939 );
or ( n1941 , n1933 , n1940 );
or ( n1942 , n1932 , n1939 );
nand ( n1943 , n1941 , n1942 );
and ( n1944 , n1696 , n1690 );
not ( n1945 , n1696 );
and ( n1946 , n1945 , n1740 );
nor ( n1947 , n1944 , n1946 );
xnor ( n1948 , n1739 , n1947 );
nor ( n1949 , n1693 , n1948 );
and ( n1950 , n1705 , n1699 );
not ( n1951 , n1705 );
and ( n1952 , n1951 , n1708 );
nor ( n1953 , n1950 , n1952 );
xnor ( n1954 , n1737 , n1953 );
nor ( n1955 , n1702 , n1954 );
and ( n1956 , n1423 , n1693 );
not ( n1957 , n1423 );
and ( n1958 , n1957 , n1429 );
nor ( n1959 , n1956 , n1958 );
not ( n1960 , n1959 );
and ( n1961 , n1515 , n1740 );
not ( n1962 , n1515 );
and ( n1963 , n1962 , n1690 );
nor ( n1964 , n1961 , n1963 );
not ( n1965 , n1964 );
or ( n1966 , n1960 , n1965 );
or ( n1967 , n1959 , n1964 );
nand ( n1968 , n1966 , n1967 );
not ( n1969 , n1461 );
xor ( n1970 , n1710 , n1714 );
xor ( n1971 , n1734 , n1970 );
nor ( n1972 , n1969 , n1971 );
and ( n1973 , n1721 , n1629 );
not ( n1974 , n1721 );
and ( n1975 , n1974 , n1716 );
nor ( n1976 , n1973 , n1975 );
and ( n1977 , n1731 , n1976 );
nor ( n1978 , n1731 , n1976 );
nor ( n1979 , n1977 , n1978 );
nor ( n1980 , n1718 , n1979 );
and ( n1981 , n1448 , n1454 );
not ( n1982 , n1448 );
and ( n1983 , n1982 , n1702 );
nor ( n1984 , n1981 , n1983 );
not ( n1985 , n1984 );
and ( n1986 , n1513 , n1708 );
not ( n1987 , n1513 );
and ( n1988 , n1987 , n1699 );
nor ( n1989 , n1986 , n1988 );
not ( n1990 , n1989 );
or ( n1991 , n1985 , n1990 );
or ( n1992 , n1984 , n1989 );
nand ( n1993 , n1991 , n1992 );
xor ( n1994 , n1730 , n1728 );
nor ( n1995 , n1500 , n1994 );
not ( n1996 , n1508 );
not ( n1997 , n1634 );
not ( n1998 , n1496 );
or ( n1999 , n1997 , n1998 );
or ( n2000 , n1634 , n1496 );
nand ( n2001 , n1999 , n2000 );
not ( n2002 , n2001 );
or ( n2003 , n1996 , n2002 );
or ( n2004 , n1508 , n2001 );
nand ( n2005 , n2003 , n2004 );
and ( n2006 , n1710 , n1461 );
not ( n2007 , n1710 );
and ( n2008 , n2007 , n1969 );
nor ( n2009 , n2006 , n2008 );
and ( n2010 , n1507 , n1325 );
not ( n2011 , n1507 );
and ( n2012 , n2011 , n1324 );
nor ( n2013 , n2010 , n2012 );
xor ( n2014 , n1801 , n1257 );
nor ( n2015 , n2014 , n653 );
xor ( n2016 , n1510 , n1476 );
xor ( n2017 , n2016 , n2009 );
endmodule
