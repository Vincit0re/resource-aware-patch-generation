module top ( g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 , g98 , g99 , g100 , g101 , g102 , g103 , g104 , g105 , g106 , g107 , g108 , g109 , g110 , g111 , g112 , g113 , g114 , g115 , g116 , g117 , g118 , g119 , g120 , g121 , g122 , g123 , g124 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g136 , g137 , g138 , g139 , g140 , g141 , g142 , g143 , g144 , g145 , g146 , g147 , g148 , g149 , g150 , g151 , g152 , g153 , g154 , g155 , g156 , g157 , g158 , g159 , g160 , g161 , g162 , g163 , g164 , g165 , g166 , g167 , g168 , g169 , g170 , g171 , g172 , g173 , g174 , g175 , g176 , g177 , g178 , g179 , g180 , g181 , g182 , g183 , g184 , g185 , g186 , g187 , g188 , g189 , g190 , g191 , g192 , g193 , g194 , g195 , g196 , g197 , g198 , g199 , g200 , g201 , g202 , g203 , g204 , g205 , g206 , g207 , g208 , g209 , g210 , g211 , g212 , g213 , g214 , g215 , g216 , g217 , g218 , g219 , g220 , g221 , g222 , g223 , g224 , g225 , g226 , g227 , g228 , g229 , g230 , g231 , g232 , g233 , g234 , g235 , g236 , g237 , g238 , g239 , g240 , g241 , g242 , g243 , g244 , g245 , g246 , g247 , g248 , g249 , g250 , g251 , g252 , g253 , g254 , g255 , g256 , g257 , g258 , g259 , g260 , g261 , g262 , g263 , g264 , g265 , g266 , g267 , g268 , g269 , g270 , g271 , g272 , g273 , g274 , g275 , g276 , g277 , g278 , g279 , g280 , g281 , g282 , g283 , g284 , g285 , g286 , g287 , g288 , g289 , g290 , g291 , g292 , g293 , g294 , g295 , g296 , g297 , g298 , g299 , g300 , g301 , g302 , g303 , g304 , g305 , g306 , g307 , g308 , g309 , g310 , g311 , g312 , g313 , g314 , g315 , g316 , g317 , g318 , g319 , g320 , g321 , g322 , g323 , g324 , g325 , g326 , g327 , g328 , g329 , g330 , g331 , g332 , g333 , g334 , g335 , g336 , g337 , g338 , g339 , g340 , g341 , g342 , g343 , g344 , g345 , g346 , g347 , g348 , g349 , g350 , g351 , g352 , g353 , g354 , g355 , g356 , g357 , g358 , g359 , g360 , g361 , g362 , g363 , g364 , g365 , g366 , g367 , g368 , g369 , g370 , g371 , g372 , g373 , g374 , g375 , g376 , g377 , g378 , g379 , g380 , g381 , g382 , g383 , g384 , g385 , g386 , g387 , g388 , g389 , g390 , g391 , g392 , g393 , g394 , g395 , g396 , g397 , g398 , g399 , g400 , g401 , g402 , g403 , g404 , g405 , g406 , g407 , g408 , g409 , g410 , g411 , g412 , g413 , g414 , g415 , g416 , g417 , g418 , g419 , g420 , g421 , g422 , g423 , g424 , g425 , g426 , g427 , g428 , g429 , g430 , g431 , g432 , g433 , g434 , g435 , g436 , g437 , g438 , g439 , g440 , g441 , g442 , g443 , g444 , g445 , g446 , g447 , g448 , g449 , g450 , g451 , g452 , g453 , g454 , g455 , g456 , g457 , g458 , g459 , g460 , g461 , g462 , g463 , g464 , g465 , g466 , g467 , g468 , g469 , g470 , g471 , g472 , g473 , g474 , g475 , g476 , g477 , g478 , g479 , g480 , g481 , g482 , g483 , g484 , g485 , g486 , g487 , g488 , g489 , g490 , g491 , g492 , g493 , g494 , g495 , g496 , g497 , g498 , g499 , g500 );
input g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 , g98 , g99 , g100 , g101 , g102 , g103 , g104 , g105 , g106 , g107 , g108 , g109 , g110 , g111 , g112 , g113 , g114 , g115 , g116 , g117 , g118 , g119 , g120 , g121 , g122 , g123 , g124 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g136 , g137 , g138 , g139 , g140 , g141 , g142 , g143 , g144 , g145 , g146 , g147 , g148 , g149 , g150 , g151 , g152 , g153 , g154 , g155 , g156 , g157 , g158 , g159 , g160 , g161 , g162 , g163 , g164 , g165 , g166 , g167 , g168 , g169 , g170 , g171 , g172 , g173 , g174 , g175 , g176 , g177 , g178 , g179 , g180 , g181 , g182 , g183 , g184 , g185 , g186 , g187 , g188 , g189 , g190 , g191 , g192 , g193 , g194 , g195 , g196 , g197 , g198 , g199 , g200 , g201 , g202 , g203 , g204 , g205 , g206 , g207 , g208 , g209 , g210 , g211 , g212 , g213 , g214 , g215 , g216 , g217 , g218 , g219 , g220 , g221 , g222 , g223 , g224 , g225 , g226 , g227 , g228 , g229 , g230 , g231 , g232 , g233 , g234 , g235 , g236 , g237 , g238 , g239 , g240 , g241 , g242 , g243 , g244 , g245 , g246 , g247 , g248 , g249 , g250 , g251 , g252 , g253 , g254 , g255 ;
output g256 , g257 , g258 , g259 , g260 , g261 , g262 , g263 , g264 , g265 , g266 , g267 , g268 , g269 , g270 , g271 , g272 , g273 , g274 , g275 , g276 , g277 , g278 , g279 , g280 , g281 , g282 , g283 , g284 , g285 , g286 , g287 , g288 , g289 , g290 , g291 , g292 , g293 , g294 , g295 , g296 , g297 , g298 , g299 , g300 , g301 , g302 , g303 , g304 , g305 , g306 , g307 , g308 , g309 , g310 , g311 , g312 , g313 , g314 , g315 , g316 , g317 , g318 , g319 , g320 , g321 , g322 , g323 , g324 , g325 , g326 , g327 , g328 , g329 , g330 , g331 , g332 , g333 , g334 , g335 , g336 , g337 , g338 , g339 , g340 , g341 , g342 , g343 , g344 , g345 , g346 , g347 , g348 , g349 , g350 , g351 , g352 , g353 , g354 , g355 , g356 , g357 , g358 , g359 , g360 , g361 , g362 , g363 , g364 , g365 , g366 , g367 , g368 , g369 , g370 , g371 , g372 , g373 , g374 , g375 , g376 , g377 , g378 , g379 , g380 , g381 , g382 , g383 , g384 , g385 , g386 , g387 , g388 , g389 , g390 , g391 , g392 , g393 , g394 , g395 , g396 , g397 , g398 , g399 , g400 , g401 , g402 , g403 , g404 , g405 , g406 , g407 , g408 , g409 , g410 , g411 , g412 , g413 , g414 , g415 , g416 , g417 , g418 , g419 , g420 , g421 , g422 , g423 , g424 , g425 , g426 , g427 , g428 , g429 , g430 , g431 , g432 , g433 , g434 , g435 , g436 , g437 , g438 , g439 , g440 , g441 , g442 , g443 , g444 , g445 , g446 , g447 , g448 , g449 , g450 , g451 , g452 , g453 , g454 , g455 , g456 , g457 , g458 , g459 , g460 , g461 , g462 , g463 , g464 , g465 , g466 , g467 , g468 , g469 , g470 , g471 , g472 , g473 , g474 , g475 , g476 , g477 , g478 , g479 , g480 , g481 , g482 , g483 , g484 , g485 , g486 , g487 , g488 , g489 , g490 , g491 , g492 , g493 , g494 , g495 , g496 , g497 , g498 , g499 , g500 ;

wire n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , 
     n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , 
     n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , 
     n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , 
     n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , 
     n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , 
     n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , 
     n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , 
     n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , 
     n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , 
     n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , 
     n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , 
     n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , 
     n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , 
     n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , 
     n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , 
     n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , 
     n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , 
     n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , 
     n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , 
     n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , 
     n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , 
     n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , 
     n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , 
     n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , 
     n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , 
     n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , 
     n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , 
     n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , 
     n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , 
     n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , 
     n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , 
     n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , 
     n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , 
     n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , 
     n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , 
     n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , 
     n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , 
     n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , 
     n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , 
     n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , 
     n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , 
     n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , 
     n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , 
     n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , 
     n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , 
     n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , 
     n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , 
     n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , 
     n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , 
     n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , 
     n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , 
     n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , 
     n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , 
     n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , 
     n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , 
     n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , 
     n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , 
     n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , 
     n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , 
     n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , 
     n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , 
     n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , 
     n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , 
     n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , 
     n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , 
     n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , 
     n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , 
     n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , 
     n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , 
     n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , 
     n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , 
     n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , 
     n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , 
     n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , 
     n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , 
     n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , 
     n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , 
     n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , 
     n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , 
     n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , 
     n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , 
     n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , 
     n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , 
     n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , 
     n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , 
     n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , 
     n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , 
     n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , 
     n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , 
     n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , 
     n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , 
     n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , 
     n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , 
     n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , 
     n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , 
     n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , 
     n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , 
     n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , 
     n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , 
     n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , 
     n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , 
     n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , 
     n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , 
     n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , 
     n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , 
     n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , 
     n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , 
     n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , 
     n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , 
     n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , 
     n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , 
     n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , 
     n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , 
     n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , 
     n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , 
     n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , 
     n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , 
     n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , 
     n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , 
     n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , 
     n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , 
     n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , 
     n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , 
     n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , 
     n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , 
     n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , 
     n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , 
     n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , 
     n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , 
     n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , 
     n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , 
     n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , 
     n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , 
     n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , 
     n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , 
     n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , 
     n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , 
     n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , 
     n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , 
     n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , 
     n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , 
     n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , 
     n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , 
     n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , 
     n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , 
     n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , 
     n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , 
     n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , 
     n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , 
     n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , 
     n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , 
     n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , 
     n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , 
     n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , 
     n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , 
     n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , 
     n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , 
     n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , 
     n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , 
     n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , 
     n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , 
     n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , 
     n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , 
     n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , 
     n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , 
     n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , 
     n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , 
     n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , 
     n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , 
     n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , 
     n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , 
     n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , 
     n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , 
     n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , 
     n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , 
     n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , 
     n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , 
     n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , 
     n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , 
     n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , 
     n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , 
     n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , 
     n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , 
     n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , 
     n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , 
     n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , 
     n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , 
     n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , 
     n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , 
     n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , 
     n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , 
     n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , 
     n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , 
     n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , 
     n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , 
     n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , 
     n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , 
     n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , 
     n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , 
     n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , 
     n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , 
     n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , 
     n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , 
     n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , 
     n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , 
     n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , 
     n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , 
     n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , 
     n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , 
     n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , 
     n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , 
     n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , 
     n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , 
     n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , 
     n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , 
     n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , 
     n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , 
     n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , 
     n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , 
     n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , 
     n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , 
     n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , 
     n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , 
     n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , 
     n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , 
     n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , 
     n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , 
     n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , 
     n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , 
     n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , 
     n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , 
     n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , 
     n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , 
     n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , 
     n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , 
     n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , 
     n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , 
     n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , 
     n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , 
     n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , 
     n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , 
     n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , 
     n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , 
     n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , 
     n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , 
     n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , 
     n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , 
     n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , 
     n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , 
     n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , 
     n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , 
     n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , 
     n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , 
     n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , 
     n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , 
     n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , 
     n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , 
     n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , 
     n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , 
     n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , 
     n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , 
     n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , 
     n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , 
     n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , 
     n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , 
     n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , 
     n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , 
     n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , 
     n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , 
     n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , 
     n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , 
     n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , 
     n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , 
     n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , 
     n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , 
     n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , 
     n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , 
     n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , 
     n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , 
     n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , 
     n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , 
     n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , 
     n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , 
     n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , 
     n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , 
     n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , 
     n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , 
     n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , 
     n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , 
     n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , 
     n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , 
     n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , 
     n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , 
     n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , 
     n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , 
     n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , 
     n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , 
     n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , 
     n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , 
     n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , 
     n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , 
     n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , 
     n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , 
     n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , 
     n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , 
     n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , 
     n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , 
     n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , 
     n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , 
     n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , 
     n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , 
     n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , 
     n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , 
     n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , 
     n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , 
     n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , 
     n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , 
     n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , 
     n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , 
     n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , 
     n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , 
     n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , 
     n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , 
     n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , 
     n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , 
     n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , 
     n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , 
     n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , 
     n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , 
     n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , 
     n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , 
     n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , 
     n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , 
     n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , 
     n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , 
     n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , 
     n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , 
     n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , 
     n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , 
     n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , 
     n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , 
     n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , 
     n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , 
     n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , 
     n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , 
     n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , 
     n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , 
     n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , 
     n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , 
     n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , 
     n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , 
     n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , 
     n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , 
     n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , 
     n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , 
     n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , 
     n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , 
     n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , 
     n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , 
     n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , 
     n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , 
     n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , 
     n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , 
     n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , 
     n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , 
     n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , 
     n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , 
     n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , 
     n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , 
     n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , 
     n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , 
     n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , 
     n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , 
     n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , 
     n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , 
     n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , 
     n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , 
     n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , 
     n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , 
     n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , 
     n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , 
     n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , 
     n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , 
     n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , 
     n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , 
     n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , 
     n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , 
     n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , 
     n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , 
     n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , 
     n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , 
     n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , 
     n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , 
     n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , 
     n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , 
     n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , 
     n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , 
     n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , 
     n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , 
     n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , 
     n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , 
     n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , 
     n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , 
     n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , 
     n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , 
     n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , 
     n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , 
     n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , 
     n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , 
     n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , 
     n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , 
     n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , 
     n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , 
     n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , 
     n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , 
     n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , 
     n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , 
     n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , 
     n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , 
     n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , 
     n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , 
     n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , 
     n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , 
     n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , 
     n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , 
     n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , 
     n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , 
     n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , 
     n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , 
     n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , 
     n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , 
     n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , 
     n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , 
     n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , 
     n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , 
     n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , 
     n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , 
     n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , 
     n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , 
     n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , 
     n4410 , n4411 , n4412 , n4413 , n4414 ;
buf ( n1  , g0 );
buf ( n2  , g1 );
buf ( n3  , g2 );
buf ( n4  , g3 );
buf ( n5  , g4 );
buf ( n6  , g5 );
buf ( n7  , g6 );
buf ( n8  , g7 );
buf ( n9  , g8 );
buf ( n10  , g9 );
buf ( n11  , g10 );
buf ( n12  , g11 );
buf ( n13  , g12 );
buf ( n14  , g13 );
buf ( n15  , g14 );
buf ( n16  , g15 );
buf ( n17  , g16 );
buf ( n18  , g17 );
buf ( n19  , g18 );
buf ( n20  , g19 );
buf ( n21  , g20 );
buf ( n22  , g21 );
buf ( n23  , g22 );
buf ( n24  , g23 );
buf ( n25  , g24 );
buf ( n26  , g25 );
buf ( n27  , g26 );
buf ( n28  , g27 );
buf ( n29  , g28 );
buf ( n30  , g29 );
buf ( n31  , g30 );
buf ( n32  , g31 );
buf ( n33  , g32 );
buf ( n34  , g33 );
buf ( n35  , g34 );
buf ( n36  , g35 );
buf ( n37  , g36 );
buf ( n38  , g37 );
buf ( n39  , g38 );
buf ( n40  , g39 );
buf ( n41  , g40 );
buf ( n42  , g41 );
buf ( n43  , g42 );
buf ( n44  , g43 );
buf ( n45  , g44 );
buf ( n46  , g45 );
buf ( n47  , g46 );
buf ( n48  , g47 );
buf ( n49  , g48 );
buf ( n50  , g49 );
buf ( n51  , g50 );
buf ( n52  , g51 );
buf ( n53  , g52 );
buf ( n54  , g53 );
buf ( n55  , g54 );
buf ( n56  , g55 );
buf ( n57  , g56 );
buf ( n58  , g57 );
buf ( n59  , g58 );
buf ( n60  , g59 );
buf ( n61  , g60 );
buf ( n62  , g61 );
buf ( n63  , g62 );
buf ( n64  , g63 );
buf ( n65  , g64 );
buf ( n66  , g65 );
buf ( n67  , g66 );
buf ( n68  , g67 );
buf ( n69  , g68 );
buf ( n70  , g69 );
buf ( n71  , g70 );
buf ( n72  , g71 );
buf ( n73  , g72 );
buf ( n74  , g73 );
buf ( n75  , g74 );
buf ( n76  , g75 );
buf ( n77  , g76 );
buf ( n78  , g77 );
buf ( n79  , g78 );
buf ( n80  , g79 );
buf ( n81  , g80 );
buf ( n82  , g81 );
buf ( n83  , g82 );
buf ( n84  , g83 );
buf ( n85  , g84 );
buf ( n86  , g85 );
buf ( n87  , g86 );
buf ( n88  , g87 );
buf ( n89  , g88 );
buf ( n90  , g89 );
buf ( n91  , g90 );
buf ( n92  , g91 );
buf ( n93  , g92 );
buf ( n94  , g93 );
buf ( n95  , g94 );
buf ( n96  , g95 );
buf ( n97  , g96 );
buf ( n98  , g97 );
buf ( n99  , g98 );
buf ( n100  , g99 );
buf ( n101  , g100 );
buf ( n102  , g101 );
buf ( n103  , g102 );
buf ( n104  , g103 );
buf ( n105  , g104 );
buf ( n106  , g105 );
buf ( n107  , g106 );
buf ( n108  , g107 );
buf ( n109  , g108 );
buf ( n110  , g109 );
buf ( n111  , g110 );
buf ( n112  , g111 );
buf ( n113  , g112 );
buf ( n114  , g113 );
buf ( n115  , g114 );
buf ( n116  , g115 );
buf ( n117  , g116 );
buf ( n118  , g117 );
buf ( n119  , g118 );
buf ( n120  , g119 );
buf ( n121  , g120 );
buf ( n122  , g121 );
buf ( n123  , g122 );
buf ( n124  , g123 );
buf ( n125  , g124 );
buf ( n126  , g125 );
buf ( n127  , g126 );
buf ( n128  , g127 );
buf ( n129  , g128 );
buf ( n130  , g129 );
buf ( n131  , g130 );
buf ( n132  , g131 );
buf ( n133  , g132 );
buf ( n134  , g133 );
buf ( n135  , g134 );
buf ( n136  , g135 );
buf ( n137  , g136 );
buf ( n138  , g137 );
buf ( n139  , g138 );
buf ( n140  , g139 );
buf ( n141  , g140 );
buf ( n142  , g141 );
buf ( n143  , g142 );
buf ( n144  , g143 );
buf ( n145  , g144 );
buf ( n146  , g145 );
buf ( n147  , g146 );
buf ( n148  , g147 );
buf ( n149  , g148 );
buf ( n150  , g149 );
buf ( n151  , g150 );
buf ( n152  , g151 );
buf ( n153  , g152 );
buf ( n154  , g153 );
buf ( n155  , g154 );
buf ( n156  , g155 );
buf ( n157  , g156 );
buf ( n158  , g157 );
buf ( n159  , g158 );
buf ( n160  , g159 );
buf ( n161  , g160 );
buf ( n162  , g161 );
buf ( n163  , g162 );
buf ( n164  , g163 );
buf ( n165  , g164 );
buf ( n166  , g165 );
buf ( n167  , g166 );
buf ( n168  , g167 );
buf ( n169  , g168 );
buf ( n170  , g169 );
buf ( n171  , g170 );
buf ( n172  , g171 );
buf ( n173  , g172 );
buf ( n174  , g173 );
buf ( n175  , g174 );
buf ( n176  , g175 );
buf ( n177  , g176 );
buf ( n178  , g177 );
buf ( n179  , g178 );
buf ( n180  , g179 );
buf ( n181  , g180 );
buf ( n182  , g181 );
buf ( n183  , g182 );
buf ( n184  , g183 );
buf ( n185  , g184 );
buf ( n186  , g185 );
buf ( n187  , g186 );
buf ( n188  , g187 );
buf ( n189  , g188 );
buf ( n190  , g189 );
buf ( n191  , g190 );
buf ( n192  , g191 );
buf ( n193  , g192 );
buf ( n194  , g193 );
buf ( n195  , g194 );
buf ( n196  , g195 );
buf ( n197  , g196 );
buf ( n198  , g197 );
buf ( n199  , g198 );
buf ( n200  , g199 );
buf ( n201  , g200 );
buf ( n202  , g201 );
buf ( n203  , g202 );
buf ( n204  , g203 );
buf ( n205  , g204 );
buf ( n206  , g205 );
buf ( n207  , g206 );
buf ( n208  , g207 );
buf ( n209  , g208 );
buf ( n210  , g209 );
buf ( n211  , g210 );
buf ( n212  , g211 );
buf ( n213  , g212 );
buf ( n214  , g213 );
buf ( n215  , g214 );
buf ( n216  , g215 );
buf ( n217  , g216 );
buf ( n218  , g217 );
buf ( n219  , g218 );
buf ( n220  , g219 );
buf ( n221  , g220 );
buf ( n222  , g221 );
buf ( n223  , g222 );
buf ( n224  , g223 );
buf ( n225  , g224 );
buf ( n226  , g225 );
buf ( n227  , g226 );
buf ( n228  , g227 );
buf ( n229  , g228 );
buf ( n230  , g229 );
buf ( n231  , g230 );
buf ( n232  , g231 );
buf ( n233  , g232 );
buf ( n234  , g233 );
buf ( n235  , g234 );
buf ( n236  , g235 );
buf ( n237  , g236 );
buf ( n238  , g237 );
buf ( n239  , g238 );
buf ( n240  , g239 );
buf ( n241  , g240 );
buf ( n242  , g241 );
buf ( n243  , g242 );
buf ( n244  , g243 );
buf ( n245  , g244 );
buf ( n246  , g245 );
buf ( n247  , g246 );
buf ( n248  , g247 );
buf ( n249  , g248 );
buf ( n250  , g249 );
buf ( n251  , g250 );
buf ( n252  , g251 );
buf ( n253  , g252 );
buf ( n254  , g253 );
buf ( n255  , g254 );
buf ( n256  , g255 );
buf ( g256 , n257  );
buf ( g257 , n258  );
buf ( g258 , n259  );
buf ( g259 , n260  );
buf ( g260 , n261  );
buf ( g261 , n262  );
buf ( g262 , n263  );
buf ( g263 , n264  );
buf ( g264 , n265  );
buf ( g265 , n266  );
buf ( g266 , n267  );
buf ( g267 , n268  );
buf ( g268 , n269  );
buf ( g269 , n270  );
buf ( g270 , n271  );
buf ( g271 , n272  );
buf ( g272 , n273  );
buf ( g273 , n274  );
buf ( g274 , n275  );
buf ( g275 , n276  );
buf ( g276 , n277  );
buf ( g277 , n278  );
buf ( g278 , n279  );
buf ( g279 , n280  );
buf ( g280 , n281  );
buf ( g281 , n282  );
buf ( g282 , n283  );
buf ( g283 , n284  );
buf ( g284 , n285  );
buf ( g285 , n286  );
buf ( g286 , n287  );
buf ( g287 , n288  );
buf ( g288 , n289  );
buf ( g289 , n290  );
buf ( g290 , n291  );
buf ( g291 , n292  );
buf ( g292 , n293  );
buf ( g293 , n294  );
buf ( g294 , n295  );
buf ( g295 , n296  );
buf ( g296 , n297  );
buf ( g297 , n298  );
buf ( g298 , n299  );
buf ( g299 , n300  );
buf ( g300 , n301  );
buf ( g301 , n302  );
buf ( g302 , n303  );
buf ( g303 , n304  );
buf ( g304 , n305  );
buf ( g305 , n306  );
buf ( g306 , n307  );
buf ( g307 , n308  );
buf ( g308 , n309  );
buf ( g309 , n310  );
buf ( g310 , n311  );
buf ( g311 , n312  );
buf ( g312 , n313  );
buf ( g313 , n314  );
buf ( g314 , n315  );
buf ( g315 , n316  );
buf ( g316 , n317  );
buf ( g317 , n318  );
buf ( g318 , n319  );
buf ( g319 , n320  );
buf ( g320 , n321  );
buf ( g321 , n322  );
buf ( g322 , n323  );
buf ( g323 , n324  );
buf ( g324 , n325  );
buf ( g325 , n326  );
buf ( g326 , n327  );
buf ( g327 , n328  );
buf ( g328 , n329  );
buf ( g329 , n330  );
buf ( g330 , n331  );
buf ( g331 , n332  );
buf ( g332 , n333  );
buf ( g333 , n334  );
buf ( g334 , n335  );
buf ( g335 , n336  );
buf ( g336 , n337  );
buf ( g337 , n338  );
buf ( g338 , n339  );
buf ( g339 , n340  );
buf ( g340 , n341  );
buf ( g341 , n342  );
buf ( g342 , n343  );
buf ( g343 , n344  );
buf ( g344 , n345  );
buf ( g345 , n346  );
buf ( g346 , n347  );
buf ( g347 , n348  );
buf ( g348 , n349  );
buf ( g349 , n350  );
buf ( g350 , n351  );
buf ( g351 , n352  );
buf ( g352 , n353  );
buf ( g353 , n354  );
buf ( g354 , n355  );
buf ( g355 , n356  );
buf ( g356 , n357  );
buf ( g357 , n358  );
buf ( g358 , n359  );
buf ( g359 , n360  );
buf ( g360 , n361  );
buf ( g361 , n362  );
buf ( g362 , n363  );
buf ( g363 , n364  );
buf ( g364 , n365  );
buf ( g365 , n366  );
buf ( g366 , n367  );
buf ( g367 , n368  );
buf ( g368 , n369  );
buf ( g369 , n370  );
buf ( g370 , n371  );
buf ( g371 , n372  );
buf ( g372 , n373  );
buf ( g373 , n374  );
buf ( g374 , n375  );
buf ( g375 , n376  );
buf ( g376 , n377  );
buf ( g377 , n378  );
buf ( g378 , n379  );
buf ( g379 , n380  );
buf ( g380 , n381  );
buf ( g381 , n382  );
buf ( g382 , n383  );
buf ( g383 , n384  );
buf ( g384 , n385  );
buf ( g385 , n386  );
buf ( g386 , n387  );
buf ( g387 , n388  );
buf ( g388 , n389  );
buf ( g389 , n390  );
buf ( g390 , n391  );
buf ( g391 , n392  );
buf ( g392 , n393  );
buf ( g393 , n394  );
buf ( g394 , n395  );
buf ( g395 , n396  );
buf ( g396 , n397  );
buf ( g397 , n398  );
buf ( g398 , n399  );
buf ( g399 , n400  );
buf ( g400 , n401  );
buf ( g401 , n402  );
buf ( g402 , n403  );
buf ( g403 , n404  );
buf ( g404 , n405  );
buf ( g405 , n406  );
buf ( g406 , n407  );
buf ( g407 , n408  );
buf ( g408 , n409  );
buf ( g409 , n410  );
buf ( g410 , n411  );
buf ( g411 , n412  );
buf ( g412 , n413  );
buf ( g413 , n414  );
buf ( g414 , n415  );
buf ( g415 , n416  );
buf ( g416 , n417  );
buf ( g417 , n418  );
buf ( g418 , n419  );
buf ( g419 , n420  );
buf ( g420 , n421  );
buf ( g421 , n422  );
buf ( g422 , n423  );
buf ( g423 , n424  );
buf ( g424 , n425  );
buf ( g425 , n426  );
buf ( g426 , n427  );
buf ( g427 , n428  );
buf ( g428 , n429  );
buf ( g429 , n430  );
buf ( g430 , n431  );
buf ( g431 , n432  );
buf ( g432 , n433  );
buf ( g433 , n434  );
buf ( g434 , n435  );
buf ( g435 , n436  );
buf ( g436 , n437  );
buf ( g437 , n438  );
buf ( g438 , n439  );
buf ( g439 , n440  );
buf ( g440 , n441  );
buf ( g441 , n442  );
buf ( g442 , n443  );
buf ( g443 , n444  );
buf ( g444 , n445  );
buf ( g445 , n446  );
buf ( g446 , n447  );
buf ( g447 , n448  );
buf ( g448 , n449  );
buf ( g449 , n450  );
buf ( g450 , n451  );
buf ( g451 , n452  );
buf ( g452 , n453  );
buf ( g453 , n454  );
buf ( g454 , n455  );
buf ( g455 , n456  );
buf ( g456 , n457  );
buf ( g457 , n458  );
buf ( g458 , n459  );
buf ( g459 , n460  );
buf ( g460 , n461  );
buf ( g461 , n462  );
buf ( g462 , n463  );
buf ( g463 , n464  );
buf ( g464 , n465  );
buf ( g465 , n466  );
buf ( g466 , n467  );
buf ( g467 , n468  );
buf ( g468 , n469  );
buf ( g469 , n470  );
buf ( g470 , n471  );
buf ( g471 , n472  );
buf ( g472 , n473  );
buf ( g473 , n474  );
buf ( g474 , n475  );
buf ( g475 , n476  );
buf ( g476 , n477  );
buf ( g477 , n478  );
buf ( g478 , n479  );
buf ( g479 , n480  );
buf ( g480 , n481  );
buf ( g481 , n482  );
buf ( g482 , n483  );
buf ( g483 , n484  );
buf ( g484 , n485  );
buf ( g485 , n486  );
buf ( g486 , n487  );
buf ( g487 , n488  );
buf ( g488 , n489  );
buf ( g489 , n490  );
buf ( g490 , n491  );
buf ( g491 , n492  );
buf ( g492 , n493  );
buf ( g493 , n494  );
buf ( g494 , n495  );
buf ( g495 , n496  );
buf ( g496 , n497  );
buf ( g497 , n498  );
buf ( g498 , n499  );
buf ( g499 , n500  );
buf ( g500 , n501  );
buf ( n257 , n3962 );
buf ( n258 , n3965 );
buf ( n259 , n3802 );
buf ( n260 , n3968 );
buf ( n261 , n3809 );
buf ( n262 , n4188 );
buf ( n263 , n3815 );
buf ( n264 , n4185 );
buf ( n265 , n3973 );
buf ( n266 , n3976 );
buf ( n267 , n3980 );
buf ( n268 , n3983 );
buf ( n269 , n3988 );
buf ( n270 , n3991 );
buf ( n271 , n3995 );
buf ( n272 , n3998 );
buf ( n273 , n4176 );
buf ( n274 , n4179 );
buf ( n275 , n4182 );
buf ( n276 , n4001 );
buf ( n277 , n4005 );
buf ( n278 , n4008 );
buf ( n279 , n4012 );
buf ( n280 , n3818 );
buf ( n281 , n4017 );
buf ( n282 , n4020 );
buf ( n283 , n4025 );
buf ( n284 , n4028 );
buf ( n285 , n4032 );
buf ( n286 , n4035 );
buf ( n287 , n4039 );
buf ( n288 , n4042 );
buf ( n289 , n4047 );
buf ( n290 , n4050 );
buf ( n291 , n4054 );
buf ( n292 , n4198 );
buf ( n293 , n4157 );
buf ( n294 , n4057 );
buf ( n295 , n4061 );
buf ( n296 , n4064 );
buf ( n297 , n4069 );
buf ( n298 , n4072 );
buf ( n299 , n3823 );
buf ( n300 , n4075 );
buf ( n301 , n4080 );
buf ( n302 , n3826 );
buf ( n303 , n4202 );
buf ( n304 , n4083 );
buf ( n305 , n4088 );
buf ( n306 , n4091 );
buf ( n307 , n4096 );
buf ( n308 , n3957 );
buf ( n309 , n4101 );
buf ( n310 , n4104 );
buf ( n311 , n4109 );
buf ( n312 , n4112 );
buf ( n313 , n2923 );
buf ( n314 , n4258 );
buf ( n315 , n2867 );
buf ( n316 , n4246 );
buf ( n317 , n2524 );
buf ( n318 , n4250 );
buf ( n319 , n2617 );
buf ( n320 , n4254 );
buf ( n321 , n2863 );
buf ( n322 , n4119 );
buf ( n323 , n2818 );
buf ( n324 , n3834 );
buf ( n325 , n2928 );
buf ( n326 , n3841 );
buf ( n327 , n676 );
buf ( n328 , n4126 );
buf ( n329 , n2465 );
buf ( n330 , n3848 );
buf ( n331 , n1924 );
buf ( n332 , n4133 );
buf ( n333 , n1650 );
buf ( n334 , n4140 );
buf ( n335 , n1898 );
buf ( n336 , n4147 );
buf ( n337 , n4410 );
buf ( n338 , n4154 );
buf ( n339 , n2094 );
buf ( n340 , n3855 );
buf ( n341 , n1683 );
buf ( n342 , n3862 );
buf ( n343 , n1730 );
buf ( n344 , n4195 );
buf ( n345 , n1587 );
buf ( n346 , n3869 );
buf ( n347 , n1041 );
buf ( n348 , n3876 );
buf ( n349 , n1088 );
buf ( n350 , n3953 );
buf ( n351 , n2549 );
buf ( n352 , n3883 );
buf ( n353 , n2425 );
buf ( n354 , n4164 );
buf ( n355 , n4414 );
buf ( n356 , n4171 );
buf ( n357 , n2301 );
buf ( n358 , n3890 );
buf ( n359 , n2244 );
buf ( n360 , n3897 );
buf ( n361 , n2658 );
buf ( n362 , n3796 );
buf ( n363 , n1308 );
buf ( n364 , n3904 );
buf ( n365 , n1152 );
buf ( n366 , n3911 );
buf ( n367 , n2329 );
buf ( n368 , n3918 );
buf ( n369 , n843 );
buf ( n370 , n3925 );
buf ( n371 , n2705 );
buf ( n372 , n3932 );
buf ( n373 , n2736 );
buf ( n374 , n3939 );
buf ( n375 , n2951 );
buf ( n376 , n3946 );
buf ( n377 , n852 );
buf ( n378 , n2740 );
buf ( n379 , n2745 );
buf ( n380 , n2358 );
buf ( n381 , n1359 );
buf ( n382 , n2770 );
buf ( n383 , n2854 );
buf ( n384 , n2955 );
buf ( n385 , n2749 );
buf ( n386 , n1365 );
buf ( n387 , n1416 );
buf ( n388 , n1433 );
buf ( n389 , n2338 );
buf ( n390 , n2343 );
buf ( n391 , n2858 );
buf ( n392 , n2790 );
buf ( n393 , n2754 );
buf ( n394 , n1421 );
buf ( n395 , n2348 );
buf ( n396 , n1426 );
buf ( n397 , n2353 );
buf ( n398 , n2333 );
buf ( n399 , n2895 );
buf ( n400 , n2758 );
buf ( n401 , n2959 );
buf ( n402 , n2363 );
buf ( n403 , n2367 );
buf ( n404 , n2762 );
buf ( n405 , n2371 );
buf ( n406 , n2375 );
buf ( n407 , n858 );
buf ( n408 , n2766 );
buf ( n409 , n4213 );
buf ( n410 , n4275 );
buf ( n411 , n4286 );
buf ( n412 , n4292 );
buf ( n413 , n4281 );
buf ( n414 , n4218 );
buf ( n415 , n4223 );
buf ( n416 , n4391 );
buf ( n417 , n4264 );
buf ( n418 , n4330 );
buf ( n419 , n4345 );
buf ( n420 , n4350 );
buf ( n421 , n4325 );
buf ( n422 , n4385 );
buf ( n423 , n4297 );
buf ( n424 , n4270 );
buf ( n425 , n4397 );
buf ( n426 , n4304 );
buf ( n427 , n4375 );
buf ( n428 , n4370 );
buf ( n429 , n4380 );
buf ( n430 , n4310 );
buf ( n431 , n4355 );
buf ( n432 , n4230 );
buf ( n433 , n4236 );
buf ( n434 , n4340 );
buf ( n435 , n4315 );
buf ( n436 , n4365 );
buf ( n437 , n4320 );
buf ( n438 , n4360 );
buf ( n439 , n4335 );
buf ( n440 , n4242 );
buf ( n441 , n4399 );
buf ( n442 , n4403 );
buf ( n443 , n4405 );
buf ( n444 , n4406 );
buf ( n445 , n3183 );
buf ( n446 , n3199 );
buf ( n447 , n3214 );
buf ( n448 , n3228 );
buf ( n449 , n3241 );
buf ( n450 , n3254 );
buf ( n451 , n3267 );
buf ( n452 , n3015 );
buf ( n453 , n3062 );
buf ( n454 , n3281 );
buf ( n455 , n3294 );
buf ( n456 , n3308 );
buf ( n457 , n3047 );
buf ( n458 , n3322 );
buf ( n459 , n3335 );
buf ( n460 , n3349 );
buf ( n461 , n3123 );
buf ( n462 , n3363 );
buf ( n463 , n3376 );
buf ( n464 , n3390 );
buf ( n465 , n3153 );
buf ( n466 , n3404 );
buf ( n467 , n3417 );
buf ( n468 , n3431 );
buf ( n469 , n3139 );
buf ( n470 , n3444 );
buf ( n471 , n3456 );
buf ( n472 , n3468 );
buf ( n473 , n3108 );
buf ( n474 , n3484 );
buf ( n475 , n3498 );
buf ( n476 , n3783 );
buf ( n477 , n3093 );
buf ( n478 , n3513 );
buf ( n479 , n3527 );
buf ( n480 , n3542 );
buf ( n481 , n3555 );
buf ( n482 , n3569 );
buf ( n483 , n3582 );
buf ( n484 , n3596 );
buf ( n485 , n3031 );
buf ( n486 , n3610 );
buf ( n487 , n3623 );
buf ( n488 , n3637 );
buf ( n489 , n3077 );
buf ( n490 , n3651 );
buf ( n491 , n3664 );
buf ( n492 , n3678 );
buf ( n493 , n3168 );
buf ( n494 , n3692 );
buf ( n495 , n3706 );
buf ( n496 , n3720 );
buf ( n497 , n3733 );
buf ( n498 , n3746 );
buf ( n499 , n3758 );
buf ( n500 , n3771 );
buf ( n501 , n4207 );
xor ( n504 , n155 , n218 );
not ( n505 , n504 );
xor ( n506 , n156 , n207 );
nor ( n507 , n505 , n506 );
buf ( n508 , n507 );
not ( n509 , n508 );
xor ( n510 , n157 , n222 );
not ( n511 , n159 );
not ( n512 , n200 );
and ( n513 , n511 , n512 );
and ( n514 , n159 , n200 );
nor ( n515 , n513 , n514 );
nand ( n516 , n510 , n515 );
not ( n517 , n516 );
xor ( n518 , n158 , n213 );
nand ( n519 , n517 , n518 );
xor ( n520 , n160 , n225 );
not ( n521 , n520 );
buf ( n522 , n521 );
nor ( n523 , n519 , n522 );
not ( n524 , n523 );
or ( n525 , n509 , n524 );
nand ( n526 , n506 , n504 );
not ( n527 , n526 );
nand ( n528 , n527 , n521 );
not ( n529 , n528 );
not ( n530 , n515 );
nand ( n531 , n530 , n518 );
not ( n532 , n510 );
nor ( n533 , n531 , n532 );
and ( n534 , n529 , n533 );
not ( n535 , n518 );
nand ( n536 , n535 , n530 , n510 );
not ( n537 , n536 );
not ( n538 , n504 );
nand ( n539 , n538 , n506 );
nor ( n540 , n539 , n520 );
and ( n541 , n537 , n540 );
nor ( n542 , n534 , n541 );
nand ( n543 , n525 , n542 );
not ( n544 , n519 );
nand ( n545 , n532 , n518 );
not ( n546 , n545 );
buf ( n547 , n515 );
not ( n548 , n547 );
nand ( n549 , n546 , n548 );
not ( n550 , n549 );
or ( n551 , n544 , n550 );
nor ( n552 , n506 , n520 );
buf ( n553 , n504 );
and ( n554 , n552 , n553 );
nand ( n555 , n551 , n554 );
not ( n556 , n531 );
nand ( n557 , n532 , n506 );
not ( n558 , n521 );
or ( n559 , n557 , n558 );
not ( n560 , n520 );
not ( n561 , n560 );
nand ( n562 , n561 , n510 , n506 );
nand ( n563 , n559 , n562 );
nand ( n564 , n556 , n563 , n553 );
buf ( n565 , n539 );
not ( n566 , n565 );
nand ( n567 , n537 , n566 );
nand ( n568 , n555 , n564 , n567 );
nor ( n569 , n543 , n568 );
not ( n570 , n553 );
and ( n571 , n552 , n570 );
nor ( n572 , n547 , n532 );
nand ( n573 , n571 , n572 , n518 );
nor ( n574 , n526 , n521 );
or ( n575 , n574 , n540 );
not ( n576 , n549 );
nand ( n577 , n575 , n576 );
nor ( n578 , n510 , n518 );
nand ( n579 , n547 , n578 );
not ( n580 , n579 );
nand ( n581 , n580 , n540 );
nand ( n582 , n573 , n577 , n581 );
not ( n583 , n582 );
nor ( n584 , n548 , n545 );
not ( n585 , n584 );
not ( n586 , n554 );
or ( n587 , n585 , n586 );
nand ( n588 , n571 , n576 );
nand ( n589 , n587 , n588 );
not ( n590 , n566 );
not ( n591 , n518 );
nand ( n592 , n517 , n591 );
nor ( n593 , n592 , n522 );
not ( n594 , n593 );
or ( n595 , n590 , n594 );
nor ( n596 , n504 , n560 );
not ( n597 , n506 );
nand ( n598 , n596 , n597 );
not ( n599 , n598 );
nand ( n600 , n599 , n537 );
nand ( n601 , n595 , n600 );
nor ( n602 , n589 , n601 );
nand ( n603 , n569 , n583 , n602 );
not ( n604 , n603 );
nand ( n605 , n537 , n507 );
not ( n606 , n515 );
nand ( n607 , n606 , n578 );
not ( n608 , n522 );
nand ( n609 , n605 , n607 , n608 );
nand ( n610 , n537 , n507 , n561 );
nand ( n611 , n610 , n565 );
nand ( n612 , n519 , n560 );
nand ( n613 , n609 , n611 , n612 );
nor ( n614 , n516 , n518 );
and ( n615 , n529 , n614 );
and ( n616 , n576 , n599 );
nor ( n617 , n615 , n616 );
and ( n618 , n613 , n617 );
not ( n619 , n507 );
nand ( n620 , n619 , n565 );
not ( n621 , n620 );
and ( n622 , n606 , n553 );
not ( n623 , n606 );
and ( n624 , n623 , n596 );
nor ( n625 , n622 , n624 );
nor ( n626 , n625 , n545 );
not ( n627 , n626 );
or ( n628 , n621 , n627 );
not ( n629 , n607 );
nand ( n630 , n629 , n552 );
nand ( n631 , n628 , n630 );
not ( n632 , n508 );
nor ( n633 , n579 , n522 );
not ( n634 , n633 );
or ( n635 , n632 , n634 );
not ( n636 , n519 );
nand ( n637 , n636 , n599 );
nand ( n638 , n635 , n637 );
nor ( n639 , n631 , n638 );
nand ( n640 , n618 , n639 );
not ( n641 , n633 );
not ( n642 , n641 );
nand ( n643 , n528 , n598 );
nand ( n644 , n643 , n537 );
not ( n645 , n644 );
or ( n646 , n642 , n645 );
nand ( n647 , n646 , n527 );
nand ( n648 , n523 , n566 );
not ( n649 , n554 );
nand ( n650 , n649 , n598 , n614 , n597 );
nand ( n651 , n647 , n648 , n650 );
nor ( n652 , n640 , n651 );
nand ( n653 , n604 , n652 );
and ( n654 , n653 , n194 );
not ( n655 , n653 );
not ( n656 , n194 );
and ( n657 , n655 , n656 );
nor ( n658 , n654 , n657 );
nand ( n659 , n196 , n197 , n198 , n199 );
not ( n660 , n659 );
buf ( n661 , n660 );
not ( n662 , n661 );
buf ( n663 , n662 );
not ( n664 , n663 );
nand ( n665 , n658 , n664 );
nand ( n666 , n659 , n199 );
buf ( n667 , n666 );
not ( n668 , n667 );
not ( n669 , n668 );
buf ( n670 , n669 );
not ( n671 , n670 );
and ( n672 , n671 , n74 );
not ( n673 , n199 );
and ( n674 , n673 , n82 );
nor ( n675 , n672 , n674 );
nand ( n676 , n665 , n675 );
xor ( n677 , n136 , n250 );
not ( n678 , n677 );
xor ( n679 , n137 , n228 );
buf ( n680 , n679 );
xor ( n681 , n135 , n231 );
not ( n682 , n681 );
not ( n683 , n682 );
nand ( n684 , n678 , n680 , n683 );
not ( n685 , n684 );
xor ( n686 , n136 , n250 );
not ( n687 , n681 );
nand ( n688 , n686 , n687 , n679 );
not ( n689 , n688 );
xor ( n690 , n139 , n235 );
not ( n691 , n690 );
nand ( n692 , n689 , n691 );
not ( n693 , n692 );
or ( n694 , n685 , n693 );
not ( n695 , n245 );
not ( n696 , n138 );
or ( n697 , n695 , n696 );
or ( n698 , n138 , n245 );
nand ( n699 , n697 , n698 );
not ( n700 , n699 );
not ( n701 , n700 );
xor ( n702 , n140 , n240 );
not ( n703 , n702 );
nor ( n704 , n701 , n703 );
nand ( n705 , n694 , n704 );
not ( n706 , n679 );
nand ( n707 , n706 , n681 );
not ( n708 , n707 );
not ( n709 , n677 );
nand ( n710 , n708 , n709 );
not ( n711 , n710 );
not ( n712 , n700 );
not ( n713 , n139 );
not ( n714 , n235 );
and ( n715 , n713 , n714 );
and ( n716 , n139 , n235 );
nor ( n717 , n715 , n716 );
xor ( n718 , n140 , n240 );
nand ( n719 , n717 , n718 );
nor ( n720 , n712 , n719 );
nand ( n721 , n711 , n720 );
not ( n722 , n686 );
nor ( n723 , n679 , n681 );
nand ( n724 , n722 , n723 );
not ( n725 , n724 );
xor ( n726 , n138 , n245 );
buf ( n727 , n726 );
not ( n728 , n727 );
not ( n729 , n728 );
nor ( n730 , n729 , n719 );
nand ( n731 , n725 , n730 );
and ( n732 , n705 , n721 , n731 );
not ( n733 , n732 );
not ( n734 , n681 );
not ( n735 , n717 );
or ( n736 , n734 , n735 );
not ( n737 , n687 );
or ( n738 , n737 , n717 );
nand ( n739 , n736 , n738 );
not ( n740 , n739 );
buf ( n741 , n740 );
and ( n742 , n733 , n741 );
not ( n743 , n725 );
nand ( n744 , n691 , n727 , n702 );
not ( n745 , n744 );
not ( n746 , n745 );
or ( n747 , n743 , n746 );
not ( n748 , n684 );
nand ( n749 , n691 , n699 , n702 );
not ( n750 , n749 );
nand ( n751 , n748 , n750 );
nand ( n752 , n747 , n751 );
not ( n753 , n752 );
nand ( n754 , n686 , n702 );
nor ( n755 , n727 , n754 );
and ( n756 , n740 , n755 );
not ( n757 , n740 );
not ( n758 , n726 );
nor ( n759 , n758 , n718 );
and ( n760 , n759 , n709 , n679 );
and ( n761 , n757 , n760 );
nor ( n762 , n756 , n761 );
not ( n763 , n759 );
nor ( n764 , n739 , n763 );
nand ( n765 , n723 , n677 );
not ( n766 , n687 );
nand ( n767 , n766 , n686 , n679 );
nand ( n768 , n765 , n767 );
nand ( n769 , n764 , n768 );
nand ( n770 , n762 , n769 );
not ( n771 , n765 );
not ( n772 , n771 );
not ( n773 , n727 );
nand ( n774 , n773 , n703 , n690 );
not ( n775 , n774 );
not ( n776 , n775 );
or ( n777 , n772 , n776 );
not ( n778 , n767 );
nand ( n779 , n720 , n778 );
nand ( n780 , n777 , n779 );
nor ( n781 , n770 , n780 );
not ( n782 , n730 );
nor ( n783 , n782 , n710 );
not ( n784 , n720 );
not ( n785 , n677 );
nand ( n786 , n785 , n680 , n682 );
nor ( n787 , n784 , n786 );
nor ( n788 , n783 , n787 );
nand ( n789 , n753 , n781 , n788 );
nor ( n790 , n742 , n789 );
not ( n791 , n719 );
nand ( n792 , n768 , n791 );
not ( n793 , n792 );
nand ( n794 , n684 , n765 );
nor ( n795 , n717 , n718 );
buf ( n796 , n795 );
nand ( n797 , n794 , n796 );
not ( n798 , n797 );
or ( n799 , n793 , n798 );
nand ( n800 , n799 , n701 );
not ( n801 , n786 );
nand ( n802 , n801 , n750 );
nand ( n803 , n800 , n802 );
not ( n804 , n803 );
buf ( n805 , n688 );
not ( n806 , n805 );
not ( n807 , n806 );
and ( n808 , n795 , n701 );
not ( n809 , n808 );
or ( n810 , n807 , n809 );
nand ( n811 , n759 , n691 );
not ( n812 , n811 );
nand ( n813 , n812 , n725 );
nand ( n814 , n810 , n813 );
nand ( n815 , n721 , n692 );
nor ( n816 , n814 , n815 );
not ( n817 , n816 );
not ( n818 , n775 );
and ( n819 , n786 , n767 );
not ( n820 , n819 );
not ( n821 , n820 );
or ( n822 , n818 , n821 );
nand ( n823 , n708 , n677 );
nor ( n824 , n823 , n763 );
not ( n825 , n728 );
not ( n826 , n677 );
nand ( n827 , n826 , n703 );
nor ( n828 , n825 , n707 , n827 );
nor ( n829 , n824 , n828 );
nand ( n830 , n822 , n829 );
nor ( n831 , n817 , n830 );
nand ( n832 , n790 , n804 , n831 );
and ( n833 , n832 , n164 );
not ( n834 , n832 );
not ( n835 , n164 );
and ( n836 , n834 , n835 );
nor ( n837 , n833 , n836 );
not ( n838 , n663 );
nand ( n839 , n837 , n838 );
and ( n840 , n671 , n116 );
and ( n841 , n673 , n124 );
nor ( n842 , n840 , n841 );
nand ( n843 , n839 , n842 );
not ( n844 , n837 );
buf ( n845 , n662 );
not ( n846 , n845 );
or ( n847 , n844 , n846 );
buf ( n848 , n661 );
not ( n849 , n848 );
not ( n850 , n2 );
or ( n851 , n849 , n850 );
nand ( n852 , n847 , n851 );
not ( n853 , n658 );
or ( n854 , n853 , n846 );
buf ( n855 , n662 );
not ( n856 , n27 );
or ( n857 , n855 , n856 );
nand ( n858 , n854 , n857 );
xor ( n859 , n163 , n252 );
not ( n860 , n859 );
xor ( n861 , n132 , n255 );
nand ( n862 , n860 , n861 );
not ( n863 , n861 );
nand ( n864 , n863 , n859 );
nand ( n865 , n862 , n864 );
xor ( n866 , n163 , n252 );
xor ( n867 , n133 , n248 );
xor ( n868 , n866 , n867 );
not ( n869 , n868 );
nor ( n870 , n865 , n869 );
buf ( n871 , n870 );
not ( n872 , n871 );
not ( n873 , n872 );
not ( n874 , n134 );
not ( n875 , n234 );
and ( n876 , n874 , n875 );
and ( n877 , n134 , n234 );
nor ( n878 , n876 , n877 );
buf ( n879 , n878 );
not ( n880 , n879 );
not ( n881 , n880 );
not ( n882 , n867 );
nor ( n883 , n866 , n861 );
nand ( n884 , n882 , n883 );
not ( n885 , n884 );
nand ( n886 , n881 , n885 );
not ( n887 , n886 );
not ( n888 , n878 );
nor ( n889 , n888 , n859 );
not ( n890 , n889 );
not ( n891 , n878 );
nand ( n892 , n891 , n859 );
nand ( n893 , n890 , n892 );
nand ( n894 , n867 , n861 );
not ( n895 , n894 );
nand ( n896 , n893 , n895 );
not ( n897 , n892 );
nor ( n898 , n896 , n897 );
not ( n899 , n898 );
not ( n900 , n899 );
or ( n901 , n887 , n900 );
xor ( n902 , n136 , n238 );
not ( n903 , n902 );
xor ( n904 , n135 , n242 );
nand ( n905 , n903 , n904 );
not ( n906 , n905 );
nand ( n907 , n901 , n906 );
not ( n908 , n907 );
or ( n909 , n873 , n908 );
not ( n910 , n897 );
nand ( n911 , n902 , n904 );
not ( n912 , n911 );
not ( n913 , n884 );
or ( n914 , n912 , n913 );
nand ( n915 , n914 , n881 );
nand ( n916 , n910 , n915 , n896 );
not ( n917 , n891 );
not ( n918 , n911 );
nand ( n919 , n917 , n918 );
nand ( n920 , n919 , n905 );
and ( n921 , n916 , n920 );
nand ( n922 , n909 , n921 );
nor ( n923 , n902 , n904 );
and ( n924 , n879 , n923 );
buf ( n925 , n867 );
not ( n926 , n925 );
nor ( n927 , n926 , n864 );
nand ( n928 , n924 , n927 );
nand ( n929 , n922 , n928 );
not ( n930 , n929 );
not ( n931 , n911 );
nand ( n932 , n925 , n883 );
not ( n933 , n932 );
or ( n934 , n931 , n933 );
nor ( n935 , n917 , n905 );
not ( n936 , n935 );
not ( n937 , n932 );
not ( n938 , n937 );
or ( n939 , n936 , n938 );
buf ( n940 , n879 );
nor ( n941 , n862 , n925 );
and ( n942 , n940 , n941 );
not ( n943 , n882 );
nor ( n944 , n864 , n943 );
nor ( n945 , n942 , n944 );
nand ( n946 , n939 , n945 );
nand ( n947 , n934 , n946 );
nand ( n948 , n870 , n923 , n897 );
buf ( n949 , n948 );
nand ( n950 , n895 , n906 );
not ( n951 , n950 );
not ( n952 , n897 );
not ( n953 , n952 );
and ( n954 , n951 , n953 );
not ( n955 , n904 );
nand ( n956 , n955 , n902 );
not ( n957 , n956 );
buf ( n958 , n888 );
and ( n959 , n957 , n958 );
and ( n960 , n959 , n941 );
nor ( n961 , n954 , n960 );
nand ( n962 , n947 , n949 , n961 );
nand ( n963 , n859 , n878 );
nor ( n964 , n963 , n894 );
not ( n965 , n964 );
not ( n966 , n965 );
not ( n967 , n886 );
or ( n968 , n966 , n967 );
nand ( n969 , n968 , n918 );
not ( n970 , n885 );
not ( n971 , n959 );
or ( n972 , n970 , n971 );
nand ( n973 , n957 , n895 , n897 );
nand ( n974 , n972 , n973 );
not ( n975 , n974 );
not ( n976 , n963 );
and ( n977 , n870 , n976 );
not ( n978 , n923 );
not ( n979 , n978 );
nand ( n980 , n977 , n979 );
nand ( n981 , n969 , n975 , n980 );
nor ( n982 , n962 , n981 );
nand ( n983 , n880 , n918 );
nand ( n984 , n906 , n879 );
nand ( n985 , n983 , n984 );
nand ( n986 , n985 , n927 );
and ( n987 , n923 , n891 );
not ( n988 , n987 );
not ( n989 , n958 );
nand ( n990 , n989 , n957 );
nand ( n991 , n988 , n990 );
nand ( n992 , n991 , n885 );
and ( n993 , n986 , n992 );
not ( n994 , n935 );
not ( n995 , n994 );
not ( n996 , n924 );
not ( n997 , n996 );
or ( n998 , n995 , n997 );
not ( n999 , n937 );
not ( n1000 , n924 );
or ( n1001 , n999 , n1000 );
not ( n1002 , n862 );
nand ( n1003 , n926 , n1002 );
nand ( n1004 , n1001 , n1003 );
nand ( n1005 , n998 , n1004 );
not ( n1006 , n902 );
and ( n1007 , n864 , n1006 );
not ( n1008 , n902 );
not ( n1009 , n861 );
not ( n1010 , n1009 );
or ( n1011 , n1008 , n1010 );
nand ( n1012 , n1011 , n958 );
nor ( n1013 , n1007 , n1012 );
or ( n1014 , n1013 , n898 );
not ( n1015 , n1012 );
or ( n1016 , n1015 , n1006 );
not ( n1017 , n904 );
nand ( n1018 , n1014 , n1016 , n1017 );
not ( n1019 , n918 );
not ( n1020 , n888 );
nor ( n1021 , n1020 , n866 , n894 );
not ( n1022 , n1021 );
or ( n1023 , n1019 , n1022 );
nand ( n1024 , n964 , n957 );
nand ( n1025 , n1023 , n1024 );
and ( n1026 , n927 , n987 );
nor ( n1027 , n1025 , n1026 );
and ( n1028 , n993 , n1005 , n1018 , n1027 );
nand ( n1029 , n930 , n982 , n1028 );
and ( n1030 , n1029 , n175 );
not ( n1031 , n1029 );
not ( n1032 , n175 );
and ( n1033 , n1031 , n1032 );
nor ( n1034 , n1030 , n1033 );
buf ( n1035 , n661 );
nand ( n1036 , n1034 , n1035 );
not ( n1037 , n669 );
and ( n1038 , n1037 , n94 );
and ( n1039 , n673 , n102 );
nor ( n1040 , n1038 , n1039 );
nand ( n1041 , n1036 , n1040 );
nand ( n1042 , n649 , n598 );
and ( n1043 , n1042 , n533 );
not ( n1044 , n567 );
nor ( n1045 , n1043 , n1044 );
nand ( n1046 , n554 , n580 );
not ( n1047 , n620 );
nand ( n1048 , n593 , n1047 );
nand ( n1049 , n571 , n584 );
and ( n1050 , n1046 , n1048 , n1049 );
not ( n1051 , n625 );
not ( n1052 , n557 );
nand ( n1053 , n1051 , n1052 );
not ( n1054 , n1053 );
nand ( n1055 , n571 , n572 );
not ( n1056 , n1055 );
or ( n1057 , n1054 , n1056 );
nand ( n1058 , n1057 , n591 );
nand ( n1059 , n1045 , n1050 , n1058 , n577 );
not ( n1060 , n527 );
not ( n1061 , n523 );
or ( n1062 , n1060 , n1061 );
nand ( n1063 , n649 , n598 , n578 , n597 );
nand ( n1064 , n1062 , n1063 );
nor ( n1065 , n1059 , n1064 );
not ( n1066 , n648 );
nor ( n1067 , n1066 , n543 );
nand ( n1068 , n643 , n584 );
not ( n1069 , n607 );
not ( n1070 , n528 );
and ( n1071 , n1069 , n1070 );
and ( n1072 , n540 , n614 );
nor ( n1073 , n1071 , n1072 );
nand ( n1074 , n1068 , n555 , n1073 );
not ( n1075 , n1074 );
and ( n1076 , n1067 , n1075 , n618 );
nand ( n1077 , n1065 , n1076 );
and ( n1078 , n1077 , n183 );
not ( n1079 , n1077 );
not ( n1080 , n183 );
and ( n1081 , n1079 , n1080 );
nor ( n1082 , n1078 , n1081 );
not ( n1083 , n663 );
nand ( n1084 , n1082 , n1083 );
and ( n1085 , n671 , n96 );
and ( n1086 , n673 , n104 );
nor ( n1087 , n1085 , n1086 );
nand ( n1088 , n1084 , n1087 );
not ( n1089 , n181 );
not ( n1090 , n1089 );
not ( n1091 , n962 );
not ( n1092 , n1003 );
not ( n1093 , n932 );
or ( n1094 , n1092 , n1093 );
not ( n1095 , n990 );
nand ( n1096 , n1094 , n1095 );
nand ( n1097 , n1096 , n996 );
and ( n1098 , n1097 , n871 );
nand ( n1099 , n898 , n957 );
nand ( n1100 , n959 , n944 );
or ( n1101 , n983 , n1003 );
nand ( n1102 , n1099 , n1100 , n1101 , n950 );
nor ( n1103 , n1098 , n1102 );
not ( n1104 , n994 );
not ( n1105 , n884 );
and ( n1106 , n1104 , n1105 );
and ( n1107 , n977 , n957 );
nor ( n1108 , n1106 , n1107 );
nand ( n1109 , n1091 , n1103 , n1108 );
not ( n1110 , n919 );
not ( n1111 , n940 );
or ( n1112 , n1110 , n1111 );
buf ( n1113 , n927 );
nand ( n1114 , n1112 , n1113 );
not ( n1115 , n1114 );
not ( n1116 , n977 );
not ( n1117 , n1116 );
or ( n1118 , n1115 , n1117 );
not ( n1119 , n1110 );
not ( n1120 , n1113 );
or ( n1121 , n1119 , n1120 );
nand ( n1122 , n1121 , n905 );
nand ( n1123 , n1118 , n1122 );
not ( n1124 , n1003 );
not ( n1125 , n886 );
or ( n1126 , n1124 , n1125 );
nand ( n1127 , n1126 , n979 );
and ( n1128 , n1127 , n975 , n928 );
not ( n1129 , n886 );
and ( n1130 , n1111 , n937 );
nor ( n1131 , n1130 , n964 );
not ( n1132 , n1131 );
or ( n1133 , n1129 , n1132 );
nand ( n1134 , n1133 , n918 );
nand ( n1135 , n959 , n927 );
nand ( n1136 , n924 , n944 );
and ( n1137 , n1135 , n1136 );
nand ( n1138 , n1134 , n1137 );
not ( n1139 , n1138 );
nand ( n1140 , n1123 , n1128 , n1139 );
nor ( n1141 , n1109 , n1140 );
not ( n1142 , n1141 );
or ( n1143 , n1090 , n1142 );
or ( n1144 , n1089 , n1141 );
nand ( n1145 , n1143 , n1144 );
buf ( n1146 , n661 );
not ( n1147 , n1146 );
or ( n1148 , n1145 , n1147 );
and ( n1149 , n1037 , n112 );
and ( n1150 , n673 , n120 );
nor ( n1151 , n1149 , n1150 );
nand ( n1152 , n1148 , n1151 );
not ( n1153 , n162 );
not ( n1154 , n217 );
and ( n1155 , n1153 , n1154 );
and ( n1156 , n162 , n217 );
nor ( n1157 , n1155 , n1156 );
not ( n1158 , n1157 );
xor ( n1159 , n132 , n214 );
nand ( n1160 , n1158 , n1159 );
not ( n1161 , n1160 );
not ( n1162 , n1159 );
nand ( n1163 , n1162 , n1157 );
not ( n1164 , n1163 );
nor ( n1165 , n1161 , n1164 );
xor ( n1166 , n161 , n204 );
not ( n1167 , n1166 );
xor ( n1168 , n160 , n227 );
not ( n1169 , n1168 );
xor ( n1170 , n159 , n223 );
and ( n1171 , n1167 , n1169 , n1170 );
nand ( n1172 , n163 , n211 );
not ( n1173 , n1172 );
nor ( n1174 , n163 , n211 );
nor ( n1175 , n1173 , n1174 );
buf ( n1176 , n1175 );
nand ( n1177 , n1165 , n1171 , n1176 );
not ( n1178 , n1159 );
and ( n1179 , n1178 , n1175 );
not ( n1180 , n1179 );
xor ( n1181 , n161 , n204 );
nand ( n1182 , n1181 , n1168 );
not ( n1183 , n1182 );
not ( n1184 , n1170 );
nor ( n1185 , n1157 , n1184 );
nand ( n1186 , n1183 , n1185 );
not ( n1187 , n1186 );
not ( n1188 , n1187 );
or ( n1189 , n1180 , n1188 );
not ( n1190 , n162 );
not ( n1191 , n217 );
and ( n1192 , n1190 , n1191 );
and ( n1193 , n162 , n217 );
nor ( n1194 , n1192 , n1193 );
not ( n1195 , n1194 );
not ( n1196 , n211 );
not ( n1197 , n163 );
or ( n1198 , n1196 , n1197 );
or ( n1199 , n163 , n211 );
nand ( n1200 , n1198 , n1199 );
nand ( n1201 , n1200 , n1159 );
nor ( n1202 , n1195 , n1201 );
nor ( n1203 , n1182 , n1170 );
nand ( n1204 , n1202 , n1203 );
nand ( n1205 , n1189 , n1204 );
not ( n1206 , n1205 );
not ( n1207 , n1181 );
nand ( n1208 , n1207 , n1184 , n1168 );
not ( n1209 , n1208 );
buf ( n1210 , n1194 );
not ( n1211 , n1210 );
nand ( n1212 , n1209 , n1211 , n1179 );
nand ( n1213 , n1177 , n1206 , n1212 );
nand ( n1214 , n1167 , n1200 );
nor ( n1215 , n1214 , n1163 );
nor ( n1216 , n1201 , n1167 );
or ( n1217 , n1215 , n1216 );
nand ( n1218 , n1170 , n1168 );
not ( n1219 , n1218 );
nor ( n1220 , n1170 , n1168 );
or ( n1221 , n1219 , n1220 );
nand ( n1222 , n1217 , n1221 );
nand ( n1223 , n1220 , n1167 );
not ( n1224 , n1223 );
and ( n1225 , n1178 , n1200 );
nand ( n1226 , n1224 , n1211 , n1225 );
nor ( n1227 , n1218 , n1166 );
buf ( n1228 , n1159 );
nor ( n1229 , n1228 , n1194 );
nand ( n1230 , n1227 , n1229 );
nand ( n1231 , n1209 , n1228 , n1210 );
nand ( n1232 , n1222 , n1226 , n1230 , n1231 );
nor ( n1233 , n1213 , n1232 );
and ( n1234 , n1159 , n1175 );
not ( n1235 , n1234 );
and ( n1236 , n1166 , n1169 , n1170 );
nand ( n1237 , n1236 , n1210 );
nand ( n1238 , n1237 , n1186 );
not ( n1239 , n1238 );
or ( n1240 , n1235 , n1239 );
nand ( n1241 , n1209 , n1164 );
not ( n1242 , n1241 );
nand ( n1243 , n1236 , n1211 );
not ( n1244 , n1243 );
or ( n1245 , n1242 , n1244 );
nand ( n1246 , n1245 , n1225 );
nand ( n1247 , n1240 , n1246 );
not ( n1248 , n1247 );
and ( n1249 , n1164 , n1175 );
and ( n1250 , n1249 , n1203 );
nand ( n1251 , n1220 , n1166 );
not ( n1252 , n1251 );
nand ( n1253 , n1252 , n1225 , n1210 );
not ( n1254 , n1253 );
nor ( n1255 , n1250 , n1254 );
nand ( n1256 , n1233 , n1248 , n1255 );
not ( n1257 , n1256 );
not ( n1258 , n1164 );
not ( n1259 , n1171 );
or ( n1260 , n1258 , n1259 );
nor ( n1261 , n1251 , n1160 );
not ( n1262 , n1261 );
nand ( n1263 , n1260 , n1262 );
nor ( n1264 , n1263 , n1176 );
not ( n1265 , n1264 );
not ( n1266 , n1160 );
not ( n1267 , n1266 );
not ( n1268 , n1171 );
or ( n1269 , n1267 , n1268 );
nand ( n1270 , n1252 , n1229 );
nand ( n1271 , n1269 , n1270 );
not ( n1272 , n1179 );
nor ( n1273 , n1218 , n1166 );
not ( n1274 , n1273 );
or ( n1275 , n1272 , n1274 );
not ( n1276 , n1182 );
and ( n1277 , n1157 , n1170 );
nand ( n1278 , n1276 , n1277 , n1228 );
nand ( n1279 , n1275 , n1278 );
nor ( n1280 , n1271 , n1279 );
nor ( n1281 , n1280 , n1229 );
not ( n1282 , n1281 );
not ( n1283 , n1282 );
or ( n1284 , n1265 , n1283 );
not ( n1285 , n1237 );
not ( n1286 , n1228 );
nand ( n1287 , n1285 , n1286 );
nand ( n1288 , n1266 , n1227 );
nand ( n1289 , n1224 , n1165 );
nand ( n1290 , n1287 , n1288 , n1289 , n1176 );
not ( n1291 , n1290 );
not ( n1292 , n1203 );
nand ( n1293 , n1292 , n1223 );
or ( n1294 , n1236 , n1293 );
nand ( n1295 , n1294 , n1266 );
nand ( n1296 , n1291 , n1295 , n1270 );
nand ( n1297 , n1284 , n1296 );
nand ( n1298 , n1257 , n1297 );
and ( n1299 , n1298 , n173 );
not ( n1300 , n1298 );
not ( n1301 , n173 );
and ( n1302 , n1300 , n1301 );
nor ( n1303 , n1299 , n1302 );
nand ( n1304 , n1303 , n1083 );
and ( n1305 , n1037 , n110 );
and ( n1306 , n673 , n118 );
nor ( n1307 , n1305 , n1306 );
nand ( n1308 , n1304 , n1307 );
not ( n1309 , n543 );
not ( n1310 , n577 );
nand ( n1311 , n1047 , n636 , n522 );
not ( n1312 , n1311 );
or ( n1313 , n1310 , n1312 );
nand ( n1314 , n1313 , n553 );
nand ( n1315 , n1309 , n1314 , n602 );
not ( n1316 , n593 );
not ( n1317 , n1316 );
not ( n1318 , n508 );
not ( n1319 , n1318 );
and ( n1320 , n1317 , n1319 );
not ( n1321 , n599 );
not ( n1322 , n580 );
or ( n1323 , n1321 , n1322 );
nand ( n1324 , n574 , n584 );
nand ( n1325 , n1323 , n1324 );
nor ( n1326 , n1320 , n1325 );
not ( n1327 , n1073 );
not ( n1328 , n620 );
nor ( n1329 , n607 , n560 );
not ( n1330 , n1329 );
or ( n1331 , n1328 , n1330 );
nand ( n1332 , n1331 , n581 );
nor ( n1333 , n1327 , n1332 );
nand ( n1334 , n549 , n536 );
nand ( n1335 , n1334 , n554 );
not ( n1336 , n519 );
not ( n1337 , n607 );
or ( n1338 , n1336 , n1337 );
nand ( n1339 , n1338 , n571 );
not ( n1340 , n563 );
nand ( n1341 , n561 , n510 );
and ( n1342 , n565 , n1341 );
nor ( n1343 , n1342 , n531 );
nand ( n1344 , n1340 , n1343 );
and ( n1345 , n1335 , n1339 , n1344 );
nand ( n1346 , n1326 , n1333 , n1345 );
nor ( n1347 , n1315 , n1346 );
and ( n1348 , n647 , n1050 , n648 );
nand ( n1349 , n1347 , n1348 );
and ( n1350 , n1349 , n168 );
not ( n1351 , n1349 );
not ( n1352 , n168 );
and ( n1353 , n1351 , n1352 );
nor ( n1354 , n1350 , n1353 );
not ( n1355 , n1354 );
or ( n1356 , n1355 , n846 );
not ( n1357 , n37 );
or ( n1358 , n855 , n1357 );
nand ( n1359 , n1356 , n1358 );
not ( n1360 , n1303 );
or ( n1361 , n1360 , n846 );
not ( n1362 , n1035 );
not ( n1363 , n63 );
or ( n1364 , n1362 , n1363 );
nand ( n1365 , n1361 , n1364 );
not ( n1366 , n691 );
nand ( n1367 , n755 , n708 );
not ( n1368 , n1367 );
not ( n1369 , n1368 );
or ( n1370 , n1366 , n1369 );
nand ( n1371 , n1370 , n769 );
nor ( n1372 , n1371 , n814 );
nand ( n1373 , n732 , n1372 );
not ( n1374 , n791 );
nand ( n1375 , n823 , n805 );
not ( n1376 , n1375 );
or ( n1377 , n1374 , n1376 );
not ( n1378 , n827 );
not ( n1379 , n691 );
nand ( n1380 , n1378 , n708 , n1379 );
nand ( n1381 , n1377 , n1380 );
nand ( n1382 , n1381 , n825 );
nand ( n1383 , n820 , n808 );
not ( n1384 , n774 );
nand ( n1385 , n1375 , n1384 );
nand ( n1386 , n1382 , n1383 , n1385 );
nor ( n1387 , n1373 , n1386 );
not ( n1388 , n803 );
not ( n1389 , n823 );
not ( n1390 , n819 );
or ( n1391 , n1389 , n1390 );
nor ( n1392 , n763 , n691 );
nand ( n1393 , n1391 , n1392 );
nand ( n1394 , n820 , n745 );
nor ( n1395 , n825 , n791 , n796 );
and ( n1396 , n711 , n1395 );
and ( n1397 , n801 , n730 );
nor ( n1398 , n1396 , n1397 );
and ( n1399 , n1393 , n1394 , n1398 );
not ( n1400 , n774 );
not ( n1401 , n724 );
and ( n1402 , n1400 , n1401 );
nor ( n1403 , n744 , n765 );
nor ( n1404 , n1402 , n1403 );
nand ( n1405 , n1387 , n1388 , n1399 , n1404 );
and ( n1406 , n1405 , n174 );
not ( n1407 , n1405 );
not ( n1408 , n174 );
and ( n1409 , n1407 , n1408 );
nor ( n1410 , n1406 , n1409 );
not ( n1411 , n1410 );
or ( n1412 , n1411 , n846 );
not ( n1413 , n1035 );
not ( n1414 , n55 );
or ( n1415 , n1413 , n1414 );
nand ( n1416 , n1412 , n1415 );
or ( n1417 , n1145 , n846 );
not ( n1418 , n1035 );
not ( n1419 , n65 );
or ( n1420 , n1418 , n1419 );
nand ( n1421 , n1417 , n1420 );
not ( n1422 , n1082 );
or ( n1423 , n1422 , n1146 );
not ( n1424 , n49 );
or ( n1425 , n855 , n1424 );
nand ( n1426 , n1423 , n1425 );
not ( n1427 , n1034 );
or ( n1428 , n1427 , n846 );
not ( n1429 , n662 );
not ( n1430 , n1429 );
not ( n1431 , n47 );
or ( n1432 , n1430 , n1431 );
nand ( n1433 , n1428 , n1432 );
not ( n1434 , n167 );
not ( n1435 , n1434 );
xor ( n1436 , n142 , n233 );
not ( n1437 , n1436 );
xor ( n1438 , n141 , n239 );
nand ( n1439 , n1437 , n1438 );
not ( n1440 , n1439 );
xor ( n1441 , n139 , n236 );
xor ( n1442 , n140 , n251 );
nand ( n1443 , n1441 , n1442 );
not ( n1444 , n1443 );
nand ( n1445 , n1440 , n1444 );
nor ( n1446 , n1436 , n1438 );
nor ( n1447 , n1441 , n1442 );
nand ( n1448 , n1446 , n1447 );
nand ( n1449 , n1445 , n1448 );
not ( n1450 , n143 );
not ( n1451 , n244 );
and ( n1452 , n1450 , n1451 );
and ( n1453 , n143 , n244 );
nor ( n1454 , n1452 , n1453 );
xor ( n1455 , n144 , n254 );
nand ( n1456 , n1454 , n1455 );
not ( n1457 , n1456 );
nand ( n1458 , n1449 , n1457 );
not ( n1459 , n1443 );
nand ( n1460 , n1446 , n1459 );
not ( n1461 , n1460 );
or ( n1462 , n1454 , n1455 );
not ( n1463 , n1462 );
nand ( n1464 , n1461 , n1463 );
nand ( n1465 , n1438 , n1436 );
not ( n1466 , n1465 );
nand ( n1467 , n1466 , n1444 );
and ( n1468 , n1458 , n1464 , n1467 );
not ( n1469 , n1455 );
buf ( n1470 , n1454 );
nand ( n1471 , n1469 , n1470 );
not ( n1472 , n1454 );
nand ( n1473 , n1472 , n1455 );
nand ( n1474 , n1471 , n1473 );
nor ( n1475 , n1468 , n1474 );
not ( n1476 , n1473 );
not ( n1477 , n1442 );
nor ( n1478 , n1477 , n1441 );
not ( n1479 , n1438 );
nand ( n1480 , n1476 , n1478 , n1479 );
not ( n1481 , n1480 );
not ( n1482 , n1436 );
and ( n1483 , n1481 , n1482 );
nor ( n1484 , n1445 , n1471 );
nor ( n1485 , n1483 , n1484 );
buf ( n1486 , n1470 );
not ( n1487 , n1486 );
not ( n1488 , n1438 );
nand ( n1489 , n1488 , n1436 );
not ( n1490 , n1489 );
nand ( n1491 , n1490 , n1459 );
nand ( n1492 , n1491 , n1469 );
nand ( n1493 , n1466 , n1447 );
not ( n1494 , n1469 );
nand ( n1495 , n1493 , n1445 , n1494 );
nand ( n1496 , n1487 , n1492 , n1495 );
or ( n1497 , n1448 , n1462 );
nand ( n1498 , n1485 , n1496 , n1497 );
nor ( n1499 , n1475 , n1498 );
and ( n1500 , n1478 , n1438 );
nand ( n1501 , n1500 , n1437 );
or ( n1502 , n1501 , n1462 );
not ( n1503 , n1471 );
nand ( n1504 , n1477 , n1441 );
or ( n1505 , n1504 , n1439 );
nand ( n1506 , n1446 , n1478 );
nand ( n1507 , n1505 , n1506 );
nand ( n1508 , n1503 , n1507 );
nand ( n1509 , n1502 , n1508 );
not ( n1510 , n1503 );
not ( n1511 , n1504 );
nand ( n1512 , n1511 , n1446 );
not ( n1513 , n1512 );
not ( n1514 , n1513 );
or ( n1515 , n1510 , n1514 );
nand ( n1516 , n1511 , n1466 );
nor ( n1517 , n1516 , n1473 );
not ( n1518 , n1517 );
nand ( n1519 , n1515 , n1518 );
nor ( n1520 , n1509 , n1519 );
and ( n1521 , n1455 , n1436 );
nand ( n1522 , n1500 , n1521 , n1486 );
not ( n1523 , n1489 );
nand ( n1524 , n1523 , n1511 );
not ( n1525 , n1524 );
not ( n1526 , n1456 );
and ( n1527 , n1525 , n1526 );
not ( n1528 , n1493 );
and ( n1529 , n1528 , n1463 );
nor ( n1530 , n1527 , n1529 );
nand ( n1531 , n1522 , n1530 );
not ( n1532 , n1461 );
not ( n1533 , n1457 );
or ( n1534 , n1532 , n1533 );
nand ( n1535 , n1490 , n1447 , n1469 );
not ( n1536 , n1535 );
nand ( n1537 , n1536 , n1486 );
nand ( n1538 , n1534 , n1537 );
nor ( n1539 , n1531 , n1538 );
nand ( n1540 , n1499 , n1520 , n1539 );
not ( n1541 , n1501 );
not ( n1542 , n1491 );
or ( n1543 , n1541 , n1542 );
nand ( n1544 , n1543 , n1476 );
not ( n1545 , n1477 );
nand ( n1546 , n1470 , n1545 );
not ( n1547 , n1546 );
not ( n1548 , n1471 );
or ( n1549 , n1547 , n1548 );
not ( n1550 , n1478 );
not ( n1551 , n1523 );
or ( n1552 , n1550 , n1551 );
nand ( n1553 , n1552 , n1493 );
nand ( n1554 , n1549 , n1553 );
not ( n1555 , n1524 );
not ( n1556 , n1462 );
and ( n1557 , n1555 , n1556 );
nand ( n1558 , n1447 , n1440 );
nor ( n1559 , n1558 , n1473 );
nor ( n1560 , n1557 , n1559 );
and ( n1561 , n1554 , n1560 );
and ( n1562 , n1479 , n1476 );
not ( n1563 , n1479 );
and ( n1564 , n1563 , n1473 );
nor ( n1565 , n1562 , n1564 );
not ( n1566 , n1470 );
not ( n1567 , n1441 );
not ( n1568 , n1567 );
and ( n1569 , n1566 , n1568 );
and ( n1570 , n1470 , n1567 );
nor ( n1571 , n1569 , n1570 );
buf ( n1572 , n1545 );
nor ( n1573 , n1565 , n1571 , n1503 , n1572 );
and ( n1574 , n1500 , n1503 );
or ( n1575 , n1573 , n1574 );
nand ( n1576 , n1575 , n1437 );
nand ( n1577 , n1544 , n1561 , n1576 );
nor ( n1578 , n1540 , n1577 );
not ( n1579 , n1578 );
or ( n1580 , n1435 , n1579 );
or ( n1581 , n1578 , n1434 );
nand ( n1582 , n1580 , n1581 );
or ( n1583 , n1582 , n855 );
and ( n1584 , n1037 , n92 );
and ( n1585 , n673 , n100 );
nor ( n1586 , n1584 , n1585 );
nand ( n1587 , n1583 , n1586 );
not ( n1588 , n185 );
not ( n1589 , n1588 );
not ( n1590 , n1512 );
not ( n1591 , n1456 );
and ( n1592 , n1590 , n1591 );
nor ( n1593 , n1592 , n1517 );
nand ( n1594 , n1593 , n1485 );
or ( n1595 , n1501 , n1474 );
nand ( n1596 , n1595 , n1560 );
not ( n1597 , n1523 );
nor ( n1598 , n1597 , n1546 , n1455 );
nor ( n1599 , n1594 , n1596 , n1598 );
not ( n1600 , n1441 );
not ( n1601 , n1439 );
or ( n1602 , n1600 , n1601 );
not ( n1603 , n1545 );
nand ( n1604 , n1469 , n1603 );
nand ( n1605 , n1602 , n1604 );
nor ( n1606 , n1523 , n1441 );
nor ( n1607 , n1605 , n1606 );
not ( n1608 , n1572 );
nand ( n1609 , n1607 , n1608 );
nor ( n1610 , n1609 , n1486 );
not ( n1611 , n1455 );
buf ( n1612 , n1611 );
or ( n1613 , n1610 , n1612 );
nand ( n1614 , n1613 , n1513 );
not ( n1615 , n1609 );
or ( n1616 , n1615 , n1612 );
and ( n1617 , n1607 , n1487 );
nand ( n1618 , n1616 , n1617 );
nand ( n1619 , n1599 , n1614 , n1618 );
not ( n1620 , n1460 );
nand ( n1621 , n1500 , n1521 );
not ( n1622 , n1621 );
or ( n1623 , n1620 , n1622 );
nand ( n1624 , n1623 , n1476 );
or ( n1625 , n1449 , n1528 );
nand ( n1626 , n1625 , n1457 );
nand ( n1627 , n1558 , n1516 );
nand ( n1628 , n1627 , n1503 );
nand ( n1629 , n1624 , n1626 , n1628 );
not ( n1630 , n1629 );
not ( n1631 , n1558 );
or ( n1632 , n1461 , n1455 );
nand ( n1633 , n1467 , n1494 );
nand ( n1634 , n1632 , n1633 );
not ( n1635 , n1634 );
or ( n1636 , n1631 , n1635 );
nand ( n1637 , n1636 , n1487 );
nand ( n1638 , n1574 , n1436 );
and ( n1639 , n1637 , n1638 );
nand ( n1640 , n1630 , n1639 , n1539 );
nor ( n1641 , n1619 , n1640 );
not ( n1642 , n1641 );
or ( n1643 , n1589 , n1642 );
or ( n1644 , n1641 , n1588 );
nand ( n1645 , n1643 , n1644 );
or ( n1646 , n1645 , n1147 );
and ( n1647 , n671 , n80 );
and ( n1648 , n673 , n88 );
nor ( n1649 , n1647 , n1648 );
nand ( n1650 , n1646 , n1649 );
nand ( n1651 , n1368 , n1379 );
not ( n1652 , n754 );
not ( n1653 , n827 );
or ( n1654 , n1652 , n1653 );
xnor ( n1655 , n699 , n687 );
nor ( n1656 , n690 , n679 );
nand ( n1657 , n1655 , n1656 );
not ( n1658 , n1657 );
nand ( n1659 , n1654 , n1658 );
nor ( n1660 , n708 , n709 );
nand ( n1661 , n1660 , n775 );
nand ( n1662 , n1651 , n792 , n1659 , n1661 );
nor ( n1663 , n1662 , n752 );
not ( n1664 , n778 );
nand ( n1665 , n1664 , n710 );
nand ( n1666 , n1665 , n808 );
nand ( n1667 , n748 , n1384 );
not ( n1668 , n763 );
nor ( n1669 , n691 , n702 );
nand ( n1670 , n1668 , n725 , n1669 );
and ( n1671 , n1666 , n1667 , n1670 );
and ( n1672 , n1663 , n816 , n1671 );
nand ( n1673 , n1672 , n1399 );
and ( n1674 , n1673 , n184 );
not ( n1675 , n1673 );
not ( n1676 , n184 );
and ( n1677 , n1675 , n1676 );
nor ( n1678 , n1674 , n1677 );
nand ( n1679 , n1678 , n664 );
and ( n1680 , n1037 , n88 );
and ( n1681 , n673 , n96 );
nor ( n1682 , n1680 , n1681 );
nand ( n1683 , n1679 , n1682 );
nand ( n1684 , n1571 , n1466 , n1572 );
not ( n1685 , n1684 );
and ( n1686 , n1685 , n1611 );
and ( n1687 , n1513 , n1463 );
nor ( n1688 , n1686 , n1687 );
not ( n1689 , n1538 );
nand ( n1690 , n1553 , n1457 );
nand ( n1691 , n1688 , n1689 , n1690 );
nor ( n1692 , n1691 , n1498 );
not ( n1693 , n1593 );
and ( n1694 , n1535 , n1516 );
nor ( n1695 , n1694 , n1462 );
nor ( n1696 , n1693 , n1695 );
nand ( n1697 , n1696 , n1502 , n1508 );
not ( n1698 , n1697 );
or ( n1699 , n1501 , n1456 );
not ( n1700 , n1521 );
not ( n1701 , n1700 );
not ( n1702 , n1684 );
or ( n1703 , n1701 , n1702 );
or ( n1704 , n1504 , n1479 );
nand ( n1705 , n1704 , n1480 );
nand ( n1706 , n1703 , n1705 );
nand ( n1707 , n1699 , n1706 );
not ( n1708 , n1448 );
not ( n1709 , n1524 );
or ( n1710 , n1708 , n1709 );
nand ( n1711 , n1710 , n1476 );
not ( n1712 , n1456 );
not ( n1713 , n1491 );
nand ( n1714 , n1713 , n1486 );
not ( n1715 , n1714 );
or ( n1716 , n1712 , n1715 );
nand ( n1717 , n1716 , n1633 );
nand ( n1718 , n1711 , n1717 );
nor ( n1719 , n1707 , n1718 );
nand ( n1720 , n1692 , n1639 , n1698 , n1719 );
and ( n1721 , n1720 , n192 );
not ( n1722 , n1720 );
not ( n1723 , n192 );
and ( n1724 , n1722 , n1723 );
or ( n1725 , n1721 , n1724 );
or ( n1726 , n1725 , n1147 );
and ( n1727 , n1037 , n90 );
and ( n1728 , n673 , n98 );
nor ( n1729 , n1727 , n1728 );
nand ( n1730 , n1726 , n1729 );
not ( n1731 , n193 );
not ( n1732 , n1731 );
xor ( n1733 , n146 , n253 );
not ( n1734 , n1733 );
not ( n1735 , n145 );
not ( n1736 , n247 );
and ( n1737 , n1735 , n1736 );
and ( n1738 , n145 , n247 );
nor ( n1739 , n1737 , n1738 );
nor ( n1740 , n1734 , n1739 );
xor ( n1741 , n144 , n237 );
not ( n1742 , n1741 );
xor ( n1743 , n143 , n229 );
nand ( n1744 , n1742 , n1743 );
not ( n1745 , n1744 );
nand ( n1746 , n1740 , n1745 );
not ( n1747 , n1746 );
xor ( n1748 , n148 , n243 );
not ( n1749 , n1748 );
xor ( n1750 , n147 , n232 );
nand ( n1751 , n1749 , n1750 );
not ( n1752 , n1751 );
and ( n1753 , n1747 , n1752 );
xor ( n1754 , n145 , n247 );
not ( n1755 , n1754 );
not ( n1756 , n1755 );
nand ( n1757 , n1743 , n1741 );
not ( n1758 , n1757 );
not ( n1759 , n1758 );
or ( n1760 , n1756 , n1759 );
nor ( n1761 , n1743 , n1741 );
nand ( n1762 , n1739 , n1733 );
not ( n1763 , n1762 );
nand ( n1764 , n1761 , n1763 );
nand ( n1765 , n1760 , n1764 );
or ( n1766 , n1750 , n1748 );
not ( n1767 , n1766 );
and ( n1768 , n1765 , n1767 );
nor ( n1769 , n1753 , n1768 );
not ( n1770 , n1733 );
nand ( n1771 , n1770 , n1739 );
not ( n1772 , n1771 );
not ( n1773 , n1741 );
nor ( n1774 , n1773 , n1743 );
not ( n1775 , n1751 );
nand ( n1776 , n1772 , n1774 , n1775 );
not ( n1777 , n1750 );
nand ( n1778 , n1777 , n1748 );
not ( n1779 , n1778 );
not ( n1780 , n1771 );
nand ( n1781 , n1779 , n1780 , n1758 );
and ( n1782 , n1776 , n1781 );
nor ( n1783 , n1742 , n1743 );
and ( n1784 , n1740 , n1783 );
not ( n1785 , n1784 );
not ( n1786 , n1785 );
not ( n1787 , n1762 );
nand ( n1788 , n1787 , n1758 );
not ( n1789 , n1788 );
or ( n1790 , n1786 , n1789 );
nand ( n1791 , n1750 , n1748 );
not ( n1792 , n1791 );
nand ( n1793 , n1790 , n1792 );
and ( n1794 , n1769 , n1782 , n1793 );
nand ( n1795 , n1780 , n1745 );
nand ( n1796 , n1740 , n1758 );
nand ( n1797 , n1774 , n1763 );
nand ( n1798 , n1795 , n1796 , n1797 );
nand ( n1799 , n1798 , n1775 );
not ( n1800 , n1799 );
not ( n1801 , n1775 );
nand ( n1802 , n1761 , n1740 );
nor ( n1803 , n1733 , n1754 );
nand ( n1804 , n1745 , n1803 );
nand ( n1805 , n1783 , n1803 );
nand ( n1806 , n1802 , n1804 , n1805 );
not ( n1807 , n1806 );
or ( n1808 , n1801 , n1807 );
nand ( n1809 , n1777 , n1748 );
not ( n1810 , n1809 );
nand ( n1811 , n1784 , n1810 );
nand ( n1812 , n1808 , n1811 );
nor ( n1813 , n1800 , n1812 );
not ( n1814 , n1802 );
not ( n1815 , n1766 );
and ( n1816 , n1814 , n1815 );
nor ( n1817 , n1764 , n1809 );
nor ( n1818 , n1816 , n1817 );
not ( n1819 , n1818 );
not ( n1820 , n1810 );
not ( n1821 , n1804 );
not ( n1822 , n1821 );
or ( n1823 , n1820 , n1822 );
not ( n1824 , n1754 );
not ( n1825 , n1743 );
not ( n1826 , n1825 );
or ( n1827 , n1824 , n1826 );
or ( n1828 , n1825 , n1754 );
nand ( n1829 , n1827 , n1828 );
not ( n1830 , n1733 );
nand ( n1831 , n1830 , n1741 );
nor ( n1832 , n1829 , n1831 );
nand ( n1833 , n1832 , n1792 );
nand ( n1834 , n1823 , n1833 );
not ( n1835 , n1829 );
not ( n1836 , n1748 );
nor ( n1837 , n1836 , n1741 );
not ( n1838 , n1837 );
or ( n1839 , n1835 , n1838 );
or ( n1840 , n1755 , n1742 );
nand ( n1841 , n1839 , n1840 );
not ( n1842 , n1825 );
buf ( n1843 , n1733 );
nor ( n1844 , n1843 , n1750 );
not ( n1845 , n1844 );
or ( n1846 , n1842 , n1845 );
nand ( n1847 , n1777 , n1743 , n1843 );
nand ( n1848 , n1846 , n1847 );
nand ( n1849 , n1841 , n1848 );
nand ( n1850 , n1745 , n1763 );
nand ( n1851 , n1778 , n1751 );
nor ( n1852 , n1850 , n1851 );
not ( n1853 , n1852 );
nand ( n1854 , n1849 , n1853 );
nor ( n1855 , n1819 , n1834 , n1854 );
nand ( n1856 , n1794 , n1813 , n1855 );
not ( n1857 , n1830 );
and ( n1858 , n1784 , n1767 );
not ( n1859 , n1843 );
nand ( n1860 , n1859 , n1837 );
nand ( n1861 , n1750 , n1825 , n1755 );
nor ( n1862 , n1860 , n1861 );
nor ( n1863 , n1858 , n1862 );
not ( n1864 , n1796 );
and ( n1865 , n1864 , n1810 );
nand ( n1866 , n1758 , n1803 );
nor ( n1867 , n1866 , n1791 );
nor ( n1868 , n1865 , n1867 );
nand ( n1869 , n1780 , n1774 );
not ( n1870 , n1869 );
not ( n1871 , n1802 );
or ( n1872 , n1870 , n1871 );
nand ( n1873 , n1872 , n1810 );
nand ( n1874 , n1863 , n1868 , n1873 );
not ( n1875 , n1874 );
or ( n1876 , n1857 , n1875 );
nand ( n1877 , n1780 , n1761 );
or ( n1878 , n1877 , n1751 );
not ( n1879 , n1878 );
not ( n1880 , n1792 );
not ( n1881 , n1869 );
not ( n1882 , n1881 );
or ( n1883 , n1880 , n1882 );
not ( n1884 , n1788 );
nand ( n1885 , n1884 , n1810 );
nand ( n1886 , n1883 , n1885 );
nor ( n1887 , n1879 , n1886 );
nand ( n1888 , n1876 , n1887 );
nor ( n1889 , n1856 , n1888 );
not ( n1890 , n1889 );
or ( n1891 , n1732 , n1890 );
or ( n1892 , n1889 , n1731 );
nand ( n1893 , n1891 , n1892 );
or ( n1894 , n1893 , n855 );
and ( n1895 , n671 , n82 );
and ( n1896 , n673 , n90 );
nor ( n1897 , n1895 , n1896 );
nand ( n1898 , n1894 , n1897 );
not ( n1899 , n177 );
nand ( n1900 , n1561 , n1544 );
nor ( n1901 , n1697 , n1900 );
nand ( n1902 , n1717 , n1638 , n1711 );
nor ( n1903 , n1629 , n1902 );
nand ( n1904 , n1467 , n1506 );
nor ( n1905 , n1904 , n1461 );
not ( n1906 , n1462 );
not ( n1907 , n1460 );
or ( n1908 , n1906 , n1907 );
nand ( n1909 , n1908 , n1611 );
nor ( n1910 , n1905 , n1909 );
or ( n1911 , n1910 , n1615 );
or ( n1912 , n1905 , n1462 );
nand ( n1913 , n1912 , n1487 );
nand ( n1914 , n1911 , n1913 );
nand ( n1915 , n1901 , n1903 , n1914 );
not ( n1916 , n1915 );
or ( n1917 , n1899 , n1916 );
or ( n1918 , n1915 , n177 );
nand ( n1919 , n1917 , n1918 );
or ( n1920 , n1919 , n1147 );
and ( n1921 , n1037 , n78 );
and ( n1922 , n673 , n86 );
nor ( n1923 , n1921 , n1922 );
nand ( n1924 , n1920 , n1923 );
not ( n1925 , n201 );
not ( n1926 , n150 );
or ( n1927 , n1925 , n1926 );
or ( n1928 , n150 , n201 );
nand ( n1929 , n1927 , n1928 );
buf ( n1930 , n1929 );
not ( n1931 , n1930 );
not ( n1932 , n147 );
not ( n1933 , n226 );
and ( n1934 , n1932 , n1933 );
and ( n1935 , n147 , n226 );
nor ( n1936 , n1934 , n1935 );
buf ( n1937 , n1936 );
xor ( n1938 , n148 , n215 );
not ( n1939 , n1938 );
not ( n1940 , n149 );
not ( n1941 , n208 );
and ( n1942 , n1940 , n1941 );
and ( n1943 , n149 , n208 );
nor ( n1944 , n1942 , n1943 );
not ( n1945 , n1944 );
and ( n1946 , n1937 , n1939 , n1945 );
not ( n1947 , n1946 );
or ( n1948 , n1931 , n1947 );
not ( n1949 , n1944 );
xor ( n1950 , n150 , n201 );
nor ( n1951 , n1949 , n1950 );
not ( n1952 , n1951 );
not ( n1953 , n1952 );
and ( n1954 , n1938 , n1936 );
nand ( n1955 , n1953 , n1954 );
nand ( n1956 , n1948 , n1955 );
xor ( n1957 , n152 , n212 );
not ( n1958 , n151 );
not ( n1959 , n221 );
and ( n1960 , n1958 , n1959 );
and ( n1961 , n151 , n221 );
nor ( n1962 , n1960 , n1961 );
nor ( n1963 , n1957 , n1962 );
buf ( n1964 , n1963 );
nand ( n1965 , n1956 , n1964 );
not ( n1966 , n1957 );
not ( n1967 , n1929 );
nand ( n1968 , n1967 , n1945 );
not ( n1969 , n1936 );
nand ( n1970 , n1969 , n1939 );
nor ( n1971 , n1968 , n1970 );
not ( n1972 , n1971 );
or ( n1973 , n1966 , n1972 );
not ( n1974 , n1962 );
and ( n1975 , n1957 , n1974 );
and ( n1976 , n1950 , n1944 );
not ( n1977 , n1970 );
nand ( n1978 , n1975 , n1976 , n1977 );
nand ( n1979 , n1973 , n1978 );
or ( n1980 , n1957 , n1974 );
not ( n1981 , n1980 );
not ( n1982 , n1981 );
not ( n1983 , n1936 );
nand ( n1984 , n1983 , n1938 );
not ( n1985 , n1984 );
nand ( n1986 , n1985 , n1951 );
not ( n1987 , n1986 );
not ( n1988 , n1987 );
or ( n1989 , n1982 , n1988 );
not ( n1990 , n1937 );
nand ( n1991 , n1929 , n1945 );
not ( n1992 , n1991 );
nand ( n1993 , n1990 , n1963 , n1992 );
nand ( n1994 , n1989 , n1993 );
nor ( n1995 , n1979 , n1994 );
not ( n1996 , n1957 );
not ( n1997 , n1996 );
nand ( n1998 , n1937 , n1950 );
not ( n1999 , n1998 );
not ( n2000 , n1999 );
or ( n2001 , n1997 , n2000 );
nor ( n2002 , n1936 , n1950 );
not ( n2003 , n2002 );
not ( n2004 , n1939 );
nand ( n2005 , n1957 , n2004 );
nor ( n2006 , n2003 , n2005 );
not ( n2007 , n2006 );
nand ( n2008 , n2001 , n2007 );
not ( n2009 , n1945 );
buf ( n2010 , n1962 );
nor ( n2011 , n2009 , n2010 );
and ( n2012 , n2008 , n2011 );
or ( n2013 , n1970 , n1991 );
not ( n2014 , n1974 );
nand ( n2015 , n2014 , n1957 );
nor ( n2016 , n2013 , n2015 );
nor ( n2017 , n2012 , n2016 );
or ( n2018 , n1968 , n1984 );
not ( n2019 , n2018 );
not ( n2020 , n1955 );
or ( n2021 , n2019 , n2020 );
or ( n2022 , n1950 , n1957 );
nand ( n2023 , n1950 , n1957 );
nand ( n2024 , n2022 , n2023 );
nor ( n2025 , n2024 , n2010 );
nand ( n2026 , n2021 , n2025 );
nand ( n2027 , n1965 , n1995 , n2017 , n2026 );
not ( n2028 , n1981 );
nand ( n2029 , n1955 , n2018 );
not ( n2030 , n2029 );
or ( n2031 , n2028 , n2030 );
not ( n2032 , n1986 );
nand ( n2033 , n1976 , n1954 );
not ( n2034 , n2033 );
or ( n2035 , n2032 , n2034 );
not ( n2036 , n2015 );
nand ( n2037 , n2035 , n2036 );
not ( n2038 , n2004 );
nand ( n2039 , n2038 , n1937 , n2009 );
not ( n2040 , n2039 );
nand ( n2041 , n2040 , n1981 , n1950 );
and ( n2042 , n1951 , n1977 );
nand ( n2043 , n2042 , n1964 );
and ( n2044 , n2037 , n2041 , n2043 );
nand ( n2045 , n2031 , n2044 );
nor ( n2046 , n2027 , n2045 );
not ( n2047 , n2002 );
nand ( n2048 , n2047 , n1998 );
nor ( n2049 , n1957 , n1938 );
not ( n2050 , n2049 );
nand ( n2051 , n2050 , n2005 );
nand ( n2052 , n2051 , n1968 );
nor ( n2053 , n2048 , n2052 );
and ( n2054 , n1952 , n2053 );
not ( n2055 , n2023 );
and ( n2056 , n1946 , n2055 );
nor ( n2057 , n2054 , n2056 );
not ( n2058 , n2057 );
not ( n2059 , n2010 );
not ( n2060 , n2059 );
and ( n2061 , n2058 , n2060 );
and ( n2062 , n1945 , n1950 );
nand ( n2063 , n2062 , n1954 );
not ( n2064 , n2063 );
nand ( n2065 , n2040 , n1930 );
not ( n2066 , n2065 );
or ( n2067 , n2064 , n2066 );
nand ( n2068 , n2067 , n2036 );
nand ( n2069 , n1992 , n1954 );
not ( n2070 , n2069 );
nand ( n2071 , n2040 , n1950 );
not ( n2072 , n2071 );
or ( n2073 , n2070 , n2072 );
nand ( n2074 , n2073 , n1975 );
not ( n2075 , n1963 );
nand ( n2076 , n2075 , n2015 );
not ( n2077 , n1984 );
nand ( n2078 , n2077 , n1976 );
nor ( n2079 , n2076 , n2078 );
nor ( n2080 , n2076 , n2069 );
nor ( n2081 , n2079 , n2080 );
nand ( n2082 , n2068 , n2074 , n2081 );
nor ( n2083 , n2061 , n2082 );
nand ( n2084 , n2046 , n2083 );
and ( n2085 , n2084 , n176 );
not ( n2086 , n2084 );
not ( n2087 , n176 );
and ( n2088 , n2086 , n2087 );
nor ( n2089 , n2085 , n2088 );
nand ( n2090 , n2089 , n838 );
and ( n2091 , n671 , n86 );
and ( n2092 , n673 , n94 );
nor ( n2093 , n2091 , n2092 );
nand ( n2094 , n2090 , n2093 );
not ( n2095 , n190 );
not ( n2096 , n2095 );
xor ( n2097 , n155 , n209 );
not ( n2098 , n2097 );
not ( n2099 , n156 );
not ( n2100 , n205 );
and ( n2101 , n2099 , n2100 );
and ( n2102 , n156 , n205 );
nor ( n2103 , n2101 , n2102 );
nand ( n2104 , n2098 , n2103 );
not ( n2105 , n2104 );
not ( n2106 , n2105 );
not ( n2107 , n154 );
not ( n2108 , n216 );
and ( n2109 , n2107 , n2108 );
and ( n2110 , n154 , n216 );
nor ( n2111 , n2109 , n2110 );
not ( n2112 , n2111 );
not ( n2113 , n2112 );
not ( n2114 , n2113 );
not ( n2115 , n2114 );
xor ( n2116 , n152 , n202 );
not ( n2117 , n151 );
not ( n2118 , n220 );
and ( n2119 , n2117 , n2118 );
and ( n2120 , n151 , n220 );
nor ( n2121 , n2119 , n2120 );
nor ( n2122 , n2116 , n2121 );
not ( n2123 , n2122 );
xor ( n2124 , n153 , n224 );
buf ( n2125 , n2124 );
or ( n2126 , n2123 , n2125 );
not ( n2127 , n2116 );
buf ( n2128 , n2121 );
nand ( n2129 , n2127 , n2128 , n2125 );
nand ( n2130 , n2126 , n2129 );
not ( n2131 , n2130 );
or ( n2132 , n2115 , n2131 );
not ( n2133 , n2125 );
nor ( n2134 , n2113 , n2133 );
not ( n2135 , n2121 );
nand ( n2136 , n2135 , n2116 );
not ( n2137 , n2136 );
nand ( n2138 , n2134 , n2137 );
nand ( n2139 , n2132 , n2138 );
not ( n2140 , n2139 );
or ( n2141 , n2106 , n2140 );
nand ( n2142 , n2116 , n2121 );
not ( n2143 , n2142 );
nand ( n2144 , n2134 , n2143 );
not ( n2145 , n2144 );
or ( n2146 , n2097 , n2103 );
not ( n2147 , n2146 );
nand ( n2148 , n2145 , n2147 );
nand ( n2149 , n2141 , n2148 );
not ( n2150 , n2149 );
and ( n2151 , n2125 , n2111 );
buf ( n2152 , n2122 );
nand ( n2153 , n2151 , n2152 );
not ( n2154 , n2124 );
nand ( n2155 , n2154 , n2111 );
not ( n2156 , n2155 );
nand ( n2157 , n2137 , n2156 );
nand ( n2158 , n2153 , n2157 );
nor ( n2159 , n2125 , n2111 );
nand ( n2160 , n2143 , n2159 );
not ( n2161 , n2160 );
nor ( n2162 , n2158 , n2161 );
not ( n2163 , n2103 );
not ( n2164 , n2163 );
or ( n2165 , n2162 , n2164 );
nand ( n2166 , n2112 , n2163 );
not ( n2167 , n2166 );
nand ( n2168 , n2167 , n2152 , n2125 );
not ( n2169 , n2168 );
nand ( n2170 , n2163 , n2097 );
nand ( n2171 , n2170 , n2104 );
nand ( n2172 , n2137 , n2151 );
nor ( n2173 , n2171 , n2172 );
nor ( n2174 , n2169 , n2173 );
nand ( n2175 , n2165 , n2174 );
nand ( n2176 , n2175 , n2098 );
nand ( n2177 , n2137 , n2159 );
and ( n2178 , n2177 , n2129 );
not ( n2179 , n2178 );
nand ( n2180 , n2143 , n2151 );
nand ( n2181 , n2138 , n2180 );
not ( n2182 , n2181 );
not ( n2183 , n2182 );
or ( n2184 , n2179 , n2183 );
buf ( n2185 , n2170 );
not ( n2186 , n2185 );
nand ( n2187 , n2184 , n2186 );
not ( n2188 , n2097 );
not ( n2189 , n2128 );
and ( n2190 , n2188 , n2189 );
and ( n2191 , n2128 , n2097 );
nor ( n2192 , n2190 , n2191 );
nand ( n2193 , n2142 , n2159 , n2192 );
nand ( n2194 , n2150 , n2176 , n2187 , n2193 );
not ( n2195 , n2160 );
not ( n2196 , n2116 );
nand ( n2197 , n2196 , n2128 , n2156 );
not ( n2198 , n2197 );
or ( n2199 , n2195 , n2198 );
not ( n2200 , n2163 );
nand ( n2201 , n2200 , n2097 );
not ( n2202 , n2201 );
nand ( n2203 , n2199 , n2202 );
nand ( n2204 , n2156 , n2122 );
not ( n2205 , n2204 );
not ( n2206 , n2201 );
and ( n2207 , n2205 , n2206 );
not ( n2208 , n2133 );
not ( n2209 , n2166 );
or ( n2210 , n2208 , n2209 );
not ( n2211 , n2116 );
nand ( n2212 , n2210 , n2211 );
nor ( n2213 , n2097 , n2125 );
nand ( n2214 , n2213 , n2128 );
nor ( n2215 , n2212 , n2214 );
nor ( n2216 , n2207 , n2215 );
or ( n2217 , n2180 , n2104 );
nand ( n2218 , n2164 , n2156 , n2143 );
and ( n2219 , n2203 , n2216 , n2217 , n2218 );
not ( n2220 , n2197 );
not ( n2221 , n2146 );
and ( n2222 , n2220 , n2221 );
and ( n2223 , n2158 , n2105 );
nor ( n2224 , n2222 , n2223 );
not ( n2225 , n2129 );
not ( n2226 , n2114 );
nand ( n2227 , n2225 , n2226 );
nand ( n2228 , n2156 , n2143 );
nand ( n2229 , n2227 , n2204 , n2228 );
nand ( n2230 , n2229 , n2186 );
nand ( n2231 , n2152 , n2159 );
nand ( n2232 , n2231 , n2144 , n2172 );
nand ( n2233 , n2232 , n2202 );
nand ( n2234 , n2219 , n2224 , n2230 , n2233 );
nor ( n2235 , n2194 , n2234 );
not ( n2236 , n2235 );
or ( n2237 , n2096 , n2236 );
or ( n2238 , n2095 , n2235 );
nand ( n2239 , n2237 , n2238 );
or ( n2240 , n2239 , n1418 );
and ( n2241 , n671 , n106 );
and ( n2242 , n673 , n114 );
nor ( n2243 , n2241 , n2242 );
nand ( n2244 , n2240 , n2243 );
not ( n2245 , n1812 );
not ( n2246 , n1802 );
nand ( n2247 , n2246 , n1792 );
nand ( n2248 , n1821 , n1767 );
nand ( n2249 , n2247 , n2248 );
nor ( n2250 , n2249 , n1886 );
nor ( n2251 , n1852 , n1862 );
and ( n2252 , n1776 , n2251 , n1781 );
not ( n2253 , n1795 );
nand ( n2254 , n2253 , n1810 );
not ( n2255 , n1877 );
nand ( n2256 , n2255 , n1792 );
nand ( n2257 , n1832 , n1767 );
and ( n2258 , n2254 , n2256 , n2257 );
nand ( n2259 , n2245 , n2250 , n2252 , n2258 );
not ( n2260 , n2259 );
nand ( n2261 , n1795 , n1764 , n1788 );
nand ( n2262 , n2261 , n1775 );
not ( n2263 , n1791 );
not ( n2264 , n1766 );
or ( n2265 , n2263 , n2264 );
not ( n2266 , n1797 );
nand ( n2267 , n2265 , n2266 );
nand ( n2268 , n1818 , n1868 , n2262 , n2267 );
not ( n2269 , n1748 );
not ( n2270 , n1844 );
not ( n2271 , n1761 );
or ( n2272 , n2270 , n2271 );
nand ( n2273 , n1758 , n1733 );
nand ( n2274 , n2272 , n2273 );
not ( n2275 , n2274 );
or ( n2276 , n2269 , n2275 );
not ( n2277 , n1847 );
nor ( n2278 , n1741 , n1748 );
nand ( n2279 , n2277 , n2278 );
nand ( n2280 , n2276 , n2279 );
nand ( n2281 , n2280 , n1755 );
nand ( n2282 , n1821 , n1748 );
not ( n2283 , n2282 );
nand ( n2284 , n2283 , n1750 );
not ( n2285 , n1877 );
not ( n2286 , n1796 );
or ( n2287 , n2285 , n2286 );
nand ( n2288 , n2287 , n1767 );
nand ( n2289 , n2281 , n2284 , n2288 );
nor ( n2290 , n2268 , n2289 );
nand ( n2291 , n2260 , n2290 );
and ( n2292 , n2291 , n182 );
not ( n2293 , n2291 );
not ( n2294 , n182 );
and ( n2295 , n2293 , n2294 );
nor ( n2296 , n2292 , n2295 );
nand ( n2297 , n2296 , n1146 );
and ( n2298 , n671 , n104 );
and ( n2299 , n673 , n112 );
nor ( n2300 , n2298 , n2299 );
nand ( n2301 , n2297 , n2300 );
and ( n2302 , n788 , n1394 , n1671 );
nand ( n2303 , n830 , n1655 );
nand ( n2304 , n794 , n720 );
nand ( n2305 , n1404 , n2304 , n1385 , n802 );
not ( n2306 , n763 );
not ( n2307 , n749 );
or ( n2308 , n2306 , n2307 );
nand ( n2309 , n2308 , n689 );
and ( n2310 , n813 , n2309 );
not ( n2311 , n1367 );
nand ( n2312 , n709 , n702 );
nor ( n2313 , n1657 , n2312 );
nor ( n2314 , n2311 , n2313 );
not ( n2315 , n811 );
nand ( n2316 , n2315 , n748 );
nand ( n2317 , n2310 , n2314 , n751 , n2316 );
nor ( n2318 , n2305 , n2317 );
nand ( n2319 , n2302 , n2303 , n2318 , n800 );
and ( n2320 , n2319 , n189 );
not ( n2321 , n2319 );
not ( n2322 , n189 );
and ( n2323 , n2321 , n2322 );
nor ( n2324 , n2320 , n2323 );
nand ( n2325 , n2324 , n664 );
and ( n2326 , n671 , n114 );
and ( n2327 , n673 , n122 );
nor ( n2328 , n2326 , n2327 );
nand ( n2329 , n2325 , n2328 );
or ( n2330 , n1645 , n846 );
not ( n2331 , n33 );
or ( n2332 , n1362 , n2331 );
nand ( n2333 , n2330 , n2332 );
not ( n2334 , n2089 );
or ( n2335 , n2334 , n846 );
not ( n2336 , n39 );
or ( n2337 , n1362 , n2336 );
nand ( n2338 , n2335 , n2337 );
not ( n2339 , n663 );
or ( n2340 , n1919 , n2339 );
not ( n2341 , n31 );
or ( n2342 , n1413 , n2341 );
nand ( n2343 , n2340 , n2342 );
not ( n2344 , n2296 );
or ( n2345 , n2344 , n846 );
not ( n2346 , n57 );
or ( n2347 , n855 , n2346 );
nand ( n2348 , n2345 , n2347 );
not ( n2349 , n1678 );
or ( n2350 , n2349 , n846 );
not ( n2351 , n41 );
or ( n2352 , n849 , n2351 );
nand ( n2353 , n2350 , n2352 );
not ( n2354 , n855 );
or ( n2355 , n1582 , n2354 );
not ( n2356 , n45 );
or ( n2357 , n1362 , n2356 );
nand ( n2358 , n2355 , n2357 );
not ( n2359 , n2324 );
or ( n2360 , n2359 , n846 );
not ( n2361 , n67 );
or ( n2362 , n1413 , n2361 );
nand ( n2363 , n2360 , n2362 );
or ( n2364 , n2239 , n846 );
not ( n2365 , n59 );
or ( n2366 , n855 , n2365 );
nand ( n2367 , n2364 , n2366 );
or ( n2368 , n1725 , n846 );
not ( n2369 , n43 );
or ( n2370 , n849 , n2369 );
nand ( n2371 , n2368 , n2370 );
or ( n2372 , n1893 , n846 );
not ( n2373 , n35 );
or ( n2374 , n1413 , n2373 );
nand ( n2375 , n2372 , n2374 );
not ( n2376 , n166 );
and ( n2377 , n2128 , n2163 , n2125 );
or ( n2378 , n2212 , n2377 );
not ( n2379 , n2378 );
or ( n2380 , n2128 , n2166 );
nand ( n2381 , n2380 , n2097 );
not ( n2382 , n2381 );
and ( n2383 , n2379 , n2382 );
nor ( n2384 , n2144 , n2185 );
nor ( n2385 , n2383 , n2384 );
nand ( n2386 , n2161 , n2105 );
and ( n2387 , n2217 , n2386 );
not ( n2388 , n2204 );
not ( n2389 , n2138 );
or ( n2390 , n2388 , n2389 );
nand ( n2391 , n2390 , n2147 );
nand ( n2392 , n2385 , n2387 , n2391 );
nand ( n2393 , n2197 , n2177 );
nand ( n2394 , n2393 , n2105 );
not ( n2395 , n2153 );
not ( n2396 , n2160 );
or ( n2397 , n2395 , n2396 );
not ( n2398 , n2171 );
nand ( n2399 , n2397 , n2398 );
or ( n2400 , n2138 , n2185 );
nand ( n2401 , n2394 , n2399 , n2400 );
nor ( n2402 , n2392 , n2401 );
nand ( n2403 , n2231 , n2180 );
not ( n2404 , n2403 );
and ( n2405 , n2404 , n2227 );
nor ( n2406 , n2405 , n2146 );
not ( n2407 , n2197 );
nor ( n2408 , n2129 , n2226 );
nor ( n2409 , n2407 , n2408 );
not ( n2410 , n2164 );
or ( n2411 , n2409 , n2410 );
nand ( n2412 , n2411 , n2157 );
or ( n2413 , n2406 , n2412 );
nand ( n2414 , n2413 , n2398 );
and ( n2415 , n2224 , n2230 , n2233 );
nand ( n2416 , n2402 , n2414 , n2415 );
not ( n2417 , n2416 );
or ( n2418 , n2376 , n2417 );
or ( n2419 , n2416 , n166 );
nand ( n2420 , n2418 , n2419 );
or ( n2421 , n2420 , n1147 );
and ( n2422 , n671 , n100 );
and ( n2423 , n673 , n108 );
nor ( n2424 , n2422 , n2423 );
nand ( n2425 , n2421 , n2424 );
not ( n2426 , n893 );
not ( n2427 , n923 );
not ( n2428 , n895 );
or ( n2429 , n2427 , n2428 );
nand ( n2430 , n868 , n957 , n1009 );
nand ( n2431 , n2429 , n2430 );
nand ( n2432 , n2426 , n2431 );
and ( n2433 , n928 , n948 , n2432 );
not ( n2434 , n937 );
not ( n2435 , n984 );
not ( n2436 , n2435 );
or ( n2437 , n2434 , n2436 );
nand ( n2438 , n2437 , n1135 );
nor ( n2439 , n974 , n2438 );
nand ( n2440 , n996 , n983 );
and ( n2441 , n2440 , n941 );
nand ( n2442 , n919 , n978 );
and ( n2443 , n2442 , n885 );
nor ( n2444 , n2441 , n2443 );
and ( n2445 , n2433 , n2439 , n2444 );
not ( n2446 , n994 );
not ( n2447 , n944 );
not ( n2448 , n2447 );
and ( n2449 , n2446 , n2448 );
not ( n2450 , n906 );
not ( n2451 , n1021 );
or ( n2452 , n2450 , n2451 );
nand ( n2453 , n882 , n866 );
or ( n2454 , n983 , n2453 );
nand ( n2455 , n2452 , n2454 );
nor ( n2456 , n2449 , n2455 );
nand ( n2457 , n2456 , n1027 , n1096 );
not ( n2458 , n2457 );
nand ( n2459 , n2445 , n1123 , n922 , n2458 );
xnor ( n2460 , n2459 , n169 );
or ( n2461 , n2460 , n1147 );
and ( n2462 , n1037 , n76 );
and ( n2463 , n673 , n84 );
nor ( n2464 , n2462 , n2463 );
nand ( n2465 , n2461 , n2464 );
not ( n2466 , n187 );
not ( n2467 , n1213 );
and ( n2468 , n1176 , n1263 );
not ( n2469 , n1176 );
and ( n2470 , n2469 , n1271 );
nor ( n2471 , n2468 , n2470 );
not ( n2472 , n1234 );
not ( n2473 , n2472 );
not ( n2474 , n1288 );
or ( n2475 , n2473 , n2474 );
and ( n2476 , n1186 , n1208 );
nand ( n2477 , n1288 , n2476 );
nand ( n2478 , n2475 , n2477 );
nand ( n2479 , n2467 , n2471 , n2478 );
not ( n2480 , n2479 );
nor ( n2481 , n1194 , n1170 );
nand ( n2482 , n2481 , n1276 );
not ( n2483 , n2482 );
not ( n2484 , n1243 );
or ( n2485 , n2483 , n2484 );
nand ( n2486 , n2485 , n1179 );
buf ( n2487 , n1200 );
not ( n2488 , n2487 );
not ( n2489 , n1261 );
or ( n2490 , n2488 , n2489 );
nand ( n2491 , n2490 , n1226 );
not ( n2492 , n1224 );
not ( n2493 , n1202 );
or ( n2494 , n2492 , n2493 );
nand ( n2495 , n1234 , n2481 , n1167 );
nand ( n2496 , n2494 , n2495 );
nor ( n2497 , n2491 , n2496 );
not ( n2498 , n1165 );
nor ( n2499 , n1219 , n1175 );
nand ( n2500 , n2498 , n2499 , n1277 );
and ( n2501 , n2486 , n2497 , n2500 );
nand ( n2502 , n1249 , n1219 );
not ( n2503 , n2502 );
nand ( n2504 , n2498 , n2499 );
not ( n2505 , n2504 );
or ( n2506 , n2503 , n2505 );
nand ( n2507 , n2506 , n1166 );
nand ( n2508 , n1227 , n1229 , n2487 );
not ( n2509 , n2508 );
nor ( n2510 , n1278 , n2487 );
nor ( n2511 , n2509 , n2510 );
nand ( n2512 , n1202 , n1273 );
nand ( n2513 , n1253 , n1241 , n2512 );
not ( n2514 , n2513 );
and ( n2515 , n2507 , n2511 , n2514 );
nand ( n2516 , n2480 , n2501 , n2515 );
not ( n2517 , n2516 );
or ( n2518 , n2466 , n2517 );
or ( n2519 , n2516 , n187 );
nand ( n2520 , n2518 , n2519 );
or ( n2521 , n2520 , n1147 );
not ( n2522 , n72 );
or ( n2523 , n2522 , n199 );
nand ( n2524 , n2521 , n2523 );
not ( n2525 , n943 );
not ( n2526 , n865 );
not ( n2527 , n2526 );
not ( n2528 , n987 );
or ( n2529 , n2527 , n2528 );
nor ( n2530 , n990 , n864 );
or ( n2531 , n2530 , n1110 );
or ( n2532 , n1002 , n1017 );
nand ( n2533 , n2531 , n2532 );
nand ( n2534 , n2529 , n2533 );
not ( n2535 , n2534 );
or ( n2536 , n2525 , n2535 );
and ( n2537 , n961 , n948 );
nand ( n2538 , n2536 , n2537 );
nor ( n2539 , n2538 , n1138 );
nand ( n2540 , n871 , n2435 );
nand ( n2541 , n993 , n1005 , n2540 );
nor ( n2542 , n2457 , n2541 );
nand ( n2543 , n2539 , n2542 , n1108 );
xnor ( n2544 , n2543 , n191 );
or ( n2545 , n2544 , n1147 );
and ( n2546 , n1037 , n98 );
and ( n2547 , n673 , n106 );
nor ( n2548 , n2546 , n2547 );
nand ( n2549 , n2545 , n2548 );
not ( n2550 , n195 );
not ( n2551 , n1956 );
not ( n2552 , n1946 );
not ( n2553 , n2552 );
not ( n2554 , n2013 );
or ( n2555 , n2553 , n2554 );
nand ( n2556 , n2555 , n1975 );
not ( n2557 , n2556 );
not ( n2558 , n2557 );
or ( n2559 , n2551 , n2558 );
not ( n2560 , n2033 );
nand ( n2561 , n2560 , n1996 );
nand ( n2562 , n1971 , n2036 );
and ( n2563 , n2561 , n1978 , n2562 );
nand ( n2564 , n2559 , n2563 );
not ( n2565 , n2036 );
not ( n2566 , n1956 );
or ( n2567 , n2565 , n2566 );
not ( n2568 , n1981 );
not ( n2569 , n1971 );
or ( n2570 , n2568 , n2569 );
nor ( n2571 , n1968 , n1984 );
nand ( n2572 , n2571 , n1975 );
nand ( n2573 , n2570 , n2572 );
not ( n2574 , n2573 );
nand ( n2575 , n2567 , n2574 );
nor ( n2576 , n2564 , n2575 );
not ( n2577 , n2082 );
not ( n2578 , n1964 );
not ( n2579 , n2053 );
or ( n2580 , n2578 , n2579 );
and ( n2581 , n2042 , n1975 );
nor ( n2582 , n2581 , n2016 );
nand ( n2583 , n2580 , n2582 );
not ( n2584 , n2010 );
not ( n2585 , n2006 );
or ( n2586 , n2584 , n2585 );
not ( n2587 , n2005 );
nand ( n2588 , n2587 , n1999 , n2059 );
nand ( n2589 , n2586 , n2588 );
not ( n2590 , n2589 );
not ( n2591 , n2038 );
not ( n2592 , n2591 );
nand ( n2593 , n2592 , n2048 , n1981 );
and ( n2594 , n2590 , n2593 );
nor ( n2595 , n2594 , n2009 );
nor ( n2596 , n2583 , n2595 );
not ( n2597 , n1964 );
nand ( n2598 , n1955 , n2063 );
not ( n2599 , n2598 );
or ( n2600 , n2597 , n2599 );
not ( n2601 , n1994 );
nand ( n2602 , n2600 , n2601 );
nand ( n2603 , n2042 , n2036 );
not ( n2604 , n2078 );
nand ( n2605 , n2604 , n1981 );
nand ( n2606 , n1987 , n1964 );
nand ( n2607 , n2603 , n2605 , n2606 );
nor ( n2608 , n2602 , n2607 );
nand ( n2609 , n2576 , n2577 , n2596 , n2608 );
not ( n2610 , n2609 );
or ( n2611 , n2550 , n2610 );
or ( n2612 , n2609 , n195 );
nand ( n2613 , n2611 , n2612 );
or ( n2614 , n2613 , n1147 );
not ( n2615 , n74 );
or ( n2616 , n2615 , n199 );
nand ( n2617 , n2614 , n2616 );
not ( n2618 , n165 );
not ( n2619 , n2471 );
nor ( n2620 , n2619 , n1281 );
not ( n2621 , n1202 );
and ( n2622 , n2621 , n2472 );
nor ( n2623 , n2622 , n1223 );
nor ( n2624 , n1205 , n2623 );
not ( n2625 , n1243 );
not ( n2626 , n2472 );
and ( n2627 , n2625 , n2626 );
and ( n2628 , n1236 , n1225 );
nor ( n2629 , n2627 , n2628 );
nand ( n2630 , n2624 , n2629 , n2514 );
nand ( n2631 , n1293 , n1249 );
not ( n2632 , n1210 );
not ( n2633 , n1252 );
or ( n2634 , n2632 , n2633 );
nand ( n2635 , n2634 , n2482 );
nand ( n2636 , n2635 , n1234 );
nand ( n2637 , n2631 , n2508 , n2636 );
nor ( n2638 , n2630 , n2637 );
not ( n2639 , n1228 );
or ( n2640 , n1208 , n1210 );
nand ( n2641 , n2640 , n1237 );
not ( n2642 , n2641 );
or ( n2643 , n2639 , n2642 );
or ( n2644 , n1277 , n2481 );
and ( n2645 , n2644 , n1276 , n1286 );
nor ( n2646 , n2645 , n1176 );
nand ( n2647 , n2643 , n2646 );
nand ( n2648 , n1290 , n2647 );
nand ( n2649 , n2620 , n2638 , n2648 );
not ( n2650 , n2649 );
or ( n2651 , n2618 , n2650 );
or ( n2652 , n2649 , n165 );
nand ( n2653 , n2651 , n2652 );
or ( n2654 , n2653 , n855 );
and ( n2655 , n671 , n108 );
and ( n2656 , n673 , n116 );
nor ( n2657 , n2655 , n2656 );
nand ( n2658 , n2654 , n2657 );
not ( n2659 , n2147 );
nand ( n2660 , n2182 , n2378 );
not ( n2661 , n2660 );
or ( n2662 , n2659 , n2661 );
nor ( n2663 , n2114 , n2104 );
and ( n2664 , n2130 , n2663 );
not ( n2665 , n2172 );
and ( n2666 , n2665 , n2186 );
nor ( n2667 , n2664 , n2666 );
nand ( n2668 , n2662 , n2667 );
nor ( n2669 , n2149 , n2668 );
not ( n2670 , n2202 );
not ( n2671 , n2181 );
or ( n2672 , n2670 , n2671 );
not ( n2673 , n2157 );
not ( n2674 , n2104 );
and ( n2675 , n2673 , n2674 );
nor ( n2676 , n2675 , n2384 );
nand ( n2677 , n2672 , n2676 );
and ( n2678 , n2231 , n2409 );
nor ( n2679 , n2678 , n2201 );
nor ( n2680 , n2677 , n2679 );
nand ( n2681 , n2218 , n2168 );
not ( n2682 , n2681 );
nand ( n2683 , n2682 , n2386 , n2217 , n2201 );
not ( n2684 , n2201 );
not ( n2685 , n2681 );
or ( n2686 , n2684 , n2685 );
nand ( n2687 , n2686 , n2162 );
nand ( n2688 , n2683 , n2687 );
not ( n2689 , n2229 );
not ( n2690 , n2689 );
nor ( n2691 , n2393 , n2161 );
not ( n2692 , n2691 );
or ( n2693 , n2690 , n2692 );
nand ( n2694 , n2693 , n2186 );
nand ( n2695 , n2669 , n2680 , n2688 , n2694 );
and ( n2696 , n2695 , n172 );
not ( n2697 , n2695 );
not ( n2698 , n172 );
and ( n2699 , n2697 , n2698 );
or ( n2700 , n2696 , n2699 );
or ( n2701 , n2700 , n1147 );
and ( n2702 , n671 , n118 );
and ( n2703 , n673 , n126 );
nor ( n2704 , n2702 , n2703 );
nand ( n2705 , n2701 , n2704 );
not ( n2706 , n2197 );
not ( n2707 , n2178 );
or ( n2708 , n2706 , n2707 );
nand ( n2709 , n2708 , n2186 );
nand ( n2710 , n2681 , n2097 );
nand ( n2711 , n2709 , n2710 , n2216 , n2391 );
nor ( n2712 , n2711 , n2401 );
not ( n2713 , n2410 );
not ( n2714 , n2227 );
or ( n2715 , n2713 , n2714 );
or ( n2716 , n2098 , n2128 );
nand ( n2717 , n2716 , n2114 , n2211 );
or ( n2718 , n2717 , n2213 );
nand ( n2719 , n2718 , n2164 );
nand ( n2720 , n2715 , n2719 );
nand ( n2721 , n2403 , n2105 );
not ( n2722 , n2173 );
nand ( n2723 , n2192 , n2156 , n2410 , n2116 );
nand ( n2724 , n2720 , n2721 , n2722 , n2723 );
nor ( n2725 , n2677 , n2724 );
nand ( n2726 , n2712 , n2725 );
and ( n2727 , n2726 , n180 );
not ( n2728 , n2726 );
not ( n2729 , n180 );
and ( n2730 , n2728 , n2729 );
nor ( n2731 , n2727 , n2730 );
nand ( n2732 , n2731 , n664 );
and ( n2733 , n671 , n120 );
and ( n2734 , n673 , n128 );
nor ( n2735 , n2733 , n2734 );
nand ( n2736 , n2732 , n2735 );
or ( n2737 , n2653 , n1146 );
not ( n2738 , n61 );
or ( n2739 , n1362 , n2738 );
nand ( n2740 , n2737 , n2739 );
or ( n2741 , n2420 , n846 );
not ( n2742 , n1429 );
not ( n2743 , n53 );
or ( n2744 , n2742 , n2743 );
nand ( n2745 , n2741 , n2744 );
or ( n2746 , n2700 , n846 );
not ( n2747 , n4 );
or ( n2748 , n1362 , n2747 );
nand ( n2749 , n2746 , n2748 );
not ( n2750 , n2731 );
or ( n2751 , n2750 , n846 );
not ( n2752 , n6 );
or ( n2753 , n1362 , n2752 );
nand ( n2754 , n2751 , n2753 );
or ( n2755 , n2520 , n846 );
not ( n2756 , n17 );
or ( n2757 , n849 , n2756 );
nand ( n2758 , n2755 , n2757 );
or ( n2759 , n2544 , n2354 );
not ( n2760 , n51 );
or ( n2761 , n1362 , n2760 );
nand ( n2762 , n2759 , n2761 );
or ( n2763 , n2613 , n1146 );
not ( n2764 , n19 );
or ( n2765 , n1430 , n2764 );
nand ( n2766 , n2763 , n2765 );
or ( n2767 , n2460 , n846 );
not ( n2768 , n29 );
or ( n2769 , n1430 , n2768 );
nand ( n2770 , n2767 , n2769 );
not ( n2771 , n179 );
not ( n2772 , n1271 );
not ( n2773 , n1279 );
not ( n2774 , n1201 );
nand ( n2775 , n2774 , n1167 , n1169 );
nand ( n2776 , n2772 , n2773 , n2775 );
nor ( n2777 , n2776 , n1247 );
and ( n2778 , n1288 , n1266 );
nor ( n2779 , n2778 , n1176 );
and ( n2780 , n2779 , n2477 );
nor ( n2781 , n2780 , n2637 );
nand ( n2782 , n2501 , n2777 , n2781 );
not ( n2783 , n2782 );
or ( n2784 , n2771 , n2783 );
or ( n2785 , n2782 , n179 );
nand ( n2786 , n2784 , n2785 );
or ( n2787 , n2786 , n846 );
not ( n2788 , n15 );
or ( n2789 , n1413 , n2788 );
nand ( n2790 , n2787 , n2789 );
not ( n2791 , n631 );
nand ( n2792 , n1326 , n2791 );
nor ( n2793 , n2792 , n1064 );
not ( n2794 , n591 );
not ( n2795 , n517 );
not ( n2796 , n554 );
or ( n2797 , n2795 , n2796 );
not ( n2798 , n547 );
nand ( n2799 , n2798 , n563 );
nand ( n2800 , n2797 , n2799 );
not ( n2801 , n2800 );
or ( n2802 , n2794 , n2801 );
nand ( n2803 , n2802 , n648 );
nor ( n2804 , n2803 , n1074 );
nand ( n2805 , n533 , n596 );
nand ( n2806 , n2805 , n1311 , n644 );
nor ( n2807 , n2806 , n582 );
nand ( n2808 , n2793 , n2804 , n2807 );
and ( n2809 , n2808 , n178 );
not ( n2810 , n2808 );
not ( n2811 , n178 );
and ( n2812 , n2810 , n2811 );
or ( n2813 , n2809 , n2812 );
or ( n2814 , n2813 , n1147 );
and ( n2815 , n671 , n70 );
and ( n2816 , n673 , n78 );
nor ( n2817 , n2815 , n2816 );
nand ( n2818 , n2814 , n2817 );
not ( n2819 , n2045 );
not ( n2820 , n1945 );
not ( n2821 , n1975 );
or ( n2822 , n2820 , n2821 );
nand ( n2823 , n2024 , n2010 );
or ( n2824 , n2823 , n1945 );
nand ( n2825 , n2822 , n2824 );
nand ( n2826 , n2825 , n1977 );
not ( n2827 , n2033 );
not ( n2828 , n1980 );
and ( n2829 , n2827 , n2828 );
nor ( n2830 , n2829 , n2056 );
nand ( n2831 , n2074 , n2826 , n2830 );
not ( n2832 , n2009 );
not ( n2833 , n2589 );
or ( n2834 , n2832 , n2833 );
not ( n2835 , n2591 );
not ( n2836 , n1992 );
or ( n2837 , n2835 , n2836 );
nand ( n2838 , n2837 , n2063 );
nand ( n2839 , n2838 , n1964 );
nand ( n2840 , n2834 , n2839 );
nor ( n2841 , n2831 , n2583 , n2840 );
not ( n2842 , n2604 );
not ( n2843 , n1964 );
or ( n2844 , n2842 , n2843 );
not ( n2845 , n2063 );
nand ( n2846 , n2845 , n1981 );
nand ( n2847 , n2844 , n2846 );
nor ( n2848 , n2575 , n2847 , n2079 );
nand ( n2849 , n2819 , n2841 , n2848 );
xnor ( n2850 , n2849 , n170 );
or ( n2851 , n2850 , n846 );
not ( n2852 , n21 );
or ( n2853 , n2742 , n2852 );
nand ( n2854 , n2851 , n2853 );
or ( n2855 , n2813 , n846 );
not ( n2856 , n23 );
or ( n2857 , n855 , n2856 );
nand ( n2858 , n2855 , n2857 );
or ( n2859 , n2850 , n1147 );
and ( n2860 , n1037 , n68 );
and ( n2861 , n673 , n76 );
nor ( n2862 , n2860 , n2861 );
nand ( n2863 , n2859 , n2862 );
or ( n2864 , n2786 , n1147 );
not ( n2865 , n70 );
or ( n2866 , n2865 , n199 );
nand ( n2867 , n2864 , n2866 );
not ( n2868 , n186 );
not ( n2869 , n2868 );
not ( n2870 , n2080 );
nand ( n2871 , n2870 , n2556 );
nor ( n2872 , n2871 , n2607 );
and ( n2873 , n2598 , n2036 );
nor ( n2874 , n2873 , n2847 );
nand ( n2875 , n2872 , n2874 , n2044 );
or ( n2876 , n1984 , n2009 );
nand ( n2877 , n2876 , n2039 );
not ( n2878 , n2877 );
not ( n2879 , n2823 );
not ( n2880 , n2879 );
or ( n2881 , n2878 , n2880 );
nand ( n2882 , n2881 , n1978 );
nor ( n2883 , n2573 , n2882 );
nand ( n2884 , n2065 , n2033 , n2013 );
nand ( n2885 , n2884 , n1964 );
nand ( n2886 , n2883 , n2017 , n2026 , n2885 );
nor ( n2887 , n2875 , n2886 );
not ( n2888 , n2887 );
or ( n2889 , n2869 , n2888 );
or ( n2890 , n2887 , n2868 );
nand ( n2891 , n2889 , n2890 );
or ( n2892 , n2891 , n846 );
not ( n2893 , n25 );
or ( n2894 , n1362 , n2893 );
nand ( n2895 , n2892 , n2894 );
not ( n2896 , n171 );
not ( n2897 , n1746 );
not ( n2898 , n1791 );
and ( n2899 , n2897 , n2898 );
nor ( n2900 , n1771 , n1757 );
and ( n2901 , n2900 , n1775 );
nor ( n2902 , n2899 , n2901 );
nand ( n2903 , n2902 , n2248 );
nand ( n2904 , n1878 , n2247 );
nor ( n2905 , n2903 , n2904 );
and ( n2906 , n1863 , n1873 );
not ( n2907 , n1805 );
not ( n2908 , n1850 );
or ( n2909 , n2907 , n2908 );
nand ( n2910 , n2909 , n1810 );
nand ( n2911 , n1835 , n1844 , n2278 );
and ( n2912 , n2282 , n2910 , n2911 );
and ( n2913 , n2905 , n2906 , n2912 );
not ( n2914 , n2268 );
nand ( n2915 , n2913 , n1794 , n2914 );
not ( n2916 , n2915 );
or ( n2917 , n2896 , n2916 );
or ( n2918 , n2915 , n171 );
nand ( n2919 , n2917 , n2918 );
or ( n2920 , n2919 , n1147 );
not ( n2921 , n68 );
or ( n2922 , n2921 , n199 );
nand ( n2923 , n2920 , n2922 );
or ( n2924 , n2891 , n1147 );
and ( n2925 , n1037 , n72 );
and ( n2926 , n673 , n80 );
nor ( n2927 , n2925 , n2926 );
nand ( n2928 , n2924 , n2927 );
not ( n2929 , n1866 );
nand ( n2930 , n1785 , n1797 , n1788 );
nand ( n2931 , n1810 , n2930 );
not ( n2932 , n2931 );
or ( n2933 , n2929 , n2932 );
nand ( n2934 , n2933 , n1777 );
not ( n2935 , n1834 );
and ( n2936 , n2258 , n1799 , n2935 );
not ( n2937 , n1874 );
nand ( n2938 , n2266 , n1792 );
not ( n2939 , n1762 );
not ( n2940 , n1861 );
or ( n2941 , n2939 , n2940 );
nand ( n2942 , n2941 , n2278 );
nand ( n2943 , n1776 , n2938 , n2942 );
nor ( n2944 , n2943 , n2903 );
nand ( n2945 , n2934 , n2936 , n2937 , n2944 );
xnor ( n2946 , n2945 , n188 );
or ( n2947 , n2946 , n1147 );
and ( n2948 , n1037 , n122 );
and ( n2949 , n673 , n130 );
nor ( n2950 , n2948 , n2949 );
nand ( n2951 , n2947 , n2950 );
or ( n2952 , n2919 , n846 );
not ( n2953 , n13 );
or ( n2954 , n1362 , n2953 );
nand ( n2955 , n2952 , n2954 );
or ( n2956 , n2946 , n846 );
not ( n2957 , n8 );
or ( n2958 , n1430 , n2957 );
nand ( n2959 , n2956 , n2958 );
and ( n2960 , n10 , n256 );
not ( n2961 , n10 );
not ( n2962 , n256 );
and ( n2963 , n2961 , n2962 );
nor ( n2964 , n2960 , n2963 );
nand ( n2965 , n660 , n2964 );
nand ( n2966 , n660 , n11 );
nand ( n2967 , n2965 , n2966 , n256 );
not ( n2968 , n2967 );
not ( n2969 , n197 );
not ( n2970 , n196 );
nand ( n2971 , n197 , n198 , n199 );
nand ( n2972 , n2970 , n2971 );
nand ( n2973 , n2972 , n198 );
not ( n2974 , n2973 );
or ( n2975 , n2969 , n2974 );
not ( n2976 , n196 );
nor ( n2977 , n198 , n199 );
nand ( n2978 , n2976 , n2977 );
not ( n2979 , n197 );
nand ( n2980 , n2978 , n2979 );
nand ( n2981 , n2975 , n2980 );
buf ( n2982 , n2981 );
nand ( n2983 , n2982 , n205 );
and ( n2984 , n2979 , n2978 );
not ( n2985 , n2979 );
and ( n2986 , n2985 , n2973 );
nor ( n2987 , n2984 , n2986 );
buf ( n2988 , n2987 );
nand ( n2989 , n2988 , n206 );
nand ( n2990 , n2968 , n2983 , n2989 );
and ( n2991 , n2966 , n2965 , n2962 );
buf ( n2992 , n2991 );
nand ( n2993 , n2982 , n209 );
nand ( n2994 , n2988 , n208 );
nand ( n2995 , n2992 , n2993 , n2994 );
nand ( n2996 , n2990 , n2995 );
nor ( n2997 , n9 , n10 );
buf ( n2998 , n2997 );
and ( n2999 , n2998 , n49 );
not ( n3000 , n9 );
nand ( n3001 , n3000 , n10 );
not ( n3002 , n3001 );
and ( n3003 , n3002 , n57 );
nor ( n3004 , n2999 , n3003 );
not ( n3005 , n3004 );
nand ( n3006 , n2966 , n3000 );
buf ( n3007 , n3006 );
not ( n3008 , n3007 );
or ( n3009 , n3005 , n3008 );
not ( n3010 , n2965 );
nand ( n3011 , n3010 , n2966 );
buf ( n3012 , n3011 );
or ( n3013 , n3012 , n207 );
nand ( n3014 , n3009 , n3013 );
nor ( n3015 , n2996 , n3014 );
nand ( n3016 , n2982 , n238 );
nand ( n3017 , n239 , n2988 );
nand ( n3018 , n2968 , n3016 , n3017 );
nand ( n3019 , n2982 , n242 );
nand ( n3020 , n2988 , n241 );
nand ( n3021 , n2992 , n3019 , n3020 );
nand ( n3022 , n3018 , n3021 );
and ( n3023 , n2998 , n3 );
and ( n3024 , n3002 , n15 );
nor ( n3025 , n3023 , n3024 );
not ( n3026 , n3025 );
not ( n3027 , n3007 );
or ( n3028 , n3026 , n3027 );
or ( n3029 , n3012 , n240 );
nand ( n3030 , n3028 , n3029 );
nor ( n3031 , n3022 , n3030 );
nand ( n3032 , n2982 , n210 );
nand ( n3033 , n211 , n2988 );
nand ( n3034 , n2968 , n3032 , n3033 );
nand ( n3035 , n2982 , n214 );
nand ( n3036 , n213 , n2988 );
nand ( n3037 , n2992 , n3035 , n3036 );
nand ( n3038 , n3034 , n3037 );
and ( n3039 , n2998 , n7 );
and ( n3040 , n3002 , n17 );
nor ( n3041 , n3039 , n3040 );
not ( n3042 , n3041 );
not ( n3043 , n3007 );
or ( n3044 , n3042 , n3043 );
or ( n3045 , n3012 , n212 );
nand ( n3046 , n3044 , n3045 );
nor ( n3047 , n3038 , n3046 );
nand ( n3048 , n2982 , n206 );
nand ( n3049 , n2988 , n207 );
nand ( n3050 , n2968 , n3048 , n3049 );
nand ( n3051 , n209 , n2988 );
nand ( n3052 , n3051 , n3032 , n2992 );
nand ( n3053 , n3050 , n3052 );
and ( n3054 , n2998 , n41 );
and ( n3055 , n3002 , n49 );
nor ( n3056 , n3054 , n3055 );
not ( n3057 , n3056 );
not ( n3058 , n3007 );
or ( n3059 , n3057 , n3058 );
or ( n3060 , n3012 , n208 );
nand ( n3061 , n3059 , n3060 );
nor ( n3062 , n3053 , n3061 );
nand ( n3063 , n243 , n2988 );
nand ( n3064 , n2968 , n3019 , n3063 );
nand ( n3065 , n2982 , n246 );
nand ( n3066 , n2988 , n245 );
nand ( n3067 , n2992 , n3065 , n3066 );
nand ( n3068 , n3064 , n3067 );
and ( n3069 , n2998 , n38 );
and ( n3070 , n3002 , n46 );
nor ( n3071 , n3069 , n3070 );
not ( n3072 , n3071 );
not ( n3073 , n3007 );
or ( n3074 , n3072 , n3073 );
or ( n3075 , n3012 , n244 );
nand ( n3076 , n3074 , n3075 );
nor ( n3077 , n3068 , n3076 );
nand ( n3078 , n2982 , n230 );
nand ( n3079 , n231 , n2988 );
nand ( n3080 , n2968 , n3078 , n3079 );
nand ( n3081 , n2982 , n234 );
nand ( n3082 , n233 , n2988 );
nand ( n3083 , n2992 , n3081 , n3082 );
nand ( n3084 , n3080 , n3083 );
and ( n3085 , n2998 , n4 );
and ( n3086 , n3002 , n48 );
nor ( n3087 , n3085 , n3086 );
not ( n3088 , n3087 );
not ( n3089 , n3007 );
or ( n3090 , n3088 , n3089 );
or ( n3091 , n3012 , n232 );
nand ( n3092 , n3090 , n3091 );
nor ( n3093 , n3084 , n3092 );
nand ( n3094 , n2982 , n254 );
nand ( n3095 , n2988 , n255 );
nand ( n3096 , n2968 , n3094 , n3095 );
nand ( n3097 , n229 , n2988 );
nand ( n3098 , n3097 , n3078 , n2992 );
nand ( n3099 , n3096 , n3098 );
and ( n3100 , n2998 , n5 );
and ( n3101 , n3002 , n13 );
nor ( n3102 , n3100 , n3101 );
not ( n3103 , n3102 );
not ( n3104 , n3007 );
or ( n3105 , n3103 , n3104 );
or ( n3106 , n3012 , n228 );
nand ( n3107 , n3105 , n3106 );
nor ( n3108 , n3099 , n3107 );
nand ( n3109 , n2988 , n215 );
nand ( n3110 , n2968 , n3035 , n3109 );
nand ( n3111 , n2982 , n218 );
nand ( n3112 , n2988 , n217 );
nand ( n3113 , n2992 , n3111 , n3112 );
nand ( n3114 , n3110 , n3113 );
and ( n3115 , n2998 , n42 );
and ( n3116 , n3002 , n50 );
nor ( n3117 , n3115 , n3116 );
not ( n3118 , n3117 );
not ( n3119 , n3007 );
or ( n3120 , n3118 , n3119 );
or ( n3121 , n3012 , n216 );
nand ( n3122 , n3120 , n3121 );
nor ( n3123 , n3114 , n3122 );
nand ( n3124 , n2988 , n223 );
nand ( n3125 , n2982 , n222 );
nand ( n3126 , n3124 , n3125 , n2968 );
nand ( n3127 , n2982 , n226 );
nand ( n3128 , n2988 , n225 );
nand ( n3129 , n2992 , n3127 , n3128 );
nand ( n3130 , n3126 , n3129 );
and ( n3131 , n2998 , n43 );
and ( n3132 , n3002 , n51 );
nor ( n3133 , n3131 , n3132 );
not ( n3134 , n3133 );
not ( n3135 , n3007 );
or ( n3136 , n3134 , n3135 );
or ( n3137 , n3012 , n224 );
nand ( n3138 , n3136 , n3137 );
nor ( n3139 , n3130 , n3138 );
nand ( n3140 , n2988 , n219 );
nand ( n3141 , n2968 , n3111 , n3140 );
nand ( n3142 , n2988 , n221 );
nand ( n3143 , n2992 , n3125 , n3142 );
nand ( n3144 , n3141 , n3143 );
and ( n3145 , n2998 , n8 );
and ( n3146 , n3002 , n18 );
nor ( n3147 , n3145 , n3146 );
not ( n3148 , n3147 );
not ( n3149 , n3007 );
or ( n3150 , n3148 , n3149 );
or ( n3151 , n3012 , n220 );
nand ( n3152 , n3150 , n3151 );
nor ( n3153 , n3144 , n3152 );
nand ( n3154 , n247 , n2988 );
nand ( n3155 , n2968 , n3065 , n3154 );
nand ( n3156 , n2982 , n250 );
nand ( n3157 , n2988 , n249 );
nand ( n3158 , n2992 , n3156 , n3157 );
nand ( n3159 , n3155 , n3158 );
and ( n3160 , n2998 , n2 );
and ( n3161 , n3002 , n14 );
nor ( n3162 , n3160 , n3161 );
not ( n3163 , n3162 );
not ( n3164 , n3007 );
or ( n3165 , n3163 , n3164 );
or ( n3166 , n3012 , n248 );
nand ( n3167 , n3165 , n3166 );
nor ( n3168 , n3159 , n3167 );
nand ( n3169 , n2988 , n227 );
nand ( n3170 , n2968 , n3127 , n3169 );
nand ( n3171 , n201 , n2988 );
nand ( n3172 , n2982 , n202 );
nand ( n3173 , n3171 , n3172 , n2992 );
nand ( n3174 , n3170 , n3173 );
and ( n3175 , n2998 , n40 );
and ( n3176 , n3002 , n19 );
nor ( n3177 , n3175 , n3176 );
not ( n3178 , n3177 );
not ( n3179 , n3007 );
or ( n3180 , n3178 , n3179 );
or ( n3181 , n3012 , n200 );
nand ( n3182 , n3180 , n3181 );
nor ( n3183 , n3174 , n3182 );
nand ( n3184 , n2982 , n227 );
nand ( n3185 , n200 , n2988 );
nand ( n3186 , n2968 , n3184 , n3185 );
nand ( n3187 , n2982 , n203 );
nand ( n3188 , n2988 , n202 );
nand ( n3189 , n2992 , n3187 , n3188 );
nand ( n3190 , n3186 , n3189 );
and ( n3191 , n2998 , n32 );
and ( n3192 , n3002 , n40 );
nor ( n3193 , n3191 , n3192 );
not ( n3194 , n3193 );
not ( n3195 , n3007 );
or ( n3196 , n3194 , n3195 );
or ( n3197 , n3012 , n201 );
nand ( n3198 , n3196 , n3197 );
nor ( n3199 , n3190 , n3198 );
nand ( n3200 , n2982 , n200 );
nand ( n3201 , n2968 , n3200 , n3171 );
nand ( n3202 , n2982 , n204 );
nand ( n3203 , n203 , n2988 );
nand ( n3204 , n2992 , n3202 , n3203 );
nand ( n3205 , n3201 , n3204 );
and ( n3206 , n2998 , n24 );
and ( n3207 , n3002 , n32 );
nor ( n3208 , n3206 , n3207 );
not ( n3209 , n3208 );
not ( n3210 , n3007 );
or ( n3211 , n3209 , n3210 );
or ( n3212 , n3012 , n202 );
nand ( n3213 , n3211 , n3212 );
nor ( n3214 , n3205 , n3213 );
nand ( n3215 , n2982 , n201 );
nand ( n3216 , n2968 , n3215 , n3188 );
nand ( n3217 , n204 , n2988 );
nand ( n3218 , n3217 , n2983 , n2992 );
nand ( n3219 , n3216 , n3218 );
and ( n3220 , n2998 , n16 );
and ( n3221 , n3002 , n24 );
nor ( n3222 , n3220 , n3221 );
not ( n3223 , n3222 );
not ( n3224 , n3007 );
or ( n3225 , n3223 , n3224 );
or ( n3226 , n3012 , n203 );
nand ( n3227 , n3225 , n3226 );
nor ( n3228 , n3219 , n3227 );
nand ( n3229 , n2968 , n3172 , n3203 );
nand ( n3230 , n2988 , n205 );
nand ( n3231 , n2992 , n3048 , n3230 );
nand ( n3232 , n3229 , n3231 );
and ( n3233 , n2998 , n6 );
and ( n3234 , n3002 , n16 );
nor ( n3235 , n3233 , n3234 );
not ( n3236 , n3235 );
not ( n3237 , n3007 );
or ( n3238 , n3236 , n3237 );
or ( n3239 , n3012 , n204 );
nand ( n3240 , n3238 , n3239 );
nor ( n3241 , n3232 , n3240 );
nand ( n3242 , n2968 , n3187 , n3217 );
nand ( n3243 , n2982 , n207 );
nand ( n3244 , n2992 , n3243 , n2989 );
nand ( n3245 , n3242 , n3244 );
and ( n3246 , n2998 , n65 );
and ( n3247 , n3002 , n6 );
nor ( n3248 , n3246 , n3247 );
not ( n3249 , n3248 );
not ( n3250 , n3007 );
or ( n3251 , n3249 , n3250 );
or ( n3252 , n3012 , n205 );
nand ( n3253 , n3251 , n3252 );
nor ( n3254 , n3245 , n3253 );
nand ( n3255 , n2968 , n3202 , n3230 );
nand ( n3256 , n2982 , n208 );
nand ( n3257 , n2992 , n3256 , n3049 );
nand ( n3258 , n3255 , n3257 );
and ( n3259 , n2998 , n57 );
and ( n3260 , n3002 , n65 );
nor ( n3261 , n3259 , n3260 );
not ( n3262 , n3261 );
not ( n3263 , n3007 );
or ( n3264 , n3262 , n3263 );
or ( n3265 , n3012 , n206 );
nand ( n3266 , n3264 , n3265 );
nor ( n3267 , n3258 , n3266 );
nand ( n3268 , n2968 , n3243 , n2994 );
nand ( n3269 , n2988 , n210 );
nand ( n3270 , n2982 , n211 );
nand ( n3271 , n3269 , n3270 , n2992 );
nand ( n3272 , n3268 , n3271 );
and ( n3273 , n2998 , n33 );
and ( n3274 , n3002 , n41 );
nor ( n3275 , n3273 , n3274 );
not ( n3276 , n3275 );
not ( n3277 , n3007 );
or ( n3278 , n3276 , n3277 );
or ( n3279 , n3012 , n209 );
nand ( n3280 , n3278 , n3279 );
nor ( n3281 , n3272 , n3280 );
nand ( n3282 , n2968 , n3256 , n3051 );
nand ( n3283 , n2982 , n212 );
nand ( n3284 , n2992 , n3283 , n3033 );
nand ( n3285 , n3282 , n3284 );
and ( n3286 , n2998 , n25 );
and ( n3287 , n3002 , n33 );
nor ( n3288 , n3286 , n3287 );
not ( n3289 , n3288 );
not ( n3290 , n3007 );
or ( n3291 , n3289 , n3290 );
or ( n3292 , n3012 , n210 );
nand ( n3293 , n3291 , n3292 );
nor ( n3294 , n3285 , n3293 );
nand ( n3295 , n2968 , n2993 , n3269 );
nand ( n3296 , n2982 , n213 );
nand ( n3297 , n212 , n2988 );
nand ( n3298 , n2992 , n3296 , n3297 );
nand ( n3299 , n3295 , n3298 );
and ( n3300 , n2998 , n17 );
and ( n3301 , n3002 , n25 );
nor ( n3302 , n3300 , n3301 );
not ( n3303 , n3302 );
not ( n3304 , n3007 );
or ( n3305 , n3303 , n3304 );
or ( n3306 , n3012 , n211 );
nand ( n3307 , n3305 , n3306 );
nor ( n3308 , n3299 , n3307 );
nand ( n3309 , n2968 , n3270 , n3297 );
nand ( n3310 , n2982 , n215 );
nand ( n3311 , n214 , n2988 );
nand ( n3312 , n2992 , n3310 , n3311 );
nand ( n3313 , n3309 , n3312 );
and ( n3314 , n2998 , n66 );
and ( n3315 , n3002 , n7 );
nor ( n3316 , n3314 , n3315 );
not ( n3317 , n3316 );
not ( n3318 , n3007 );
or ( n3319 , n3317 , n3318 );
or ( n3320 , n3012 , n213 );
nand ( n3321 , n3319 , n3320 );
nor ( n3322 , n3313 , n3321 );
nand ( n3323 , n2968 , n3283 , n3036 );
nand ( n3324 , n2982 , n216 );
nand ( n3325 , n2992 , n3324 , n3109 );
nand ( n3326 , n3323 , n3325 );
and ( n3327 , n2998 , n58 );
and ( n3328 , n3002 , n66 );
nor ( n3329 , n3327 , n3328 );
not ( n3330 , n3329 );
not ( n3331 , n3007 );
or ( n3332 , n3330 , n3331 );
or ( n3333 , n3012 , n214 );
nand ( n3334 , n3332 , n3333 );
nor ( n3335 , n3326 , n3334 );
nand ( n3336 , n2968 , n3296 , n3311 );
nand ( n3337 , n2982 , n217 );
nand ( n3338 , n216 , n2988 );
nand ( n3339 , n2992 , n3337 , n3338 );
nand ( n3340 , n3336 , n3339 );
and ( n3341 , n2998 , n50 );
and ( n3342 , n3002 , n58 );
nor ( n3343 , n3341 , n3342 );
not ( n3344 , n3343 );
not ( n3345 , n3007 );
or ( n3346 , n3344 , n3345 );
or ( n3347 , n3012 , n215 );
nand ( n3348 , n3346 , n3347 );
nor ( n3349 , n3340 , n3348 );
nand ( n3350 , n2968 , n3310 , n3338 );
nand ( n3351 , n2982 , n219 );
nand ( n3352 , n2988 , n218 );
nand ( n3353 , n2992 , n3351 , n3352 );
nand ( n3354 , n3350 , n3353 );
and ( n3355 , n2998 , n34 );
and ( n3356 , n3002 , n42 );
nor ( n3357 , n3355 , n3356 );
not ( n3358 , n3357 );
not ( n3359 , n3007 );
or ( n3360 , n3358 , n3359 );
or ( n3361 , n3012 , n217 );
nand ( n3362 , n3360 , n3361 );
nor ( n3363 , n3354 , n3362 );
nand ( n3364 , n2968 , n3324 , n3112 );
nand ( n3365 , n2982 , n220 );
nand ( n3366 , n2992 , n3365 , n3140 );
nand ( n3367 , n3364 , n3366 );
and ( n3368 , n2998 , n26 );
and ( n3369 , n3002 , n34 );
nor ( n3370 , n3368 , n3369 );
not ( n3371 , n3370 );
not ( n3372 , n3007 );
or ( n3373 , n3371 , n3372 );
or ( n3374 , n3012 , n218 );
nand ( n3375 , n3373 , n3374 );
nor ( n3376 , n3367 , n3375 );
nand ( n3377 , n2968 , n3337 , n3352 );
nand ( n3378 , n220 , n2988 );
nand ( n3379 , n2982 , n221 );
nand ( n3380 , n3378 , n3379 , n2992 );
nand ( n3381 , n3377 , n3380 );
and ( n3382 , n2998 , n18 );
and ( n3383 , n3002 , n26 );
nor ( n3384 , n3382 , n3383 );
not ( n3385 , n3384 );
not ( n3386 , n3007 );
or ( n3387 , n3385 , n3386 );
or ( n3388 , n3012 , n219 );
nand ( n3389 , n3387 , n3388 );
nor ( n3390 , n3381 , n3389 );
nand ( n3391 , n2968 , n3351 , n3378 );
nand ( n3392 , n2982 , n223 );
nand ( n3393 , n2988 , n222 );
nand ( n3394 , n2992 , n3392 , n3393 );
nand ( n3395 , n3391 , n3394 );
and ( n3396 , n2998 , n67 );
and ( n3397 , n3002 , n8 );
nor ( n3398 , n3396 , n3397 );
not ( n3399 , n3398 );
not ( n3400 , n3007 );
or ( n3401 , n3399 , n3400 );
or ( n3402 , n3012 , n221 );
nand ( n3403 , n3401 , n3402 );
nor ( n3404 , n3395 , n3403 );
nand ( n3405 , n2968 , n3365 , n3142 );
nand ( n3406 , n2982 , n224 );
nand ( n3407 , n2992 , n3406 , n3124 );
nand ( n3408 , n3405 , n3407 );
and ( n3409 , n2998 , n59 );
and ( n3410 , n3002 , n67 );
nor ( n3411 , n3409 , n3410 );
not ( n3412 , n3411 );
not ( n3413 , n3007 );
or ( n3414 , n3412 , n3413 );
or ( n3415 , n3012 , n222 );
nand ( n3416 , n3414 , n3415 );
nor ( n3417 , n3408 , n3416 );
nand ( n3418 , n2968 , n3379 , n3393 );
nand ( n3419 , n224 , n2988 );
nand ( n3420 , n2982 , n225 );
nand ( n3421 , n3419 , n3420 , n2992 );
nand ( n3422 , n3418 , n3421 );
and ( n3423 , n2998 , n51 );
and ( n3424 , n3002 , n59 );
nor ( n3425 , n3423 , n3424 );
not ( n3426 , n3425 );
not ( n3427 , n3007 );
or ( n3428 , n3426 , n3427 );
or ( n3429 , n3012 , n223 );
nand ( n3430 , n3428 , n3429 );
nor ( n3431 , n3422 , n3430 );
nand ( n3432 , n2968 , n3392 , n3419 );
nand ( n3433 , n2988 , n226 );
nand ( n3434 , n2992 , n3184 , n3433 );
nand ( n3435 , n3432 , n3434 );
and ( n3436 , n2998 , n35 );
and ( n3437 , n3002 , n43 );
nor ( n3438 , n3436 , n3437 );
not ( n3439 , n3438 );
not ( n3440 , n3007 );
or ( n3441 , n3439 , n3440 );
or ( n3442 , n3012 , n225 );
nand ( n3443 , n3441 , n3442 );
nor ( n3444 , n3435 , n3443 );
nand ( n3445 , n2968 , n3406 , n3128 );
nand ( n3446 , n2992 , n3200 , n3169 );
nand ( n3447 , n3445 , n3446 );
and ( n3448 , n2998 , n27 );
and ( n3449 , n3002 , n35 );
nor ( n3450 , n3448 , n3449 );
not ( n3451 , n3450 );
not ( n3452 , n3007 );
or ( n3453 , n3451 , n3452 );
or ( n3454 , n3012 , n226 );
nand ( n3455 , n3453 , n3454 );
nor ( n3456 , n3447 , n3455 );
nand ( n3457 , n2968 , n3420 , n3433 );
nand ( n3458 , n3185 , n3215 , n2992 );
nand ( n3459 , n3457 , n3458 );
and ( n3460 , n2998 , n19 );
and ( n3461 , n3002 , n27 );
nor ( n3462 , n3460 , n3461 );
not ( n3463 , n3462 );
not ( n3464 , n3007 );
or ( n3465 , n3463 , n3464 );
or ( n3466 , n3012 , n227 );
nand ( n3467 , n3465 , n3466 );
nor ( n3468 , n3459 , n3467 );
nand ( n3469 , n2982 , n255 );
nand ( n3470 , n228 , n2988 );
nand ( n3471 , n2968 , n3469 , n3470 );
nand ( n3472 , n2982 , n231 );
nand ( n3473 , n2988 , n230 );
nand ( n3474 , n2992 , n3472 , n3473 );
nand ( n3475 , n3471 , n3474 );
and ( n3476 , n2998 , n64 );
and ( n3477 , n3002 , n5 );
nor ( n3478 , n3476 , n3477 );
not ( n3479 , n3478 );
not ( n3480 , n3007 );
or ( n3481 , n3479 , n3480 );
or ( n3482 , n3012 , n229 );
nand ( n3483 , n3481 , n3482 );
nor ( n3484 , n3475 , n3483 );
nand ( n3485 , n2982 , n228 );
nand ( n3486 , n2968 , n3485 , n3097 );
nand ( n3487 , n2982 , n232 );
nand ( n3488 , n2992 , n3487 , n3079 );
nand ( n3489 , n3486 , n3488 );
and ( n3490 , n2998 , n56 );
and ( n3491 , n3002 , n64 );
nor ( n3492 , n3490 , n3491 );
not ( n3493 , n3492 );
not ( n3494 , n3007 );
or ( n3495 , n3493 , n3494 );
or ( n3496 , n3012 , n230 );
nand ( n3497 , n3495 , n3496 );
nor ( n3498 , n3489 , n3497 );
nand ( n3499 , n232 , n2988 );
nand ( n3500 , n2968 , n3472 , n3499 );
nand ( n3501 , n2982 , n235 );
nand ( n3502 , n234 , n2988 );
nand ( n3503 , n2992 , n3501 , n3502 );
nand ( n3504 , n3500 , n3503 );
and ( n3505 , n2998 , n63 );
and ( n3506 , n3002 , n4 );
nor ( n3507 , n3505 , n3506 );
not ( n3508 , n3507 );
not ( n3509 , n3007 );
or ( n3510 , n3508 , n3509 );
or ( n3511 , n3012 , n233 );
nand ( n3512 , n3510 , n3511 );
nor ( n3513 , n3504 , n3512 );
nand ( n3514 , n2968 , n3487 , n3082 );
nand ( n3515 , n2982 , n236 );
nand ( n3516 , n235 , n2988 );
nand ( n3517 , n2992 , n3515 , n3516 );
nand ( n3518 , n3514 , n3517 );
and ( n3519 , n2998 , n55 );
and ( n3520 , n3002 , n63 );
nor ( n3521 , n3519 , n3520 );
not ( n3522 , n3521 );
not ( n3523 , n3007 );
or ( n3524 , n3522 , n3523 );
or ( n3525 , n3012 , n234 );
nand ( n3526 , n3524 , n3525 );
nor ( n3527 , n3518 , n3526 );
nand ( n3528 , n2982 , n233 );
nand ( n3529 , n2968 , n3528 , n3502 );
nand ( n3530 , n2982 , n237 );
nand ( n3531 , n2988 , n236 );
nand ( n3532 , n2992 , n3530 , n3531 );
nand ( n3533 , n3529 , n3532 );
and ( n3534 , n2998 , n47 );
and ( n3535 , n3002 , n55 );
nor ( n3536 , n3534 , n3535 );
not ( n3537 , n3536 );
not ( n3538 , n3007 );
or ( n3539 , n3537 , n3538 );
or ( n3540 , n3012 , n235 );
nand ( n3541 , n3539 , n3540 );
nor ( n3542 , n3533 , n3541 );
nand ( n3543 , n2968 , n3081 , n3516 );
nand ( n3544 , n237 , n2988 );
nand ( n3545 , n2992 , n3016 , n3544 );
nand ( n3546 , n3543 , n3545 );
and ( n3547 , n2998 , n39 );
and ( n3548 , n3002 , n47 );
nor ( n3549 , n3547 , n3548 );
not ( n3550 , n3549 );
not ( n3551 , n3007 );
or ( n3552 , n3550 , n3551 );
or ( n3553 , n3012 , n236 );
nand ( n3554 , n3552 , n3553 );
nor ( n3555 , n3546 , n3554 );
nand ( n3556 , n2968 , n3501 , n3531 );
nand ( n3557 , n2982 , n239 );
nand ( n3558 , n238 , n2988 );
nand ( n3559 , n3557 , n3558 , n2992 );
nand ( n3560 , n3556 , n3559 );
and ( n3561 , n2998 , n31 );
and ( n3562 , n3002 , n39 );
nor ( n3563 , n3561 , n3562 );
not ( n3564 , n3563 );
not ( n3565 , n3007 );
or ( n3566 , n3564 , n3565 );
or ( n3567 , n3012 , n237 );
nand ( n3568 , n3566 , n3567 );
nor ( n3569 , n3560 , n3568 );
nand ( n3570 , n2968 , n3515 , n3544 );
nand ( n3571 , n2982 , n240 );
nand ( n3572 , n2992 , n3571 , n3017 );
nand ( n3573 , n3570 , n3572 );
and ( n3574 , n2998 , n23 );
and ( n3575 , n3002 , n31 );
nor ( n3576 , n3574 , n3575 );
not ( n3577 , n3576 );
not ( n3578 , n3007 );
or ( n3579 , n3577 , n3578 );
or ( n3580 , n3012 , n238 );
nand ( n3581 , n3579 , n3580 );
nor ( n3582 , n3573 , n3581 );
nand ( n3583 , n2968 , n3530 , n3558 );
nand ( n3584 , n2982 , n241 );
nand ( n3585 , n2988 , n240 );
nand ( n3586 , n2992 , n3584 , n3585 );
nand ( n3587 , n3583 , n3586 );
and ( n3588 , n2998 , n15 );
and ( n3589 , n3002 , n23 );
nor ( n3590 , n3588 , n3589 );
not ( n3591 , n3590 );
not ( n3592 , n3007 );
or ( n3593 , n3591 , n3592 );
or ( n3594 , n3012 , n239 );
nand ( n3595 , n3593 , n3594 );
nor ( n3596 , n3587 , n3595 );
nand ( n3597 , n2968 , n3557 , n3585 );
nand ( n3598 , n2982 , n243 );
nand ( n3599 , n2988 , n242 );
nand ( n3600 , n2992 , n3598 , n3599 );
nand ( n3601 , n3597 , n3600 );
and ( n3602 , n2998 , n62 );
and ( n3603 , n3002 , n3 );
nor ( n3604 , n3602 , n3603 );
not ( n3605 , n3604 );
not ( n3606 , n3007 );
or ( n3607 , n3605 , n3606 );
or ( n3608 , n3012 , n241 );
nand ( n3609 , n3607 , n3608 );
nor ( n3610 , n3601 , n3609 );
nand ( n3611 , n2968 , n3571 , n3020 );
nand ( n3612 , n2982 , n244 );
nand ( n3613 , n2992 , n3612 , n3063 );
nand ( n3614 , n3611 , n3613 );
and ( n3615 , n2998 , n54 );
and ( n3616 , n3002 , n62 );
nor ( n3617 , n3615 , n3616 );
not ( n3618 , n3617 );
not ( n3619 , n3007 );
or ( n3620 , n3618 , n3619 );
or ( n3621 , n3012 , n242 );
nand ( n3622 , n3620 , n3621 );
nor ( n3623 , n3614 , n3622 );
nand ( n3624 , n2968 , n3584 , n3599 );
nand ( n3625 , n2982 , n245 );
nand ( n3626 , n2988 , n244 );
nand ( n3627 , n2992 , n3625 , n3626 );
nand ( n3628 , n3624 , n3627 );
and ( n3629 , n2998 , n46 );
and ( n3630 , n3002 , n54 );
nor ( n3631 , n3629 , n3630 );
not ( n3632 , n3631 );
not ( n3633 , n3007 );
or ( n3634 , n3632 , n3633 );
or ( n3635 , n3012 , n243 );
nand ( n3636 , n3634 , n3635 );
nor ( n3637 , n3628 , n3636 );
nand ( n3638 , n2968 , n3598 , n3626 );
nand ( n3639 , n2982 , n247 );
nand ( n3640 , n2988 , n246 );
nand ( n3641 , n2992 , n3639 , n3640 );
nand ( n3642 , n3638 , n3641 );
and ( n3643 , n2998 , n30 );
and ( n3644 , n3002 , n38 );
nor ( n3645 , n3643 , n3644 );
not ( n3646 , n3645 );
not ( n3647 , n3007 );
or ( n3648 , n3646 , n3647 );
or ( n3649 , n3012 , n245 );
nand ( n3650 , n3648 , n3649 );
nor ( n3651 , n3642 , n3650 );
nand ( n3652 , n2968 , n3612 , n3066 );
nand ( n3653 , n2982 , n248 );
nand ( n3654 , n3154 , n3653 , n2992 );
nand ( n3655 , n3652 , n3654 );
and ( n3656 , n2998 , n22 );
and ( n3657 , n3002 , n30 );
nor ( n3658 , n3656 , n3657 );
not ( n3659 , n3658 );
not ( n3660 , n3007 );
or ( n3661 , n3659 , n3660 );
or ( n3662 , n3012 , n246 );
nand ( n3663 , n3661 , n3662 );
nor ( n3664 , n3655 , n3663 );
nand ( n3665 , n2968 , n3625 , n3640 );
nand ( n3666 , n2982 , n249 );
nand ( n3667 , n248 , n2988 );
nand ( n3668 , n3666 , n3667 , n2992 );
nand ( n3669 , n3665 , n3668 );
and ( n3670 , n2998 , n14 );
and ( n3671 , n3002 , n22 );
nor ( n3672 , n3670 , n3671 );
not ( n3673 , n3672 );
not ( n3674 , n3007 );
or ( n3675 , n3673 , n3674 );
or ( n3676 , n3012 , n247 );
nand ( n3677 , n3675 , n3676 );
nor ( n3678 , n3669 , n3677 );
nand ( n3679 , n2968 , n3639 , n3667 );
nand ( n3680 , n2982 , n251 );
nand ( n3681 , n2988 , n250 );
nand ( n3682 , n2992 , n3680 , n3681 );
nand ( n3683 , n3679 , n3682 );
and ( n3684 , n2998 , n61 );
and ( n3685 , n3002 , n2 );
nor ( n3686 , n3684 , n3685 );
not ( n3687 , n3686 );
not ( n3688 , n3007 );
or ( n3689 , n3687 , n3688 );
or ( n3690 , n3012 , n249 );
nand ( n3691 , n3689 , n3690 );
nor ( n3692 , n3683 , n3691 );
nand ( n3693 , n2968 , n3653 , n3157 );
nand ( n3694 , n2982 , n252 );
nand ( n3695 , n251 , n2988 );
nand ( n3696 , n2992 , n3694 , n3695 );
nand ( n3697 , n3693 , n3696 );
and ( n3698 , n2998 , n53 );
and ( n3699 , n3002 , n61 );
nor ( n3700 , n3698 , n3699 );
not ( n3701 , n3700 );
not ( n3702 , n3007 );
or ( n3703 , n3701 , n3702 );
or ( n3704 , n3012 , n250 );
nand ( n3705 , n3703 , n3704 );
nor ( n3706 , n3697 , n3705 );
nand ( n3707 , n2968 , n3666 , n3681 );
nand ( n3708 , n2982 , n253 );
nand ( n3709 , n2988 , n252 );
nand ( n3710 , n2992 , n3708 , n3709 );
nand ( n3711 , n3707 , n3710 );
and ( n3712 , n2998 , n45 );
and ( n3713 , n3002 , n53 );
nor ( n3714 , n3712 , n3713 );
not ( n3715 , n3714 );
not ( n3716 , n3007 );
or ( n3717 , n3715 , n3716 );
or ( n3718 , n3012 , n251 );
nand ( n3719 , n3717 , n3718 );
nor ( n3720 , n3711 , n3719 );
nand ( n3721 , n2968 , n3156 , n3695 );
nand ( n3722 , n2988 , n253 );
nand ( n3723 , n2992 , n3094 , n3722 );
nand ( n3724 , n3721 , n3723 );
and ( n3725 , n2998 , n37 );
and ( n3726 , n3002 , n45 );
nor ( n3727 , n3725 , n3726 );
not ( n3728 , n3727 );
not ( n3729 , n3007 );
or ( n3730 , n3728 , n3729 );
or ( n3731 , n3012 , n252 );
nand ( n3732 , n3730 , n3731 );
nor ( n3733 , n3724 , n3732 );
nand ( n3734 , n2968 , n3680 , n3709 );
nand ( n3735 , n254 , n2988 );
nand ( n3736 , n3735 , n3469 , n2992 );
nand ( n3737 , n3734 , n3736 );
and ( n3738 , n2998 , n29 );
and ( n3739 , n3002 , n37 );
nor ( n3740 , n3738 , n3739 );
not ( n3741 , n3740 );
not ( n3742 , n3007 );
or ( n3743 , n3741 , n3742 );
or ( n3744 , n3012 , n253 );
nand ( n3745 , n3743 , n3744 );
nor ( n3746 , n3737 , n3745 );
nand ( n3747 , n2968 , n3694 , n3722 );
nand ( n3748 , n2992 , n3485 , n3095 );
nand ( n3749 , n3747 , n3748 );
and ( n3750 , n2998 , n21 );
and ( n3751 , n3002 , n29 );
nor ( n3752 , n3750 , n3751 );
not ( n3753 , n3752 );
not ( n3754 , n3007 );
or ( n3755 , n3753 , n3754 );
or ( n3756 , n3012 , n254 );
nand ( n3757 , n3755 , n3756 );
nor ( n3758 , n3749 , n3757 );
nand ( n3759 , n2968 , n3708 , n3735 );
nand ( n3760 , n2982 , n229 );
nand ( n3761 , n2992 , n3760 , n3470 );
nand ( n3762 , n3759 , n3761 );
and ( n3763 , n2998 , n13 );
and ( n3764 , n3002 , n21 );
nor ( n3765 , n3763 , n3764 );
not ( n3766 , n3765 );
not ( n3767 , n3007 );
or ( n3768 , n3766 , n3767 );
or ( n3769 , n3012 , n255 );
nand ( n3770 , n3768 , n3769 );
nor ( n3771 , n3762 , n3770 );
nand ( n3772 , n2968 , n3760 , n3473 );
nand ( n3773 , n2992 , n3528 , n3499 );
nand ( n3774 , n3772 , n3773 );
and ( n3775 , n2998 , n48 );
and ( n3776 , n3002 , n56 );
nor ( n3777 , n3775 , n3776 );
not ( n3778 , n3777 );
not ( n3779 , n3007 );
or ( n3780 , n3778 , n3779 );
or ( n3781 , n3012 , n231 );
nand ( n3782 , n3780 , n3781 );
nor ( n3783 , n3774 , n3782 );
and ( n3784 , n671 , n102 );
and ( n3785 , n673 , n110 );
nor ( n3786 , n3784 , n3785 );
and ( n3787 , n671 , n84 );
and ( n3788 , n673 , n92 );
nor ( n3789 , n3787 , n3788 );
not ( n3790 , n109 );
not ( n3791 , n668 );
or ( n3792 , n3790 , n3791 );
and ( n3793 , n1146 , n133 );
and ( n3794 , n673 , n117 );
nor ( n3795 , n3793 , n3794 );
nand ( n3796 , n3792 , n3795 );
not ( n3797 , n14 );
not ( n3798 , n673 );
or ( n3799 , n3797 , n3798 );
not ( n3800 , n22 );
or ( n3801 , n669 , n3800 );
nand ( n3802 , n3799 , n3801 );
not ( n3803 , n16 );
not ( n3804 , n673 );
or ( n3805 , n3803 , n3804 );
not ( n3806 , n668 );
not ( n3807 , n24 );
or ( n3808 , n3806 , n3807 );
nand ( n3809 , n3805 , n3808 );
not ( n3810 , n18 );
not ( n3811 , n673 );
or ( n3812 , n3810 , n3811 );
not ( n3813 , n26 );
or ( n3814 , n3806 , n3813 );
nand ( n3815 , n3812 , n3814 );
or ( n3816 , n3806 , n2369 );
or ( n3817 , n2373 , n199 );
nand ( n3818 , n3816 , n3817 );
not ( n3819 , n62 );
or ( n3820 , n669 , n3819 );
not ( n3821 , n54 );
or ( n3822 , n3821 , n199 );
nand ( n3823 , n3820 , n3822 );
or ( n3824 , n3806 , n1419 );
or ( n3825 , n2346 , n199 );
nand ( n3826 , n3824 , n3825 );
not ( n3827 , n71 );
not ( n3828 , n667 );
not ( n3829 , n3828 );
or ( n3830 , n3827 , n3829 );
and ( n3831 , n848 , n146 );
and ( n3832 , n673 , n79 );
nor ( n3833 , n3831 , n3832 );
nand ( n3834 , n3830 , n3833 );
not ( n3835 , n73 );
not ( n3836 , n3828 );
or ( n3837 , n3835 , n3836 );
and ( n3838 , n848 , n154 );
and ( n3839 , n673 , n81 );
nor ( n3840 , n3838 , n3839 );
nand ( n3841 , n3837 , n3840 );
not ( n3842 , n77 );
not ( n3843 , n3828 );
or ( n3844 , n3842 , n3843 );
and ( n3845 , n1146 , n137 );
and ( n3846 , n673 , n85 );
nor ( n3847 , n3845 , n3846 );
nand ( n3848 , n3844 , n3847 );
not ( n3849 , n87 );
not ( n3850 , n3828 );
or ( n3851 , n3849 , n3850 );
and ( n3852 , n848 , n144 );
and ( n3853 , n673 , n95 );
nor ( n3854 , n3852 , n3853 );
nand ( n3855 , n3851 , n3854 );
not ( n3856 , n89 );
not ( n3857 , n668 );
or ( n3858 , n3856 , n3857 );
and ( n3859 , n1146 , n152 );
and ( n3860 , n673 , n97 );
nor ( n3861 , n3859 , n3860 );
nand ( n3862 , n3858 , n3861 );
not ( n3863 , n93 );
not ( n3864 , n668 );
or ( n3865 , n3863 , n3864 );
and ( n3866 , n1146 , n135 );
and ( n3867 , n673 , n101 );
nor ( n3868 , n3866 , n3867 );
nand ( n3869 , n3865 , n3868 );
not ( n3870 , n95 );
not ( n3871 , n3828 );
or ( n3872 , n3870 , n3871 );
and ( n3873 , n848 , n143 );
and ( n3874 , n673 , n103 );
nor ( n3875 , n3873 , n3874 );
nand ( n3876 , n3872 , n3875 );
not ( n3877 , n99 );
not ( n3878 , n668 );
or ( n3879 , n3877 , n3878 );
and ( n3880 , n1146 , n159 );
and ( n3881 , n673 , n107 );
nor ( n3882 , n3880 , n3881 );
nand ( n3883 , n3879 , n3882 );
not ( n3884 , n105 );
not ( n3885 , n3828 );
or ( n3886 , n3884 , n3885 );
and ( n3887 , n1146 , n150 );
and ( n3888 , n673 , n113 );
nor ( n3889 , n3887 , n3888 );
nand ( n3890 , n3886 , n3889 );
not ( n3891 , n107 );
not ( n3892 , n668 );
or ( n3893 , n3891 , n3892 );
and ( n3894 , n848 , n158 );
and ( n3895 , n673 , n115 );
nor ( n3896 , n3894 , n3895 );
nand ( n3897 , n3893 , n3896 );
not ( n3898 , n111 );
not ( n3899 , n668 );
or ( n3900 , n3898 , n3899 );
and ( n3901 , n848 , n141 );
and ( n3902 , n673 , n119 );
nor ( n3903 , n3901 , n3902 );
nand ( n3904 , n3900 , n3903 );
not ( n3905 , n113 );
not ( n3906 , n3828 );
or ( n3907 , n3905 , n3906 );
and ( n3908 , n1146 , n149 );
and ( n3909 , n673 , n121 );
nor ( n3910 , n3908 , n3909 );
nand ( n3911 , n3907 , n3910 );
not ( n3912 , n115 );
not ( n3913 , n668 );
or ( n3914 , n3912 , n3913 );
and ( n3915 , n1429 , n157 );
and ( n3916 , n673 , n123 );
nor ( n3917 , n3915 , n3916 );
nand ( n3918 , n3914 , n3917 );
not ( n3919 , n117 );
not ( n3920 , n668 );
or ( n3921 , n3919 , n3920 );
and ( n3922 , n848 , n132 );
and ( n3923 , n673 , n125 );
nor ( n3924 , n3922 , n3923 );
nand ( n3925 , n3921 , n3924 );
not ( n3926 , n119 );
not ( n3927 , n668 );
or ( n3928 , n3926 , n3927 );
and ( n3929 , n848 , n140 );
and ( n3930 , n673 , n127 );
nor ( n3931 , n3929 , n3930 );
nand ( n3932 , n3928 , n3931 );
not ( n3933 , n121 );
not ( n3934 , n668 );
or ( n3935 , n3933 , n3934 );
and ( n3936 , n1146 , n148 );
and ( n3937 , n673 , n129 );
nor ( n3938 , n3936 , n3937 );
nand ( n3939 , n3935 , n3938 );
not ( n3940 , n123 );
not ( n3941 , n668 );
or ( n3942 , n3940 , n3941 );
and ( n3943 , n848 , n156 );
and ( n3944 , n673 , n131 );
nor ( n3945 , n3943 , n3944 );
nand ( n3946 , n3942 , n3945 );
not ( n3947 , n97 );
not ( n3948 , n3828 );
or ( n3949 , n3947 , n3948 );
and ( n3950 , n848 , n151 );
and ( n3951 , n673 , n105 );
nor ( n3952 , n3950 , n3951 );
nand ( n3953 , n3949 , n3952 );
buf ( n3954 , n667 );
or ( n3955 , n3954 , n2747 );
or ( n3956 , n1363 , n199 );
nand ( n3957 , n3955 , n3956 );
not ( n3958 , n20 );
not ( n3959 , n668 );
or ( n3960 , n3958 , n3959 );
nand ( n3961 , n673 , n12 );
nand ( n3962 , n3960 , n3961 );
or ( n3963 , n3954 , n2852 );
or ( n3964 , n2953 , n199 );
nand ( n3965 , n3963 , n3964 );
or ( n3966 , n3954 , n2856 );
or ( n3967 , n2788 , n199 );
nand ( n3968 , n3966 , n3967 );
not ( n3969 , n28 );
not ( n3970 , n3828 );
or ( n3971 , n3969 , n3970 );
nand ( n3972 , n673 , n20 );
nand ( n3973 , n3971 , n3972 );
or ( n3974 , n3954 , n2768 );
or ( n3975 , n2852 , n199 );
nand ( n3976 , n3974 , n3975 );
not ( n3977 , n30 );
or ( n3978 , n3954 , n3977 );
or ( n3979 , n3800 , n199 );
nand ( n3980 , n3978 , n3979 );
or ( n3981 , n3954 , n2341 );
or ( n3982 , n2856 , n199 );
nand ( n3983 , n3981 , n3982 );
buf ( n3984 , n667 );
not ( n3985 , n32 );
or ( n3986 , n3984 , n3985 );
or ( n3987 , n3807 , n199 );
nand ( n3988 , n3986 , n3987 );
or ( n3989 , n3954 , n2331 );
or ( n3990 , n2893 , n199 );
nand ( n3991 , n3989 , n3990 );
not ( n3992 , n34 );
or ( n3993 , n3954 , n3992 );
or ( n3994 , n3813 , n199 );
nand ( n3995 , n3993 , n3994 );
or ( n3996 , n3954 , n2373 );
or ( n3997 , n856 , n199 );
nand ( n3998 , n3996 , n3997 );
or ( n3999 , n3984 , n2336 );
or ( n4000 , n2341 , n199 );
nand ( n4001 , n3999 , n4000 );
not ( n4002 , n40 );
or ( n4003 , n3984 , n4002 );
or ( n4004 , n3985 , n199 );
nand ( n4005 , n4003 , n4004 );
or ( n4006 , n3984 , n2351 );
or ( n4007 , n2331 , n199 );
nand ( n4008 , n4006 , n4007 );
not ( n4009 , n42 );
or ( n4010 , n3954 , n4009 );
or ( n4011 , n3992 , n199 );
nand ( n4012 , n4010 , n4011 );
not ( n4013 , n44 );
not ( n4014 , n3828 );
or ( n4015 , n4013 , n4014 );
nand ( n4016 , n673 , n36 );
nand ( n4017 , n4015 , n4016 );
or ( n4018 , n3954 , n2356 );
or ( n4019 , n1357 , n199 );
nand ( n4020 , n4018 , n4019 );
not ( n4021 , n46 );
or ( n4022 , n3954 , n4021 );
not ( n4023 , n38 );
or ( n4024 , n4023 , n199 );
nand ( n4025 , n4022 , n4024 );
or ( n4026 , n3984 , n1431 );
or ( n4027 , n2336 , n199 );
nand ( n4028 , n4026 , n4027 );
not ( n4029 , n48 );
or ( n4030 , n3984 , n4029 );
or ( n4031 , n4002 , n199 );
nand ( n4032 , n4030 , n4031 );
or ( n4033 , n3954 , n1424 );
or ( n4034 , n2351 , n199 );
nand ( n4035 , n4033 , n4034 );
not ( n4036 , n50 );
or ( n4037 , n3954 , n4036 );
or ( n4038 , n4009 , n199 );
nand ( n4039 , n4037 , n4038 );
or ( n4040 , n3954 , n2760 );
or ( n4041 , n2369 , n199 );
nand ( n4042 , n4040 , n4041 );
not ( n4043 , n52 );
not ( n4044 , n3828 );
or ( n4045 , n4043 , n4044 );
nand ( n4046 , n673 , n44 );
nand ( n4047 , n4045 , n4046 );
or ( n4048 , n3954 , n2743 );
or ( n4049 , n2356 , n199 );
nand ( n4050 , n4048 , n4049 );
buf ( n4051 , n667 );
or ( n4052 , n4051 , n3821 );
or ( n4053 , n4021 , n199 );
nand ( n4054 , n4052 , n4053 );
or ( n4055 , n4051 , n2346 );
or ( n4056 , n1424 , n199 );
nand ( n4057 , n4055 , n4056 );
not ( n4058 , n58 );
or ( n4059 , n4051 , n4058 );
or ( n4060 , n4036 , n199 );
nand ( n4061 , n4059 , n4060 );
or ( n4062 , n4051 , n2365 );
or ( n4063 , n2760 , n199 );
nand ( n4064 , n4062 , n4063 );
not ( n4065 , n60 );
not ( n4066 , n668 );
or ( n4067 , n4065 , n4066 );
nand ( n4068 , n673 , n52 );
nand ( n4069 , n4067 , n4068 );
or ( n4070 , n4051 , n2738 );
or ( n4071 , n2743 , n199 );
nand ( n4072 , n4070 , n4071 );
or ( n4073 , n3984 , n1363 );
or ( n4074 , n1414 , n199 );
nand ( n4075 , n4073 , n4074 );
not ( n4076 , n64 );
or ( n4077 , n4051 , n4076 );
not ( n4078 , n56 );
or ( n4079 , n4078 , n199 );
nand ( n4080 , n4077 , n4079 );
or ( n4081 , n3984 , n2361 );
or ( n4082 , n2365 , n199 );
nand ( n4083 , n4081 , n4082 );
not ( n4084 , n1 );
not ( n4085 , n3828 );
or ( n4086 , n4084 , n4085 );
nand ( n4087 , n673 , n60 );
nand ( n4088 , n4086 , n4087 );
or ( n4089 , n4051 , n850 );
or ( n4090 , n2738 , n199 );
nand ( n4091 , n4089 , n4090 );
not ( n4092 , n3 );
not ( n4093 , n3828 );
or ( n4094 , n4092 , n4093 );
nand ( n4095 , n673 , n62 );
nand ( n4096 , n4094 , n4095 );
not ( n4097 , n5 );
not ( n4098 , n668 );
or ( n4099 , n4097 , n4098 );
nand ( n4100 , n673 , n64 );
nand ( n4101 , n4099 , n4100 );
or ( n4102 , n4051 , n2752 );
or ( n4103 , n1419 , n199 );
nand ( n4104 , n4102 , n4103 );
not ( n4105 , n7 );
not ( n4106 , n668 );
or ( n4107 , n4105 , n4106 );
nand ( n4108 , n673 , n66 );
nand ( n4109 , n4107 , n4108 );
or ( n4110 , n4051 , n2957 );
or ( n4111 , n2361 , n199 );
nand ( n4112 , n4110 , n4111 );
not ( n4113 , n69 );
not ( n4114 , n3828 );
or ( n4115 , n4113 , n4114 );
and ( n4116 , n1146 , n138 );
and ( n4117 , n673 , n77 );
nor ( n4118 , n4116 , n4117 );
nand ( n4119 , n4115 , n4118 );
not ( n4120 , n75 );
not ( n4121 , n668 );
or ( n4122 , n4120 , n4121 );
and ( n4123 , n1146 , n162 );
and ( n4124 , n673 , n83 );
nor ( n4125 , n4123 , n4124 );
nand ( n4126 , n4122 , n4125 );
not ( n4127 , n79 );
not ( n4128 , n3828 );
or ( n4129 , n4127 , n4128 );
and ( n4130 , n1146 , n145 );
and ( n4131 , n673 , n87 );
nor ( n4132 , n4130 , n4131 );
nand ( n4133 , n4129 , n4132 );
not ( n4134 , n81 );
not ( n4135 , n668 );
or ( n4136 , n4134 , n4135 );
and ( n4137 , n1146 , n153 );
and ( n4138 , n673 , n89 );
nor ( n4139 , n4137 , n4138 );
nand ( n4140 , n4136 , n4139 );
not ( n4141 , n83 );
not ( n4142 , n668 );
or ( n4143 , n4141 , n4142 );
and ( n4144 , n1035 , n161 );
and ( n4145 , n673 , n91 );
nor ( n4146 , n4144 , n4145 );
nand ( n4147 , n4143 , n4146 );
not ( n4148 , n85 );
not ( n4149 , n668 );
or ( n4150 , n4148 , n4149 );
and ( n4151 , n1146 , n136 );
and ( n4152 , n673 , n93 );
nor ( n4153 , n4151 , n4152 );
nand ( n4154 , n4150 , n4153 );
or ( n4155 , n4051 , n4078 );
or ( n4156 , n4029 , n199 );
nand ( n4157 , n4155 , n4156 );
not ( n4158 , n101 );
not ( n4159 , n668 );
or ( n4160 , n4158 , n4159 );
and ( n4161 , n1146 , n134 );
and ( n4162 , n673 , n109 );
nor ( n4163 , n4161 , n4162 );
nand ( n4164 , n4160 , n4163 );
not ( n4165 , n103 );
not ( n4166 , n3828 );
or ( n4167 , n4165 , n4166 );
and ( n4168 , n1146 , n142 );
and ( n4169 , n673 , n111 );
nor ( n4170 , n4168 , n4169 );
nand ( n4171 , n4167 , n4170 );
not ( n4172 , n36 );
not ( n4173 , n668 );
or ( n4174 , n4172 , n4173 );
nand ( n4175 , n673 , n28 );
nand ( n4176 , n4174 , n4175 );
or ( n4177 , n4051 , n1357 );
or ( n4178 , n2768 , n199 );
nand ( n4179 , n4177 , n4178 );
or ( n4180 , n4051 , n4023 );
or ( n4181 , n3977 , n199 );
nand ( n4182 , n4180 , n4181 );
or ( n4183 , n4051 , n856 );
or ( n4184 , n2764 , n199 );
nand ( n4185 , n4183 , n4184 );
or ( n4186 , n4051 , n2893 );
or ( n4187 , n2756 , n199 );
nand ( n4188 , n4186 , n4187 );
not ( n4189 , n91 );
not ( n4190 , n668 );
or ( n4191 , n4189 , n4190 );
and ( n4192 , n1146 , n160 );
and ( n4193 , n673 , n99 );
nor ( n4194 , n4192 , n4193 );
nand ( n4195 , n4191 , n4194 );
or ( n4196 , n4051 , n1414 );
or ( n4197 , n1431 , n199 );
nand ( n4198 , n4196 , n4197 );
not ( n4199 , n66 );
or ( n4200 , n4051 , n4199 );
or ( n4201 , n4058 , n199 );
nand ( n4202 , n4200 , n4201 );
not ( n4203 , n10 );
not ( n4204 , n1035 );
or ( n4205 , n4203 , n4204 );
or ( n4206 , n2339 , n2962 );
nand ( n4207 , n4205 , n4206 );
not ( n4208 , n1 );
not ( n4209 , n1035 );
or ( n4210 , n4208 , n4209 );
not ( n4211 , n132 );
or ( n4212 , n838 , n4211 );
nand ( n4213 , n4210 , n4212 );
not ( n4214 , n28 );
not ( n4215 , n1429 );
or ( n4216 , n4214 , n4215 );
nand ( n4217 , n845 , n137 );
nand ( n4218 , n4216 , n4217 );
not ( n4219 , n20 );
not ( n4220 , n1429 );
or ( n4221 , n4219 , n4220 );
nand ( n4222 , n845 , n138 );
nand ( n4223 , n4221 , n4222 );
not ( n4224 , n16 );
not ( n4225 , n1146 );
or ( n4226 , n4224 , n4225 );
not ( n4227 , n663 );
not ( n4228 , n155 );
or ( n4229 , n4227 , n4228 );
nand ( n4230 , n4226 , n4229 );
not ( n4231 , n7 );
not ( n4232 , n1035 );
or ( n4233 , n4231 , n4232 );
not ( n4234 , n156 );
or ( n4235 , n838 , n4234 );
nand ( n4236 , n4233 , n4235 );
not ( n4237 , n18 );
not ( n4238 , n1035 );
or ( n4239 , n4237 , n4238 );
not ( n4240 , n163 );
or ( n4241 , n4227 , n4240 );
nand ( n4242 , n4239 , n4241 );
and ( n4243 , n1035 , n147 );
and ( n4244 , n673 , n71 );
nor ( n4245 , n4243 , n4244 );
not ( n4246 , n4245 );
and ( n4247 , n1035 , n155 );
and ( n4248 , n673 , n73 );
nor ( n4249 , n4247 , n4248 );
not ( n4250 , n4249 );
and ( n4251 , n1429 , n163 );
and ( n4252 , n673 , n75 );
nor ( n4253 , n4251 , n4252 );
not ( n4254 , n4253 );
and ( n4255 , n1429 , n139 );
and ( n4256 , n673 , n69 );
nor ( n4257 , n4255 , n4256 );
not ( n4258 , n4257 );
not ( n4259 , n3 );
not ( n4260 , n1035 );
or ( n4261 , n4259 , n4260 );
not ( n4262 , n140 );
or ( n4263 , n4227 , n4262 );
nand ( n4264 , n4261 , n4263 );
not ( n4265 , n14 );
not ( n4266 , n1146 );
or ( n4267 , n4265 , n4266 );
not ( n4268 , n147 );
or ( n4269 , n2339 , n4268 );
nand ( n4270 , n4267 , n4269 );
not ( n4271 , n60 );
not ( n4272 , n1146 );
or ( n4273 , n4271 , n4272 );
nand ( n4274 , n855 , n133 );
nand ( n4275 , n4273 , n4274 );
not ( n4276 , n36 );
not ( n4277 , n1035 );
or ( n4278 , n4276 , n4277 );
not ( n4279 , n136 );
or ( n4280 , n2339 , n4279 );
nand ( n4281 , n4278 , n4280 );
not ( n4282 , n52 );
not ( n4283 , n1146 );
or ( n4284 , n4282 , n4283 );
nand ( n4285 , n855 , n134 );
nand ( n4286 , n4284 , n4285 );
not ( n4287 , n44 );
not ( n4288 , n1035 );
or ( n4289 , n4287 , n4288 );
not ( n4290 , n135 );
or ( n4291 , n4227 , n4290 );
nand ( n4292 , n4289 , n4291 );
not ( n4293 , n146 );
not ( n4294 , n663 );
or ( n4295 , n4293 , n4294 );
or ( n4296 , n855 , n3800 );
nand ( n4297 , n4295 , n4296 );
not ( n4298 , n1429 );
not ( n4299 , n4298 );
not ( n4300 , n149 );
or ( n4301 , n4299 , n4300 );
not ( n4302 , n1035 );
or ( n4303 , n4302 , n4076 );
nand ( n4304 , n4301 , n4303 );
not ( n4305 , n153 );
not ( n4306 , n848 );
not ( n4307 , n4306 );
or ( n4308 , n4305 , n4307 );
or ( n4309 , n1362 , n3985 );
nand ( n4310 , n4308 , n4309 );
not ( n4311 , n4298 );
not ( n4312 , n158 );
or ( n4313 , n4311 , n4312 );
or ( n4314 , n1362 , n4058 );
nand ( n4315 , n4313 , n4314 );
not ( n4316 , n160 );
not ( n4317 , n855 );
or ( n4318 , n4316 , n4317 );
or ( n4319 , n4306 , n4009 );
nand ( n4320 , n4318 , n4319 );
not ( n4321 , n144 );
not ( n4322 , n845 );
or ( n4323 , n4321 , n4322 );
or ( n4324 , n4302 , n4023 );
nand ( n4325 , n4323 , n4324 );
not ( n4326 , n141 );
not ( n4327 , n4298 );
or ( n4328 , n4326 , n4327 );
or ( n4329 , n4306 , n3819 );
nand ( n4330 , n4328 , n4329 );
not ( n4331 , n162 );
not ( n4332 , n855 );
or ( n4333 , n4331 , n4332 );
or ( n4334 , n1362 , n3813 );
nand ( n4335 , n4333 , n4334 );
not ( n4336 , n157 );
not ( n4337 , n855 );
or ( n4338 , n4336 , n4337 );
or ( n4339 , n1362 , n4199 );
nand ( n4340 , n4338 , n4339 );
not ( n4341 , n142 );
not ( n4342 , n4306 );
or ( n4343 , n4341 , n4342 );
or ( n4344 , n4302 , n3821 );
nand ( n4345 , n4343 , n4344 );
not ( n4346 , n143 );
not ( n4347 , n855 );
or ( n4348 , n4346 , n4347 );
or ( n4349 , n1418 , n4021 );
nand ( n4350 , n4348 , n4349 );
not ( n4351 , n154 );
not ( n4352 , n855 );
or ( n4353 , n4351 , n4352 );
or ( n4354 , n1362 , n3807 );
nand ( n4355 , n4353 , n4354 );
not ( n4356 , n4298 );
not ( n4357 , n161 );
or ( n4358 , n4356 , n4357 );
or ( n4359 , n1418 , n3992 );
nand ( n4360 , n4358 , n4359 );
not ( n4361 , n159 );
not ( n4362 , n4306 );
or ( n4363 , n4361 , n4362 );
or ( n4364 , n4306 , n4036 );
nand ( n4365 , n4363 , n4364 );
not ( n4366 , n151 );
not ( n4367 , n855 );
or ( n4368 , n4366 , n4367 );
or ( n4369 , n855 , n4029 );
nand ( n4370 , n4368 , n4369 );
not ( n4371 , n150 );
not ( n4372 , n4306 );
or ( n4373 , n4371 , n4372 );
or ( n4374 , n4302 , n4078 );
nand ( n4375 , n4373 , n4374 );
not ( n4376 , n152 );
not ( n4377 , n855 );
or ( n4378 , n4376 , n4377 );
or ( n4379 , n1362 , n4002 );
nand ( n4380 , n4378 , n4379 );
not ( n4381 , n145 );
not ( n4382 , n855 );
or ( n4383 , n4381 , n4382 );
or ( n4384 , n4306 , n3977 );
nand ( n4385 , n4383 , n4384 );
not ( n4386 , n12 );
not ( n4387 , n1035 );
or ( n4388 , n4386 , n4387 );
not ( n4389 , n139 );
or ( n4390 , n2339 , n4389 );
nand ( n4391 , n4388 , n4390 );
not ( n4392 , n5 );
not ( n4393 , n1035 );
or ( n4394 , n4392 , n4393 );
not ( n4395 , n148 );
or ( n4396 , n2339 , n4395 );
nand ( n4397 , n4394 , n4396 );
not ( n4398 , n2972 );
nor ( n4399 , n1146 , n4398 , n9 );
nand ( n4400 , n198 , n199 );
and ( n4401 , n4400 , n2979 );
not ( n4402 , n2971 );
nor ( n4403 , n4401 , n4402 , n9 );
not ( n4404 , n4400 );
nor ( n4405 , n4404 , n2977 , n9 );
nor ( n4406 , n9 , n199 );
not ( n4407 , n1354 );
not ( n4408 , n1146 );
or ( n4409 , n4407 , n4408 );
nand ( n4410 , n4409 , n3789 );
not ( n4411 , n1410 );
not ( n4412 , n2339 );
or ( n4413 , n4411 , n4412 );
nand ( n4414 , n4413 , n3786 );
endmodule
