module top ( g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 , g98 , g99 , g100 , g101 , g102 , g103 , g104 , g105 , g106 , g107 , g108 , g109 , g110 , g111 , g112 , g113 , g114 , g115 , g116 , g117 , g118 , g119 , g120 , g121 , g122 , g123 , g124 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g136 , g137 , g138 , g139 , g140 , g141 , g142 , g143 , g144 , g145 , g146 , g147 , g148 , g149 , g150 , g151 , g152 , g153 , g154 , g155 , g156 , g157 , g158 , g159 , g160 );
input g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 ;
output g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 , g98 , g99 , g100 , g101 , g102 , g103 , g104 , g105 , g106 , g107 , g108 , g109 , g110 , g111 , g112 , g113 , g114 , g115 , g116 , g117 , g118 , g119 , g120 , g121 , g122 , g123 , g124 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g136 , g137 , g138 , g139 , g140 , g141 , g142 , g143 , g144 , g145 , g146 , g147 , g148 , g149 , g150 , g151 , g152 , g153 , g154 , g155 , g156 , g157 , g158 , g159 , g160 ;

wire n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , 
     n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , 
     n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , 
     n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , 
     n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , 
     n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , 
     n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , 
     n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , 
     n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , 
     n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , 
     n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , 
     n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , 
     n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , 
     n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , 
     n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , 
     n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , 
     n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , 
     n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , 
     n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , 
     n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , 
     n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , 
     n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , 
     n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , 
     n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , 
     n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , 
     n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , 
     n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , 
     n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , 
     n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , 
     n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , 
     n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , 
     n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , 
     n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , 
     n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , 
     n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , 
     n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , 
     n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , 
     n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , 
     n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , 
     n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , 
     n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , 
     n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , 
     n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , 
     n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , 
     n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , 
     n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , 
     n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , 
     n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , 
     n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , 
     n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , 
     n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , 
     n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , 
     n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , 
     n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , 
     n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , 
     n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , 
     n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , 
     n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , 
     n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , 
     n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , 
     n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , 
     n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , 
     n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , 
     n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , 
     n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , 
     n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , 
     n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , 
     n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , 
     n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , 
     n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , 
     n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , 
     n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , 
     n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , 
     n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , 
     n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , 
     n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , 
     n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , 
     n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , 
     n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , 
     n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , 
     n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , 
     n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , 
     n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , 
     n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , 
     n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , 
     n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , 
     n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , 
     n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , 
     n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , 
     n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , 
     n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , 
     n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , 
     n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , 
     n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , 
     n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , 
     n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , 
     n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , 
     n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , 
     n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , 
     n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , 
     n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , 
     n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , 
     n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , 
     n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , 
     n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , 
     n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , 
     n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , 
     n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , 
     n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , 
     n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , 
     n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , 
     n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , 
     n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , 
     n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , 
     n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , 
     n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , 
     n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , 
     n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , 
     n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , 
     n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , 
     n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , 
     n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , 
     n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , 
     n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , 
     n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , 
     n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , 
     n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , 
     n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , 
     n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , 
     n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , 
     n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , 
     n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , 
     n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , 
     n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , 
     n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , 
     n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , 
     n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , 
     n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , 
     n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , 
     n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , 
     n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , 
     n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , 
     n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , 
     n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , 
     n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , 
     n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , 
     n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , 
     n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , 
     n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , 
     n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , 
     n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , 
     n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , 
     n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , 
     n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , 
     n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , 
     n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , g349 , 
     g350 , g351 , g352 , g353 , g354 , g355 , g356 , g357 ;
wire t_0 , t_1 ;
buf ( g349  , g0 );
buf ( g350  , g1 );
buf ( g351  , g2 );
buf ( g352  , g3 );
buf ( g353  , g4 );
buf ( g354  , g5 );
buf ( g355  , g6 );
buf ( g356  , g7 );
buf ( g357  , g8 );
buf ( n28  , g9 );
buf ( n29  , g10 );
buf ( n30  , g11 );
buf ( n31  , g12 );
buf ( n32  , g13 );
buf ( n33  , g14 );
buf ( n34  , g15 );
buf ( n35  , g16 );
buf ( n36  , g17 );
buf ( n37  , g18 );
buf ( n38  , g19 );
buf ( n39  , g20 );
buf ( n40  , g21 );
buf ( n41  , g22 );
buf ( n42  , g23 );
buf ( n43  , g24 );
buf ( n44  , g25 );
buf ( n45  , g26 );
buf ( n46  , g27 );
buf ( n47  , g28 );
buf ( n48  , g29 );
buf ( n49  , g30 );
buf ( n50  , g31 );
buf ( g32 , n51  );
buf ( g33 , n52  );
buf ( g34 , n53  );
buf ( g35 , n54  );
buf ( g36 , n55  );
buf ( g37 , n56  );
buf ( g38 , n57  );
buf ( g39 , n58  );
buf ( g40 , n59  );
buf ( g41 , n60  );
buf ( g42 , n61  );
buf ( g43 , n62  );
buf ( g44 , n63  );
buf ( g45 , n64  );
buf ( g46 , n65  );
buf ( g47 , n66  );
buf ( g48 , n67  );
buf ( g49 , n68  );
buf ( g50 , n69  );
buf ( g51 , n70  );
buf ( g52 , n71  );
buf ( g53 , n72  );
buf ( g54 , n73  );
buf ( g55 , n74  );
buf ( g56 , n75  );
buf ( g57 , n76  );
buf ( g58 , n77  );
buf ( g59 , n78  );
buf ( g60 , n79  );
buf ( g61 , n80  );
buf ( g62 , n81  );
buf ( g63 , n82  );
buf ( g64 , n83  );
buf ( g65 , n84  );
buf ( g66 , n85  );
buf ( g67 , n86  );
buf ( g68 , n87  );
buf ( g69 , n88  );
buf ( g70 , n89  );
buf ( g71 , n90  );
buf ( g72 , n91  );
buf ( g73 , n92  );
buf ( g74 , n93  );
buf ( g75 , n94  );
buf ( g76 , n95  );
buf ( g77 , n96  );
buf ( g78 , n97  );
buf ( g79 , n98  );
buf ( g80 , n99  );
buf ( g81 , n100  );
buf ( g82 , n101  );
buf ( g83 , n102  );
buf ( g84 , n103  );
buf ( g85 , n104  );
buf ( g86 , n105  );
buf ( g87 , n106  );
buf ( g88 , n107  );
buf ( g89 , n108  );
buf ( g90 , n109  );
buf ( g91 , n110  );
buf ( g92 , n111  );
buf ( g93 , n112  );
buf ( g94 , n113  );
buf ( g95 , n114  );
buf ( g96 , n115  );
buf ( g97 , n116  );
buf ( g98 , n117  );
buf ( g99 , n118  );
buf ( g100 , n119  );
buf ( g101 , n120  );
buf ( g102 , n121  );
buf ( g103 , n122  );
buf ( g104 , n123  );
buf ( g105 , n124  );
buf ( g106 , n125  );
buf ( g107 , n126  );
buf ( g108 , n127  );
buf ( g109 , n128  );
buf ( g110 , n129  );
buf ( g111 , n130  );
buf ( g112 , n131  );
buf ( g113 , n132  );
buf ( g114 , n133  );
buf ( g115 , n134  );
buf ( g116 , n135  );
buf ( g117 , n136  );
buf ( g118 , n137  );
buf ( g119 , n138  );
buf ( g120 , n139  );
buf ( g121 , n140  );
buf ( g122 , n141  );
buf ( g123 , n142  );
buf ( g124 , n143  );
buf ( g125 , n144  );
buf ( g126 , n145  );
buf ( g127 , n146  );
buf ( g128 , n147  );
buf ( g129 , n148  );
buf ( g130 , n149  );
buf ( g131 , n150  );
buf ( g132 , n151  );
buf ( g133 , n152  );
buf ( g134 , n153  );
buf ( g135 , n154  );
buf ( g136 , n155  );
buf ( g137 , n156  );
buf ( g138 , n157  );
buf ( g139 , n158  );
buf ( g140 , n159  );
buf ( g141 , n160  );
buf ( g142 , n161  );
buf ( g143 , n162  );
buf ( g144 , n163  );
buf ( g145 , n164  );
buf ( g146 , n165  );
buf ( g147 , n166  );
buf ( g148 , n167  );
buf ( g149 , n168  );
buf ( g150 , n169  );
buf ( g151 , n170  );
buf ( g152 , n171  );
buf ( g153 , n172  );
buf ( g154 , n173  );
buf ( g155 , n174  );
buf ( g156 , n175  );
buf ( g157 , n176  );
buf ( g158 , n177  );
buf ( g159 , n178  );
buf ( g160 , n179  );
buf ( n51 , 1'b0 );
buf ( n52 , 1'b0 );
buf ( n53 , 1'b0 );
buf ( n54 , 1'b0 );
buf ( n55 , 1'b0 );
buf ( n56 , 1'b0 );
buf ( n57 , 1'b0 );
buf ( n58 , 1'b0 );
buf ( n59 , 1'b0 );
buf ( n60 , 1'b0 );
buf ( n61 , 1'b0 );
buf ( n62 , 1'b0 );
buf ( n63 , 1'b0 );
buf ( n64 , 1'b0 );
buf ( n65 , 1'b0 );
buf ( n66 , 1'b0 );
buf ( n67 , 1'b0 );
buf ( n68 , 1'b0 );
buf ( n69 , 1'b0 );
buf ( n70 , 1'b0 );
buf ( n71 , 1'b0 );
buf ( n72 , 1'b0 );
buf ( n73 , 1'b0 );
buf ( n74 , 1'b0 );
buf ( n75 , 1'b0 );
buf ( n76 , 1'b0 );
buf ( n77 , 1'b0 );
buf ( n78 , 1'b0 );
buf ( n79 , 1'b0 );
buf ( n80 , 1'b0 );
buf ( n81 , 1'b0 );
buf ( n82 , 1'b0 );
buf ( n83 , 1'b0 );
buf ( n84 , 1'b0 );
buf ( n85 , 1'b0 );
buf ( n86 , 1'b0 );
buf ( n87 , 1'b0 );
buf ( n88 , 1'b0 );
buf ( n89 , 1'b0 );
buf ( n90 , 1'b0 );
buf ( n91 , 1'b0 );
buf ( n92 , 1'b0 );
buf ( n93 , 1'b0 );
buf ( n94 , 1'b0 );
buf ( n95 , 1'b0 );
buf ( n96 , 1'b0 );
buf ( n97 , 1'b0 );
buf ( n98 , 1'b0 );
buf ( n99 , n1518 );
buf ( n100 , n1520 );
buf ( n101 , n1522 );
buf ( n102 , n1524 );
buf ( n103 , n1526 );
buf ( n104 , n1528 );
buf ( n105 , n1530 );
buf ( n106 , n1532 );
buf ( n107 , n1535 );
buf ( n108 , n1538 );
buf ( n109 , n1541 );
buf ( n110 , n1544 );
buf ( n111 , n1547 );
buf ( n112 , n1550 );
buf ( n113 , n1553 );
buf ( n114 , n1556 );
buf ( n115 , n1558 );
buf ( n116 , 1'b0 );
buf ( n117 , 1'b0 );
buf ( n118 , 1'b0 );
buf ( n119 , 1'b0 );
buf ( n120 , 1'b0 );
buf ( n121 , 1'b0 );
buf ( n122 , 1'b0 );
buf ( n123 , 1'b0 );
buf ( n124 , 1'b0 );
buf ( n125 , 1'b0 );
buf ( n126 , 1'b0 );
buf ( n127 , 1'b0 );
buf ( n128 , 1'b0 );
buf ( n129 , 1'b0 );
buf ( n130 , 1'b0 );
buf ( n131 , 1'b0 );
buf ( n132 , 1'b0 );
buf ( n133 , 1'b0 );
buf ( n134 , 1'b0 );
buf ( n135 , 1'b0 );
buf ( n136 , 1'b0 );
buf ( n137 , 1'b0 );
buf ( n138 , 1'b0 );
buf ( n139 , 1'b0 );
buf ( n140 , 1'b0 );
buf ( n141 , 1'b0 );
buf ( n142 , 1'b0 );
buf ( n143 , 1'b0 );
buf ( n144 , 1'b0 );
buf ( n145 , 1'b0 );
buf ( n146 , 1'b0 );
buf ( n147 , 1'b0 );
buf ( n148 , 1'b0 );
buf ( n149 , 1'b0 );
buf ( n150 , 1'b0 );
buf ( n151 , 1'b0 );
buf ( n152 , 1'b0 );
buf ( n153 , 1'b0 );
buf ( n154 , 1'b0 );
buf ( n155 , 1'b0 );
buf ( n156 , 1'b0 );
buf ( n157 , 1'b0 );
buf ( n158 , 1'b0 );
buf ( n159 , 1'b0 );
buf ( n160 , 1'b0 );
buf ( n161 , 1'b0 );
buf ( n162 , 1'b0 );
buf ( n163 , n1413 );
buf ( n164 , n1415 );
buf ( n165 , n1417 );
buf ( n166 , n1419 );
buf ( n167 , n1421 );
buf ( n168 , n1423 );
buf ( n169 , n1425 );
buf ( n170 , n1427 );
buf ( n171 , n1430 );
buf ( n172 , n1433 );
buf ( n173 , n1436 );
buf ( n174 , n1439 );
buf ( n175 , n1442 );
buf ( n176 , n1445 );
buf ( n177 , n1448 );
buf ( n178 , n1451 );
buf ( n179 , n1453 );
buf ( n298 , n42 );
buf ( n299 , n50 );
xor ( n300 , n298 , n299 );
buf ( n301 , n300 );
buf ( n302 , g356 );
buf ( n303 , n34 );
xor ( n304 , n302 , n303 );
buf ( n305 , n304 );
buf ( n306 , g356 );
buf ( n307 , n36 );
and ( n308 , n306 , n307 );
buf ( n309 , g355 );
buf ( n310 , n37 );
and ( n311 , n309 , n310 );
and ( n312 , n308 , n311 );
buf ( n313 , g354 );
buf ( n314 , n38 );
and ( n315 , n313 , n314 );
and ( n316 , n311 , n315 );
and ( n317 , n308 , n315 );
or ( n318 , n312 , n316 , n317 );
buf ( n319 , n40 );
and ( n320 , n313 , n319 );
buf ( n321 , g353 );
buf ( n322 , n41 );
and ( n323 , n321 , n322 );
and ( n324 , n320 , n323 );
buf ( n325 , g352 );
buf ( n326 , n42 );
and ( n327 , n325 , n326 );
and ( n328 , n323 , n327 );
and ( n329 , n320 , n327 );
or ( n330 , n324 , n328 , n329 );
and ( n331 , n321 , n319 );
and ( n332 , n330 , n331 );
and ( n333 , n325 , n322 );
buf ( n334 , g351 );
and ( n335 , n334 , n326 );
xor ( n336 , n333 , n335 );
and ( n337 , n331 , n336 );
and ( n338 , n330 , n336 );
or ( n339 , n332 , n337 , n338 );
xor ( n340 , n308 , n311 );
xor ( n341 , n340 , n315 );
and ( n342 , n339 , n341 );
and ( n343 , n333 , n335 );
buf ( n344 , n39 );
and ( n345 , n321 , n344 );
xor ( n346 , n343 , n345 );
and ( n347 , n325 , n319 );
and ( n348 , n334 , n322 );
xor ( n349 , n347 , n348 );
buf ( n350 , g350 );
and ( n351 , n350 , n326 );
xor ( n352 , n349 , n351 );
xor ( n353 , n346 , n352 );
and ( n354 , n341 , n353 );
and ( n355 , n339 , n353 );
or ( n356 , n342 , n354 , n355 );
xor ( n357 , n318 , n356 );
and ( n358 , n343 , n345 );
and ( n359 , n345 , n352 );
and ( n360 , n343 , n352 );
or ( n361 , n358 , n359 , n360 );
and ( n362 , n347 , n348 );
and ( n363 , n348 , n351 );
and ( n364 , n347 , n351 );
or ( n365 , n362 , n363 , n364 );
and ( n366 , n309 , n307 );
and ( n367 , n313 , n310 );
xor ( n368 , n366 , n367 );
and ( n369 , n321 , n314 );
xor ( n370 , n368 , n369 );
xor ( n371 , n365 , n370 );
and ( n372 , n325 , n344 );
and ( n373 , n334 , n319 );
xor ( n374 , n372 , n373 );
and ( n375 , n350 , n322 );
xor ( n376 , n374 , n375 );
xor ( n377 , n371 , n376 );
xor ( n378 , n361 , n377 );
not ( n379 , n306 );
buf ( n380 , n35 );
not ( n381 , n380 );
and ( n382 , n381 , n306 );
nor ( n383 , n379 , n382 );
buf ( n384 , g349 );
not ( n385 , n384 );
and ( n386 , n385 , n326 );
not ( n387 , n326 );
nor ( n388 , n386 , n387 );
xor ( n389 , n383 , n388 );
xor ( n390 , n378 , n389 );
xor ( n391 , n357 , n390 );
and ( n392 , n309 , n314 );
and ( n393 , n313 , n344 );
and ( n394 , n392 , n393 );
and ( n395 , n309 , n319 );
and ( n396 , n313 , n322 );
and ( n397 , n395 , n396 );
and ( n398 , n321 , n326 );
and ( n399 , n396 , n398 );
and ( n400 , n395 , n398 );
or ( n401 , n397 , n399 , n400 );
and ( n402 , n309 , n344 );
and ( n403 , n401 , n402 );
xor ( n404 , n320 , n323 );
xor ( n405 , n404 , n327 );
and ( n406 , n402 , n405 );
and ( n407 , n401 , n405 );
or ( n408 , n403 , n406 , n407 );
xor ( n409 , n392 , n393 );
and ( n410 , n408 , n409 );
xor ( n411 , n330 , n331 );
xor ( n412 , n411 , n336 );
and ( n413 , n409 , n412 );
and ( n414 , n408 , n412 );
or ( n415 , n410 , n413 , n414 );
and ( n416 , n394 , n415 );
xor ( n417 , n339 , n341 );
xor ( n418 , n417 , n353 );
and ( n419 , n415 , n418 );
and ( n420 , n394 , n418 );
or ( n421 , n416 , n419 , n420 );
xor ( n422 , n391 , n421 );
xor ( n423 , n394 , n415 );
xor ( n424 , n423 , n418 );
and ( n425 , n306 , n319 );
and ( n426 , n309 , n322 );
and ( n427 , n425 , n426 );
and ( n428 , n313 , n326 );
and ( n429 , n426 , n428 );
and ( n430 , n425 , n428 );
or ( n431 , n427 , n429 , n430 );
and ( n432 , n306 , n344 );
and ( n433 , n431 , n432 );
xor ( n434 , n395 , n396 );
xor ( n435 , n434 , n398 );
and ( n436 , n432 , n435 );
and ( n437 , n431 , n435 );
or ( n438 , n433 , n436 , n437 );
and ( n439 , n306 , n314 );
and ( n440 , n438 , n439 );
xor ( n441 , n401 , n402 );
xor ( n442 , n441 , n405 );
and ( n443 , n439 , n442 );
and ( n444 , n438 , n442 );
or ( n445 , n440 , n443 , n444 );
xor ( n446 , n408 , n409 );
xor ( n447 , n446 , n412 );
and ( n448 , n445 , n447 );
and ( n449 , n424 , n448 );
xor ( n450 , n424 , n448 );
and ( n451 , n306 , n310 );
xor ( n452 , n445 , n447 );
and ( n453 , n451 , n452 );
xor ( n454 , n451 , n452 );
xor ( n455 , n438 , n439 );
xor ( n456 , n455 , n442 );
xor ( n457 , n431 , n432 );
xor ( n458 , n457 , n435 );
xor ( n459 , n425 , n426 );
xor ( n460 , n459 , n428 );
and ( n461 , n306 , n322 );
and ( n462 , n309 , n326 );
and ( n463 , n461 , n462 );
and ( n464 , n460 , n463 );
and ( n465 , n458 , n464 );
and ( n466 , n456 , n465 );
and ( n467 , n454 , n466 );
or ( n468 , n453 , n467 );
and ( n469 , n450 , n468 );
or ( n470 , n449 , n469 );
buf ( n471 , n34 );
buf ( n472 , n44 );
and ( n473 , n471 , n472 );
buf ( n474 , n33 );
buf ( n475 , n45 );
and ( n476 , n474 , n475 );
and ( n477 , n473 , n476 );
buf ( n478 , n32 );
buf ( n479 , n46 );
and ( n480 , n478 , n479 );
and ( n481 , n476 , n480 );
and ( n482 , n473 , n480 );
or ( n483 , n477 , n481 , n482 );
buf ( n484 , n48 );
and ( n485 , n478 , n484 );
buf ( n486 , n31 );
buf ( n487 , n49 );
and ( n488 , n486 , n487 );
and ( n489 , n485 , n488 );
buf ( n490 , n30 );
buf ( n491 , n50 );
and ( n492 , n490 , n491 );
and ( n493 , n488 , n492 );
and ( n494 , n485 , n492 );
or ( n495 , n489 , n493 , n494 );
and ( n496 , n486 , n484 );
and ( n497 , n495 , n496 );
and ( n498 , n490 , n487 );
buf ( n499 , n29 );
and ( n500 , n499 , n491 );
xor ( n501 , n498 , n500 );
and ( n502 , n496 , n501 );
and ( n503 , n495 , n501 );
or ( n504 , n497 , n502 , n503 );
xor ( n505 , n473 , n476 );
xor ( n506 , n505 , n480 );
and ( n507 , n504 , n506 );
and ( n508 , n498 , n500 );
buf ( n509 , n47 );
and ( n510 , n486 , n509 );
xor ( n511 , n508 , n510 );
and ( n512 , n490 , n484 );
and ( n513 , n499 , n487 );
xor ( n514 , n512 , n513 );
buf ( n515 , n28 );
and ( n516 , n515 , n491 );
xor ( n517 , n514 , n516 );
xor ( n518 , n511 , n517 );
and ( n519 , n506 , n518 );
and ( n520 , n504 , n518 );
or ( n521 , n507 , n519 , n520 );
xor ( n522 , n483 , n521 );
and ( n523 , n508 , n510 );
and ( n524 , n510 , n517 );
and ( n525 , n508 , n517 );
or ( n526 , n523 , n524 , n525 );
and ( n527 , n512 , n513 );
and ( n528 , n513 , n516 );
and ( n529 , n512 , n516 );
or ( n530 , n527 , n528 , n529 );
and ( n531 , n474 , n472 );
and ( n532 , n478 , n475 );
xor ( n533 , n531 , n532 );
and ( n534 , n486 , n479 );
xor ( n535 , n533 , n534 );
xor ( n536 , n530 , n535 );
and ( n537 , n490 , n509 );
and ( n538 , n499 , n484 );
xor ( n539 , n537 , n538 );
and ( n540 , n515 , n487 );
xor ( n541 , n539 , n540 );
xor ( n542 , n536 , n541 );
xor ( n543 , n526 , n542 );
not ( n544 , n471 );
buf ( n545 , n43 );
not ( n546 , n545 );
and ( n547 , n546 , n471 );
nor ( n548 , n544 , n547 );
buf ( n549 , g357 );
not ( n550 , n549 );
and ( n551 , n550 , n491 );
not ( n552 , n491 );
nor ( n553 , n551 , n552 );
xor ( n554 , n548 , n553 );
xor ( n555 , n543 , n554 );
xor ( n556 , n522 , n555 );
and ( n557 , n474 , n479 );
and ( n558 , n478 , n509 );
and ( n559 , n557 , n558 );
and ( n560 , n474 , n484 );
and ( n561 , n478 , n487 );
and ( n562 , n560 , n561 );
and ( n563 , n486 , n491 );
and ( n564 , n561 , n563 );
and ( n565 , n560 , n563 );
or ( n566 , n562 , n564 , n565 );
and ( n567 , n474 , n509 );
and ( n568 , n566 , n567 );
xor ( n569 , n485 , n488 );
xor ( n570 , n569 , n492 );
and ( n571 , n567 , n570 );
and ( n572 , n566 , n570 );
or ( n573 , n568 , n571 , n572 );
xor ( n574 , n557 , n558 );
and ( n575 , n573 , n574 );
xor ( n576 , n495 , n496 );
xor ( n577 , n576 , n501 );
and ( n578 , n574 , n577 );
and ( n579 , n573 , n577 );
or ( n580 , n575 , n578 , n579 );
and ( n581 , n559 , n580 );
xor ( n582 , n504 , n506 );
xor ( n583 , n582 , n518 );
and ( n584 , n580 , n583 );
and ( n585 , n559 , n583 );
or ( n586 , n581 , n584 , n585 );
xor ( n587 , n556 , n586 );
xor ( n588 , n559 , n580 );
xor ( n589 , n588 , n583 );
and ( n590 , n471 , n484 );
and ( n591 , n474 , n487 );
and ( n592 , n590 , n591 );
and ( n593 , n478 , n491 );
and ( n594 , n591 , n593 );
and ( n595 , n590 , n593 );
or ( n596 , n592 , n594 , n595 );
and ( n597 , n471 , n509 );
and ( n598 , n596 , n597 );
xor ( n599 , n560 , n561 );
xor ( n600 , n599 , n563 );
and ( n601 , n597 , n600 );
and ( n602 , n596 , n600 );
or ( n603 , n598 , n601 , n602 );
and ( n604 , n471 , n479 );
and ( n605 , n603 , n604 );
xor ( n606 , n566 , n567 );
xor ( n607 , n606 , n570 );
and ( n608 , n604 , n607 );
and ( n609 , n603 , n607 );
or ( n610 , n605 , n608 , n609 );
xor ( n611 , n573 , n574 );
xor ( n612 , n611 , n577 );
and ( n613 , n610 , n612 );
and ( n614 , n589 , n613 );
xor ( n615 , n589 , n613 );
and ( n616 , n471 , n475 );
xor ( n617 , n610 , n612 );
and ( n618 , n616 , n617 );
xor ( n619 , n616 , n617 );
xor ( n620 , n603 , n604 );
xor ( n621 , n620 , n607 );
xor ( n622 , n596 , n597 );
xor ( n623 , n622 , n600 );
xor ( n624 , n590 , n591 );
xor ( n625 , n624 , n593 );
and ( n626 , n471 , n487 );
and ( n627 , n474 , n491 );
and ( n628 , n626 , n627 );
and ( n629 , n625 , n628 );
and ( n630 , n623 , n629 );
and ( n631 , n621 , n630 );
and ( n632 , n619 , n631 );
or ( n633 , n618 , n632 );
and ( n634 , n615 , n633 );
or ( n635 , n614 , n634 );
xor ( n636 , n587 , n635 );
buf ( n637 , n636 );
xor ( n638 , n450 , n468 );
buf ( n639 , n638 );
buf ( n640 , n639 );
xor ( n641 , n615 , n633 );
buf ( n642 , n641 );
buf ( n643 , n642 );
and ( n644 , n640 , n643 );
xor ( n645 , n454 , n466 );
buf ( n646 , n645 );
buf ( n647 , n646 );
xor ( n648 , n619 , n631 );
buf ( n649 , n648 );
buf ( n650 , n649 );
and ( n651 , n647 , n650 );
xor ( n652 , n456 , n465 );
buf ( n653 , n652 );
buf ( n654 , n653 );
xor ( n655 , n621 , n630 );
buf ( n656 , n655 );
buf ( n657 , n656 );
and ( n658 , n654 , n657 );
xor ( n659 , n458 , n464 );
buf ( n660 , n659 );
buf ( n661 , n660 );
xor ( n662 , n623 , n629 );
buf ( n663 , n662 );
buf ( n664 , n663 );
and ( n665 , n661 , n664 );
xor ( n666 , n460 , n463 );
buf ( n667 , n666 );
buf ( n668 , n667 );
xor ( n669 , n625 , n628 );
buf ( n670 , n669 );
buf ( n671 , n670 );
and ( n672 , n668 , n671 );
xor ( n673 , n461 , n462 );
buf ( n674 , n673 );
buf ( n675 , n674 );
xor ( n676 , n626 , n627 );
buf ( n677 , n676 );
buf ( n678 , n677 );
and ( n679 , n675 , n678 );
and ( n680 , n306 , n326 );
buf ( n681 , n680 );
buf ( n682 , n681 );
and ( n683 , n471 , n491 );
buf ( n684 , n683 );
buf ( n685 , n684 );
and ( n686 , n682 , n685 );
and ( n687 , n678 , n686 );
and ( n688 , n675 , n686 );
or ( n689 , n679 , n687 , n688 );
and ( n690 , n671 , n689 );
and ( n691 , n668 , n689 );
or ( n692 , n672 , n690 , n691 );
and ( n693 , n664 , n692 );
and ( n694 , n661 , n692 );
or ( n695 , n665 , n693 , n694 );
and ( n696 , n657 , n695 );
and ( n697 , n654 , n695 );
or ( n698 , n658 , n696 , n697 );
and ( n699 , n650 , n698 );
and ( n700 , n647 , n698 );
or ( n701 , n651 , n699 , n700 );
and ( n702 , n643 , n701 );
and ( n703 , n640 , n701 );
or ( n704 , n644 , n702 , n703 );
xor ( n705 , t_0 , n704 );
buf ( n706 , n705 );
not ( n1 , n706 );
and ( n2 , n1 , n301 );
and ( n3 , n305 , n706 );
or ( n707 , n2 , n3 );
buf ( n708 , n41 );
buf ( n709 , n49 );
xor ( n710 , n708 , n709 );
and ( n711 , n298 , n299 );
xor ( n712 , n710 , n711 );
buf ( n713 , n712 );
buf ( n714 , g355 );
buf ( n715 , n33 );
xor ( n716 , n714 , n715 );
and ( n717 , n302 , n303 );
xor ( n718 , n716 , n717 );
buf ( n719 , n718 );
not ( n4 , n706 );
and ( n5 , n4 , n713 );
and ( n6 , n719 , n706 );
or ( n720 , n5 , n6 );
buf ( n721 , n40 );
buf ( n722 , n48 );
xor ( n723 , n721 , n722 );
and ( n724 , n708 , n709 );
and ( n725 , n709 , n711 );
and ( n726 , n708 , n711 );
or ( n727 , n724 , n725 , n726 );
xor ( n728 , n723 , n727 );
buf ( n729 , n728 );
buf ( n730 , g354 );
buf ( n731 , n32 );
xor ( n732 , n730 , n731 );
and ( n733 , n714 , n715 );
and ( n734 , n715 , n717 );
and ( n735 , n714 , n717 );
or ( n736 , n733 , n734 , n735 );
xor ( n737 , n732 , n736 );
buf ( n738 , n737 );
not ( n7 , n706 );
and ( n8 , n7 , n729 );
and ( n9 , n738 , n706 );
or ( n739 , n8 , n9 );
buf ( n740 , n39 );
buf ( n741 , n47 );
xor ( n742 , n740 , n741 );
and ( n743 , n721 , n722 );
and ( n744 , n722 , n727 );
and ( n745 , n721 , n727 );
or ( n746 , n743 , n744 , n745 );
xor ( n747 , n742 , n746 );
buf ( n748 , n747 );
buf ( n749 , g353 );
buf ( n750 , n31 );
xor ( n751 , n749 , n750 );
and ( n752 , n730 , n731 );
and ( n753 , n731 , n736 );
and ( n754 , n730 , n736 );
or ( n755 , n752 , n753 , n754 );
xor ( n756 , n751 , n755 );
buf ( n757 , n756 );
not ( n10 , n706 );
and ( n11 , n10 , n748 );
and ( n12 , n757 , n706 );
or ( n758 , n11 , n12 );
buf ( n759 , n38 );
buf ( n760 , n46 );
xor ( n761 , n759 , n760 );
and ( n762 , n740 , n741 );
and ( n763 , n741 , n746 );
and ( n764 , n740 , n746 );
or ( n765 , n762 , n763 , n764 );
xor ( n766 , n761 , n765 );
buf ( n767 , n766 );
buf ( n768 , g352 );
buf ( n769 , n30 );
xor ( n770 , n768 , n769 );
and ( n771 , n749 , n750 );
and ( n772 , n750 , n755 );
and ( n773 , n749 , n755 );
or ( n774 , n771 , n772 , n773 );
xor ( n775 , n770 , n774 );
buf ( n776 , n775 );
not ( n13 , n706 );
and ( n14 , n13 , n767 );
and ( n15 , n776 , n706 );
or ( n777 , n14 , n15 );
buf ( n778 , n37 );
buf ( n779 , n45 );
xor ( n780 , n778 , n779 );
and ( n781 , n759 , n760 );
and ( n782 , n760 , n765 );
and ( n783 , n759 , n765 );
or ( n784 , n781 , n782 , n783 );
xor ( n785 , n780 , n784 );
buf ( n786 , n785 );
buf ( n787 , g351 );
buf ( n788 , n29 );
xor ( n789 , n787 , n788 );
and ( n790 , n768 , n769 );
and ( n791 , n769 , n774 );
and ( n792 , n768 , n774 );
or ( n793 , n790 , n791 , n792 );
xor ( n794 , n789 , n793 );
buf ( n795 , n794 );
not ( n16 , n706 );
and ( n17 , n16 , n786 );
and ( n18 , n795 , n706 );
or ( n796 , n17 , n18 );
buf ( n797 , n36 );
buf ( n798 , n44 );
xor ( n799 , n797 , n798 );
and ( n800 , n778 , n779 );
and ( n801 , n779 , n784 );
and ( n802 , n778 , n784 );
or ( n803 , n800 , n801 , n802 );
xor ( n804 , n799 , n803 );
buf ( n805 , n804 );
buf ( n806 , g350 );
buf ( n807 , n28 );
xor ( n808 , n806 , n807 );
and ( n809 , n787 , n788 );
and ( n810 , n788 , n793 );
and ( n811 , n787 , n793 );
or ( n812 , n809 , n810 , n811 );
xor ( n813 , n808 , n812 );
buf ( n814 , n813 );
not ( n19 , n706 );
and ( n20 , n19 , n805 );
and ( n21 , n814 , n706 );
or ( n815 , n20 , n21 );
buf ( n816 , n35 );
buf ( n817 , n43 );
xor ( n818 , n816 , n817 );
and ( n819 , n797 , n798 );
and ( n820 , n798 , n803 );
and ( n821 , n797 , n803 );
or ( n822 , n819 , n820 , n821 );
xor ( n823 , n818 , n822 );
buf ( n824 , n823 );
buf ( n825 , g349 );
buf ( n826 , g357 );
xor ( n827 , n825 , n826 );
and ( n828 , n806 , n807 );
and ( n829 , n807 , n812 );
and ( n830 , n806 , n812 );
or ( n831 , n828 , n829 , n830 );
xor ( n832 , n827 , n831 );
buf ( n833 , n832 );
not ( n22 , n706 );
and ( n23 , n22 , n824 );
and ( n24 , n833 , n706 );
or ( n834 , n23 , n24 );
and ( n835 , n816 , n817 );
and ( n836 , n817 , n822 );
and ( n837 , n816 , n822 );
or ( n838 , n835 , n836 , n837 );
buf ( n839 , n838 );
and ( n840 , n825 , n826 );
and ( n841 , n826 , n831 );
and ( n842 , n825 , n831 );
or ( n843 , n840 , n841 , n842 );
buf ( n844 , n843 );
not ( n25 , n706 );
and ( n26 , n25 , n839 );
and ( n27 , n844 , n706 );
or ( n845 , n26 , n27 );
xor ( n846 , n640 , n643 );
xor ( n847 , n846 , n701 );
buf ( n848 , n847 );
xor ( n849 , n647 , n650 );
xor ( n850 , n849 , n698 );
buf ( n851 , n850 );
xor ( n852 , n654 , n657 );
xor ( n853 , n852 , n695 );
buf ( n854 , n853 );
xor ( n855 , n661 , n664 );
xor ( n856 , n855 , n692 );
buf ( n857 , n856 );
xor ( n858 , n668 , n671 );
xor ( n859 , n858 , n689 );
buf ( n860 , n859 );
xor ( n861 , n675 , n678 );
xor ( n862 , n861 , n686 );
buf ( n863 , n862 );
xor ( n864 , n682 , n685 );
buf ( n865 , n864 );
and ( n866 , n549 , n545 );
not ( n867 , n490 );
and ( n868 , n546 , n490 );
nor ( n869 , n867 , n868 );
and ( n870 , n499 , n472 );
and ( n871 , n869 , n870 );
and ( n872 , n515 , n475 );
and ( n873 , n870 , n872 );
and ( n874 , n869 , n872 );
or ( n875 , n871 , n873 , n874 );
not ( n876 , n499 );
and ( n877 , n546 , n499 );
nor ( n878 , n876 , n877 );
and ( n879 , n875 , n878 );
and ( n880 , n515 , n472 );
and ( n881 , n878 , n880 );
and ( n882 , n875 , n880 );
or ( n883 , n879 , n881 , n882 );
not ( n884 , n515 );
and ( n885 , n546 , n515 );
nor ( n886 , n884 , n885 );
and ( n887 , n883 , n886 );
and ( n888 , n550 , n472 );
not ( n889 , n472 );
nor ( n890 , n888 , n889 );
and ( n891 , n886 , n890 );
and ( n892 , n883 , n890 );
or ( n893 , n887 , n891 , n892 );
and ( n894 , n866 , n893 );
xor ( n895 , n866 , n893 );
xor ( n896 , n883 , n886 );
xor ( n897 , n896 , n890 );
not ( n898 , n486 );
and ( n899 , n546 , n486 );
nor ( n900 , n898 , n899 );
and ( n901 , n490 , n472 );
and ( n902 , n900 , n901 );
and ( n903 , n550 , n509 );
not ( n904 , n509 );
nor ( n905 , n903 , n904 );
and ( n906 , n901 , n905 );
and ( n907 , n900 , n905 );
or ( n908 , n902 , n906 , n907 );
and ( n909 , n490 , n475 );
and ( n910 , n499 , n479 );
and ( n911 , n909 , n910 );
and ( n912 , n515 , n509 );
and ( n913 , n910 , n912 );
and ( n914 , n909 , n912 );
or ( n915 , n911 , n913 , n914 );
and ( n916 , n499 , n475 );
and ( n917 , n915 , n916 );
and ( n918 , n515 , n479 );
and ( n919 , n916 , n918 );
and ( n920 , n915 , n918 );
or ( n921 , n917 , n919 , n920 );
and ( n922 , n908 , n921 );
xor ( n923 , n869 , n870 );
xor ( n924 , n923 , n872 );
and ( n925 , n921 , n924 );
and ( n926 , n908 , n924 );
or ( n927 , n922 , n925 , n926 );
and ( n928 , n550 , n475 );
not ( n929 , n475 );
nor ( n930 , n928 , n929 );
and ( n931 , n927 , n930 );
xor ( n932 , n875 , n878 );
xor ( n933 , n932 , n880 );
and ( n934 , n930 , n933 );
and ( n935 , n927 , n933 );
or ( n936 , n931 , n934 , n935 );
and ( n937 , n897 , n936 );
xor ( n938 , n897 , n936 );
xor ( n939 , n927 , n930 );
xor ( n940 , n939 , n933 );
and ( n941 , n490 , n479 );
and ( n942 , n499 , n509 );
and ( n943 , n941 , n942 );
and ( n944 , n515 , n484 );
and ( n945 , n942 , n944 );
and ( n946 , n941 , n944 );
or ( n947 , n943 , n945 , n946 );
and ( n948 , n478 , n472 );
and ( n949 , n486 , n475 );
and ( n950 , n948 , n949 );
and ( n951 , n947 , n950 );
xor ( n952 , n909 , n910 );
xor ( n953 , n952 , n912 );
and ( n954 , n950 , n953 );
and ( n955 , n947 , n953 );
or ( n956 , n951 , n954 , n955 );
xor ( n957 , n900 , n901 );
xor ( n958 , n957 , n905 );
and ( n959 , n956 , n958 );
xor ( n960 , n915 , n916 );
xor ( n961 , n960 , n918 );
and ( n962 , n958 , n961 );
and ( n963 , n956 , n961 );
or ( n964 , n959 , n962 , n963 );
and ( n965 , n550 , n479 );
not ( n966 , n479 );
nor ( n967 , n965 , n966 );
and ( n968 , n964 , n967 );
xor ( n969 , n908 , n921 );
xor ( n970 , n969 , n924 );
and ( n971 , n967 , n970 );
and ( n972 , n964 , n970 );
or ( n973 , n968 , n971 , n972 );
and ( n974 , n940 , n973 );
xor ( n975 , n940 , n973 );
xor ( n976 , n964 , n967 );
xor ( n977 , n976 , n970 );
not ( n978 , n478 );
and ( n979 , n546 , n478 );
nor ( n980 , n978 , n979 );
and ( n981 , n486 , n472 );
and ( n982 , n980 , n981 );
and ( n983 , n550 , n484 );
not ( n984 , n484 );
nor ( n985 , n983 , n984 );
and ( n986 , n981 , n985 );
and ( n987 , n980 , n985 );
or ( n988 , n982 , n986 , n987 );
and ( n989 , n537 , n538 );
and ( n990 , n538 , n540 );
and ( n991 , n537 , n540 );
or ( n992 , n989 , n990 , n991 );
xor ( n993 , n941 , n942 );
xor ( n994 , n993 , n944 );
and ( n995 , n992 , n994 );
xor ( n996 , n948 , n949 );
and ( n997 , n994 , n996 );
and ( n998 , n992 , n996 );
or ( n999 , n995 , n997 , n998 );
xor ( n1000 , n980 , n981 );
xor ( n1001 , n1000 , n985 );
and ( n1002 , n999 , n1001 );
xor ( n1003 , n947 , n950 );
xor ( n1004 , n1003 , n953 );
and ( n1005 , n1001 , n1004 );
and ( n1006 , n999 , n1004 );
or ( n1007 , n1002 , n1005 , n1006 );
and ( n1008 , n988 , n1007 );
xor ( n1009 , n956 , n958 );
xor ( n1010 , n1009 , n961 );
and ( n1011 , n1007 , n1010 );
and ( n1012 , n988 , n1010 );
or ( n1013 , n1008 , n1011 , n1012 );
and ( n1014 , n977 , n1013 );
xor ( n1015 , n977 , n1013 );
xor ( n1016 , n988 , n1007 );
xor ( n1017 , n1016 , n1010 );
and ( n1018 , n531 , n532 );
and ( n1019 , n532 , n534 );
and ( n1020 , n531 , n534 );
or ( n1021 , n1018 , n1019 , n1020 );
not ( n1022 , n474 );
and ( n1023 , n546 , n474 );
nor ( n1024 , n1022 , n1023 );
and ( n1025 , n1021 , n1024 );
and ( n1026 , n550 , n487 );
not ( n1027 , n487 );
nor ( n1028 , n1026 , n1027 );
and ( n1029 , n1024 , n1028 );
and ( n1030 , n1021 , n1028 );
or ( n1031 , n1025 , n1029 , n1030 );
and ( n1032 , n530 , n535 );
and ( n1033 , n535 , n541 );
and ( n1034 , n530 , n541 );
or ( n1035 , n1032 , n1033 , n1034 );
xor ( n1036 , n1021 , n1024 );
xor ( n1037 , n1036 , n1028 );
and ( n1038 , n1035 , n1037 );
xor ( n1039 , n992 , n994 );
xor ( n1040 , n1039 , n996 );
and ( n1041 , n1037 , n1040 );
and ( n1042 , n1035 , n1040 );
or ( n1043 , n1038 , n1041 , n1042 );
and ( n1044 , n1031 , n1043 );
xor ( n1045 , n999 , n1001 );
xor ( n1046 , n1045 , n1004 );
and ( n1047 , n1043 , n1046 );
and ( n1048 , n1031 , n1046 );
or ( n1049 , n1044 , n1047 , n1048 );
and ( n1050 , n1017 , n1049 );
xor ( n1051 , n1017 , n1049 );
xor ( n1052 , n1031 , n1043 );
xor ( n1053 , n1052 , n1046 );
and ( n1054 , n548 , n553 );
and ( n1055 , n526 , n542 );
and ( n1056 , n542 , n554 );
and ( n1057 , n526 , n554 );
or ( n1058 , n1055 , n1056 , n1057 );
and ( n1059 , n1054 , n1058 );
xor ( n1060 , n1035 , n1037 );
xor ( n1061 , n1060 , n1040 );
and ( n1062 , n1058 , n1061 );
and ( n1063 , n1054 , n1061 );
or ( n1064 , n1059 , n1062 , n1063 );
and ( n1065 , n1053 , n1064 );
xor ( n1066 , n1053 , n1064 );
xor ( n1067 , n1054 , n1058 );
xor ( n1068 , n1067 , n1061 );
and ( n1069 , n483 , n521 );
and ( n1070 , n521 , n555 );
and ( n1071 , n483 , n555 );
or ( n1072 , n1069 , n1070 , n1071 );
and ( n1073 , n1068 , n1072 );
xor ( n1074 , n1068 , n1072 );
and ( n1075 , n556 , n586 );
and ( n1076 , n587 , n635 );
or ( n1077 , n1075 , n1076 );
and ( n1078 , n1074 , n1077 );
or ( n1079 , n1073 , n1078 );
and ( n1080 , n1066 , n1079 );
or ( n1081 , n1065 , n1080 );
and ( n1082 , n1051 , n1081 );
or ( n1083 , n1050 , n1082 );
and ( n1084 , n1015 , n1083 );
or ( n1085 , n1014 , n1084 );
and ( n1086 , n975 , n1085 );
or ( n1087 , n974 , n1086 );
and ( n1088 , n938 , n1087 );
or ( n1089 , n937 , n1088 );
and ( n1090 , n895 , n1089 );
or ( n1091 , n894 , n1090 );
buf ( n1092 , n1091 );
xor ( n1093 , n895 , n1089 );
buf ( n1094 , n1093 );
xor ( n1095 , n938 , n1087 );
buf ( n1096 , n1095 );
xor ( n1097 , n975 , n1085 );
buf ( n1098 , n1097 );
xor ( n1099 , n1015 , n1083 );
buf ( n1100 , n1099 );
xor ( n1101 , n1051 , n1081 );
buf ( n1102 , n1101 );
xor ( n1103 , n1066 , n1079 );
buf ( n1104 , n1103 );
xor ( n1105 , n1074 , n1077 );
buf ( n1106 , n1105 );
and ( n1107 , n384 , n380 );
not ( n1108 , n325 );
and ( n1109 , n381 , n325 );
nor ( n1110 , n1108 , n1109 );
and ( n1111 , n334 , n307 );
and ( n1112 , n1110 , n1111 );
and ( n1113 , n350 , n310 );
and ( n1114 , n1111 , n1113 );
and ( n1115 , n1110 , n1113 );
or ( n1116 , n1112 , n1114 , n1115 );
not ( n1117 , n334 );
and ( n1118 , n381 , n334 );
nor ( n1119 , n1117 , n1118 );
and ( n1120 , n1116 , n1119 );
and ( n1121 , n350 , n307 );
and ( n1122 , n1119 , n1121 );
and ( n1123 , n1116 , n1121 );
or ( n1124 , n1120 , n1122 , n1123 );
not ( n1125 , n350 );
and ( n1126 , n381 , n350 );
nor ( n1127 , n1125 , n1126 );
and ( n1128 , n1124 , n1127 );
and ( n1129 , n385 , n307 );
not ( n1130 , n307 );
nor ( n1131 , n1129 , n1130 );
and ( n1132 , n1127 , n1131 );
and ( n1133 , n1124 , n1131 );
or ( n1134 , n1128 , n1132 , n1133 );
and ( n1135 , n1107 , n1134 );
xor ( n1136 , n1107 , n1134 );
xor ( n1137 , n1124 , n1127 );
xor ( n1138 , n1137 , n1131 );
not ( n1139 , n321 );
and ( n1140 , n381 , n321 );
nor ( n1141 , n1139 , n1140 );
and ( n1142 , n325 , n307 );
and ( n1143 , n1141 , n1142 );
and ( n1144 , n385 , n344 );
not ( n1145 , n344 );
nor ( n1146 , n1144 , n1145 );
and ( n1147 , n1142 , n1146 );
and ( n1148 , n1141 , n1146 );
or ( n1149 , n1143 , n1147 , n1148 );
and ( n1150 , n325 , n310 );
and ( n1151 , n334 , n314 );
and ( n1152 , n1150 , n1151 );
and ( n1153 , n350 , n344 );
and ( n1154 , n1151 , n1153 );
and ( n1155 , n1150 , n1153 );
or ( n1156 , n1152 , n1154 , n1155 );
and ( n1157 , n334 , n310 );
and ( n1158 , n1156 , n1157 );
and ( n1159 , n350 , n314 );
and ( n1160 , n1157 , n1159 );
and ( n1161 , n1156 , n1159 );
or ( n1162 , n1158 , n1160 , n1161 );
and ( n1163 , n1149 , n1162 );
xor ( n1164 , n1110 , n1111 );
xor ( n1165 , n1164 , n1113 );
and ( n1166 , n1162 , n1165 );
and ( n1167 , n1149 , n1165 );
or ( n1168 , n1163 , n1166 , n1167 );
and ( n1169 , n385 , n310 );
not ( n1170 , n310 );
nor ( n1171 , n1169 , n1170 );
and ( n1172 , n1168 , n1171 );
xor ( n1173 , n1116 , n1119 );
xor ( n1174 , n1173 , n1121 );
and ( n1175 , n1171 , n1174 );
and ( n1176 , n1168 , n1174 );
or ( n1177 , n1172 , n1175 , n1176 );
and ( n1178 , n1138 , n1177 );
xor ( n1179 , n1138 , n1177 );
xor ( n1180 , n1168 , n1171 );
xor ( n1181 , n1180 , n1174 );
and ( n1182 , n325 , n314 );
and ( n1183 , n334 , n344 );
and ( n1184 , n1182 , n1183 );
and ( n1185 , n350 , n319 );
and ( n1186 , n1183 , n1185 );
and ( n1187 , n1182 , n1185 );
or ( n1188 , n1184 , n1186 , n1187 );
and ( n1189 , n313 , n307 );
and ( n1190 , n321 , n310 );
and ( n1191 , n1189 , n1190 );
and ( n1192 , n1188 , n1191 );
xor ( n1193 , n1150 , n1151 );
xor ( n1194 , n1193 , n1153 );
and ( n1195 , n1191 , n1194 );
and ( n1196 , n1188 , n1194 );
or ( n1197 , n1192 , n1195 , n1196 );
xor ( n1198 , n1141 , n1142 );
xor ( n1199 , n1198 , n1146 );
and ( n1200 , n1197 , n1199 );
xor ( n1201 , n1156 , n1157 );
xor ( n1202 , n1201 , n1159 );
and ( n1203 , n1199 , n1202 );
and ( n1204 , n1197 , n1202 );
or ( n1205 , n1200 , n1203 , n1204 );
and ( n1206 , n385 , n314 );
not ( n1207 , n314 );
nor ( n1208 , n1206 , n1207 );
and ( n1209 , n1205 , n1208 );
xor ( n1210 , n1149 , n1162 );
xor ( n1211 , n1210 , n1165 );
and ( n1212 , n1208 , n1211 );
and ( n1213 , n1205 , n1211 );
or ( n1214 , n1209 , n1212 , n1213 );
and ( n1215 , n1181 , n1214 );
xor ( n1216 , n1181 , n1214 );
xor ( n1217 , n1205 , n1208 );
xor ( n1218 , n1217 , n1211 );
not ( n1219 , n313 );
and ( n1220 , n381 , n313 );
nor ( n1221 , n1219 , n1220 );
and ( n1222 , n321 , n307 );
and ( n1223 , n1221 , n1222 );
and ( n1224 , n385 , n319 );
not ( n1225 , n319 );
nor ( n1226 , n1224 , n1225 );
and ( n1227 , n1222 , n1226 );
and ( n1228 , n1221 , n1226 );
or ( n1229 , n1223 , n1227 , n1228 );
and ( n1230 , n372 , n373 );
and ( n1231 , n373 , n375 );
and ( n1232 , n372 , n375 );
or ( n1233 , n1230 , n1231 , n1232 );
xor ( n1234 , n1182 , n1183 );
xor ( n1235 , n1234 , n1185 );
and ( n1236 , n1233 , n1235 );
xor ( n1237 , n1189 , n1190 );
and ( n1238 , n1235 , n1237 );
and ( n1239 , n1233 , n1237 );
or ( n1240 , n1236 , n1238 , n1239 );
xor ( n1241 , n1221 , n1222 );
xor ( n1242 , n1241 , n1226 );
and ( n1243 , n1240 , n1242 );
xor ( n1244 , n1188 , n1191 );
xor ( n1245 , n1244 , n1194 );
and ( n1246 , n1242 , n1245 );
and ( n1247 , n1240 , n1245 );
or ( n1248 , n1243 , n1246 , n1247 );
and ( n1249 , n1229 , n1248 );
xor ( n1250 , n1197 , n1199 );
xor ( n1251 , n1250 , n1202 );
and ( n1252 , n1248 , n1251 );
and ( n1253 , n1229 , n1251 );
or ( n1254 , n1249 , n1252 , n1253 );
and ( n1255 , n1218 , n1254 );
xor ( n1256 , n1218 , n1254 );
xor ( n1257 , n1229 , n1248 );
xor ( n1258 , n1257 , n1251 );
and ( n1259 , n366 , n367 );
and ( n1260 , n367 , n369 );
and ( n1261 , n366 , n369 );
or ( n1262 , n1259 , n1260 , n1261 );
not ( n1263 , n309 );
and ( n1264 , n381 , n309 );
nor ( n1265 , n1263 , n1264 );
and ( n1266 , n1262 , n1265 );
and ( n1267 , n385 , n322 );
not ( n1268 , n322 );
nor ( n1269 , n1267 , n1268 );
and ( n1270 , n1265 , n1269 );
and ( n1271 , n1262 , n1269 );
or ( n1272 , n1266 , n1270 , n1271 );
and ( n1273 , n365 , n370 );
and ( n1274 , n370 , n376 );
and ( n1275 , n365 , n376 );
or ( n1276 , n1273 , n1274 , n1275 );
xor ( n1277 , n1262 , n1265 );
xor ( n1278 , n1277 , n1269 );
and ( n1279 , n1276 , n1278 );
xor ( n1280 , n1233 , n1235 );
xor ( n1281 , n1280 , n1237 );
and ( n1282 , n1278 , n1281 );
and ( n1283 , n1276 , n1281 );
or ( n1284 , n1279 , n1282 , n1283 );
and ( n1285 , n1272 , n1284 );
xor ( n1286 , n1240 , n1242 );
xor ( n1287 , n1286 , n1245 );
and ( n1288 , n1284 , n1287 );
and ( n1289 , n1272 , n1287 );
or ( n1290 , n1285 , n1288 , n1289 );
and ( n1291 , n1258 , n1290 );
xor ( n1292 , n1258 , n1290 );
xor ( n1293 , n1272 , n1284 );
xor ( n1294 , n1293 , n1287 );
and ( n1295 , n383 , n388 );
and ( n1296 , n361 , n377 );
and ( n1297 , n377 , n389 );
and ( n1298 , n361 , n389 );
or ( n1299 , n1296 , n1297 , n1298 );
and ( n1300 , n1295 , n1299 );
xor ( n1301 , n1276 , n1278 );
xor ( n1302 , n1301 , n1281 );
and ( n1303 , n1299 , n1302 );
and ( n1304 , n1295 , n1302 );
or ( n1305 , n1300 , n1303 , n1304 );
and ( n1306 , n1294 , n1305 );
xor ( n1307 , n1294 , n1305 );
xor ( n1308 , n1295 , n1299 );
xor ( n1309 , n1308 , n1302 );
and ( n1310 , n318 , n356 );
and ( n1311 , n356 , n390 );
and ( n1312 , n318 , n390 );
or ( n1313 , n1310 , n1311 , n1312 );
and ( n1314 , n1309 , n1313 );
xor ( n1315 , n1309 , n1313 );
and ( n1316 , n391 , n421 );
and ( n1317 , n422 , n470 );
or ( n1318 , n1316 , n1317 );
and ( n1319 , n1315 , n1318 );
or ( n1320 , n1314 , n1319 );
and ( n1321 , n1307 , n1320 );
or ( n1322 , n1306 , n1321 );
and ( n1323 , n1292 , n1322 );
or ( n1324 , n1291 , n1323 );
and ( n1325 , n1256 , n1324 );
or ( n1326 , n1255 , n1325 );
and ( n1327 , n1216 , n1326 );
or ( n1328 , n1215 , n1327 );
and ( n1329 , n1179 , n1328 );
or ( n1330 , n1178 , n1329 );
and ( n1331 , n1136 , n1330 );
or ( n1332 , n1135 , n1331 );
buf ( n1333 , n1332 );
xor ( n1334 , n1136 , n1330 );
buf ( n1335 , n1334 );
xor ( n1336 , n1179 , n1328 );
buf ( n1337 , n1336 );
xor ( n1338 , n1216 , n1326 );
buf ( n1339 , n1338 );
xor ( n1340 , n1256 , n1324 );
buf ( n1341 , n1340 );
xor ( n1342 , n1292 , n1322 );
buf ( n1343 , n1342 );
xor ( n1344 , n1307 , n1320 );
buf ( n1345 , n1344 );
xor ( n1346 , n1315 , n1318 );
buf ( n1347 , n1346 );
buf ( n1348 , n845 );
buf ( n1349 , n834 );
buf ( n1350 , n815 );
buf ( n1351 , n796 );
buf ( n1352 , n777 );
buf ( n1353 , n758 );
buf ( n1354 , n739 );
buf ( n1355 , n720 );
buf ( n1356 , n707 );
buf ( n1357 , n1092 );
buf ( n1358 , n1094 );
buf ( n1359 , n1096 );
buf ( n1360 , n1098 );
buf ( n1361 , n1100 );
buf ( n1362 , n1102 );
buf ( n1363 , n1104 );
buf ( n1364 , n1106 );
buf ( n1365 , n637 );
buf ( n1366 , n642 );
buf ( n1367 , n649 );
buf ( n1368 , n656 );
buf ( n1369 , n663 );
buf ( n1370 , n670 );
buf ( n1371 , n677 );
buf ( n1372 , n684 );
and ( n1373 , n1348 , n1364 );
and ( n1374 , n1349 , n1365 );
and ( n1375 , n1350 , n1366 );
and ( n1376 , n1351 , n1367 );
and ( n1377 , n1352 , n1368 );
and ( n1378 , n1353 , n1369 );
and ( n1379 , n1354 , n1370 );
and ( n1380 , n1355 , n1371 );
and ( n1381 , n1356 , n1372 );
and ( n1382 , n1371 , n1381 );
and ( n1383 , n1355 , n1381 );
or ( n1384 , n1380 , n1382 , n1383 );
and ( n1385 , n1370 , n1384 );
and ( n1386 , n1354 , n1384 );
or ( n1387 , n1379 , n1385 , n1386 );
and ( n1388 , n1369 , n1387 );
and ( n1389 , n1353 , n1387 );
or ( n1390 , n1378 , n1388 , n1389 );
and ( n1391 , n1368 , n1390 );
and ( n1392 , n1352 , n1390 );
or ( n1393 , n1377 , n1391 , n1392 );
and ( n1394 , n1367 , n1393 );
and ( n1395 , n1351 , n1393 );
or ( n1396 , n1376 , n1394 , n1395 );
and ( n1397 , n1366 , n1396 );
and ( n1398 , n1350 , n1396 );
or ( n1399 , n1375 , n1397 , n1398 );
and ( n1400 , n1365 , n1399 );
and ( n1401 , n1349 , n1399 );
or ( n1402 , n1374 , n1400 , n1401 );
and ( n1403 , n1364 , n1402 );
and ( n1404 , n1348 , n1402 );
or ( n1405 , n1373 , n1403 , n1404 );
and ( n1406 , n1363 , n1405 );
and ( n1407 , n1362 , n1406 );
and ( n1408 , n1361 , n1407 );
and ( n1409 , n1360 , n1408 );
and ( n1410 , n1359 , n1409 );
and ( n1411 , n1358 , n1410 );
and ( n1412 , n1357 , n1411 );
buf ( n1413 , n1412 );
xor ( n1414 , n1357 , n1411 );
buf ( n1415 , n1414 );
xor ( n1416 , n1358 , n1410 );
buf ( n1417 , n1416 );
xor ( n1418 , n1359 , n1409 );
buf ( n1419 , n1418 );
xor ( n1420 , n1360 , n1408 );
buf ( n1421 , n1420 );
xor ( n1422 , n1361 , n1407 );
buf ( n1423 , n1422 );
xor ( n1424 , n1362 , n1406 );
buf ( n1425 , n1424 );
xor ( n1426 , n1363 , n1405 );
buf ( n1427 , n1426 );
xor ( n1428 , n1348 , n1364 );
xor ( n1429 , n1428 , n1402 );
buf ( n1430 , n1429 );
xor ( n1431 , n1349 , n1365 );
xor ( n1432 , n1431 , n1399 );
buf ( n1433 , n1432 );
xor ( n1434 , n1350 , n1366 );
xor ( n1435 , n1434 , n1396 );
buf ( n1436 , n1435 );
xor ( n1437 , n1351 , n1367 );
xor ( n1438 , n1437 , n1393 );
buf ( n1439 , n1438 );
xor ( n1440 , n1352 , n1368 );
xor ( n1441 , n1440 , n1390 );
buf ( n1442 , n1441 );
xor ( n1443 , n1353 , n1369 );
xor ( n1444 , n1443 , n1387 );
buf ( n1445 , n1444 );
xor ( n1446 , n1354 , n1370 );
xor ( n1447 , n1446 , n1384 );
buf ( n1448 , n1447 );
xor ( n1449 , n1355 , n1371 );
xor ( n1450 , n1449 , n1381 );
buf ( n1451 , n1450 );
xor ( n1452 , n1356 , n1372 );
buf ( n1453 , n1452 );
buf ( n1454 , n845 );
buf ( n1455 , n834 );
buf ( n1456 , n815 );
buf ( n1457 , n796 );
buf ( n1458 , n777 );
buf ( n1459 , n758 );
buf ( n1460 , n739 );
buf ( n1461 , n720 );
buf ( n1462 , n707 );
buf ( n1463 , n1333 );
buf ( n1464 , n1335 );
buf ( n1465 , n1337 );
buf ( n1466 , n1339 );
buf ( n1467 , n1341 );
buf ( n1468 , n1343 );
buf ( n1469 , n1345 );
buf ( n1470 , n1347 );
buf ( n1471 , n639 );
buf ( n1472 , n646 );
buf ( n1473 , n653 );
buf ( n1474 , n660 );
buf ( n1475 , n667 );
buf ( n1476 , n674 );
buf ( n1477 , n681 );
and ( n1478 , n1454 , n1470 );
and ( n1479 , n1455 , t_1 );
and ( n1480 , n1456 , n1471 );
and ( n1481 , n1457 , n1472 );
and ( n1482 , n1458 , n1473 );
and ( n1483 , n1459 , n1474 );
and ( n1484 , n1460 , n1475 );
and ( n1485 , n1461 , n1476 );
and ( n1486 , n1462 , n1477 );
and ( n1487 , n1476 , n1486 );
and ( n1488 , n1461 , n1486 );
or ( n1489 , n1485 , n1487 , n1488 );
and ( n1490 , n1475 , n1489 );
and ( n1491 , n1460 , n1489 );
or ( n1492 , n1484 , n1490 , n1491 );
and ( n1493 , n1474 , n1492 );
and ( n1494 , n1459 , n1492 );
or ( n1495 , n1483 , n1493 , n1494 );
and ( n1496 , n1473 , n1495 );
and ( n1497 , n1458 , n1495 );
or ( n1498 , n1482 , n1496 , n1497 );
and ( n1499 , n1472 , n1498 );
and ( n1500 , n1457 , n1498 );
or ( n1501 , n1481 , n1499 , n1500 );
and ( n1502 , n1471 , n1501 );
and ( n1503 , n1456 , n1501 );
or ( n1504 , n1480 , n1502 , n1503 );
and ( n1505 , t_1 , n1504 );
and ( n1506 , n1455 , n1504 );
or ( n1507 , n1479 , n1505 , n1506 );
and ( n1508 , n1470 , n1507 );
and ( n1509 , n1454 , n1507 );
or ( n1510 , n1478 , n1508 , n1509 );
and ( n1511 , n1469 , n1510 );
and ( n1512 , n1468 , n1511 );
and ( n1513 , n1467 , n1512 );
and ( n1514 , n1466 , n1513 );
and ( n1515 , n1465 , n1514 );
and ( n1516 , n1464 , n1515 );
and ( n1517 , n1463 , n1516 );
buf ( n1518 , n1517 );
xor ( n1519 , n1463 , n1516 );
buf ( n1520 , n1519 );
xor ( n1521 , n1464 , n1515 );
buf ( n1522 , n1521 );
xor ( n1523 , n1465 , n1514 );
buf ( n1524 , n1523 );
xor ( n1525 , n1466 , n1513 );
buf ( n1526 , n1525 );
xor ( n1527 , n1467 , n1512 );
buf ( n1528 , n1527 );
xor ( n1529 , n1468 , n1511 );
buf ( n1530 , n1529 );
xor ( n1531 , n1469 , n1510 );
buf ( n1532 , n1531 );
xor ( n1533 , n1454 , n1470 );
xor ( n1534 , n1533 , n1507 );
buf ( n1535 , n1534 );
xor ( n1536 , n1455 , t_1 );
xor ( n1537 , n1536 , n1504 );
buf ( n1538 , n1537 );
xor ( n1539 , n1456 , n1471 );
xor ( n1540 , n1539 , n1501 );
buf ( n1541 , n1540 );
xor ( n1542 , n1457 , n1472 );
xor ( n1543 , n1542 , n1498 );
buf ( n1544 , n1543 );
xor ( n1545 , n1458 , n1473 );
xor ( n1546 , n1545 , n1495 );
buf ( n1547 , n1546 );
xor ( n1548 , n1459 , n1474 );
xor ( n1549 , n1548 , n1492 );
buf ( n1550 , n1549 );
xor ( n1551 , n1460 , n1475 );
xor ( n1552 , n1551 , n1489 );
buf ( n1553 , n1552 );
xor ( n1554 , n1461 , n1476 );
xor ( n1555 , n1554 , n1486 );
buf ( n1556 , n1555 );
xor ( n1557 , n1462 , n1477 );
buf ( n1558 , n1557 );
endmodule
