module top ( g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 , g98 , g99 , g100 , g101 , g102 , g103 , g104 , g105 , g106 , g107 , g108 , g109 , g110 , g111 , g112 , g113 , g114 , g115 , g116 , g117 , g118 , g119 , g120 , g121 , g122 , g123 , g124 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g136 , g137 , g138 , g139 , g140 , g141 , g142 , g143 , g144 , g145 , g146 , g147 , g148 , g149 , g150 , g151 , g152 , g153 , g154 , g155 , g156 , g157 , g158 , g159 , g160 );
input g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 ;
output g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 , g98 , g99 , g100 , g101 , g102 , g103 , g104 , g105 , g106 , g107 , g108 , g109 , g110 , g111 , g112 , g113 , g114 , g115 , g116 , g117 , g118 , g119 , g120 , g121 , g122 , g123 , g124 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g136 , g137 , g138 , g139 , g140 , g141 , g142 , g143 , g144 , g145 , g146 , g147 , g148 , g149 , g150 , g151 , g152 , g153 , g154 , g155 , g156 , g157 , g158 , g159 , g160 ;

wire n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , 
     n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , 
     n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , 
     n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , 
     n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , 
     n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , 
     n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , 
     n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , 
     n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , 
     n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , 
     n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , 
     n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , 
     n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , 
     n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , 
     n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , 
     n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , 
     n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , 
     n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , 
     n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , 
     n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , 
     n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , 
     n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , 
     n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , 
     n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , 
     n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , 
     n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , 
     n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , 
     n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , 
     n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , 
     n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , 
     n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , 
     n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , 
     n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , 
     n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , 
     n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , 
     n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , 
     n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , 
     n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , 
     n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , 
     n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , 
     n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , 
     n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , 
     n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , 
     n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , 
     n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , 
     n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , 
     n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , 
     n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , 
     n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , 
     n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , 
     n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , 
     n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , 
     n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , 
     n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , 
     n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , 
     n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , 
     n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , 
     n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , 
     n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , 
     n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , 
     n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , 
     n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , 
     n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , 
     n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , 
     n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , 
     n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , 
     n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , 
     n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , 
     n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , 
     n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , 
     n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , 
     n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , 
     n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , 
     n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , 
     n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , 
     n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , 
     n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , 
     n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , 
     n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , 
     n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , 
     n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , 
     n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , 
     n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , 
     n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , 
     n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , 
     n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , 
     n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , 
     n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , 
     n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , 
     n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , 
     n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , 
     n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , 
     n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , 
     n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , 
     n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , 
     n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , 
     n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , 
     n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , 
     n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , 
     n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , 
     n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , 
     n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , 
     n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , 
     n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , 
     n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , 
     n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , 
     n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , 
     n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , 
     n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , 
     n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , 
     n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , 
     n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , 
     n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , 
     n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , 
     n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , 
     n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , 
     n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , 
     n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , 
     n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , 
     n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , 
     n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , 
     n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , 
     n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , 
     n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , 
     n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , 
     n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , 
     n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , 
     n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , 
     n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , 
     n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , 
     n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , 
     n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , 
     n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , 
     n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , 
     n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , 
     n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , 
     n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , 
     n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , 
     n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , 
     n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , 
     n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , 
     n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , 
     n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , 
     n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , 
     n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , 
     n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , 
     n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , 
     n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , 
     n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , 
     n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , 
     n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , 
     n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , 
     n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , 
     n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , 
     n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , 
     n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , 
     n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , 
     n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , 
     n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , 
     n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , 
     n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , 
     n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , 
     n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , 
     n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , 
     n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , 
     n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , 
     n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , 
     n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , 
     n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , 
     n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , 
     n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , 
     n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , 
     n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , 
     n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , 
     n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , 
     n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , 
     n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , 
     n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , 
     n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , 
     n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , 
     n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , 
     n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , 
     n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , 
     n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , 
     n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , 
     n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , 
     n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , 
     n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , 
     n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , 
     n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , 
     n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , 
     n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , 
     n1920 , n1921 , n1922 , n1923 , n1924 , n1925 ;
buf ( n1  , g0 );
buf ( n2  , g1 );
buf ( n3  , g2 );
buf ( n4  , g3 );
buf ( n5  , g4 );
buf ( n6  , g5 );
buf ( n7  , g6 );
buf ( n8  , g7 );
buf ( n9  , g8 );
buf ( n10  , g9 );
buf ( n11  , g10 );
buf ( n12  , g11 );
buf ( n13  , g12 );
buf ( n14  , g13 );
buf ( n15  , g14 );
buf ( n16  , g15 );
buf ( n17  , g16 );
buf ( n18  , g17 );
buf ( n19  , g18 );
buf ( n20  , g19 );
buf ( n21  , g20 );
buf ( n22  , g21 );
buf ( n23  , g22 );
buf ( n24  , g23 );
buf ( n25  , g24 );
buf ( n26  , g25 );
buf ( n27  , g26 );
buf ( n28  , g27 );
buf ( n29  , g28 );
buf ( n30  , g29 );
buf ( n31  , g30 );
buf ( n32  , g31 );
buf ( g32 , n33  );
buf ( g33 , n34  );
buf ( g34 , n35  );
buf ( g35 , n36  );
buf ( g36 , n37  );
buf ( g37 , n38  );
buf ( g38 , n39  );
buf ( g39 , n40  );
buf ( g40 , n41  );
buf ( g41 , n42  );
buf ( g42 , n43  );
buf ( g43 , n44  );
buf ( g44 , n45  );
buf ( g45 , n46  );
buf ( g46 , n47  );
buf ( g47 , n48  );
buf ( g48 , n49  );
buf ( g49 , n50  );
buf ( g50 , n51  );
buf ( g51 , n52  );
buf ( g52 , n53  );
buf ( g53 , n54  );
buf ( g54 , n55  );
buf ( g55 , n56  );
buf ( g56 , n57  );
buf ( g57 , n58  );
buf ( g58 , n59  );
buf ( g59 , n60  );
buf ( g60 , n61  );
buf ( g61 , n62  );
buf ( g62 , n63  );
buf ( g63 , n64  );
buf ( g64 , n65  );
buf ( g65 , n66  );
buf ( g66 , n67  );
buf ( g67 , n68  );
buf ( g68 , n69  );
buf ( g69 , n70  );
buf ( g70 , n71  );
buf ( g71 , n72  );
buf ( g72 , n73  );
buf ( g73 , n74  );
buf ( g74 , n75  );
buf ( g75 , n76  );
buf ( g76 , n77  );
buf ( g77 , n78  );
buf ( g78 , n79  );
buf ( g79 , n80  );
buf ( g80 , n81  );
buf ( g81 , n82  );
buf ( g82 , n83  );
buf ( g83 , n84  );
buf ( g84 , n85  );
buf ( g85 , n86  );
buf ( g86 , n87  );
buf ( g87 , n88  );
buf ( g88 , n89  );
buf ( g89 , n90  );
buf ( g90 , n91  );
buf ( g91 , n92  );
buf ( g92 , n93  );
buf ( g93 , n94  );
buf ( g94 , n95  );
buf ( g95 , n96  );
buf ( g96 , n97  );
buf ( g97 , n98  );
buf ( g98 , n99  );
buf ( g99 , n100  );
buf ( g100 , n101  );
buf ( g101 , n102  );
buf ( g102 , n103  );
buf ( g103 , n104  );
buf ( g104 , n105  );
buf ( g105 , n106  );
buf ( g106 , n107  );
buf ( g107 , n108  );
buf ( g108 , n109  );
buf ( g109 , n110  );
buf ( g110 , n111  );
buf ( g111 , n112  );
buf ( g112 , n113  );
buf ( g113 , n114  );
buf ( g114 , n115  );
buf ( g115 , n116  );
buf ( g116 , n117  );
buf ( g117 , n118  );
buf ( g118 , n119  );
buf ( g119 , n120  );
buf ( g120 , n121  );
buf ( g121 , n122  );
buf ( g122 , n123  );
buf ( g123 , n124  );
buf ( g124 , n125  );
buf ( g125 , n126  );
buf ( g126 , n127  );
buf ( g127 , n128  );
buf ( g128 , n129  );
buf ( g129 , n130  );
buf ( g130 , n131  );
buf ( g131 , n132  );
buf ( g132 , n133  );
buf ( g133 , n134  );
buf ( g134 , n135  );
buf ( g135 , n136  );
buf ( g136 , n137  );
buf ( g137 , n138  );
buf ( g138 , n139  );
buf ( g139 , n140  );
buf ( g140 , n141  );
buf ( g141 , n142  );
buf ( g142 , n143  );
buf ( g143 , n144  );
buf ( g144 , n145  );
buf ( g145 , n146  );
buf ( g146 , n147  );
buf ( g147 , n148  );
buf ( g148 , n149  );
buf ( g149 , n150  );
buf ( g150 , n151  );
buf ( g151 , n152  );
buf ( g152 , n153  );
buf ( g153 , n154  );
buf ( g154 , n155  );
buf ( g155 , n156  );
buf ( g156 , n157  );
buf ( g157 , n158  );
buf ( g158 , n159  );
buf ( g159 , n160  );
buf ( g160 , n161  );
buf ( n33 , 1'b0 );
buf ( n34 , 1'b0 );
buf ( n35 , 1'b0 );
buf ( n36 , 1'b0 );
buf ( n37 , 1'b0 );
buf ( n38 , 1'b0 );
buf ( n39 , 1'b0 );
buf ( n40 , 1'b0 );
buf ( n41 , 1'b0 );
buf ( n42 , 1'b0 );
buf ( n43 , 1'b0 );
buf ( n44 , 1'b0 );
buf ( n45 , 1'b0 );
buf ( n46 , 1'b0 );
buf ( n47 , 1'b0 );
buf ( n48 , 1'b0 );
buf ( n49 , 1'b0 );
buf ( n50 , 1'b0 );
buf ( n51 , 1'b0 );
buf ( n52 , 1'b0 );
buf ( n53 , 1'b0 );
buf ( n54 , 1'b0 );
buf ( n55 , 1'b0 );
buf ( n56 , 1'b0 );
buf ( n57 , 1'b0 );
buf ( n58 , 1'b0 );
buf ( n59 , 1'b0 );
buf ( n60 , 1'b0 );
buf ( n61 , 1'b0 );
buf ( n62 , 1'b0 );
buf ( n63 , 1'b0 );
buf ( n64 , 1'b0 );
buf ( n65 , 1'b0 );
buf ( n66 , 1'b0 );
buf ( n67 , 1'b0 );
buf ( n68 , 1'b0 );
buf ( n69 , 1'b0 );
buf ( n70 , 1'b0 );
buf ( n71 , 1'b0 );
buf ( n72 , 1'b0 );
buf ( n73 , 1'b0 );
buf ( n74 , 1'b0 );
buf ( n75 , 1'b0 );
buf ( n76 , 1'b0 );
buf ( n77 , 1'b0 );
buf ( n78 , 1'b0 );
buf ( n79 , 1'b0 );
buf ( n80 , 1'b0 );
buf ( n81 , 1'b0 );
buf ( n82 , n1630 );
buf ( n83 , n1635 );
buf ( n84 , n1919 );
buf ( n85 , n1274 );
buf ( n86 , n1280 );
buf ( n87 , n1286 );
buf ( n88 , n1925 );
buf ( n89 , n1675 );
buf ( n90 , n1805 );
buf ( n91 , n1698 );
buf ( n92 , n1811 );
buf ( n93 , n1846 );
buf ( n94 , n1860 );
buf ( n95 , n1871 );
buf ( n96 , n1907 );
buf ( n97 , n1913 );
buf ( n98 , 1'b0 );
buf ( n99 , 1'b0 );
buf ( n100 , 1'b0 );
buf ( n101 , 1'b0 );
buf ( n102 , 1'b0 );
buf ( n103 , 1'b0 );
buf ( n104 , 1'b0 );
buf ( n105 , 1'b0 );
buf ( n106 , 1'b0 );
buf ( n107 , 1'b0 );
buf ( n108 , 1'b0 );
buf ( n109 , 1'b0 );
buf ( n110 , 1'b0 );
buf ( n111 , 1'b0 );
buf ( n112 , 1'b0 );
buf ( n113 , 1'b0 );
buf ( n114 , 1'b0 );
buf ( n115 , 1'b0 );
buf ( n116 , 1'b0 );
buf ( n117 , 1'b0 );
buf ( n118 , 1'b0 );
buf ( n119 , 1'b0 );
buf ( n120 , 1'b0 );
buf ( n121 , 1'b0 );
buf ( n122 , 1'b0 );
buf ( n123 , 1'b0 );
buf ( n124 , 1'b0 );
buf ( n125 , 1'b0 );
buf ( n126 , 1'b0 );
buf ( n127 , 1'b0 );
buf ( n128 , 1'b0 );
buf ( n129 , 1'b0 );
buf ( n130 , 1'b0 );
buf ( n131 , 1'b0 );
buf ( n132 , 1'b0 );
buf ( n133 , 1'b0 );
buf ( n134 , 1'b0 );
buf ( n135 , 1'b0 );
buf ( n136 , 1'b0 );
buf ( n137 , 1'b0 );
buf ( n138 , 1'b0 );
buf ( n139 , 1'b0 );
buf ( n140 , 1'b0 );
buf ( n141 , 1'b0 );
buf ( n142 , 1'b0 );
buf ( n143 , 1'b0 );
buf ( n144 , 1'b0 );
buf ( n145 , 1'b0 );
buf ( n146 , n1761 );
buf ( n147 , n1755 );
buf ( n148 , n1771 );
buf ( n149 , n1571 );
buf ( n150 , n1665 );
buf ( n151 , n1641 );
buf ( n152 , n1766 );
buf ( n153 , n1777 );
buf ( n154 , n1924 );
buf ( n155 , n1796 );
buf ( n156 , n1822 );
buf ( n157 , n1837 );
buf ( n158 , n1880 );
buf ( n159 , n1890 );
buf ( n160 , n1899 );
buf ( n161 , n1918 );
nand ( n261 , n15 , n27 );
nand ( n262 , n14 , n28 );
xor ( n263 , n261 , n262 );
nand ( n264 , n16 , n26 );
and ( n265 , n263 , n264 );
and ( n266 , n261 , n262 );
or ( n267 , n265 , n266 );
not ( n268 , n267 );
nand ( n269 , n10 , n32 );
not ( n270 , n269 );
nand ( n271 , n12 , n30 );
not ( n272 , n271 );
and ( n273 , n11 , n31 );
and ( n274 , n272 , n273 );
not ( n275 , n272 );
nand ( n276 , n11 , n31 );
and ( n277 , n275 , n276 );
nor ( n278 , n274 , n277 );
not ( n279 , n278 );
or ( n280 , n270 , n279 );
or ( n281 , n269 , n278 );
nand ( n282 , n280 , n281 );
not ( n283 , n282 );
nand ( n284 , n11 , n32 );
nand ( n285 , n12 , n31 );
nor ( n286 , n284 , n285 );
not ( n287 , n286 );
nand ( n288 , n13 , n29 );
not ( n289 , n288 );
and ( n290 , n287 , n289 );
nand ( n291 , n11 , n32 );
nand ( n292 , n12 , n31 );
nor ( n293 , n291 , n292 );
and ( n294 , n293 , n288 );
nor ( n295 , n290 , n294 );
not ( n296 , n295 );
and ( n297 , n283 , n296 );
and ( n298 , n282 , n295 );
nor ( n299 , n297 , n298 );
not ( n300 , n299 );
xor ( n301 , n261 , n262 );
xor ( n302 , n301 , n264 );
not ( n303 , n302 );
or ( n304 , n300 , n303 );
and ( n305 , n13 , n30 );
not ( n306 , n291 );
not ( n307 , n292 );
not ( n308 , n307 );
or ( n309 , n306 , n308 );
not ( n310 , n285 );
or ( n311 , n284 , n310 );
nand ( n312 , n309 , n311 );
xor ( n313 , n305 , n312 );
nand ( n314 , n14 , n30 );
nand ( n315 , n13 , n31 );
nand ( n316 , n314 , n315 );
not ( n317 , n316 );
nand ( n318 , n12 , n32 );
not ( n319 , n318 );
not ( n320 , n319 );
or ( n321 , n317 , n320 );
nand ( n322 , n13 , n14 , n30 , n31 );
nand ( n323 , n321 , n322 );
and ( n324 , n313 , n323 );
and ( n325 , n305 , n312 );
or ( n326 , n324 , n325 );
buf ( n327 , n326 );
nand ( n328 , n304 , n327 );
not ( n329 , n302 );
nand ( n330 , n329 , n300 );
nand ( n331 , n328 , n330 );
not ( n332 , n331 );
or ( n333 , n268 , n332 );
or ( n334 , n331 , n267 );
nand ( n335 , n333 , n334 );
not ( n336 , n16 );
not ( n337 , n25 );
nor ( n338 , n336 , n337 );
not ( n339 , n338 );
nand ( n340 , n9 , n32 );
not ( n341 , n340 );
and ( n342 , n339 , n341 );
and ( n343 , n338 , n340 );
nor ( n344 , n342 , n343 );
buf ( n345 , n282 );
not ( n346 , n293 );
nand ( n347 , n346 , n288 );
and ( n348 , n345 , n347 );
not ( n349 , n293 );
nor ( n350 , n349 , n288 );
nor ( n351 , n348 , n350 );
xor ( n352 , n344 , n351 );
nand ( n353 , n10 , n32 );
nand ( n354 , n276 , n353 );
and ( n355 , n354 , n272 );
nor ( n356 , n353 , n276 );
nor ( n357 , n355 , n356 );
nand ( n358 , n14 , n27 );
nand ( n359 , n13 , n28 );
xor ( n360 , n358 , n359 );
nand ( n361 , n15 , n26 );
xor ( n362 , n360 , n361 );
xor ( n363 , n357 , n362 );
nand ( n364 , n11 , n30 );
nand ( n365 , n10 , n31 );
xor ( n366 , n364 , n365 );
nand ( n367 , n12 , n29 );
xor ( n368 , n366 , n367 );
xor ( n369 , n363 , n368 );
xor ( n370 , n352 , n369 );
not ( n371 , n370 );
and ( n372 , n335 , n371 );
not ( n373 , n335 );
and ( n374 , n373 , n370 );
nor ( n375 , n372 , n374 );
nand ( n376 , n14 , n29 );
not ( n377 , n376 );
and ( n378 , n15 , n28 );
nand ( n379 , n377 , n378 );
xor ( n380 , n302 , n326 );
xnor ( n381 , n380 , n299 );
xor ( n382 , n379 , n381 );
not ( n383 , n378 );
not ( n384 , n376 );
and ( n385 , n383 , n384 );
and ( n386 , n376 , n378 );
nor ( n387 , n385 , n386 );
buf ( n388 , n387 );
xor ( n389 , n305 , n312 );
xor ( n390 , n389 , n323 );
not ( n391 , n390 );
nand ( n392 , n388 , n391 );
nand ( n393 , n13 , n31 );
xor ( n394 , n393 , n314 );
and ( n395 , n394 , n318 );
not ( n396 , n394 );
and ( n397 , n396 , n319 );
nor ( n398 , n395 , n397 );
not ( n399 , n398 );
nand ( n400 , n15 , n29 );
not ( n401 , n400 );
or ( n402 , n399 , n401 );
nand ( n403 , n13 , n32 );
not ( n404 , n403 );
not ( n405 , n404 );
nand ( n406 , n15 , n30 );
not ( n407 , n406 );
not ( n408 , n407 );
or ( n409 , n405 , n408 );
not ( n410 , n403 );
not ( n411 , n406 );
or ( n412 , n410 , n411 );
and ( n413 , n14 , n31 );
nand ( n414 , n412 , n413 );
nand ( n415 , n409 , n414 );
buf ( n416 , n415 );
nand ( n417 , n402 , n416 );
nand ( n418 , n399 , n401 );
nand ( n419 , n417 , n418 );
buf ( n420 , n419 );
and ( n421 , n392 , n420 );
nor ( n422 , n391 , n388 );
nor ( n423 , n421 , n422 );
and ( n424 , n382 , n423 );
and ( n425 , n379 , n381 );
or ( n426 , n424 , n425 );
xor ( n427 , n375 , n426 );
not ( n428 , n427 );
xor ( n429 , n379 , n381 );
xor ( n430 , n429 , n423 );
and ( n431 , n16 , n28 );
not ( n432 , n431 );
not ( n433 , n432 );
xor ( n434 , n400 , n415 );
xnor ( n435 , n434 , n398 );
not ( n436 , n435 );
or ( n437 , n433 , n436 );
nand ( n438 , n16 , n29 );
not ( n439 , n438 );
nand ( n440 , n14 , n31 );
not ( n441 , n440 );
not ( n442 , n407 );
or ( n443 , n441 , n442 );
not ( n444 , n406 );
or ( n445 , n440 , n444 );
nand ( n446 , n443 , n445 );
and ( n447 , n446 , n404 );
not ( n448 , n446 );
not ( n449 , n404 );
and ( n450 , n448 , n449 );
nor ( n451 , n447 , n450 );
nor ( n452 , n439 , n451 );
nand ( n453 , n15 , n31 );
not ( n454 , n453 );
nand ( n455 , n16 , n30 );
not ( n456 , n455 );
or ( n457 , n454 , n456 );
nand ( n458 , n14 , n32 );
not ( n459 , n458 );
nand ( n460 , n457 , n459 );
not ( n461 , n455 );
not ( n462 , n453 );
nand ( n463 , n461 , n462 );
nand ( n464 , n460 , n463 );
not ( n465 , n464 );
or ( n466 , n452 , n465 );
nand ( n467 , n451 , n439 );
nand ( n468 , n466 , n467 );
nand ( n469 , n437 , n468 );
not ( n470 , n435 );
nand ( n471 , n470 , n431 );
nand ( n472 , n469 , n471 );
not ( n473 , n472 );
not ( n474 , n473 );
xor ( n475 , n387 , n419 );
xnor ( n476 , n475 , n390 );
nand ( n477 , n474 , n476 );
nand ( n478 , n430 , n477 );
not ( n479 , n478 );
not ( n480 , n16 );
not ( n481 , n27 );
nor ( n482 , n480 , n481 );
xor ( n483 , n431 , n435 );
not ( n484 , n468 );
xnor ( n485 , n483 , n484 );
xor ( n486 , n438 , n464 );
not ( n487 , n451 );
xnor ( n488 , n486 , n487 );
not ( n489 , n488 );
not ( n490 , n453 );
not ( n491 , n461 );
or ( n492 , n490 , n491 );
or ( n493 , n453 , n461 );
nand ( n494 , n492 , n493 );
and ( n495 , n494 , n459 );
not ( n496 , n494 );
and ( n497 , n496 , n458 );
nor ( n498 , n495 , n497 );
and ( n499 , n15 , n32 );
and ( n500 , n16 , n31 );
and ( n501 , n499 , n500 );
and ( n502 , n498 , n501 );
nand ( n503 , n489 , n502 );
nor ( n504 , n485 , n503 );
xor ( n505 , n482 , n504 );
not ( n506 , n473 );
not ( n507 , n476 );
or ( n508 , n506 , n507 );
or ( n509 , n473 , n476 );
nand ( n510 , n508 , n509 );
and ( n511 , n505 , n510 );
and ( n512 , n482 , n504 );
or ( n513 , n511 , n512 );
not ( n514 , n513 );
or ( n515 , n479 , n514 );
not ( n516 , n430 );
not ( n517 , n477 );
nand ( n518 , n516 , n517 );
nand ( n519 , n515 , n518 );
not ( n520 , n519 );
or ( n521 , n428 , n520 );
not ( n522 , n517 );
not ( n523 , n430 );
or ( n524 , n522 , n523 );
or ( n525 , n517 , n430 );
nand ( n526 , n524 , n525 );
not ( n527 , n526 );
not ( n528 , n513 );
or ( n529 , n527 , n528 );
not ( n530 , n518 );
nor ( n531 , n427 , n530 );
nand ( n532 , n529 , n531 );
nand ( n533 , n521 , n532 );
nand ( n534 , n6 , n21 );
nand ( n535 , n7 , n20 );
or ( n536 , n534 , n535 );
not ( n537 , n536 );
nand ( n538 , n8 , n18 );
nand ( n539 , n7 , n19 );
xor ( n540 , n538 , n539 );
nand ( n541 , n6 , n20 );
xor ( n542 , n540 , n541 );
nand ( n543 , n5 , n22 );
nand ( n544 , n4 , n23 );
not ( n545 , n544 );
nand ( n546 , n3 , n24 );
and ( n547 , n545 , n546 );
not ( n548 , n545 );
and ( n549 , n3 , n24 );
and ( n550 , n548 , n549 );
nor ( n551 , n547 , n550 );
xor ( n552 , n543 , n551 );
nand ( n553 , n6 , n22 );
nand ( n554 , n4 , n24 );
xor ( n555 , n553 , n554 );
nand ( n556 , n5 , n23 );
and ( n557 , n555 , n556 );
and ( n558 , n553 , n554 );
or ( n559 , n557 , n558 );
and ( n560 , n552 , n559 );
and ( n561 , n543 , n551 );
or ( n562 , n560 , n561 );
xor ( n563 , n542 , n562 );
nand ( n564 , n4 , n22 );
nand ( n565 , n3 , n23 );
xor ( n566 , n564 , n565 );
nand ( n567 , n2 , n24 );
xor ( n568 , n566 , n567 );
nand ( n569 , n5 , n21 );
not ( n570 , n569 );
not ( n571 , n545 );
nor ( n572 , n571 , n546 );
xor ( n573 , n570 , n572 );
xor ( n574 , n568 , n573 );
xor ( n575 , n563 , n574 );
not ( n576 , n575 );
or ( n577 , n537 , n576 );
not ( n578 , n535 );
not ( n579 , n578 );
not ( n580 , n534 );
and ( n581 , n579 , n580 );
and ( n582 , n534 , n578 );
nor ( n583 , n581 , n582 );
not ( n584 , n583 );
xor ( n585 , n543 , n551 );
xor ( n586 , n585 , n559 );
not ( n587 , n586 );
or ( n588 , n584 , n587 );
nand ( n589 , n7 , n21 );
not ( n590 , n589 );
not ( n591 , n590 );
nand ( n592 , n6 , n23 );
not ( n593 , n592 );
nand ( n594 , n7 , n22 );
not ( n595 , n594 );
or ( n596 , n593 , n595 );
and ( n597 , n5 , n24 );
nand ( n598 , n596 , n597 );
not ( n599 , n592 );
not ( n600 , n594 );
nand ( n601 , n599 , n600 );
nand ( n602 , n598 , n601 );
not ( n603 , n602 );
or ( n604 , n591 , n603 );
not ( n605 , n589 );
not ( n606 , n602 );
not ( n607 , n606 );
or ( n608 , n605 , n607 );
xor ( n609 , n553 , n554 );
xor ( n610 , n609 , n556 );
not ( n611 , n610 );
nand ( n612 , n608 , n611 );
nand ( n613 , n604 , n612 );
nand ( n614 , n588 , n613 );
not ( n615 , n583 );
not ( n616 , n586 );
nand ( n617 , n615 , n616 );
nand ( n618 , n614 , n617 );
nand ( n619 , n577 , n618 );
or ( n620 , n575 , n536 );
and ( n621 , n619 , n620 );
xor ( n622 , n538 , n539 );
and ( n623 , n622 , n541 );
and ( n624 , n538 , n539 );
or ( n625 , n623 , n624 );
xor ( n626 , n542 , n562 );
and ( n627 , n626 , n574 );
and ( n628 , n542 , n562 );
or ( n629 , n627 , n628 );
xor ( n630 , n625 , n629 );
nand ( n631 , n8 , n17 );
nand ( n632 , n1 , n24 );
xnor ( n633 , n631 , n632 );
not ( n634 , n568 );
not ( n635 , n572 );
nand ( n636 , n635 , n569 );
and ( n637 , n634 , n636 );
and ( n638 , n570 , n572 );
nor ( n639 , n637 , n638 );
xor ( n640 , n633 , n639 );
xor ( n641 , n564 , n565 );
and ( n642 , n641 , n567 );
and ( n643 , n564 , n565 );
or ( n644 , n642 , n643 );
nand ( n645 , n7 , n18 );
nand ( n646 , n6 , n19 );
xor ( n647 , n645 , n646 );
nand ( n648 , n5 , n20 );
xor ( n649 , n647 , n648 );
xor ( n650 , n644 , n649 );
nand ( n651 , n4 , n21 );
nand ( n652 , n3 , n22 );
xor ( n653 , n651 , n652 );
nand ( n654 , n2 , n23 );
xor ( n655 , n653 , n654 );
xor ( n656 , n650 , n655 );
xor ( n657 , n640 , n656 );
xor ( n658 , n630 , n657 );
xnor ( n659 , n621 , n658 );
not ( n660 , n659 );
not ( n661 , n660 );
nand ( n662 , n8 , n19 );
nand ( n663 , n8 , n20 );
not ( n664 , n663 );
and ( n665 , n8 , n21 );
nand ( n666 , n7 , n23 );
not ( n667 , n666 );
nand ( n668 , n8 , n22 );
not ( n669 , n668 );
or ( n670 , n667 , n669 );
nand ( n671 , n6 , n24 );
not ( n672 , n671 );
nand ( n673 , n670 , n672 );
or ( n674 , n666 , n668 );
nand ( n675 , n673 , n674 );
xor ( n676 , n665 , n675 );
nand ( n677 , n6 , n23 );
xor ( n678 , n677 , n600 );
xnor ( n679 , n678 , n597 );
and ( n680 , n676 , n679 );
and ( n681 , n665 , n675 );
or ( n682 , n680 , n681 );
xor ( n683 , n664 , n682 );
xor ( n684 , n590 , n606 );
xnor ( n685 , n684 , n610 );
xnor ( n686 , n683 , n685 );
xor ( n687 , n665 , n675 );
xor ( n688 , n687 , n679 );
and ( n689 , n8 , n23 );
not ( n690 , n689 );
nand ( n691 , n7 , n24 );
nor ( n692 , n690 , n691 );
not ( n693 , n692 );
xor ( n694 , n668 , n666 );
and ( n695 , n694 , n671 );
not ( n696 , n694 );
and ( n697 , n696 , n672 );
nor ( n698 , n695 , n697 );
nor ( n699 , n693 , n698 );
and ( n700 , n688 , n699 );
nand ( n701 , n686 , n700 );
xor ( n702 , n662 , n701 );
xor ( n703 , n583 , n613 );
xnor ( n704 , n703 , n586 );
not ( n705 , n664 );
nand ( n706 , n705 , n685 );
and ( n707 , n706 , n682 );
nor ( n708 , n685 , n663 );
nor ( n709 , n707 , n708 );
and ( n710 , n704 , n709 );
not ( n711 , n704 );
not ( n712 , n709 );
and ( n713 , n711 , n712 );
or ( n714 , n710 , n713 );
and ( n715 , n702 , n714 );
and ( n716 , n662 , n701 );
or ( n717 , n715 , n716 );
not ( n718 , n717 );
not ( n719 , n718 );
not ( n720 , n704 );
and ( n721 , n720 , n712 );
not ( n722 , n721 );
xor ( n723 , n536 , n618 );
xnor ( n724 , n723 , n575 );
nand ( n725 , n722 , n724 );
not ( n726 , n725 );
or ( n727 , n719 , n726 );
not ( n728 , n724 );
nand ( n729 , n728 , n721 );
nand ( n730 , n727 , n729 );
not ( n731 , n730 );
not ( n732 , n731 );
or ( n733 , n661 , n732 );
nand ( n734 , n730 , n659 );
nand ( n735 , n733 , n734 );
xor ( n736 , n533 , n735 );
not ( n737 , n513 );
xnor ( n738 , n737 , n526 );
not ( n739 , n738 );
xnor ( n740 , n502 , n488 );
not ( n741 , n689 );
not ( n742 , n691 );
and ( n743 , n741 , n742 );
and ( n744 , n691 , n689 );
nor ( n745 , n743 , n744 );
nand ( n746 , n16 , n32 );
not ( n747 , n746 );
nand ( n748 , n8 , n24 );
not ( n749 , n748 );
nand ( n750 , n747 , n749 );
nand ( n751 , n745 , n750 );
xor ( n752 , n499 , n500 );
and ( n753 , n751 , n752 );
nor ( n754 , n745 , n750 );
nor ( n755 , n753 , n754 );
not ( n756 , n755 );
xnor ( n757 , n501 , n498 );
not ( n758 , n757 );
or ( n759 , n756 , n758 );
xnor ( n760 , n692 , n698 );
nand ( n761 , n759 , n760 );
or ( n762 , n755 , n757 );
nand ( n763 , n761 , n762 );
nor ( n764 , n740 , n763 );
xnor ( n765 , n688 , n699 );
or ( n766 , n764 , n765 );
nand ( n767 , n740 , n763 );
nand ( n768 , n766 , n767 );
not ( n769 , n768 );
xnor ( n770 , n686 , n700 );
nand ( n771 , n769 , n770 );
not ( n772 , n503 );
not ( n773 , n772 );
buf ( n774 , n485 );
not ( n775 , n774 );
or ( n776 , n773 , n775 );
or ( n777 , n774 , n772 );
nand ( n778 , n776 , n777 );
and ( n779 , n771 , n778 );
nor ( n780 , n769 , n770 );
nor ( n781 , n779 , n780 );
not ( n782 , n781 );
xor ( n783 , n662 , n701 );
xor ( n784 , n783 , n714 );
not ( n785 , n784 );
or ( n786 , n782 , n785 );
xor ( n787 , n482 , n504 );
xor ( n788 , n787 , n510 );
nand ( n789 , n786 , n788 );
xor ( n790 , n721 , n724 );
xnor ( n791 , n790 , n717 );
not ( n792 , n784 );
not ( n793 , n781 );
nand ( n794 , n792 , n793 );
nand ( n795 , n789 , n791 , n794 );
not ( n796 , n795 );
or ( n797 , n739 , n796 );
not ( n798 , n794 );
not ( n799 , n789 );
or ( n800 , n798 , n799 );
not ( n801 , n791 );
nand ( n802 , n800 , n801 );
nand ( n803 , n797 , n802 );
xnor ( n804 , n736 , n803 );
not ( n805 , n804 );
not ( n806 , n805 );
nand ( n807 , n8 , n16 );
not ( n808 , n807 );
xnor ( n809 , n15 , n7 );
not ( n810 , n809 );
or ( n811 , n808 , n810 );
or ( n812 , n809 , n807 );
nand ( n813 , n811 , n812 );
nor ( n814 , n806 , n813 );
not ( n815 , n814 );
not ( n816 , n805 );
xor ( n817 , n31 , n23 );
not ( n818 , n24 );
not ( n819 , n32 );
nor ( n820 , n818 , n819 );
xor ( n821 , n817 , n820 );
nand ( n822 , n816 , n821 );
nand ( n823 , n815 , n822 );
and ( n824 , n819 , n24 );
and ( n825 , n818 , n32 );
nor ( n826 , n824 , n825 );
or ( n827 , n826 , n805 );
not ( n828 , n8 );
or ( n829 , n828 , n16 );
or ( n830 , n480 , n8 );
nand ( n831 , n829 , n830 );
nand ( n832 , n805 , n831 );
nand ( n833 , n827 , n832 );
nand ( n834 , n833 , n749 );
not ( n835 , n834 );
nand ( n836 , n823 , n835 );
buf ( n837 , n765 );
not ( n838 , n837 );
xor ( n839 , n13 , n5 );
xor ( n840 , n14 , n6 );
not ( n841 , n15 );
not ( n842 , n7 );
or ( n843 , n841 , n842 );
nor ( n844 , n7 , n15 );
or ( n845 , n844 , n807 );
nand ( n846 , n843 , n845 );
and ( n847 , n840 , n846 );
and ( n848 , n14 , n6 );
or ( n849 , n847 , n848 );
xor ( n850 , n839 , n849 );
not ( n851 , n850 );
not ( n852 , n804 );
not ( n853 , n852 );
or ( n854 , n851 , n853 );
not ( n855 , n30 );
not ( n856 , n22 );
or ( n857 , n855 , n856 );
or ( n858 , n22 , n30 );
xor ( n859 , n31 , n23 );
and ( n860 , n859 , n820 );
and ( n861 , n31 , n23 );
or ( n862 , n860 , n861 );
nand ( n863 , n858 , n862 );
nand ( n864 , n857 , n863 );
xnor ( n865 , n29 , n21 );
xnor ( n866 , n864 , n865 );
nand ( n867 , n866 , n804 );
nand ( n868 , n854 , n867 );
nand ( n869 , n838 , n868 );
xor ( n870 , n14 , n6 );
xor ( n871 , n870 , n846 );
not ( n872 , n871 );
not ( n873 , n816 );
not ( n874 , n873 );
or ( n875 , n872 , n874 );
xnor ( n876 , n30 , n22 );
or ( n877 , n862 , n876 );
not ( n878 , n877 );
nand ( n879 , n862 , n876 );
not ( n880 , n879 );
or ( n881 , n878 , n880 );
not ( n882 , n852 );
nand ( n883 , n881 , n882 );
nand ( n884 , n875 , n883 );
nand ( n885 , n884 , n760 );
and ( n886 , n836 , n869 , n885 );
not ( n887 , n886 );
xor ( n888 , n11 , n3 );
xor ( n889 , n12 , n4 );
xor ( n890 , n13 , n5 );
and ( n891 , n890 , n849 );
and ( n892 , n13 , n5 );
or ( n893 , n891 , n892 );
and ( n894 , n889 , n893 );
and ( n895 , n12 , n4 );
or ( n896 , n894 , n895 );
xor ( n897 , n888 , n896 );
not ( n898 , n897 );
not ( n899 , n852 );
or ( n900 , n898 , n899 );
not ( n901 , n882 );
xor ( n902 , n28 , n20 );
not ( n903 , n29 );
not ( n904 , n21 );
or ( n905 , n903 , n904 );
or ( n906 , n21 , n29 );
nand ( n907 , n906 , n864 );
nand ( n908 , n905 , n907 );
and ( n909 , n902 , n908 );
and ( n910 , n28 , n20 );
or ( n911 , n909 , n910 );
and ( n912 , n19 , n481 );
not ( n913 , n19 );
and ( n914 , n913 , n27 );
nor ( n915 , n912 , n914 );
xor ( n916 , n911 , n915 );
or ( n917 , n901 , n916 );
nand ( n918 , n900 , n917 );
not ( n919 , n918 );
buf ( n920 , n784 );
nand ( n921 , n919 , n920 );
xor ( n922 , n11 , n3 );
and ( n923 , n922 , n896 );
and ( n924 , n11 , n3 );
or ( n925 , n923 , n924 );
xnor ( n926 , n10 , n2 );
xnor ( n927 , n925 , n926 );
not ( n928 , n927 );
not ( n929 , n852 );
or ( n930 , n928 , n929 );
xor ( n931 , n26 , n18 );
not ( n932 , n27 );
not ( n933 , n19 );
or ( n934 , n932 , n933 );
or ( n935 , n19 , n27 );
nand ( n936 , n935 , n911 );
nand ( n937 , n934 , n936 );
xor ( n938 , n931 , n937 );
nand ( n939 , n882 , n938 );
nand ( n940 , n930 , n939 );
not ( n941 , n940 );
not ( n942 , n801 );
nand ( n943 , n941 , n942 );
nand ( n944 , n921 , n943 );
not ( n945 , n944 );
not ( n946 , n884 );
not ( n947 , n760 );
nand ( n948 , n946 , n947 );
not ( n949 , n948 );
and ( n950 , n949 , n869 );
xor ( n951 , n12 , n4 );
xor ( n952 , n951 , n893 );
not ( n953 , n952 );
not ( n954 , n852 );
or ( n955 , n953 , n954 );
xor ( n956 , n28 , n20 );
xor ( n957 , n956 , n908 );
nand ( n958 , n806 , n957 );
nand ( n959 , n955 , n958 );
not ( n960 , n959 );
buf ( n961 , n770 );
nand ( n962 , n960 , n961 );
not ( n963 , n868 );
nand ( n964 , n963 , n837 );
nand ( n965 , n962 , n964 );
nor ( n966 , n950 , n965 );
nand ( n967 , n887 , n945 , n966 );
not ( n968 , n967 );
not ( n969 , n968 );
xor ( n970 , n9 , n1 );
not ( n971 , n10 );
not ( n972 , n2 );
or ( n973 , n971 , n972 );
or ( n974 , n2 , n10 );
nand ( n975 , n974 , n925 );
nand ( n976 , n973 , n975 );
and ( n977 , n970 , n976 );
and ( n978 , n9 , n1 );
or ( n979 , n977 , n978 );
not ( n980 , n979 );
buf ( n981 , n816 );
not ( n982 , n981 );
not ( n983 , n982 );
or ( n984 , n980 , n983 );
not ( n985 , n981 );
xor ( n986 , n26 , n18 );
and ( n987 , n986 , n937 );
and ( n988 , n26 , n18 );
or ( n989 , n987 , n988 );
not ( n990 , n17 );
nand ( n991 , n990 , n337 );
and ( n992 , n989 , n991 );
and ( n993 , n17 , n25 );
nor ( n994 , n992 , n993 );
or ( n995 , n985 , n994 );
nand ( n996 , n984 , n995 );
not ( n997 , n730 );
not ( n998 , n660 );
or ( n999 , n997 , n998 );
or ( n1000 , n658 , n621 );
nand ( n1001 , n999 , n1000 );
xor ( n1002 , n633 , n639 );
and ( n1003 , n1002 , n656 );
and ( n1004 , n633 , n639 );
or ( n1005 , n1003 , n1004 );
or ( n1006 , n632 , n631 );
xor ( n1007 , n1005 , n1006 );
nand ( n1008 , n6 , n18 );
nand ( n1009 , n5 , n19 );
xnor ( n1010 , n1008 , n1009 );
xor ( n1011 , n651 , n652 );
and ( n1012 , n1011 , n654 );
and ( n1013 , n651 , n652 );
or ( n1014 , n1012 , n1013 );
xor ( n1015 , n1010 , n1014 );
nand ( n1016 , n4 , n20 );
nand ( n1017 , n3 , n21 );
xor ( n1018 , n1016 , n1017 );
nand ( n1019 , n2 , n22 );
xor ( n1020 , n1018 , n1019 );
xor ( n1021 , n1015 , n1020 );
nand ( n1022 , n7 , n17 );
nand ( n1023 , n1 , n23 );
xor ( n1024 , n1022 , n1023 );
xor ( n1025 , n645 , n646 );
and ( n1026 , n1025 , n648 );
and ( n1027 , n645 , n646 );
or ( n1028 , n1026 , n1027 );
xor ( n1029 , n1024 , n1028 );
xor ( n1030 , n1021 , n1029 );
xor ( n1031 , n644 , n649 );
and ( n1032 , n1031 , n655 );
and ( n1033 , n644 , n649 );
or ( n1034 , n1032 , n1033 );
xor ( n1035 , n1030 , n1034 );
xor ( n1036 , n1007 , n1035 );
xor ( n1037 , n625 , n629 );
and ( n1038 , n1037 , n657 );
and ( n1039 , n625 , n629 );
or ( n1040 , n1038 , n1039 );
xor ( n1041 , n1036 , n1040 );
xor ( n1042 , n1001 , n1041 );
nand ( n1043 , n996 , n1042 );
not ( n1044 , n1043 );
buf ( n1045 , n735 );
not ( n1046 , n1045 );
xor ( n1047 , n9 , n1 );
xor ( n1048 , n1047 , n976 );
and ( n1049 , n852 , n1048 );
not ( n1050 , n852 );
and ( n1051 , n337 , n17 );
and ( n1052 , n990 , n25 );
nor ( n1053 , n1051 , n1052 );
xnor ( n1054 , n1053 , n989 );
and ( n1055 , n1050 , n1054 );
or ( n1056 , n1049 , n1055 );
not ( n1057 , n1056 );
nand ( n1058 , n1046 , n1057 );
nor ( n1059 , n1044 , n1058 );
not ( n1060 , n1042 );
nor ( n1061 , n1059 , n1060 );
not ( n1062 , n1061 );
or ( n1063 , n969 , n1062 );
buf ( n1064 , n996 );
and ( n1065 , n1064 , n1058 );
nand ( n1066 , n968 , n1065 );
nand ( n1067 , n1063 , n1066 );
not ( n1068 , n1065 );
nand ( n1069 , n948 , n964 );
nor ( n1070 , n1069 , n944 );
not ( n1071 , n834 );
not ( n1072 , n823 );
not ( n1073 , n1072 );
or ( n1074 , n1071 , n1073 );
not ( n1075 , n745 );
nand ( n1076 , n1074 , n1075 );
not ( n1077 , n962 );
nor ( n1078 , n1076 , n1077 );
nand ( n1079 , n1070 , n1078 );
not ( n1080 , n1079 );
not ( n1081 , n1080 );
or ( n1082 , n1068 , n1081 );
buf ( n1083 , n959 );
not ( n1084 , n961 );
and ( n1085 , n1083 , n1084 );
not ( n1086 , n1085 );
not ( n1087 , n945 );
or ( n1088 , n1086 , n1087 );
not ( n1089 , n919 );
not ( n1090 , n920 );
and ( n1091 , n1089 , n1090 );
and ( n1092 , n1091 , n943 );
not ( n1093 , n801 );
nor ( n1094 , n1093 , n941 );
nor ( n1095 , n1092 , n1094 );
nand ( n1096 , n1088 , n1095 );
nand ( n1097 , n1096 , n1061 );
nand ( n1098 , n1082 , n1097 );
nor ( n1099 , n1067 , n1098 );
not ( n1100 , n1078 );
not ( n1101 , n1070 );
or ( n1102 , n1100 , n1101 );
nand ( n1103 , n1056 , n1045 );
and ( n1104 , n1103 , n1043 );
nand ( n1105 , n1102 , n1104 );
and ( n1106 , n1105 , n1061 );
not ( n1107 , n1096 );
not ( n1108 , n1065 );
or ( n1109 , n1107 , n1108 );
not ( n1110 , n1103 );
nand ( n1111 , n1064 , n1110 );
nand ( n1112 , n1109 , n1111 );
nor ( n1113 , n1106 , n1112 );
nand ( n1114 , n1099 , n1113 );
nand ( n1115 , n5 , n18 );
nand ( n1116 , n6 , n17 );
xor ( n1117 , n1115 , n1116 );
nand ( n1118 , n1 , n22 );
and ( n1119 , n1117 , n1118 );
and ( n1120 , n1115 , n1116 );
or ( n1121 , n1119 , n1120 );
nand ( n1122 , n3 , n19 );
nand ( n1123 , n2 , n20 );
xor ( n1124 , n1122 , n1123 );
nand ( n1125 , n3 , n20 );
nand ( n1126 , n4 , n19 );
xor ( n1127 , n1125 , n1126 );
nand ( n1128 , n2 , n21 );
and ( n1129 , n1127 , n1128 );
and ( n1130 , n1125 , n1126 );
or ( n1131 , n1129 , n1130 );
xor ( n1132 , n1124 , n1131 );
nand ( n1133 , n4 , n18 );
nand ( n1134 , n5 , n17 );
xor ( n1135 , n1133 , n1134 );
nand ( n1136 , n1 , n21 );
xor ( n1137 , n1135 , n1136 );
xor ( n1138 , n1132 , n1137 );
xor ( n1139 , n1016 , n1017 );
and ( n1140 , n1139 , n1019 );
and ( n1141 , n1016 , n1017 );
or ( n1142 , n1140 , n1141 );
or ( n1143 , n1009 , n1008 );
xor ( n1144 , n1142 , n1143 );
xor ( n1145 , n1125 , n1126 );
xor ( n1146 , n1145 , n1128 );
and ( n1147 , n1144 , n1146 );
and ( n1148 , n1142 , n1143 );
or ( n1149 , n1147 , n1148 );
xor ( n1150 , n1138 , n1149 );
and ( n1151 , n1121 , n1150 );
xor ( n1152 , n1142 , n1143 );
xor ( n1153 , n1152 , n1146 );
xor ( n1154 , n1115 , n1116 );
xor ( n1155 , n1154 , n1118 );
xor ( n1156 , n1153 , n1155 );
xor ( n1157 , n1010 , n1014 );
and ( n1158 , n1157 , n1020 );
and ( n1159 , n1010 , n1014 );
or ( n1160 , n1158 , n1159 );
and ( n1161 , n1156 , n1160 );
and ( n1162 , n1153 , n1155 );
or ( n1163 , n1161 , n1162 );
xor ( n1164 , n1132 , n1137 );
xor ( n1165 , n1164 , n1149 );
and ( n1166 , n1163 , n1165 );
and ( n1167 , n1121 , n1163 );
or ( n1168 , n1151 , n1166 , n1167 );
nand ( n1169 , n2 , n19 );
nand ( n1170 , n3 , n18 );
xor ( n1171 , n1169 , n1170 );
nand ( n1172 , n4 , n17 );
xor ( n1173 , n1171 , n1172 );
xor ( n1174 , n1133 , n1134 );
and ( n1175 , n1174 , n1136 );
and ( n1176 , n1133 , n1134 );
or ( n1177 , n1175 , n1176 );
xor ( n1178 , n1173 , n1177 );
xor ( n1179 , n1122 , n1123 );
and ( n1180 , n1179 , n1131 );
and ( n1181 , n1122 , n1123 );
or ( n1182 , n1180 , n1181 );
xor ( n1183 , n1178 , n1182 );
nand ( n1184 , n1 , n20 );
xor ( n1185 , n1132 , n1137 );
and ( n1186 , n1185 , n1149 );
and ( n1187 , n1132 , n1137 );
or ( n1188 , n1186 , n1187 );
xor ( n1189 , n1184 , n1188 );
xor ( n1190 , n1183 , n1189 );
xor ( n1191 , n1168 , n1190 );
xor ( n1192 , n1153 , n1155 );
xor ( n1193 , n1192 , n1160 );
xor ( n1194 , n1022 , n1023 );
and ( n1195 , n1194 , n1028 );
and ( n1196 , n1022 , n1023 );
or ( n1197 , n1195 , n1196 );
xor ( n1198 , n1193 , n1197 );
xor ( n1199 , n1021 , n1029 );
and ( n1200 , n1199 , n1034 );
and ( n1201 , n1021 , n1029 );
or ( n1202 , n1200 , n1201 );
and ( n1203 , n1198 , n1202 );
and ( n1204 , n1193 , n1197 );
or ( n1205 , n1203 , n1204 );
xor ( n1206 , n1132 , n1137 );
xor ( n1207 , n1206 , n1149 );
xor ( n1208 , n1121 , n1163 );
xor ( n1209 , n1207 , n1208 );
xor ( n1210 , n1205 , n1209 );
not ( n1211 , n1210 );
xor ( n1212 , n1193 , n1197 );
xor ( n1213 , n1212 , n1202 );
xor ( n1214 , n1005 , n1006 );
and ( n1215 , n1214 , n1035 );
and ( n1216 , n1005 , n1006 );
or ( n1217 , n1215 , n1216 );
xor ( n1218 , n1213 , n1217 );
not ( n1219 , n1218 );
not ( n1220 , n1041 );
not ( n1221 , n1001 );
or ( n1222 , n1220 , n1221 );
or ( n1223 , n1036 , n1040 );
nand ( n1224 , n1222 , n1223 );
not ( n1225 , n1224 );
or ( n1226 , n1219 , n1225 );
or ( n1227 , n1213 , n1217 );
nand ( n1228 , n1226 , n1227 );
not ( n1229 , n1228 );
or ( n1230 , n1211 , n1229 );
or ( n1231 , n1205 , n1209 );
nand ( n1232 , n1230 , n1231 );
xor ( n1233 , n1191 , n1232 );
xor ( n1234 , n1228 , n1210 );
xor ( n1235 , n1224 , n1218 );
and ( n1236 , n1234 , n1235 );
nand ( n1237 , n1233 , n1236 );
not ( n1238 , n1237 );
nand ( n1239 , n1114 , n1238 );
xor ( n1240 , n1173 , n1177 );
xor ( n1241 , n1240 , n1182 );
and ( n1242 , n1184 , n1241 );
xor ( n1243 , n1173 , n1177 );
xor ( n1244 , n1243 , n1182 );
and ( n1245 , n1188 , n1244 );
and ( n1246 , n1184 , n1188 );
or ( n1247 , n1242 , n1245 , n1246 );
nand ( n1248 , n3 , n17 );
nand ( n1249 , n2 , n18 );
xor ( n1250 , n1248 , n1249 );
xor ( n1251 , n1169 , n1170 );
and ( n1252 , n1251 , n1172 );
and ( n1253 , n1169 , n1170 );
or ( n1254 , n1252 , n1253 );
xor ( n1255 , n1250 , n1254 );
nand ( n1256 , n1 , n19 );
xor ( n1257 , n1173 , n1177 );
and ( n1258 , n1257 , n1182 );
and ( n1259 , n1173 , n1177 );
or ( n1260 , n1258 , n1259 );
xor ( n1261 , n1256 , n1260 );
xor ( n1262 , n1255 , n1261 );
xor ( n1263 , n1247 , n1262 );
not ( n1264 , n1191 );
not ( n1265 , n1232 );
or ( n1266 , n1264 , n1265 );
or ( n1267 , n1168 , n1190 );
nand ( n1268 , n1266 , n1267 );
xor ( n1269 , n1263 , n1268 );
not ( n1270 , n1269 );
and ( n1271 , n1239 , n1270 );
not ( n1272 , n1239 );
and ( n1273 , n1272 , n1269 );
nor ( n1274 , n1271 , n1273 );
nand ( n1275 , n1114 , n1236 );
not ( n1276 , n1233 );
and ( n1277 , n1275 , n1276 );
not ( n1278 , n1275 );
and ( n1279 , n1278 , n1233 );
nor ( n1280 , n1277 , n1279 );
nand ( n1281 , n1114 , n1235 );
not ( n1282 , n1234 );
and ( n1283 , n1281 , n1282 );
not ( n1284 , n1281 );
and ( n1285 , n1284 , n1234 );
nor ( n1286 , n1283 , n1285 );
buf ( n1287 , n533 );
nand ( n1288 , n1056 , n1287 );
not ( n1289 , n1288 );
nor ( n1290 , n918 , n788 );
buf ( n1291 , n738 );
nor ( n1292 , n940 , n1291 );
nor ( n1293 , n1290 , n1292 );
not ( n1294 , n1293 );
buf ( n1295 , n740 );
nand ( n1296 , n868 , n1295 );
buf ( n1297 , n778 );
nor ( n1298 , n959 , n1297 );
or ( n1299 , n1296 , n1298 );
nand ( n1300 , n959 , n1297 );
nand ( n1301 , n1299 , n1300 );
not ( n1302 , n1301 );
or ( n1303 , n1294 , n1302 );
nand ( n1304 , n918 , n788 );
not ( n1305 , n1304 );
not ( n1306 , n1292 );
and ( n1307 , n1305 , n1306 );
and ( n1308 , n940 , n1291 );
nor ( n1309 , n1307 , n1308 );
nand ( n1310 , n1303 , n1309 );
not ( n1311 , n1287 );
nand ( n1312 , n1311 , n1057 );
nand ( n1313 , n1310 , n1312 );
not ( n1314 , n1313 );
or ( n1315 , n1289 , n1314 );
not ( n1316 , n427 );
buf ( n1317 , n519 );
nand ( n1318 , n1316 , n1317 );
not ( n1319 , n375 );
or ( n1320 , n1319 , n426 );
nand ( n1321 , n1318 , n1320 );
not ( n1322 , n340 );
nand ( n1323 , n1322 , n338 );
xor ( n1324 , n344 , n351 );
and ( n1325 , n1324 , n369 );
and ( n1326 , n344 , n351 );
or ( n1327 , n1325 , n1326 );
xor ( n1328 , n1323 , n1327 );
nand ( n1329 , n15 , n25 );
nand ( n1330 , n9 , n31 );
xor ( n1331 , n1329 , n1330 );
xor ( n1332 , n358 , n359 );
and ( n1333 , n1332 , n361 );
and ( n1334 , n358 , n359 );
or ( n1335 , n1333 , n1334 );
xor ( n1336 , n1331 , n1335 );
and ( n1337 , n14 , n26 );
not ( n1338 , n1337 );
nand ( n1339 , n13 , n27 );
not ( n1340 , n1339 );
and ( n1341 , n1338 , n1340 );
and ( n1342 , n1337 , n1339 );
nor ( n1343 , n1341 , n1342 );
xor ( n1344 , n364 , n365 );
and ( n1345 , n1344 , n367 );
and ( n1346 , n364 , n365 );
or ( n1347 , n1345 , n1346 );
xor ( n1348 , n1343 , n1347 );
nand ( n1349 , n11 , n29 );
nand ( n1350 , n10 , n30 );
xor ( n1351 , n1349 , n1350 );
nand ( n1352 , n12 , n28 );
xor ( n1353 , n1351 , n1352 );
xor ( n1354 , n1348 , n1353 );
xor ( n1355 , n1336 , n1354 );
xor ( n1356 , n357 , n362 );
and ( n1357 , n1356 , n368 );
and ( n1358 , n357 , n362 );
or ( n1359 , n1357 , n1358 );
xor ( n1360 , n1355 , n1359 );
xor ( n1361 , n1328 , n1360 );
not ( n1362 , n370 );
not ( n1363 , n267 );
and ( n1364 , n1362 , n1363 );
nand ( n1365 , n370 , n267 );
and ( n1366 , n1365 , n331 );
nor ( n1367 , n1364 , n1366 );
xor ( n1368 , n1361 , n1367 );
xor ( n1369 , n1321 , n1368 );
nor ( n1370 , n1369 , n996 );
not ( n1371 , n1370 );
nand ( n1372 , n1315 , n1371 );
buf ( n1373 , n757 );
nand ( n1374 , n946 , n1373 );
not ( n1375 , n1374 );
not ( n1376 , n746 );
nand ( n1377 , n1376 , n833 );
not ( n1378 , n752 );
nand ( n1379 , n822 , n1378 );
nor ( n1380 , n1379 , n814 );
or ( n1381 , n1377 , n1380 );
nand ( n1382 , n823 , n752 );
nand ( n1383 , n1381 , n1382 );
not ( n1384 , n1383 );
or ( n1385 , n1375 , n1384 );
not ( n1386 , n946 );
not ( n1387 , n1373 );
nand ( n1388 , n1386 , n1387 );
nand ( n1389 , n1385 , n1388 );
not ( n1390 , n1293 );
not ( n1391 , n1298 );
or ( n1392 , n868 , n1295 );
nand ( n1393 , n1391 , n1392 );
nor ( n1394 , n1390 , n1393 );
not ( n1395 , n1312 );
nor ( n1396 , n1395 , n1370 );
nand ( n1397 , n1389 , n1394 , n1396 );
not ( n1398 , n1369 );
not ( n1399 , n1398 );
nand ( n1400 , n1399 , n1064 );
and ( n1401 , n1372 , n1397 , n1400 );
not ( n1402 , n1401 );
nand ( n1403 , n11 , n27 );
nand ( n1404 , n10 , n28 );
xor ( n1405 , n1403 , n1404 );
nand ( n1406 , n11 , n28 );
nand ( n1407 , n10 , n29 );
xor ( n1408 , n1406 , n1407 );
nand ( n1409 , n12 , n27 );
and ( n1410 , n1408 , n1409 );
and ( n1411 , n1406 , n1407 );
or ( n1412 , n1410 , n1411 );
xor ( n1413 , n1405 , n1412 );
nand ( n1414 , n9 , n29 );
nand ( n1415 , n12 , n26 );
xor ( n1416 , n1414 , n1415 );
nand ( n1417 , n13 , n25 );
xor ( n1418 , n1416 , n1417 );
xor ( n1419 , n1413 , n1418 );
not ( n1420 , n1339 );
nand ( n1421 , n1420 , n1337 );
xor ( n1422 , n1349 , n1350 );
and ( n1423 , n1422 , n1352 );
and ( n1424 , n1349 , n1350 );
or ( n1425 , n1423 , n1424 );
xor ( n1426 , n1421 , n1425 );
xor ( n1427 , n1406 , n1407 );
xor ( n1428 , n1427 , n1409 );
and ( n1429 , n1426 , n1428 );
and ( n1430 , n1421 , n1425 );
or ( n1431 , n1429 , n1430 );
xor ( n1432 , n1419 , n1431 );
nand ( n1433 , n9 , n30 );
nand ( n1434 , n13 , n26 );
xor ( n1435 , n1433 , n1434 );
nand ( n1436 , n14 , n25 );
and ( n1437 , n1435 , n1436 );
and ( n1438 , n1433 , n1434 );
or ( n1439 , n1437 , n1438 );
xor ( n1440 , n1433 , n1434 );
xor ( n1441 , n1440 , n1436 );
xor ( n1442 , n1421 , n1425 );
xor ( n1443 , n1442 , n1428 );
xor ( n1444 , n1441 , n1443 );
xor ( n1445 , n1343 , n1347 );
and ( n1446 , n1445 , n1353 );
and ( n1447 , n1343 , n1347 );
or ( n1448 , n1446 , n1447 );
and ( n1449 , n1444 , n1448 );
and ( n1450 , n1441 , n1443 );
or ( n1451 , n1449 , n1450 );
xor ( n1452 , n1439 , n1451 );
xor ( n1453 , n1432 , n1452 );
xor ( n1454 , n1329 , n1330 );
and ( n1455 , n1454 , n1335 );
and ( n1456 , n1329 , n1330 );
or ( n1457 , n1455 , n1456 );
xor ( n1458 , n1441 , n1443 );
xor ( n1459 , n1458 , n1448 );
and ( n1460 , n1457 , n1459 );
xor ( n1461 , n1336 , n1354 );
and ( n1462 , n1461 , n1359 );
and ( n1463 , n1336 , n1354 );
or ( n1464 , n1462 , n1463 );
xor ( n1465 , n1441 , n1443 );
xor ( n1466 , n1465 , n1448 );
and ( n1467 , n1464 , n1466 );
and ( n1468 , n1457 , n1464 );
or ( n1469 , n1460 , n1467 , n1468 );
xor ( n1470 , n1453 , n1469 );
not ( n1471 , n1470 );
xor ( n1472 , n1441 , n1443 );
xor ( n1473 , n1472 , n1448 );
xor ( n1474 , n1457 , n1464 );
xor ( n1475 , n1473 , n1474 );
xor ( n1476 , n1323 , n1327 );
and ( n1477 , n1476 , n1360 );
and ( n1478 , n1323 , n1327 );
or ( n1479 , n1477 , n1478 );
xor ( n1480 , n1475 , n1479 );
not ( n1481 , n1480 );
not ( n1482 , n1368 );
not ( n1483 , n1321 );
or ( n1484 , n1482 , n1483 );
or ( n1485 , n1361 , n1367 );
nand ( n1486 , n1484 , n1485 );
not ( n1487 , n1486 );
or ( n1488 , n1481 , n1487 );
or ( n1489 , n1479 , n1475 );
nand ( n1490 , n1488 , n1489 );
not ( n1491 , n1490 );
or ( n1492 , n1471 , n1491 );
or ( n1493 , n1469 , n1453 );
nand ( n1494 , n1492 , n1493 );
xor ( n1495 , n1413 , n1418 );
xor ( n1496 , n1495 , n1431 );
and ( n1497 , n1439 , n1496 );
xor ( n1498 , n1413 , n1418 );
xor ( n1499 , n1498 , n1431 );
and ( n1500 , n1451 , n1499 );
and ( n1501 , n1439 , n1451 );
or ( n1502 , n1497 , n1500 , n1501 );
nand ( n1503 , n10 , n27 );
nand ( n1504 , n11 , n26 );
xor ( n1505 , n1503 , n1504 );
nand ( n1506 , n12 , n25 );
xor ( n1507 , n1505 , n1506 );
xor ( n1508 , n1414 , n1415 );
and ( n1509 , n1508 , n1417 );
and ( n1510 , n1414 , n1415 );
or ( n1511 , n1509 , n1510 );
xor ( n1512 , n1507 , n1511 );
xor ( n1513 , n1403 , n1404 );
and ( n1514 , n1513 , n1412 );
and ( n1515 , n1403 , n1404 );
or ( n1516 , n1514 , n1515 );
xor ( n1517 , n1512 , n1516 );
nand ( n1518 , n9 , n28 );
xor ( n1519 , n1413 , n1418 );
and ( n1520 , n1519 , n1431 );
and ( n1521 , n1413 , n1418 );
or ( n1522 , n1520 , n1521 );
xor ( n1523 , n1518 , n1522 );
xor ( n1524 , n1517 , n1523 );
xor ( n1525 , n1502 , n1524 );
and ( n1526 , n1494 , n1525 );
not ( n1527 , n1494 );
not ( n1528 , n1525 );
and ( n1529 , n1527 , n1528 );
nor ( n1530 , n1526 , n1529 );
xor ( n1531 , n1470 , n1490 );
xor ( n1532 , n1486 , n1480 );
and ( n1533 , n1531 , n1532 );
nand ( n1534 , n1530 , n1533 );
not ( n1535 , n1534 );
nand ( n1536 , n1402 , n1535 );
xor ( n1537 , n1507 , n1511 );
xor ( n1538 , n1537 , n1516 );
and ( n1539 , n1518 , n1538 );
xor ( n1540 , n1507 , n1511 );
xor ( n1541 , n1540 , n1516 );
and ( n1542 , n1522 , n1541 );
and ( n1543 , n1518 , n1522 );
or ( n1544 , n1539 , n1542 , n1543 );
nand ( n1545 , n11 , n25 );
nand ( n1546 , n10 , n26 );
xor ( n1547 , n1545 , n1546 );
xor ( n1548 , n1503 , n1504 );
and ( n1549 , n1548 , n1506 );
and ( n1550 , n1503 , n1504 );
or ( n1551 , n1549 , n1550 );
xor ( n1552 , n1547 , n1551 );
nand ( n1553 , n9 , n27 );
xor ( n1554 , n1507 , n1511 );
and ( n1555 , n1554 , n1516 );
and ( n1556 , n1507 , n1511 );
or ( n1557 , n1555 , n1556 );
xor ( n1558 , n1553 , n1557 );
xor ( n1559 , n1552 , n1558 );
xor ( n1560 , n1544 , n1559 );
not ( n1561 , n1525 );
not ( n1562 , n1494 );
or ( n1563 , n1561 , n1562 );
or ( n1564 , n1502 , n1524 );
nand ( n1565 , n1563 , n1564 );
xor ( n1566 , n1560 , n1565 );
not ( n1567 , n1566 );
and ( n1568 , n1536 , n1567 );
not ( n1569 , n1536 );
and ( n1570 , n1569 , n1566 );
nor ( n1571 , n1568 , n1570 );
not ( n1572 , n1064 );
not ( n1573 , n1042 );
and ( n1574 , n1572 , n1573 );
nor ( n1575 , n1574 , n1237 );
and ( n1576 , n1575 , n1269 , n1058 );
not ( n1577 , n1576 );
not ( n1578 , n1096 );
nand ( n1579 , n1079 , n967 , n1578 );
not ( n1580 , n1579 );
or ( n1581 , n1577 , n1580 );
nand ( n1582 , n1044 , n1238 );
not ( n1583 , n1582 );
nand ( n1584 , n1575 , n1110 );
not ( n1585 , n1584 );
or ( n1586 , n1583 , n1585 );
nand ( n1587 , n1586 , n1269 );
nand ( n1588 , n1581 , n1587 );
not ( n1589 , n1263 );
not ( n1590 , n1268 );
or ( n1591 , n1589 , n1590 );
or ( n1592 , n1247 , n1262 );
nand ( n1593 , n1591 , n1592 );
xor ( n1594 , n1248 , n1249 );
xor ( n1595 , n1594 , n1254 );
and ( n1596 , n1256 , n1595 );
xor ( n1597 , n1248 , n1249 );
xor ( n1598 , n1597 , n1254 );
and ( n1599 , n1260 , n1598 );
and ( n1600 , n1256 , n1260 );
or ( n1601 , n1596 , n1599 , n1600 );
nand ( n1602 , n2 , n17 );
nand ( n1603 , n1 , n18 );
xor ( n1604 , n1602 , n1603 );
xor ( n1605 , n1248 , n1249 );
and ( n1606 , n1605 , n1254 );
and ( n1607 , n1248 , n1249 );
or ( n1608 , n1606 , n1607 );
xor ( n1609 , n1604 , n1608 );
xor ( n1610 , n1601 , n1609 );
xor ( n1611 , n1593 , n1610 );
nand ( n1612 , n1588 , n1611 );
not ( n1613 , n1610 );
not ( n1614 , n1593 );
or ( n1615 , n1613 , n1614 );
or ( n1616 , n1601 , n1609 );
nand ( n1617 , n1615 , n1616 );
xor ( n1618 , n1602 , n1603 );
and ( n1619 , n1618 , n1608 );
and ( n1620 , n1602 , n1603 );
or ( n1621 , n1619 , n1620 );
nand ( n1622 , n1 , n17 );
xnor ( n1623 , n1621 , n1622 );
xor ( n1624 , n1617 , n1623 );
or ( n1625 , n1612 , n1624 );
not ( n1626 , n1623 );
and ( n1627 , n1617 , n1626 );
nor ( n1628 , n1621 , n1622 );
nor ( n1629 , n1627 , n1628 );
nand ( n1630 , n1625 , n1629 );
and ( n1631 , n1612 , n1624 );
not ( n1632 , n1612 );
not ( n1633 , n1624 );
and ( n1634 , n1632 , n1633 );
nor ( n1635 , n1631 , n1634 );
nand ( n1636 , n1402 , n1532 );
not ( n1637 , n1531 );
and ( n1638 , n1636 , n1637 );
not ( n1639 , n1636 );
and ( n1640 , n1639 , n1531 );
nor ( n1641 , n1638 , n1640 );
not ( n1642 , n1533 );
nor ( n1643 , n1642 , n1370 );
not ( n1644 , n1643 );
not ( n1645 , n1312 );
not ( n1646 , n1389 );
not ( n1647 , n1394 );
or ( n1648 , n1646 , n1647 );
not ( n1649 , n1310 );
nand ( n1650 , n1648 , n1649 );
not ( n1651 , n1650 );
or ( n1652 , n1645 , n1651 );
not ( n1653 , n1288 );
not ( n1654 , n1653 );
nand ( n1655 , n1652 , n1654 );
not ( n1656 , n1655 );
or ( n1657 , n1644 , n1656 );
not ( n1658 , n1400 );
nand ( n1659 , n1658 , n1533 );
nand ( n1660 , n1657 , n1659 );
and ( n1661 , n1660 , n1530 );
not ( n1662 , n1660 );
not ( n1663 , n1530 );
and ( n1664 , n1662 , n1663 );
nor ( n1665 , n1661 , n1664 );
not ( n1666 , n1058 );
not ( n1667 , n1579 );
or ( n1668 , n1666 , n1667 );
nand ( n1669 , n1668 , n1103 );
xor ( n1670 , n1060 , n1064 );
not ( n1671 , n1670 );
and ( n1672 , n1669 , n1671 );
not ( n1673 , n1669 );
and ( n1674 , n1673 , n1670 );
nor ( n1675 , n1672 , n1674 );
not ( n1676 , n1069 );
nand ( n1677 , n1076 , n836 );
nand ( n1678 , n1676 , n1677 );
not ( n1679 , n885 );
nand ( n1680 , n1679 , n964 );
and ( n1681 , n1678 , n1680 , n869 );
not ( n1682 , n1681 );
not ( n1683 , n1077 );
and ( n1684 , n1682 , n1683 );
nor ( n1685 , n1684 , n1085 );
not ( n1686 , n921 );
or ( n1687 , n1685 , n1686 );
not ( n1688 , n1091 );
nand ( n1689 , n1687 , n1688 );
and ( n1690 , n801 , n941 );
not ( n1691 , n801 );
and ( n1692 , n1691 , n940 );
nor ( n1693 , n1690 , n1692 );
not ( n1694 , n1693 );
and ( n1695 , n1689 , n1694 );
not ( n1696 , n1689 );
and ( n1697 , n1696 , n1693 );
nor ( n1698 , n1695 , n1697 );
nor ( n1699 , n1534 , n1370 );
and ( n1700 , n1699 , n1566 , n1312 );
not ( n1701 , n1700 );
not ( n1702 , n1650 );
or ( n1703 , n1701 , n1702 );
nand ( n1704 , n1658 , n1535 );
not ( n1705 , n1704 );
nand ( n1706 , n1699 , n1653 );
not ( n1707 , n1706 );
or ( n1708 , n1705 , n1707 );
nand ( n1709 , n1708 , n1566 );
nand ( n1710 , n1703 , n1709 );
not ( n1711 , n1565 );
not ( n1712 , n1560 );
or ( n1713 , n1711 , n1712 );
or ( n1714 , n1544 , n1559 );
nand ( n1715 , n1713 , n1714 );
xor ( n1716 , n1545 , n1546 );
xor ( n1717 , n1716 , n1551 );
and ( n1718 , n1553 , n1717 );
xor ( n1719 , n1545 , n1546 );
xor ( n1720 , n1719 , n1551 );
and ( n1721 , n1557 , n1720 );
and ( n1722 , n1553 , n1557 );
or ( n1723 , n1718 , n1721 , n1722 );
nand ( n1724 , n10 , n25 );
nand ( n1725 , n9 , n26 );
xor ( n1726 , n1724 , n1725 );
xor ( n1727 , n1545 , n1546 );
and ( n1728 , n1727 , n1551 );
and ( n1729 , n1545 , n1546 );
or ( n1730 , n1728 , n1729 );
xor ( n1731 , n1726 , n1730 );
xor ( n1732 , n1723 , n1731 );
xor ( n1733 , n1715 , n1732 );
nand ( n1734 , n1710 , n1733 );
not ( n1735 , n1732 );
not ( n1736 , n1715 );
or ( n1737 , n1735 , n1736 );
or ( n1738 , n1723 , n1731 );
nand ( n1739 , n1737 , n1738 );
not ( n1740 , n1739 );
xor ( n1741 , n1724 , n1725 );
and ( n1742 , n1741 , n1730 );
and ( n1743 , n1724 , n1725 );
or ( n1744 , n1742 , n1743 );
nand ( n1745 , n9 , n25 );
xnor ( n1746 , n1744 , n1745 );
not ( n1747 , n1746 );
and ( n1748 , n1740 , n1747 );
and ( n1749 , n1739 , n1746 );
nor ( n1750 , n1748 , n1749 );
and ( n1751 , n1734 , n1750 );
not ( n1752 , n1734 );
not ( n1753 , n1750 );
and ( n1754 , n1752 , n1753 );
nor ( n1755 , n1751 , n1754 );
or ( n1756 , n1734 , n1750 );
not ( n1757 , n1746 );
and ( n1758 , n1739 , n1757 );
nor ( n1759 , n1744 , n1745 );
nor ( n1760 , n1758 , n1759 );
nand ( n1761 , n1756 , n1760 );
not ( n1762 , n1532 );
not ( n1763 , n1401 );
or ( n1764 , n1762 , n1763 );
or ( n1765 , n1401 , n1532 );
nand ( n1766 , n1764 , n1765 );
and ( n1767 , n1710 , n1733 );
not ( n1768 , n1710 );
not ( n1769 , n1733 );
and ( n1770 , n1768 , n1769 );
nor ( n1771 , n1767 , n1770 );
xor ( n1772 , n1398 , n1064 );
not ( n1773 , n1772 );
and ( n1774 , n1655 , n1773 );
not ( n1775 , n1655 );
and ( n1776 , n1775 , n1772 );
nor ( n1777 , n1774 , n1776 );
not ( n1778 , n1290 );
not ( n1779 , n1778 );
not ( n1780 , n1383 );
not ( n1781 , n1374 );
nor ( n1782 , n1781 , n1393 );
not ( n1783 , n1782 );
or ( n1784 , n1780 , n1783 );
nor ( n1785 , n1388 , n1393 );
nor ( n1786 , n1785 , n1301 );
nand ( n1787 , n1784 , n1786 );
not ( n1788 , n1787 );
or ( n1789 , n1779 , n1788 );
nand ( n1790 , n1789 , n1304 );
xor ( n1791 , n941 , n1291 );
not ( n1792 , n1791 );
and ( n1793 , n1790 , n1792 );
not ( n1794 , n1790 );
and ( n1795 , n1794 , n1791 );
nor ( n1796 , n1793 , n1795 );
and ( n1797 , n1045 , n1057 );
not ( n1798 , n1045 );
and ( n1799 , n1798 , n1056 );
nor ( n1800 , n1797 , n1799 );
not ( n1801 , n1800 );
and ( n1802 , n1579 , n1801 );
not ( n1803 , n1579 );
and ( n1804 , n1803 , n1800 );
nor ( n1805 , n1802 , n1804 );
xnor ( n1806 , n1089 , n1090 );
and ( n1807 , n1685 , n1806 );
not ( n1808 , n1685 );
not ( n1809 , n1806 );
and ( n1810 , n1808 , n1809 );
nor ( n1811 , n1807 , n1810 );
not ( n1812 , n788 );
not ( n1813 , n1812 );
not ( n1814 , n1089 );
or ( n1815 , n1813 , n1814 );
or ( n1816 , n1812 , n1089 );
nand ( n1817 , n1815 , n1816 );
and ( n1818 , n1787 , n1817 );
not ( n1819 , n1787 );
not ( n1820 , n1817 );
and ( n1821 , n1819 , n1820 );
nor ( n1822 , n1818 , n1821 );
not ( n1823 , n1392 );
not ( n1824 , n1389 );
or ( n1825 , n1823 , n1824 );
nand ( n1826 , n1825 , n1296 );
not ( n1827 , n1083 );
not ( n1828 , n1297 );
not ( n1829 , n1828 );
and ( n1830 , n1827 , n1829 );
and ( n1831 , n1083 , n1828 );
nor ( n1832 , n1830 , n1831 );
not ( n1833 , n1832 );
and ( n1834 , n1826 , n1833 );
not ( n1835 , n1826 );
and ( n1836 , n1835 , n1832 );
nor ( n1837 , n1834 , n1836 );
and ( n1838 , n1083 , n961 );
not ( n1839 , n1083 );
and ( n1840 , n1839 , n1084 );
nor ( n1841 , n1838 , n1840 );
and ( n1842 , n1681 , n1841 );
not ( n1843 , n1681 );
not ( n1844 , n1841 );
and ( n1845 , n1843 , n1844 );
nor ( n1846 , n1842 , n1845 );
not ( n1847 , n948 );
not ( n1848 , n1677 );
or ( n1849 , n1847 , n1848 );
not ( n1850 , n1679 );
nand ( n1851 , n1849 , n1850 );
and ( n1852 , n837 , n868 );
not ( n1853 , n837 );
and ( n1854 , n1853 , n963 );
nor ( n1855 , n1852 , n1854 );
not ( n1856 , n1855 );
and ( n1857 , n1851 , n1856 );
not ( n1858 , n1851 );
and ( n1859 , n1858 , n1855 );
nor ( n1860 , n1857 , n1859 );
not ( n1861 , n1386 );
not ( n1862 , n947 );
and ( n1863 , n1861 , n1862 );
not ( n1864 , n946 );
and ( n1865 , n1864 , n947 );
nor ( n1866 , n1863 , n1865 );
not ( n1867 , n1866 );
and ( n1868 , n1677 , n1867 );
not ( n1869 , n1677 );
and ( n1870 , n1869 , n1866 );
nor ( n1871 , n1868 , n1870 );
and ( n1872 , n1295 , n963 );
not ( n1873 , n1295 );
and ( n1874 , n1873 , n868 );
nor ( n1875 , n1872 , n1874 );
not ( n1876 , n1875 );
and ( n1877 , n1389 , n1876 );
not ( n1878 , n1389 );
and ( n1879 , n1878 , n1875 );
nor ( n1880 , n1877 , n1879 );
not ( n1881 , n1386 );
not ( n1882 , n1373 );
and ( n1883 , n1881 , n1882 );
and ( n1884 , n1864 , n1373 );
nor ( n1885 , n1883 , n1884 );
not ( n1886 , n1383 );
and ( n1887 , n1885 , n1886 );
not ( n1888 , n1885 );
and ( n1889 , n1888 , n1383 );
nor ( n1890 , n1887 , n1889 );
and ( n1891 , n823 , n752 );
not ( n1892 , n823 );
and ( n1893 , n1892 , n1378 );
nor ( n1894 , n1891 , n1893 );
not ( n1895 , n1377 );
and ( n1896 , n1894 , n1895 );
not ( n1897 , n1894 );
and ( n1898 , n1897 , n1377 );
nor ( n1899 , n1896 , n1898 );
and ( n1900 , n823 , n1075 );
not ( n1901 , n823 );
and ( n1902 , n1901 , n745 );
nor ( n1903 , n1900 , n1902 );
and ( n1904 , n1903 , n835 );
not ( n1905 , n1903 );
and ( n1906 , n1905 , n834 );
nor ( n1907 , n1904 , n1906 );
not ( n1908 , n748 );
buf ( n1909 , n833 );
not ( n1910 , n1909 );
or ( n1911 , n1908 , n1910 );
or ( n1912 , n748 , n1909 );
nand ( n1913 , n1911 , n1912 );
not ( n1914 , n746 );
not ( n1915 , n1909 );
or ( n1916 , n1914 , n1915 );
or ( n1917 , n1909 , n746 );
nand ( n1918 , n1916 , n1917 );
xor ( n1919 , n1588 , n1611 );
and ( n1920 , n1287 , n1057 );
not ( n1921 , n1287 );
and ( n1922 , n1921 , n1056 );
nor ( n1923 , n1920 , n1922 );
xnor ( n1924 , n1650 , n1923 );
xor ( n1925 , n1235 , n1114 );
endmodule
