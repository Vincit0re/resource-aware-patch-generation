module top ( g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 , g98 , g99 , g100 , g101 , g102 , g103 , g104 , g105 , g106 , g107 , g108 , g109 , g110 , g111 , g112 , g113 , g114 , g115 , g116 , g117 , g118 , g119 , g120 , g121 , g122 , g123 , g124 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g136 , g137 , g138 , g139 , g140 , g141 , g142 , g143 , g144 , g145 , g146 , g147 , g148 , g149 , g150 , g151 , g152 , g153 , g154 , g155 , g156 , g157 , g158 , g159 , g160 , g161 , g162 , g163 , g164 , g165 , g166 , g167 , g168 , g169 , g170 , g171 , g172 , g173 , g174 , g175 , g176 , g177 , g178 , g179 , g180 , g181 , g182 , g183 , g184 , g185 , g186 , g187 , g188 , g189 , g190 , g191 , g192 , g193 , g194 , g195 , g196 , g197 , g198 , g199 , g200 , g201 , g202 , g203 , g204 , g205 , g206 , g207 , g208 , g209 , g210 , g211 , g212 , g213 , g214 , g215 , g216 , g217 , g218 , g219 , g220 , g221 , g222 , g223 , g224 , g225 , g226 , g227 , g228 , g229 , g230 , g231 , g232 , g233 , g234 , g235 , g236 , g237 , g238 , g239 , g240 , g241 , g242 , g243 , g244 , g245 , g246 , g247 , g248 , g249 , g250 , g251 , g252 , g253 , g254 , g255 , g256 , g257 , g258 , g259 , g260 , g261 , g262 , g263 , g264 , g265 , g266 , g267 , g268 , g269 , g270 , g271 , g272 , g273 , g274 , g275 , g276 , g277 , g278 , g279 , g280 , g281 , g282 , g283 , g284 , g285 , g286 , g287 , g288 , g289 , g290 , g291 , g292 , g293 , g294 , g295 , g296 , g297 , g298 , g299 , g300 , g301 , g302 , g303 , g304 , g305 , g306 , g307 , g308 , g309 , g310 , g311 , g312 , g313 , g314 , g315 , g316 , g317 , g318 , g319 , g320 , g321 , g322 , g323 , g324 , g325 , g326 , g327 , g328 , g329 , g330 , g331 , g332 , g333 , g334 , g335 , g336 , g337 , g338 , g339 , g340 , g341 , g342 , g343 , g344 , g345 , g346 , g347 , g348 , g349 , g350 , g351 , g352 , g353 , g354 , g355 , g356 , g357 , g358 , g359 , g360 , g361 , g362 , g363 , g364 , g365 , g366 , g367 , g368 , g369 , g370 , g371 , g372 , g373 , g374 , g375 , g376 , g377 , g378 , g379 , g380 , g381 , g382 , g383 , g384 , g385 , g386 , g387 , g388 , g389 , g390 , g391 , g392 , g393 , g394 , g395 , g396 , g397 , g398 , g399 , g400 , g401 , g402 , g403 , g404 , g405 , g406 , g407 , g408 , g409 , g410 , g411 , g412 , g413 , g414 , g415 , g416 , g417 , g418 , g419 , g420 , g421 , g422 , g423 , g424 , g425 , g426 , g427 , g428 , g429 , g430 , g431 , g432 , g433 , g434 , g435 , g436 , g437 , g438 , g439 , g440 , g441 , g442 , g443 , g444 , g445 , g446 , g447 , g448 , g449 , g450 , g451 , g452 , g453 , g454 , g455 , g456 , g457 , g458 , g459 , g460 , g461 , g462 , g463 , g464 , g465 , g466 , g467 , g468 , g469 , g470 , g471 , g472 , g473 , g474 , g475 , g476 , g477 , g478 , g479 , g480 , g481 , g482 , g483 , g484 , g485 , g486 , g487 , g488 , g489 , g490 , g491 , g492 , g493 , g494 , g495 , g496 , g497 , g498 , g499 , g500 , g501 , g502 , g503 , g504 , g505 , g506 , g507 , g508 , g509 , g510 , g511 , g512 , g513 , g514 , g515 , g516 , g517 , g518 , g519 , g520 , g521 , g522 , g523 , g524 , g525 , g526 , g527 , g528 , g529 , g530 , g531 , g532 , g533 , g534 , g535 , g536 , g537 , g538 , g539 , g540 , g541 , g542 , g543 , g544 , g545 , g546 , g547 , g548 , g549 , g550 , g551 , g552 , g553 , g554 , g555 , g556 , g557 , g558 , g559 , g560 , g561 , g562 , g563 , g564 , g565 , g566 , g567 , g568 , g569 , g570 , g571 , g572 , g573 , g574 , g575 , g576 , g577 , g578 , g579 , g580 , g581 , g582 , g583 , g584 , g585 , g586 , g587 , g588 , g589 , g590 , g591 , g592 , g593 , g594 , g595 , g596 , g597 , g598 , g599 , g600 , g601 , g602 , g603 , g604 , g605 , g606 , g607 , g608 , g609 , g610 , g611 , g612 , g613 , g614 , g615 , g616 , g617 , g618 , g619 , g620 , g621 , g622 , g623 , g624 , g625 , g626 , g627 , g628 , g629 , g630 , g631 , g632 , g633 , g634 , g635 , g636 , g637 , g638 , g639 , g640 , g641 , g642 , g643 , g644 , g645 , g646 , g647 , g648 , g649 , g650 , g651 , g652 , g653 , g654 , g655 , g656 , g657 , g658 , g659 , g660 , g661 , g662 , g663 , g664 , g665 , g666 , g667 , g668 , g669 , g670 , g671 , g672 , g673 , g674 , g675 , g676 , g677 , g678 , g679 , g680 , g681 , g682 , g683 , g684 , g685 , g686 , g687 , g688 , g689 , g690 , g691 , g692 , g693 , g694 , g695 , g696 , g697 , g698 , g699 , g700 , g701 , g702 , g703 , g704 , g705 , g706 , g707 , g708 , g709 , g710 , g711 , g712 , g713 , g714 , g715 , g716 , g717 , g718 , g719 , g720 , g721 , g722 , g723 , g724 , g725 , g726 , g727 , g728 , g729 , g730 , g731 , g732 , g733 , g734 , g735 , g736 , g737 , g738 , g739 , g740 , g741 , g742 , g743 , g744 , g745 , g746 , g747 , g748 , g749 , g750 , g751 , g752 , g753 , g754 , g755 , g756 , g757 , g758 , g759 , g760 , g761 , g762 , g763 , g764 , g765 , g766 , g767 , g768 , g769 , g770 , g771 , g772 , g773 , g774 , g775 , g776 , g777 , g778 , g779 , g780 , g781 , g782 , g783 , g784 , g785 , g786 , g787 , g788 , g789 , g790 , g791 , g792 , g793 , g794 , g795 , g796 , g797 , g798 , g799 , g800 , g801 , g802 , g803 , g804 , g805 , g806 , g807 , g808 , g809 , g810 , g811 , g812 , g813 , g814 , g815 , g816 , g817 , g818 , g819 , g820 , g821 , g822 , g823 , g824 , g825 , g826 , g827 , g828 , g829 , g830 , g831 , g832 , g833 , g834 , g835 , g836 , g837 , g838 , g839 , g840 , g841 , g842 , g843 , g844 , g845 , g846 , g847 , g848 , g849 , g850 , g851 , g852 , g853 , g854 , g855 , g856 , g857 , g858 , g859 , g860 , g861 , g862 , g863 , g864 , g865 , g866 , g867 , g868 , g869 , g870 , g871 , g872 , g873 , g874 , g875 , g876 , g877 , g878 , g879 , g880 , g881 , g882 , g883 , g884 , g885 , g886 , g887 , g888 , g889 , g890 , g891 , g892 , g893 , g894 , g895 , g896 , g897 , g898 , g899 , g900 , g901 , g902 , g903 , g904 , g905 , g906 , g907 , g908 , g909 , g910 , g911 , g912 , g913 , g914 , g915 , g916 , g917 , g918 , g919 , g920 , g921 , g922 , g923 , g924 , g925 , g926 , g927 , g928 , g929 , g930 , g931 , g932 , g933 , g934 , g935 , g936 , g937 , g938 , g939 , g940 , g941 , g942 , g943 , g944 , g945 , g946 , g947 , g948 , g949 , g950 , g951 , g952 , g953 , g954 , g955 , g956 , g957 , g958 , g959 , g960 , g961 , g962 , g963 , g964 , g965 , g966 , g967 , g968 , g969 , g970 , g971 , g972 , g973 , g974 , g975 , g976 , g977 , g978 , g979 , g980 , g981 , g982 , g983 , g984 , g985 , g986 , g987 , g988 , g989 , g990 , g991 , g992 , g993 , g994 , g995 , g996 , g997 , g998 , g999 , g1000 , g1001 , g1002 , g1003 , g1004 , g1005 , g1006 , g1007 , g1008 , g1009 , g1010 , g1011 , g1012 , g1013 , g1014 , g1015 , g1016 , g1017 , g1018 , g1019 , g1020 , g1021 , g1022 , g1023 , g1024 , g1025 , g1026 , g1027 , g1028 , g1029 , g1030 , g1031 , g1032 , g1033 , g1034 , g1035 , g1036 , g1037 , g1038 , g1039 , g1040 , g1041 , g1042 , g1043 , g1044 , g1045 , g1046 , g1047 , g1048 , g1049 , g1050 , g1051 , g1052 , g1053 , g1054 , g1055 , g1056 , g1057 , g1058 , g1059 , g1060 , g1061 , g1062 , g1063 , g1064 , g1065 , g1066 , g1067 , g1068 , g1069 , g1070 , g1071 , g1072 , g1073 , g1074 , g1075 , g1076 , g1077 , g1078 , g1079 , g1080 , g1081 , g1082 , g1083 , g1084 , g1085 , g1086 , g1087 , g1088 , g1089 , g1090 , g1091 , g1092 , g1093 , g1094 , g1095 , g1096 , g1097 , g1098 , g1099 , g1100 , g1101 , g1102 , g1103 , g1104 , g1105 , g1106 , g1107 , g1108 , g1109 , g1110 , g1111 , g1112 , g1113 , g1114 , g1115 , g1116 , g1117 , g1118 , g1119 , g1120 , g1121 , g1122 , g1123 , g1124 , g1125 , g1126 , g1127 , g1128 , g1129 , g1130 , g1131 , g1132 , g1133 , g1134 , g1135 , g1136 , g1137 , g1138 , g1139 , g1140 , g1141 , g1142 , g1143 , g1144 , g1145 , g1146 , g1147 , g1148 , g1149 , g1150 , g1151 , g1152 , g1153 , g1154 , g1155 , g1156 , g1157 , g1158 , g1159 , g1160 , g1161 , g1162 , g1163 , g1164 , g1165 , g1166 , g1167 , g1168 , g1169 , g1170 , g1171 , g1172 , g1173 , g1174 , g1175 , g1176 , g1177 , g1178 , g1179 , g1180 , g1181 , g1182 , g1183 , g1184 , g1185 , g1186 , g1187 , g1188 , g1189 , g1190 , g1191 , g1192 , g1193 , g1194 , g1195 , g1196 , g1197 , g1198 , g1199 , g1200 , g1201 , g1202 , g1203 , g1204 , g1205 , g1206 , g1207 , g1208 , g1209 , g1210 , g1211 , g1212 , g1213 , g1214 , g1215 , g1216 , g1217 , g1218 , g1219 , g1220 , g1221 , g1222 , g1223 , g1224 , g1225 , g1226 , g1227 , g1228 , g1229 , g1230 , g1231 , g1232 , g1233 , g1234 , g1235 , g1236 , g1237 , g1238 , g1239 , g1240 , g1241 , g1242 , g1243 , g1244 , g1245 , g1246 , g1247 , g1248 , g1249 , g1250 , g1251 , g1252 , g1253 , g1254 , g1255 , g1256 , g1257 , g1258 , g1259 , g1260 , g1261 , g1262 , g1263 , g1264 , g1265 , g1266 , g1267 , g1268 , g1269 , g1270 , g1271 , g1272 , g1273 , g1274 , g1275 , g1276 , g1277 , g1278 , g1279 , g1280 , g1281 , g1282 , g1283 , g1284 , g1285 , g1286 , g1287 , g1288 , g1289 , g1290 , g1291 , g1292 , g1293 , g1294 , g1295 , g1296 , g1297 , g1298 , g1299 , g1300 , g1301 , g1302 , g1303 , g1304 , g1305 , g1306 , g1307 , g1308 , g1309 , g1310 , g1311 , g1312 , g1313 , g1314 , g1315 , g1316 , g1317 , g1318 , g1319 , g1320 , g1321 , g1322 , g1323 , g1324 , g1325 , g1326 , g1327 , g1328 , g1329 , g1330 , g1331 , g1332 , g1333 , g1334 , g1335 , g1336 , g1337 , g1338 , g1339 , g1340 , g1341 , g1342 , g1343 , g1344 , g1345 , g1346 , g1347 , g1348 , g1349 , g1350 , g1351 , g1352 , g1353 , g1354 , g1355 , g1356 , g1357 , g1358 , g1359 , g1360 , g1361 , g1362 , g1363 , g1364 , g1365 , g1366 , g1367 , g1368 , g1369 , g1370 , g1371 , g1372 , g1373 , g1374 , g1375 , g1376 , g1377 , g1378 , g1379 , g1380 , g1381 , g1382 , g1383 , g1384 , g1385 , g1386 , g1387 , g1388 , g1389 , g1390 , g1391 , g1392 , g1393 , g1394 , g1395 , g1396 , g1397 , g1398 , g1399 , g1400 , g1401 , g1402 , g1403 , g1404 , g1405 , g1406 , g1407 , g1408 , g1409 , g1410 , g1411 , g1412 , g1413 , g1414 , g1415 , g1416 , g1417 , g1418 , g1419 , g1420 , g1421 , g1422 , g1423 , g1424 , g1425 , g1426 , g1427 , g1428 , g1429 , g1430 , g1431 , g1432 , g1433 , g1434 , g1435 , g1436 , g1437 , g1438 , g1439 , g1440 , g1441 , g1442 , g1443 , g1444 , g1445 , g1446 , g1447 , g1448 , g1449 , g1450 , g1451 , g1452 , g1453 , g1454 , g1455 , g1456 , g1457 , g1458 , g1459 , g1460 , g1461 , g1462 , g1463 , g1464 , g1465 , g1466 , g1467 , g1468 , g1469 , g1470 , g1471 , g1472 , g1473 , g1474 , g1475 , g1476 , g1477 , g1478 , g1479 , g1480 , g1481 , g1482 , g1483 , g1484 , g1485 , g1486 , g1487 , g1488 , g1489 , g1490 , g1491 , g1492 , g1493 , g1494 , g1495 , g1496 , g1497 , g1498 , g1499 , g1500 , g1501 , g1502 , g1503 , g1504 , g1505 , g1506 , g1507 , g1508 , g1509 , g1510 , g1511 , g1512 , g1513 , g1514 , g1515 , g1516 , g1517 , g1518 , g1519 , g1520 , g1521 , g1522 , g1523 , g1524 , g1525 , g1526 , g1527 , g1528 , g1529 , g1530 , g1531 , g1532 , g1533 , g1534 , g1535 , g1536 , g1537 , g1538 , g1539 , g1540 , g1541 , g1542 , g1543 , g1544 , g1545 , g1546 , g1547 , g1548 , g1549 , g1550 , g1551 , g1552 , g1553 , g1554 , g1555 , g1556 , g1557 , g1558 , g1559 , g1560 , g1561 , g1562 , g1563 , g1564 , g1565 , g1566 , g1567 , g1568 , g1569 , g1570 , g1571 , g1572 , g1573 , g1574 , g1575 , g1576 , g1577 , g1578 , g1579 , g1580 , g1581 , g1582 , g1583 , g1584 , g1585 , g1586 , g1587 , g1588 , g1589 , g1590 , g1591 , g1592 , g1593 , g1594 , g1595 , g1596 , g1597 , g1598 , g1599 , g1600 , g1601 , g1602 , g1603 , g1604 , g1605 , g1606 , g1607 , g1608 , g1609 , g1610 , g1611 , g1612 , g1613 , g1614 , g1615 , g1616 , g1617 , g1618 , g1619 , g1620 , g1621 , g1622 , g1623 , g1624 , g1625 , g1626 , g1627 , g1628 , g1629 , g1630 , g1631 , g1632 , g1633 , g1634 , g1635 , g1636 , g1637 , g1638 , g1639 , g1640 , g1641 , g1642 , g1643 , g1644 , g1645 , g1646 , g1647 , g1648 , g1649 , g1650 , g1651 , g1652 , g1653 , g1654 , g1655 , g1656 , g1657 , g1658 , g1659 , g1660 , g1661 , g1662 , g1663 , g1664 , g1665 , g1666 , g1667 , g1668 , g1669 , g1670 , g1671 , g1672 , g1673 , g1674 , g1675 , g1676 , g1677 , g1678 , g1679 , g1680 , g1681 , g1682 , g1683 , g1684 , g1685 , g1686 , g1687 , g1688 , g1689 , g1690 , g1691 , g1692 , g1693 , g1694 , g1695 , g1696 , g1697 , g1698 , g1699 , g1700 , g1701 , g1702 , g1703 , g1704 , g1705 , g1706 , g1707 , g1708 , g1709 , g1710 , g1711 , g1712 , g1713 , g1714 , g1715 , g1716 , g1717 , g1718 , g1719 , g1720 , g1721 , g1722 , g1723 , g1724 , g1725 , g1726 , g1727 , g1728 , g1729 , g1730 , g1731 , g1732 , g1733 , g1734 , g1735 , g1736 , g1737 , g1738 , g1739 , g1740 , g1741 , g1742 , g1743 , g1744 , g1745 , g1746 , g1747 , g1748 , g1749 , g1750 , g1751 , g1752 , g1753 , g1754 , g1755 , g1756 , g1757 , g1758 , g1759 , g1760 , g1761 , g1762 , g1763 , g1764 , g1765 , g1766 , g1767 , g1768 , g1769 , g1770 , g1771 , g1772 , g1773 , g1774 , g1775 , g1776 , g1777 , g1778 , g1779 , g1780 , g1781 , g1782 , g1783 , g1784 , g1785 , g1786 , g1787 , g1788 , g1789 , g1790 , g1791 , g1792 , g1793 , g1794 , g1795 , g1796 , g1797 , g1798 , g1799 , g1800 , g1801 , g1802 , g1803 , g1804 , g1805 , g1806 , g1807 , g1808 , g1809 , g1810 , g1811 , g1812 , g1813 , g1814 , g1815 , g1816 , g1817 , g1818 , g1819 , g1820 , g1821 , g1822 , g1823 , g1824 , g1825 , g1826 , g1827 , g1828 , g1829 , g1830 , g1831 , g1832 , g1833 , g1834 , g1835 , g1836 , g1837 , g1838 , g1839 , g1840 , g1841 , g1842 , g1843 , g1844 , g1845 , g1846 , g1847 , g1848 , g1849 , g1850 , g1851 , g1852 , g1853 , g1854 , g1855 , g1856 , g1857 , g1858 , g1859 , g1860 , g1861 , g1862 , g1863 , g1864 , g1865 , g1866 , g1867 , g1868 , g1869 , g1870 , g1871 , g1872 , g1873 , g1874 , g1875 , g1876 , g1877 , g1878 , g1879 , g1880 , g1881 , g1882 , g1883 , g1884 , g1885 , g1886 , g1887 , g1888 , g1889 , g1890 , g1891 , g1892 , g1893 , g1894 , g1895 , g1896 , g1897 , g1898 , g1899 , g1900 , g1901 , g1902 , g1903 , g1904 , g1905 , g1906 , g1907 , g1908 , g1909 , g1910 , g1911 , g1912 , g1913 , g1914 , g1915 , g1916 , g1917 , g1918 , g1919 , g1920 , g1921 , g1922 , g1923 , g1924 , g1925 , g1926 , g1927 , g1928 , g1929 , g1930 , g1931 , g1932 , g1933 , g1934 , g1935 , g1936 , g1937 , g1938 , g1939 , g1940 , g1941 , g1942 , g1943 , g1944 , g1945 , g1946 , g1947 , g1948 , g1949 , g1950 , g1951 , g1952 , g1953 , g1954 , g1955 , g1956 , g1957 , g1958 , g1959 , g1960 , g1961 , g1962 , g1963 , g1964 , g1965 , g1966 , g1967 , g1968 , g1969 , g1970 , g1971 , g1972 , g1973 , g1974 , g1975 , g1976 , g1977 , g1978 , g1979 , g1980 , g1981 , g1982 , g1983 , g1984 , g1985 , g1986 , g1987 , g1988 , g1989 , g1990 , g1991 , g1992 , g1993 , g1994 , g1995 , g1996 , g1997 , g1998 , g1999 , g2000 , g2001 , g2002 , g2003 , g2004 , g2005 , g2006 , g2007 , g2008 , g2009 , g2010 , g2011 , g2012 , g2013 , g2014 , g2015 , g2016 , g2017 , g2018 , g2019 , g2020 , g2021 , g2022 , g2023 , g2024 , g2025 , g2026 , g2027 , g2028 , g2029 , g2030 , g2031 , g2032 , g2033 , g2034 , g2035 , g2036 , g2037 , g2038 , g2039 , g2040 , g2041 , g2042 , g2043 , g2044 , g2045 , g2046 , g2047 , g2048 , g2049 , g2050 , g2051 , g2052 , g2053 , g2054 , g2055 , g2056 , g2057 , g2058 , g2059 , g2060 , g2061 , g2062 , g2063 , g2064 , g2065 , g2066 , g2067 , g2068 , g2069 , g2070 , g2071 , g2072 , g2073 , g2074 , g2075 , g2076 , g2077 , g2078 , g2079 , g2080 , g2081 , g2082 , g2083 , g2084 , g2085 , g2086 , g2087 , g2088 , g2089 , g2090 , g2091 , g2092 , g2093 , g2094 , g2095 , g2096 , g2097 , g2098 , g2099 , g2100 , g2101 , g2102 , g2103 , g2104 , g2105 , g2106 , g2107 , g2108 , g2109 , g2110 , g2111 , g2112 , g2113 , g2114 , g2115 , g2116 , g2117 , g2118 , g2119 , g2120 , g2121 , g2122 , g2123 , g2124 , g2125 , g2126 , g2127 , g2128 , g2129 , g2130 , g2131 , g2132 , g2133 , g2134 , g2135 , g2136 , g2137 , g2138 , g2139 , g2140 , g2141 , g2142 , g2143 , g2144 , g2145 , g2146 , g2147 , g2148 , g2149 , g2150 , g2151 , g2152 , g2153 , g2154 , g2155 , g2156 , g2157 , g2158 , g2159 , g2160 , g2161 , g2162 , g2163 , g2164 , g2165 , g2166 , g2167 , g2168 , g2169 , g2170 , g2171 , g2172 , g2173 , g2174 , g2175 , g2176 , g2177 , g2178 , g2179 , g2180 , g2181 , g2182 , g2183 , g2184 , g2185 , g2186 , g2187 , g2188 , g2189 , g2190 , g2191 , g2192 , g2193 , g2194 , g2195 , g2196 , g2197 , g2198 , g2199 , g2200 , g2201 , g2202 , g2203 , g2204 , g2205 , g2206 , g2207 , g2208 , g2209 , g2210 , g2211 , g2212 , g2213 , g2214 , g2215 , g2216 , g2217 , g2218 , g2219 , g2220 , g2221 , g2222 , g2223 , g2224 , g2225 , g2226 , g2227 , g2228 , g2229 , g2230 , g2231 , g2232 , g2233 , g2234 , g2235 , g2236 , g2237 , g2238 , g2239 , g2240 , g2241 , g2242 , g2243 , g2244 , g2245 , g2246 , g2247 , g2248 , g2249 , g2250 , g2251 , g2252 , g2253 , g2254 , g2255 , g2256 , g2257 , g2258 , g2259 , g2260 , g2261 , g2262 , g2263 , g2264 , g2265 , g2266 , g2267 , g2268 , g2269 , g2270 , g2271 , g2272 , g2273 , g2274 , g2275 , g2276 , g2277 , g2278 , g2279 , g2280 , g2281 , g2282 , g2283 , g2284 , g2285 , g2286 , g2287 , g2288 , g2289 , g2290 , g2291 , g2292 , g2293 , g2294 , g2295 , g2296 , g2297 , g2298 , g2299 , g2300 , g2301 , g2302 , g2303 , g2304 , g2305 , g2306 , g2307 , g2308 , g2309 , g2310 , g2311 , g2312 , g2313 , g2314 , g2315 , g2316 , g2317 , g2318 , g2319 , g2320 , g2321 , g2322 , g2323 , g2324 , g2325 , g2326 , g2327 , g2328 , g2329 , g2330 , g2331 , g2332 , g2333 , g2334 , g2335 , g2336 , g2337 , g2338 , g2339 , g2340 , g2341 , g2342 , g2343 , g2344 , g2345 , g2346 , g2347 , g2348 , g2349 , g2350 , g2351 , g2352 , g2353 , g2354 , g2355 , g2356 , g2357 , g2358 , g2359 , g2360 , g2361 , g2362 , g2363 , g2364 , g2365 , g2366 , g2367 , g2368 , g2369 , g2370 , g2371 , g2372 , g2373 , g2374 , g2375 , g2376 , g2377 , g2378 , g2379 , g2380 , g2381 , g2382 , g2383 , g2384 , g2385 , g2386 , g2387 , g2388 , g2389 , g2390 , g2391 , g2392 , g2393 , g2394 , g2395 , g2396 , g2397 , g2398 , g2399 , g2400 , g2401 , g2402 , g2403 , g2404 , g2405 , g2406 , g2407 , g2408 , g2409 , g2410 , g2411 , g2412 , g2413 , g2414 , g2415 , g2416 , g2417 , g2418 , g2419 , g2420 , g2421 , g2422 , g2423 , g2424 , g2425 , g2426 , g2427 , g2428 , g2429 , g2430 , g2431 , g2432 , g2433 , g2434 , g2435 , g2436 , g2437 , g2438 , g2439 , g2440 , g2441 , g2442 , g2443 , g2444 , g2445 , g2446 , g2447 , g2448 , g2449 , g2450 , g2451 , g2452 , g2453 , g2454 , g2455 , g2456 , g2457 , g2458 , g2459 , g2460 , g2461 , g2462 , g2463 , g2464 , g2465 , g2466 , g2467 , g2468 , g2469 , g2470 , g2471 , g2472 , g2473 , g2474 , g2475 , g2476 , g2477 , g2478 , g2479 , g2480 , g2481 , g2482 , g2483 , g2484 , g2485 , g2486 , g2487 , g2488 , g2489 , g2490 , g2491 , g2492 , g2493 , g2494 , g2495 , g2496 , g2497 , g2498 , g2499 , g2500 , g2501 , g2502 , g2503 , g2504 , g2505 , g2506 , g2507 , g2508 , g2509 , g2510 , g2511 , g2512 , g2513 , g2514 , g2515 , g2516 , g2517 , g2518 , g2519 , g2520 , g2521 , g2522 , g2523 , g2524 , g2525 , g2526 , g2527 , g2528 , g2529 , g2530 , g2531 , g2532 , g2533 , g2534 , g2535 , g2536 , g2537 , g2538 , g2539 , g2540 , g2541 , g2542 , g2543 , g2544 , g2545 , g2546 , g2547 , g2548 , g2549 , g2550 , g2551 , g2552 , g2553 , g2554 , g2555 , g2556 , g2557 , g2558 , g2559 , g2560 , g2561 , g2562 , g2563 , g2564 , g2565 , g2566 , g2567 , g2568 , g2569 , g2570 , g2571 , g2572 , g2573 , g2574 , g2575 , g2576 , g2577 , g2578 , g2579 , g2580 , g2581 , g2582 , g2583 , g2584 , g2585 , g2586 , g2587 , g2588 , g2589 , g2590 , g2591 , g2592 , g2593 , g2594 , g2595 , g2596 , g2597 , g2598 , g2599 , g2600 , g2601 , g2602 , g2603 , g2604 , g2605 , g2606 , g2607 , g2608 , g2609 , g2610 , g2611 , g2612 , g2613 , g2614 , g2615 , g2616 , g2617 , g2618 , g2619 , g2620 , g2621 , g2622 , g2623 , g2624 , g2625 , g2626 , g2627 , g2628 , g2629 , g2630 , g2631 , g2632 , g2633 , g2634 , g2635 , g2636 , g2637 , g2638 , g2639 , g2640 , g2641 , g2642 , g2643 , g2644 , g2645 , g2646 , g2647 , g2648 , g2649 , g2650 , g2651 , g2652 , g2653 , g2654 , g2655 , g2656 , g2657 , g2658 , g2659 , g2660 , g2661 , g2662 , g2663 , g2664 , g2665 , g2666 , g2667 , g2668 , g2669 , g2670 , g2671 , g2672 , g2673 , g2674 , g2675 , g2676 , g2677 , g2678 , g2679 , g2680 , g2681 , g2682 , g2683 , g2684 , g2685 , g2686 , g2687 , g2688 , g2689 , g2690 , g2691 , g2692 , g2693 , g2694 , g2695 , g2696 , g2697 , g2698 , g2699 , g2700 , g2701 , g2702 , g2703 , g2704 , g2705 , g2706 , g2707 , g2708 , g2709 , g2710 , g2711 , g2712 , g2713 , g2714 , g2715 , g2716 , g2717 , g2718 , g2719 , g2720 , g2721 , g2722 , g2723 , g2724 , g2725 , g2726 , g2727 , g2728 , g2729 , g2730 , g2731 , g2732 , g2733 , g2734 , g2735 , g2736 , g2737 , g2738 , g2739 , g2740 , g2741 , g2742 , g2743 , g2744 , g2745 , g2746 , g2747 , g2748 , g2749 , g2750 , g2751 , g2752 , g2753 , g2754 , g2755 , g2756 , g2757 , g2758 , g2759 , g2760 , g2761 , g2762 , g2763 , g2764 , g2765 , g2766 , g2767 , g2768 , g2769 , g2770 , g2771 , g2772 , g2773 , g2774 , g2775 , g2776 , g2777 , g2778 , g2779 , g2780 , g2781 , g2782 , g2783 , g2784 , g2785 , g2786 , g2787 , g2788 , g2789 , g2790 , g2791 , g2792 , g2793 , g2794 , g2795 , g2796 , g2797 , g2798 , g2799 , g2800 , g2801 , g2802 , g2803 , g2804 , g2805 , g2806 , g2807 , g2808 , g2809 , g2810 , g2811 , g2812 , g2813 , g2814 , g2815 , g2816 , g2817 , g2818 , g2819 , g2820 , g2821 , g2822 , g2823 , g2824 , g2825 , g2826 , g2827 , g2828 , g2829 , g2830 , g2831 , g2832 , g2833 , g2834 , g2835 , g2836 , g2837 , g2838 , g2839 , g2840 , g2841 , g2842 , g2843 , g2844 , g2845 , g2846 , g2847 , g2848 , g2849 , g2850 , g2851 , g2852 , g2853 , g2854 , g2855 , g2856 , g2857 , g2858 , g2859 , g2860 , g2861 , g2862 , g2863 , g2864 , g2865 , g2866 , g2867 , g2868 , g2869 , g2870 , g2871 , g2872 , g2873 , g2874 , g2875 , g2876 , g2877 , g2878 , g2879 , g2880 , g2881 , g2882 , g2883 , g2884 , g2885 , g2886 , g2887 , g2888 , g2889 , g2890 , g2891 , g2892 , g2893 , g2894 , g2895 , g2896 , g2897 , g2898 , g2899 , g2900 , g2901 , g2902 , g2903 , g2904 , g2905 , g2906 , g2907 , g2908 , g2909 , g2910 , g2911 , g2912 , g2913 , g2914 , g2915 , g2916 , g2917 , g2918 , g2919 , g2920 , g2921 , g2922 , g2923 , g2924 , g2925 , g2926 , g2927 , g2928 , g2929 , g2930 , g2931 , g2932 , g2933 , g2934 , g2935 , g2936 , g2937 , g2938 , g2939 , g2940 , g2941 , g2942 , g2943 , g2944 , g2945 , g2946 , g2947 , g2948 , g2949 , g2950 , g2951 , g2952 , g2953 , g2954 , g2955 , g2956 , g2957 , g2958 , g2959 , g2960 , g2961 , g2962 , g2963 , g2964 , g2965 , g2966 , g2967 , g2968 , g2969 , g2970 , g2971 , g2972 , g2973 , g2974 , g2975 , g2976 , g2977 , g2978 , g2979 , g2980 , g2981 , g2982 , g2983 , g2984 , g2985 , g2986 , g2987 , g2988 , g2989 , g2990 , g2991 , g2992 , g2993 , g2994 , g2995 , g2996 , g2997 , g2998 , g2999 , g3000 , g3001 , g3002 , g3003 , g3004 , g3005 , g3006 , g3007 , g3008 , g3009 , g3010 , g3011 , g3012 , g3013 , g3014 , g3015 , g3016 , g3017 , g3018 , g3019 , g3020 , g3021 , g3022 , g3023 , g3024 , g3025 , g3026 , g3027 , g3028 , g3029 , g3030 , g3031 , g3032 , g3033 , g3034 , g3035 , g3036 , g3037 , g3038 , g3039 , g3040 , g3041 , g3042 , g3043 , g3044 , g3045 , g3046 , g3047 , g3048 , g3049 , g3050 , g3051 , g3052 , g3053 , g3054 , g3055 , g3056 , g3057 , g3058 , g3059 , g3060 , g3061 , g3062 , g3063 , g3064 , g3065 , g3066 , g3067 , g3068 , g3069 , g3070 , g3071 , g3072 , g3073 , g3074 , g3075 , g3076 , g3077 , g3078 , g3079 , g3080 , g3081 , g3082 , g3083 , g3084 , g3085 , g3086 , g3087 , g3088 , g3089 , g3090 , g3091 , g3092 , g3093 , g3094 , g3095 , g3096 , g3097 , g3098 , g3099 , g3100 , g3101 , g3102 , g3103 , g3104 , g3105 , g3106 , g3107 , g3108 , g3109 , g3110 , g3111 , g3112 , g3113 , g3114 , g3115 , g3116 , g3117 , g3118 , g3119 , g3120 , g3121 , g3122 , g3123 , g3124 , g3125 , g3126 , g3127 , g3128 , g3129 , g3130 , g3131 , g3132 , g3133 , g3134 , g3135 , g3136 , g3137 , g3138 , g3139 , g3140 , g3141 , g3142 , g3143 , g3144 , g3145 , g3146 , g3147 , g3148 , g3149 , g3150 , g3151 , g3152 , g3153 , g3154 , g3155 , g3156 , g3157 , g3158 , g3159 , g3160 , g3161 , g3162 , g3163 , g3164 , g3165 , g3166 , g3167 , g3168 , g3169 , g3170 , g3171 , g3172 , g3173 , g3174 , g3175 , g3176 , g3177 , g3178 , g3179 , g3180 , g3181 , g3182 , g3183 , g3184 , g3185 , g3186 , g3187 , g3188 , g3189 , g3190 , g3191 , g3192 , g3193 , g3194 , g3195 , g3196 , g3197 , g3198 , g3199 , g3200 , g3201 , g3202 , g3203 , g3204 , g3205 , g3206 , g3207 , g3208 , g3209 , g3210 , g3211 , g3212 , g3213 , g3214 , g3215 , g3216 , g3217 , g3218 , g3219 , g3220 , g3221 , g3222 , g3223 , g3224 , g3225 , g3226 , g3227 , g3228 , g3229 , g3230 , g3231 , g3232 , g3233 , g3234 , g3235 , g3236 , g3237 , g3238 , g3239 , g3240 , g3241 , g3242 , g3243 , g3244 , g3245 , g3246 , g3247 , g3248 , g3249 , g3250 , g3251 , g3252 , g3253 , g3254 , g3255 , g3256 , g3257 , g3258 , g3259 , g3260 , g3261 , g3262 , g3263 , g3264 , g3265 , g3266 , g3267 , g3268 , g3269 , g3270 , g3271 , g3272 , g3273 , g3274 , g3275 , g3276 , g3277 , g3278 , g3279 , g3280 , g3281 , g3282 , g3283 , g3284 , g3285 , g3286 , g3287 , g3288 , g3289 , g3290 , g3291 , g3292 , g3293 , g3294 , g3295 , g3296 , g3297 , g3298 , g3299 , g3300 , g3301 , g3302 , g3303 , g3304 , g3305 , g3306 , g3307 , g3308 , g3309 , g3310 , g3311 , g3312 , g3313 , g3314 , g3315 , g3316 , g3317 , g3318 , g3319 , g3320 , g3321 , g3322 , g3323 , g3324 , g3325 , g3326 , g3327 , g3328 , g3329 , g3330 , g3331 , g3332 , g3333 , g3334 , g3335 , g3336 , g3337 , g3338 , g3339 , g3340 , g3341 , g3342 , g3343 , g3344 , g3345 , g3346 , g3347 , g3348 , g3349 , g3350 , g3351 , g3352 , g3353 , g3354 , g3355 , g3356 , g3357 , g3358 , g3359 , g3360 , g3361 , g3362 , g3363 , g3364 , g3365 , g3366 , g3367 , g3368 , g3369 , g3370 , g3371 , g3372 , g3373 , g3374 , g3375 , g3376 , g3377 , g3378 , g3379 , g3380 , g3381 , g3382 , g3383 , g3384 , g3385 , g3386 , g3387 , g3388 , g3389 , g3390 , g3391 , g3392 , g3393 , g3394 , g3395 , g3396 , g3397 , g3398 , g3399 , g3400 , g3401 , g3402 , g3403 , g3404 , g3405 , g3406 , g3407 , g3408 , g3409 , g3410 , g3411 , g3412 , g3413 , g3414 , g3415 , g3416 , g3417 , g3418 , g3419 , g3420 , g3421 , g3422 , g3423 , g3424 , g3425 , g3426 , g3427 , g3428 , g3429 , g3430 , g3431 , g3432 , g3433 , g3434 , g3435 , g3436 , g3437 , g3438 , g3439 , g3440 , g3441 , g3442 , g3443 , g3444 , g3445 , g3446 , g3447 , g3448 , g3449 , g3450 , g3451 , g3452 , g3453 , g3454 , g3455 , g3456 , g3457 , g3458 , g3459 , g3460 , g3461 , g3462 , g3463 , g3464 , g3465 , g3466 , g3467 , g3468 , g3469 , g3470 , g3471 , g3472 , g3473 , g3474 , g3475 , g3476 , g3477 , g3478 , g3479 , g3480 , g3481 , g3482 , g3483 , g3484 , g3485 , g3486 , g3487 , g3488 , g3489 , g3490 , g3491 , g3492 , g3493 , g3494 , g3495 , g3496 , g3497 , g3498 , g3499 , g3500 , g3501 , g3502 , g3503 , g3504 , g3505 , g3506 , g3507 , g3508 , g3509 , g3510 , g3511 , g3512 , g3513 , g3514 , g3515 , g3516 , g3517 , g3518 , g3519 , g3520 , g3521 , g3522 , g3523 , g3524 , g3525 , g3526 , g3527 , g3528 , g3529 , g3530 , g3531 , g3532 , g3533 , g3534 , g3535 , g3536 , g3537 , g3538 , g3539 , g3540 , g3541 , g3542 , g3543 , g3544 , g3545 , g3546 , g3547 , g3548 , g3549 , g3550 , g3551 , g3552 , g3553 , g3554 , g3555 , g3556 , g3557 , g3558 , g3559 , g3560 , g3561 , g3562 , g3563 , g3564 , g3565 , g3566 , g3567 , g3568 , g3569 , g3570 , g3571 , g3572 , g3573 , g3574 , g3575 , g3576 , g3577 , g3578 , g3579 , g3580 , g3581 , g3582 , g3583 , g3584 , g3585 , g3586 , g3587 , g3588 , g3589 , g3590 , g3591 , g3592 , g3593 , g3594 , g3595 , g3596 , g3597 , g3598 , g3599 , g3600 , g3601 , g3602 , g3603 , g3604 , g3605 , g3606 , g3607 , g3608 , g3609 , g3610 , g3611 , g3612 , g3613 , g3614 , g3615 , g3616 , g3617 , g3618 , g3619 , g3620 , g3621 , g3622 , g3623 , g3624 , g3625 , g3626 , g3627 , g3628 , g3629 , g3630 , g3631 , g3632 , g3633 , g3634 , g3635 , g3636 , g3637 , g3638 , g3639 , g3640 , g3641 , g3642 , g3643 , g3644 , g3645 , g3646 , g3647 , g3648 , g3649 , g3650 , g3651 , g3652 , g3653 , g3654 , g3655 , g3656 , g3657 , g3658 , g3659 , g3660 , g3661 , g3662 , g3663 , g3664 , g3665 , g3666 , g3667 , g3668 , g3669 , g3670 , g3671 , g3672 , g3673 , g3674 , g3675 , g3676 , g3677 , g3678 , g3679 , g3680 , g3681 , g3682 , g3683 , g3684 , g3685 , g3686 , g3687 , g3688 , g3689 , g3690 , g3691 , g3692 , g3693 , g3694 , g3695 , g3696 , g3697 , g3698 , g3699 , g3700 , g3701 , g3702 , g3703 , g3704 , g3705 , g3706 , g3707 , g3708 , g3709 , g3710 , g3711 , g3712 , g3713 , g3714 , g3715 , g3716 , g3717 , g3718 , g3719 , g3720 , g3721 , g3722 , g3723 , g3724 , g3725 , g3726 , g3727 , g3728 , g3729 , g3730 , g3731 , g3732 , g3733 , g3734 , g3735 , g3736 , g3737 , g3738 , g3739 , g3740 , g3741 , g3742 , g3743 , g3744 , g3745 , g3746 , g3747 , g3748 , g3749 , g3750 , g3751 , g3752 , g3753 , g3754 , g3755 , g3756 , g3757 , g3758 , g3759 , g3760 , g3761 , g3762 , g3763 , g3764 , g3765 , g3766 , g3767 , g3768 , g3769 , g3770 , g3771 , g3772 , g3773 , g3774 , g3775 , g3776 , g3777 , g3778 , g3779 , g3780 , g3781 , g3782 , g3783 , g3784 , g3785 , g3786 , g3787 , g3788 , g3789 , g3790 , g3791 , g3792 , g3793 , g3794 , g3795 , g3796 , g3797 , g3798 , g3799 , g3800 , g3801 , g3802 , g3803 , g3804 , g3805 , g3806 , g3807 , g3808 , g3809 , g3810 , g3811 , g3812 , g3813 , g3814 , g3815 , g3816 , g3817 , g3818 , g3819 , g3820 , g3821 , g3822 , g3823 , g3824 , g3825 , g3826 , g3827 , g3828 , g3829 , g3830 , g3831 , g3832 , g3833 , g3834 , g3835 , g3836 , g3837 , g3838 , g3839 , g3840 , g3841 , g3842 , g3843 , g3844 , g3845 , g3846 , g3847 , g3848 , g3849 , g3850 , g3851 , g3852 , g3853 , g3854 , g3855 , g3856 , g3857 , g3858 , g3859 , g3860 , g3861 , g3862 , g3863 , g3864 , g3865 , g3866 , g3867 , g3868 , g3869 , g3870 , g3871 , g3872 , g3873 , g3874 , g3875 , g3876 , g3877 , g3878 , g3879 , g3880 , g3881 , g3882 , g3883 , g3884 , g3885 , g3886 , g3887 , g3888 , g3889 , g3890 , g3891 , g3892 , g3893 , g3894 , g3895 , g3896 , g3897 , g3898 , g3899 , g3900 , g3901 , g3902 , g3903 , g3904 , g3905 , g3906 , g3907 , g3908 , g3909 , g3910 , g3911 , g3912 , g3913 , g3914 , g3915 , g3916 , g3917 , g3918 , g3919 , g3920 , g3921 , g3922 , g3923 , g3924 , g3925 , g3926 , g3927 , g3928 , g3929 , g3930 , g3931 , g3932 , g3933 , g3934 , g3935 , g3936 , g3937 , g3938 , g3939 , g3940 , g3941 , g3942 , g3943 , g3944 , g3945 , g3946 , g3947 , g3948 , g3949 , g3950 , g3951 , g3952 , g3953 , g3954 , g3955 , g3956 , g3957 , g3958 , g3959 , g3960 , g3961 , g3962 , g3963 , g3964 , g3965 , g3966 , g3967 , g3968 , g3969 , g3970 , g3971 , g3972 , g3973 , g3974 , g3975 , g3976 , g3977 , g3978 , g3979 , g3980 , g3981 , g3982 , g3983 , g3984 , g3985 , g3986 , g3987 , g3988 , g3989 , g3990 , g3991 , g3992 , g3993 , g3994 , g3995 , g3996 , g3997 , g3998 , g3999 , g4000 , g4001 , g4002 , g4003 , g4004 , g4005 , g4006 , g4007 , g4008 , g4009 , g4010 , g4011 , g4012 , g4013 , g4014 , g4015 , g4016 , g4017 , g4018 , g4019 , g4020 , g4021 , g4022 , g4023 , g4024 , g4025 , g4026 , g4027 , g4028 , g4029 , g4030 , g4031 , g4032 , g4033 , g4034 , g4035 , g4036 , g4037 , g4038 , g4039 , g4040 , g4041 , g4042 , g4043 , g4044 , g4045 , g4046 , g4047 , g4048 , g4049 , g4050 , g4051 , g4052 , g4053 , g4054 , g4055 , g4056 , g4057 , g4058 , g4059 , g4060 , g4061 , g4062 , g4063 , g4064 , g4065 , g4066 , g4067 , g4068 , g4069 , g4070 , g4071 , g4072 , g4073 , g4074 , g4075 , g4076 , g4077 , g4078 , g4079 , g4080 , g4081 , g4082 , g4083 , g4084 , g4085 , g4086 , g4087 , g4088 , g4089 , g4090 , g4091 , g4092 , g4093 , g4094 , g4095 , g4096 , g4097 , g4098 , g4099 , g4100 , g4101 , g4102 , g4103 , g4104 , g4105 , g4106 , g4107 , g4108 , g4109 , g4110 , g4111 , g4112 , g4113 , g4114 , g4115 , g4116 , g4117 , g4118 , g4119 , g4120 , g4121 , g4122 , g4123 , g4124 , g4125 , g4126 , g4127 , g4128 , g4129 , g4130 , g4131 , g4132 , g4133 , g4134 , g4135 , g4136 , g4137 , g4138 , g4139 , g4140 , g4141 , g4142 , g4143 , g4144 , g4145 , g4146 , g4147 , g4148 , g4149 , g4150 , g4151 , g4152 , g4153 , g4154 , g4155 , g4156 , g4157 , g4158 , g4159 , g4160 , g4161 , g4162 , g4163 , g4164 , g4165 , g4166 , g4167 , g4168 , g4169 , g4170 , g4171 , g4172 , g4173 , g4174 , g4175 , g4176 , g4177 , g4178 , g4179 , g4180 , g4181 , g4182 , g4183 , g4184 , g4185 , g4186 , g4187 , g4188 , g4189 , g4190 , g4191 , g4192 , g4193 , g4194 , g4195 , g4196 , g4197 , g4198 , g4199 , g4200 , g4201 , g4202 , g4203 , g4204 , g4205 , g4206 , g4207 , g4208 , g4209 , g4210 , g4211 , g4212 , g4213 , g4214 , g4215 , g4216 , g4217 , g4218 , g4219 , g4220 , g4221 , g4222 , g4223 , g4224 , g4225 , g4226 , g4227 , g4228 , g4229 , g4230 , g4231 , g4232 , g4233 , g4234 , g4235 , g4236 , g4237 , g4238 , g4239 , g4240 , g4241 , g4242 , g4243 , g4244 , g4245 , g4246 , g4247 , g4248 , g4249 , g4250 , g4251 , g4252 , g4253 , g4254 , g4255 , g4256 , g4257 , g4258 , g4259 , g4260 , g4261 , g4262 , g4263 , g4264 , g4265 , g4266 , g4267 , g4268 , g4269 , g4270 , g4271 , g4272 , g4273 , g4274 , g4275 , g4276 , g4277 , g4278 , g4279 , g4280 , g4281 , g4282 , g4283 , g4284 , g4285 , g4286 , g4287 , g4288 , g4289 , g4290 , g4291 , g4292 , g4293 , g4294 , g4295 , g4296 , g4297 , g4298 , g4299 , g4300 , g4301 , g4302 , g4303 , g4304 , g4305 , g4306 , g4307 , g4308 , g4309 , g4310 , g4311 , g4312 , g4313 , g4314 , g4315 , g4316 , g4317 , g4318 , g4319 , g4320 , g4321 , g4322 , g4323 , g4324 , g4325 , g4326 , g4327 , g4328 , g4329 , g4330 , g4331 , g4332 , g4333 , g4334 , g4335 , g4336 , g4337 , g4338 , g4339 , g4340 , g4341 , g4342 , g4343 , g4344 , g4345 , g4346 , g4347 , g4348 , g4349 , g4350 , g4351 , g4352 , g4353 , g4354 , g4355 , g4356 , g4357 , g4358 , g4359 , g4360 , g4361 , g4362 , g4363 , g4364 , g4365 , g4366 , g4367 , g4368 , g4369 , g4370 , g4371 , g4372 , g4373 , g4374 , g4375 , g4376 , g4377 , g4378 , g4379 , g4380 , g4381 , g4382 , g4383 , g4384 , g4385 , g4386 , g4387 , g4388 , g4389 , g4390 , g4391 , g4392 , g4393 , g4394 , g4395 , g4396 , g4397 , g4398 , g4399 , g4400 , g4401 , g4402 , g4403 , g4404 , g4405 , g4406 , g4407 , g4408 , g4409 , g4410 , g4411 , g4412 , g4413 , g4414 , g4415 , g4416 , g4417 , g4418 , g4419 , g4420 , g4421 , g4422 , g4423 , g4424 , g4425 , g4426 , g4427 , g4428 , g4429 , g4430 , g4431 , g4432 , g4433 , g4434 , g4435 , g4436 , g4437 , g4438 , g4439 , g4440 , g4441 , g4442 , g4443 , g4444 , g4445 , g4446 , g4447 , g4448 , g4449 , g4450 , g4451 , g4452 , g4453 , g4454 , g4455 , g4456 , g4457 , g4458 , g4459 , g4460 , g4461 , g4462 , g4463 , g4464 , g4465 , g4466 , g4467 , g4468 , g4469 , g4470 , g4471 , g4472 , g4473 , g4474 , g4475 , g4476 , g4477 , g4478 , g4479 , g4480 , g4481 , g4482 , g4483 , g4484 , g4485 , g4486 , g4487 , g4488 , g4489 , g4490 , g4491 , g4492 , g4493 , g4494 , g4495 , g4496 , g4497 , g4498 , g4499 , g4500 , g4501 , g4502 , g4503 , g4504 , g4505 , g4506 , g4507 , g4508 , g4509 , g4510 , g4511 , g4512 , g4513 , g4514 , g4515 , g4516 , g4517 , g4518 , g4519 , g4520 , g4521 , g4522 , g4523 , g4524 , g4525 , g4526 , g4527 , g4528 , g4529 , g4530 , g4531 , g4532 , g4533 , g4534 , g4535 , g4536 , g4537 , g4538 , g4539 , g4540 , g4541 , g4542 , g4543 , g4544 , g4545 , g4546 , g4547 , g4548 , g4549 , g4550 , g4551 , g4552 , g4553 , g4554 , g4555 , g4556 , g4557 , g4558 , g4559 , g4560 , g4561 , g4562 , g4563 , g4564 , g4565 , g4566 , g4567 , g4568 , g4569 , g4570 , g4571 , g4572 , g4573 , g4574 , g4575 , g4576 , g4577 , g4578 , g4579 , g4580 , g4581 , g4582 , g4583 , g4584 , g4585 , g4586 , g4587 , g4588 , g4589 , g4590 , g4591 , g4592 , g4593 , g4594 , g4595 , g4596 , g4597 , g4598 , g4599 , g4600 , g4601 , g4602 , g4603 , g4604 , g4605 , g4606 , g4607 , g4608 , g4609 , g4610 , g4611 , g4612 , g4613 , g4614 , g4615 , g4616 , g4617 , g4618 , g4619 , g4620 , g4621 , g4622 , g4623 , g4624 , g4625 , g4626 , g4627 , g4628 , g4629 , g4630 , g4631 , g4632 , g4633 , g4634 , g4635 , g4636 , g4637 , g4638 , g4639 , g4640 , g4641 , g4642 , g4643 , g4644 , g4645 , g4646 , g4647 , g4648 , g4649 , g4650 , g4651 , g4652 , g4653 , g4654 , g4655 , g4656 , g4657 , g4658 , g4659 , g4660 , g4661 , g4662 , g4663 , g4664 , g4665 , g4666 , g4667 , g4668 , g4669 , g4670 , g4671 , g4672 , g4673 , g4674 , g4675 , g4676 , g4677 , g4678 , g4679 , g4680 , g4681 , g4682 , g4683 , g4684 , g4685 , g4686 , g4687 , g4688 , g4689 , g4690 , g4691 , g4692 , g4693 , g4694 , g4695 , g4696 , g4697 , g4698 , g4699 , g4700 , g4701 , g4702 , g4703 , g4704 , g4705 , g4706 , g4707 , g4708 , g4709 , g4710 , g4711 , g4712 , g4713 , g4714 , g4715 , g4716 , g4717 , g4718 , g4719 , g4720 , g4721 , g4722 , g4723 , g4724 , g4725 , g4726 , g4727 , g4728 , g4729 , g4730 , g4731 , g4732 , g4733 , g4734 , g4735 , g4736 , g4737 , g4738 , g4739 , g4740 , g4741 , g4742 , g4743 , g4744 , g4745 , g4746 , g4747 , g4748 , g4749 , g4750 , g4751 , g4752 , g4753 , g4754 , g4755 , g4756 , g4757 , g4758 , g4759 , g4760 , g4761 , g4762 , g4763 , g4764 , g4765 , g4766 , g4767 , g4768 , g4769 , g4770 , g4771 , g4772 , g4773 , g4774 , g4775 , g4776 , g4777 , g4778 , g4779 , g4780 , g4781 , g4782 , g4783 , g4784 , g4785 , g4786 , g4787 , g4788 , g4789 , g4790 , g4791 , g4792 , g4793 , g4794 , g4795 , g4796 , g4797 , g4798 , g4799 , g4800 , g4801 , g4802 , g4803 , g4804 , g4805 , g4806 , g4807 , g4808 , g4809 , g4810 , g4811 , g4812 , g4813 , g4814 , g4815 , g4816 , g4817 , g4818 , g4819 , g4820 , g4821 , g4822 , g4823 , g4824 , g4825 , g4826 , g4827 , g4828 , g4829 , g4830 , g4831 , g4832 , g4833 , g4834 , g4835 , g4836 , g4837 , g4838 , g4839 , g4840 , g4841 , g4842 , g4843 , g4844 , g4845 , g4846 , g4847 , g4848 , g4849 , g4850 , g4851 , g4852 , g4853 , g4854 , g4855 , g4856 , g4857 , g4858 , g4859 , g4860 , g4861 , g4862 , g4863 , g4864 , g4865 , g4866 , g4867 , g4868 , g4869 , g4870 , g4871 , g4872 , g4873 , g4874 , g4875 , g4876 , g4877 , g4878 , g4879 , g4880 , g4881 , g4882 , g4883 , g4884 , g4885 , g4886 , g4887 , g4888 , g4889 , g4890 , g4891 , g4892 , g4893 , g4894 , g4895 , g4896 , g4897 , g4898 , g4899 , g4900 , g4901 , g4902 , g4903 , g4904 , g4905 , g4906 , g4907 , g4908 , g4909 , g4910 , g4911 , g4912 , g4913 , g4914 , g4915 , g4916 , g4917 , g4918 , g4919 , g4920 , g4921 , g4922 , g4923 , g4924 , g4925 , g4926 , g4927 , g4928 , g4929 , g4930 , g4931 , g4932 , g4933 , g4934 , g4935 , g4936 , g4937 , g4938 , g4939 , g4940 , g4941 , g4942 , g4943 , g4944 , g4945 , g4946 , g4947 , g4948 , g4949 , g4950 , g4951 , g4952 , g4953 , g4954 , g4955 , g4956 , g4957 , g4958 , g4959 , g4960 , g4961 , g4962 , g4963 , g4964 , g4965 , g4966 , g4967 , g4968 , g4969 , g4970 , g4971 , g4972 , g4973 , g4974 , g4975 , g4976 , g4977 , g4978 , g4979 , g4980 , g4981 , g4982 , g4983 , g4984 , g4985 , g4986 , g4987 , g4988 , g4989 , g4990 , g4991 , g4992 , g4993 , g4994 , g4995 , g4996 , g4997 , g4998 , g4999 , g5000 , g5001 , g5002 , g5003 , g5004 , g5005 , g5006 , g5007 , g5008 , g5009 , g5010 , g5011 , g5012 , g5013 , g5014 , g5015 , g5016 , g5017 , g5018 , g5019 , g5020 , g5021 , g5022 , g5023 , g5024 , g5025 , g5026 , g5027 , g5028 , g5029 , g5030 , g5031 , g5032 , g5033 , g5034 , g5035 , g5036 , g5037 , g5038 , g5039 , g5040 , g5041 , g5042 , g5043 , g5044 , g5045 , g5046 , g5047 , g5048 , g5049 , g5050 , g5051 , g5052 , g5053 , g5054 , g5055 , g5056 , g5057 , g5058 , g5059 , g5060 , g5061 , g5062 , g5063 , g5064 , g5065 , g5066 , g5067 , g5068 , g5069 , g5070 , g5071 , g5072 , g5073 , g5074 , g5075 , g5076 , g5077 , g5078 , g5079 , g5080 , g5081 , g5082 , g5083 , g5084 , g5085 , g5086 , g5087 , g5088 , g5089 , g5090 , g5091 , g5092 , g5093 , g5094 , g5095 , g5096 , g5097 , g5098 , g5099 , g5100 , g5101 , g5102 , g5103 , g5104 , g5105 , g5106 , g5107 , g5108 , g5109 , g5110 , g5111 , g5112 , g5113 , g5114 , g5115 , g5116 , g5117 , g5118 , g5119 , g5120 , g5121 , g5122 , g5123 , g5124 , g5125 , g5126 , g5127 , g5128 , g5129 , g5130 , g5131 , g5132 , g5133 , g5134 , g5135 , g5136 , g5137 , g5138 , g5139 , g5140 , g5141 , g5142 , g5143 , g5144 , g5145 , g5146 , g5147 , g5148 , g5149 , g5150 , g5151 , g5152 , g5153 , g5154 , g5155 , g5156 , g5157 , g5158 , g5159 , g5160 , g5161 , g5162 , g5163 , g5164 , g5165 , g5166 , g5167 , g5168 , g5169 , g5170 , g5171 , g5172 , g5173 , g5174 , g5175 , g5176 , g5177 , g5178 , g5179 , g5180 , g5181 , g5182 , g5183 , g5184 , g5185 , g5186 , g5187 , g5188 , g5189 , g5190 , g5191 , g5192 , g5193 , g5194 , g5195 , g5196 , g5197 , g5198 , g5199 , g5200 , g5201 , g5202 , g5203 , g5204 , g5205 , g5206 , g5207 , g5208 , g5209 , g5210 , g5211 , g5212 , g5213 , g5214 , g5215 , g5216 , g5217 , g5218 , g5219 , g5220 , g5221 , g5222 , g5223 , g5224 , g5225 , g5226 , g5227 , g5228 , g5229 , g5230 , g5231 , g5232 , g5233 , g5234 , g5235 , g5236 , g5237 , g5238 , g5239 , g5240 , g5241 , g5242 , g5243 , g5244 , g5245 , g5246 , g5247 , g5248 , g5249 , g5250 , g5251 , g5252 , g5253 , g5254 , g5255 , g5256 , g5257 , g5258 , g5259 , g5260 , g5261 , g5262 , g5263 , g5264 , g5265 , g5266 , g5267 , g5268 , g5269 , g5270 , g5271 , g5272 , g5273 , g5274 , g5275 , g5276 , g5277 , g5278 , g5279 , g5280 , g5281 , g5282 , g5283 , g5284 , g5285 , g5286 , g5287 , g5288 , g5289 , g5290 , g5291 , g5292 , g5293 , g5294 , g5295 , g5296 , g5297 , g5298 , g5299 , g5300 , g5301 , g5302 , g5303 , g5304 , g5305 , g5306 , g5307 , g5308 , g5309 , g5310 , g5311 , g5312 , g5313 , g5314 , g5315 , g5316 , g5317 , g5318 , g5319 , g5320 , g5321 , g5322 , g5323 , g5324 , g5325 , g5326 , g5327 , g5328 , g5329 , g5330 , g5331 , g5332 , g5333 , g5334 , g5335 , g5336 , g5337 , g5338 , g5339 , g5340 , g5341 , g5342 , g5343 , g5344 , g5345 , g5346 , g5347 , g5348 , g5349 , g5350 , g5351 , g5352 , g5353 , g5354 , g5355 , g5356 , g5357 , g5358 , g5359 , g5360 , g5361 , g5362 , g5363 , g5364 , g5365 , g5366 , g5367 , g5368 , g5369 , g5370 , g5371 , g5372 , g5373 , g5374 , g5375 , g5376 , g5377 , g5378 , g5379 , g5380 , g5381 , g5382 , g5383 , g5384 , g5385 , g5386 , g5387 , g5388 , g5389 , g5390 , g5391 , g5392 , g5393 , g5394 , g5395 , g5396 , g5397 , g5398 , g5399 , g5400 , g5401 , g5402 , g5403 , g5404 , g5405 , g5406 , g5407 , g5408 , g5409 , g5410 , g5411 , g5412 , g5413 , g5414 , g5415 , g5416 , g5417 , g5418 , g5419 , g5420 , g5421 , g5422 , g5423 , g5424 , g5425 , g5426 , g5427 , g5428 , g5429 , g5430 , g5431 , g5432 , g5433 , g5434 , g5435 , g5436 , g5437 , g5438 , g5439 , g5440 , g5441 , g5442 , g5443 , g5444 , g5445 , g5446 , g5447 , g5448 , g5449 , g5450 , g5451 , g5452 , g5453 , g5454 , g5455 , g5456 , g5457 , g5458 , g5459 , g5460 , g5461 , g5462 , g5463 , g5464 , g5465 , g5466 , g5467 , g5468 , g5469 , g5470 , g5471 , g5472 , g5473 , g5474 , g5475 , g5476 , g5477 , g5478 , g5479 , g5480 , g5481 , g5482 , g5483 , g5484 , g5485 , g5486 , g5487 , g5488 , g5489 , g5490 , g5491 , g5492 , g5493 , g5494 , g5495 , g5496 , g5497 , g5498 , g5499 , g5500 , g5501 , g5502 , g5503 , g5504 , g5505 , g5506 , g5507 , g5508 , g5509 , g5510 , g5511 , g5512 , g5513 , g5514 , g5515 , g5516 , g5517 , g5518 , g5519 , g5520 , g5521 , g5522 , g5523 , g5524 , g5525 , g5526 , g5527 , g5528 , g5529 , g5530 , g5531 , g5532 , g5533 , g5534 , g5535 , g5536 , g5537 , g5538 , g5539 , g5540 , g5541 , g5542 , g5543 , g5544 , g5545 , g5546 , g5547 , g5548 , g5549 , g5550 , g5551 , g5552 , g5553 , g5554 , g5555 , g5556 , g5557 , g5558 , g5559 , g5560 , g5561 , g5562 , g5563 , g5564 , g5565 , g5566 , g5567 , g5568 , g5569 , g5570 , g5571 , g5572 , g5573 , g5574 , g5575 , g5576 , g5577 , g5578 , g5579 , g5580 , g5581 , g5582 , g5583 , g5584 , g5585 , g5586 , g5587 , g5588 , g5589 , g5590 , g5591 , g5592 , g5593 , g5594 , g5595 , g5596 , g5597 , g5598 , g5599 , g5600 , g5601 , g5602 , g5603 , g5604 , g5605 , g5606 , g5607 , g5608 , g5609 , g5610 , g5611 , g5612 , g5613 , g5614 , g5615 , g5616 , g5617 , g5618 , g5619 , g5620 , g5621 , g5622 , g5623 , g5624 , g5625 , g5626 , g5627 , g5628 , g5629 , g5630 , g5631 , g5632 , g5633 , g5634 , g5635 , g5636 , g5637 , g5638 , g5639 , g5640 , g5641 , g5642 , g5643 , g5644 , g5645 , g5646 , g5647 , g5648 , g5649 , g5650 , g5651 , g5652 , g5653 , g5654 , g5655 , g5656 , g5657 , g5658 , g5659 , g5660 , g5661 , g5662 , g5663 , g5664 , g5665 , g5666 , g5667 , g5668 , g5669 , g5670 , g5671 , g5672 , g5673 , g5674 , g5675 , g5676 , g5677 , g5678 , g5679 , g5680 , g5681 , g5682 , g5683 , g5684 , g5685 , g5686 , g5687 , g5688 , g5689 , g5690 , g5691 , g5692 , g5693 , g5694 , g5695 , g5696 , g5697 , g5698 , g5699 , g5700 , g5701 , g5702 , g5703 , g5704 , g5705 , g5706 , g5707 , g5708 , g5709 , g5710 , g5711 , g5712 , g5713 , g5714 , g5715 , g5716 , g5717 , g5718 , g5719 , g5720 , g5721 , g5722 , g5723 , g5724 , g5725 , g5726 , g5727 , g5728 , g5729 , g5730 , g5731 , g5732 , g5733 , g5734 , g5735 , g5736 , g5737 , g5738 , g5739 , g5740 , g5741 , g5742 , g5743 , g5744 , g5745 , g5746 , g5747 , g5748 , g5749 , g5750 , g5751 , g5752 , g5753 , g5754 , g5755 , g5756 , g5757 , g5758 , g5759 , g5760 , g5761 , g5762 , g5763 , g5764 , g5765 , g5766 , g5767 , g5768 , g5769 , g5770 , g5771 , g5772 , g5773 , g5774 , g5775 , g5776 , g5777 , g5778 , g5779 , g5780 , g5781 , g5782 , g5783 , g5784 , g5785 , g5786 , g5787 , g5788 , g5789 , g5790 , g5791 , g5792 , g5793 , g5794 , g5795 , g5796 , g5797 , g5798 , g5799 , g5800 , g5801 , g5802 , g5803 , g5804 , g5805 , g5806 , g5807 , g5808 , g5809 , g5810 , g5811 , g5812 , g5813 , g5814 , g5815 , g5816 , g5817 , g5818 , g5819 , g5820 , g5821 , g5822 , g5823 , g5824 , g5825 , g5826 , g5827 , g5828 , g5829 , g5830 , g5831 , g5832 , g5833 , g5834 , g5835 , g5836 , g5837 , g5838 , g5839 , g5840 , g5841 , g5842 , g5843 , g5844 , g5845 , g5846 , g5847 , g5848 , g5849 , g5850 , g5851 , g5852 , g5853 , g5854 , g5855 , g5856 , g5857 , g5858 , g5859 , g5860 , g5861 , g5862 , g5863 , g5864 , g5865 , g5866 , g5867 , g5868 , g5869 , g5870 , g5871 , g5872 , g5873 , g5874 , g5875 , g5876 , g5877 , g5878 , g5879 , g5880 , g5881 , g5882 , g5883 , g5884 , g5885 , g5886 , g5887 , g5888 , g5889 , g5890 , g5891 , g5892 , g5893 , g5894 , g5895 , g5896 , g5897 , g5898 , g5899 , g5900 , g5901 , g5902 , g5903 , g5904 , g5905 , g5906 , g5907 , g5908 , g5909 , g5910 , g5911 , g5912 , g5913 , g5914 , g5915 , g5916 , g5917 , g5918 , g5919 , g5920 , g5921 , g5922 , g5923 , g5924 , g5925 , g5926 , g5927 , g5928 , g5929 , g5930 , g5931 , g5932 , g5933 , g5934 , g5935 , g5936 , g5937 , g5938 , g5939 , g5940 , g5941 , g5942 , g5943 , g5944 , g5945 , g5946 , g5947 , g5948 , g5949 , g5950 , g5951 , g5952 , g5953 , g5954 , g5955 , g5956 , g5957 , g5958 , g5959 , g5960 , g5961 , g5962 , g5963 , g5964 , g5965 , g5966 , g5967 , g5968 , g5969 , g5970 , g5971 , g5972 , g5973 , g5974 , g5975 , g5976 , g5977 , g5978 , g5979 , g5980 , g5981 , g5982 , g5983 , g5984 , g5985 , g5986 , g5987 , g5988 , g5989 , g5990 , g5991 , g5992 , g5993 , g5994 , g5995 , g5996 , g5997 , g5998 , g5999 , g6000 , g6001 , g6002 , g6003 , g6004 , g6005 , g6006 , g6007 , g6008 , g6009 , g6010 , g6011 , g6012 , g6013 , g6014 , g6015 , g6016 , g6017 , g6018 , g6019 , g6020 , g6021 , g6022 , g6023 , g6024 , g6025 , g6026 , g6027 , g6028 , g6029 , g6030 , g6031 , g6032 , g6033 , g6034 , g6035 , g6036 , g6037 , g6038 , g6039 , g6040 , g6041 , g6042 , g6043 , g6044 , g6045 , g6046 , g6047 , g6048 , g6049 , g6050 , g6051 , g6052 , g6053 , g6054 , g6055 , g6056 , g6057 , g6058 , g6059 , g6060 , g6061 , g6062 , g6063 , g6064 , g6065 , g6066 , g6067 , g6068 , g6069 , g6070 , g6071 , g6072 , g6073 , g6074 , g6075 , g6076 , g6077 , g6078 , g6079 , g6080 , g6081 , g6082 , g6083 , g6084 , g6085 , g6086 , g6087 , g6088 , g6089 , g6090 , g6091 , g6092 , g6093 , g6094 , g6095 , g6096 , g6097 , g6098 , g6099 , g6100 , g6101 , g6102 , g6103 , g6104 , g6105 , g6106 , g6107 , g6108 , g6109 , g6110 , g6111 , g6112 , g6113 , g6114 , g6115 , g6116 , g6117 , g6118 , g6119 , g6120 , g6121 , g6122 , g6123 , g6124 , g6125 , g6126 , g6127 , g6128 , g6129 , g6130 , g6131 , g6132 , g6133 , g6134 , g6135 , g6136 , g6137 , g6138 , g6139 , g6140 , g6141 , g6142 , g6143 , g6144 , g6145 , g6146 , g6147 , g6148 , g6149 , g6150 , g6151 , g6152 , g6153 , g6154 , g6155 , g6156 , g6157 , g6158 , g6159 , g6160 , g6161 , g6162 , g6163 , g6164 , g6165 , g6166 , g6167 , g6168 , g6169 , g6170 , g6171 , g6172 , g6173 , g6174 , g6175 , g6176 , g6177 , g6178 , g6179 , g6180 , g6181 , g6182 , g6183 , g6184 , g6185 , g6186 , g6187 , g6188 , g6189 , g6190 , g6191 , g6192 , g6193 , g6194 , g6195 , g6196 , g6197 , g6198 , g6199 , g6200 , g6201 , g6202 , g6203 , g6204 , g6205 , g6206 , g6207 , g6208 , g6209 , g6210 , g6211 , g6212 , g6213 , g6214 , g6215 , g6216 , g6217 , g6218 , g6219 , g6220 , g6221 , g6222 , g6223 , g6224 , g6225 , g6226 , g6227 , g6228 , g6229 , g6230 , g6231 , g6232 , g6233 , g6234 , g6235 , g6236 , g6237 , g6238 , g6239 , g6240 , g6241 , g6242 , g6243 , g6244 , g6245 , g6246 , g6247 , g6248 , g6249 , g6250 , g6251 , g6252 , g6253 , g6254 , g6255 , g6256 , g6257 , g6258 , g6259 , g6260 , g6261 , g6262 , g6263 , g6264 , g6265 , g6266 , g6267 , g6268 , g6269 , g6270 , g6271 , g6272 , g6273 , g6274 , g6275 , g6276 , g6277 , g6278 , g6279 , g6280 , g6281 , g6282 , g6283 , g6284 , g6285 , g6286 , g6287 , g6288 , g6289 , g6290 , g6291 , g6292 , g6293 , g6294 , g6295 , g6296 , g6297 , g6298 , g6299 , g6300 , g6301 , g6302 , g6303 , g6304 , g6305 , g6306 , g6307 , g6308 , g6309 , g6310 , g6311 , g6312 , g6313 , g6314 , g6315 , g6316 , g6317 , g6318 , g6319 , g6320 , g6321 , g6322 , g6323 , g6324 , g6325 , g6326 , g6327 , g6328 , g6329 , g6330 , g6331 , g6332 , g6333 , g6334 , g6335 , g6336 , g6337 , g6338 , g6339 , g6340 , g6341 , g6342 , g6343 , g6344 , g6345 , g6346 , g6347 , g6348 , g6349 , g6350 , g6351 , g6352 , g6353 , g6354 , g6355 , g6356 , g6357 , g6358 , g6359 , g6360 , g6361 , g6362 , g6363 , g6364 , g6365 , g6366 , g6367 , g6368 , g6369 , g6370 , g6371 , g6372 , g6373 , g6374 , g6375 , g6376 , g6377 , g6378 , g6379 , g6380 , g6381 , g6382 , g6383 , g6384 , g6385 , g6386 , g6387 , g6388 , g6389 , g6390 , g6391 , g6392 , g6393 , g6394 , g6395 , g6396 , g6397 , g6398 , g6399 , g6400 , g6401 , g6402 , g6403 , g6404 , g6405 , g6406 , g6407 , g6408 , g6409 , g6410 , g6411 , g6412 , g6413 , g6414 , g6415 , g6416 , g6417 , g6418 , g6419 , g6420 , g6421 , g6422 , g6423 , g6424 , g6425 , g6426 , g6427 , g6428 , g6429 , g6430 , g6431 , g6432 , g6433 , g6434 , g6435 , g6436 , g6437 , g6438 , g6439 , g6440 , g6441 , g6442 , g6443 , g6444 , g6445 , g6446 , g6447 , g6448 , g6449 , g6450 , g6451 , g6452 , g6453 , g6454 , g6455 , g6456 , g6457 , g6458 , g6459 , g6460 , g6461 , g6462 , g6463 , g6464 , g6465 , g6466 , g6467 , g6468 , g6469 , g6470 , g6471 , g6472 , g6473 , g6474 , g6475 , g6476 , g6477 , g6478 , g6479 , g6480 , g6481 , g6482 , g6483 , g6484 , g6485 , g6486 , g6487 , g6488 , g6489 , g6490 , g6491 , g6492 , g6493 , g6494 , g6495 , g6496 , g6497 , g6498 , g6499 , g6500 , g6501 , g6502 , g6503 , g6504 , g6505 , g6506 , g6507 , g6508 , g6509 , g6510 , g6511 , g6512 , g6513 , g6514 , g6515 , g6516 , g6517 , g6518 , g6519 , g6520 , g6521 , g6522 , g6523 , g6524 , g6525 , g6526 , g6527 , g6528 , g6529 , g6530 , g6531 , g6532 , g6533 , g6534 , g6535 , g6536 , g6537 , g6538 , g6539 , g6540 , g6541 , g6542 , g6543 , g6544 , g6545 , g6546 , g6547 , g6548 , g6549 , g6550 , g6551 , g6552 , g6553 , g6554 , g6555 , g6556 , g6557 , g6558 , g6559 , g6560 , g6561 , g6562 , g6563 , g6564 , g6565 , g6566 , g6567 , g6568 , g6569 , g6570 , g6571 , g6572 , g6573 , g6574 , g6575 , g6576 , g6577 , g6578 , g6579 , g6580 , g6581 , g6582 , g6583 , g6584 , g6585 , g6586 , g6587 , g6588 , g6589 , g6590 , g6591 , g6592 , g6593 , g6594 , g6595 , g6596 , g6597 , g6598 , g6599 , g6600 , g6601 , g6602 , g6603 , g6604 , g6605 , g6606 , g6607 , g6608 , g6609 , g6610 , g6611 , g6612 , g6613 , g6614 , g6615 , g6616 , g6617 , g6618 , g6619 , g6620 , g6621 , g6622 , g6623 , g6624 , g6625 , g6626 , g6627 , g6628 , g6629 , g6630 , g6631 , g6632 , g6633 , g6634 , g6635 , g6636 , g6637 , g6638 , g6639 , g6640 , g6641 , g6642 , g6643 , g6644 , g6645 , g6646 , g6647 , g6648 , g6649 , g6650 , g6651 , g6652 , g6653 , g6654 , g6655 , g6656 , g6657 , g6658 , g6659 , g6660 , g6661 , g6662 , g6663 , g6664 , g6665 , g6666 , g6667 , g6668 , g6669 , g6670 , g6671 , g6672 , g6673 , g6674 , g6675 , g6676 , g6677 , g6678 , g6679 , g6680 , g6681 , g6682 , g6683 , g6684 , g6685 , g6686 , g6687 , g6688 , g6689 , g6690 , g6691 , g6692 , g6693 , g6694 , g6695 , g6696 , g6697 , g6698 , g6699 , g6700 , g6701 , g6702 , g6703 , g6704 , g6705 , g6706 , g6707 , g6708 , g6709 , g6710 , g6711 , g6712 , g6713 , g6714 , g6715 , g6716 , g6717 , g6718 , g6719 , g6720 , g6721 , g6722 , g6723 , g6724 , g6725 , g6726 , g6727 , g6728 , g6729 , g6730 , g6731 , g6732 , g6733 , g6734 , g6735 , g6736 , g6737 , g6738 , g6739 , g6740 , g6741 , g6742 , g6743 , g6744 , g6745 , g6746 , g6747 , g6748 , g6749 , g6750 , g6751 , g6752 , g6753 , g6754 , g6755 , g6756 , g6757 , g6758 , g6759 , g6760 , g6761 , g6762 , g6763 , g6764 , g6765 , g6766 , g6767 , g6768 , g6769 , g6770 , g6771 , g6772 , g6773 , g6774 , g6775 , g6776 , g6777 , g6778 , g6779 , g6780 , g6781 , g6782 , g6783 , g6784 , g6785 , g6786 , g6787 , g6788 , g6789 , g6790 , g6791 , g6792 , g6793 , g6794 , g6795 , g6796 , g6797 , g6798 , g6799 , g6800 , g6801 , g6802 , g6803 , g6804 , g6805 , g6806 , g6807 , g6808 , g6809 , g6810 , g6811 , g6812 , g6813 , g6814 , g6815 , g6816 , g6817 , g6818 , g6819 , g6820 , g6821 , g6822 , g6823 , g6824 , g6825 , g6826 , g6827 , g6828 , g6829 , g6830 , g6831 , g6832 , g6833 , g6834 , g6835 , g6836 , g6837 , g6838 , g6839 , g6840 , g6841 , g6842 , g6843 , g6844 , g6845 , g6846 , g6847 , g6848 , g6849 , g6850 , g6851 , g6852 , g6853 , g6854 , g6855 , g6856 , g6857 , g6858 , g6859 , g6860 , g6861 , g6862 , g6863 , g6864 , g6865 , g6866 , g6867 , g6868 , g6869 , g6870 , g6871 , g6872 , g6873 , g6874 , g6875 , g6876 , g6877 , g6878 , g6879 , g6880 , g6881 , g6882 , g6883 , g6884 , g6885 , g6886 , g6887 , g6888 , g6889 , g6890 , g6891 , g6892 , g6893 , g6894 , g6895 , g6896 , g6897 , g6898 , g6899 , g6900 , g6901 , g6902 , g6903 , g6904 , g6905 , g6906 , g6907 , g6908 , g6909 , g6910 , g6911 , g6912 , g6913 , g6914 , g6915 , g6916 , g6917 , g6918 , g6919 , g6920 , g6921 , g6922 , g6923 , g6924 , g6925 , g6926 , g6927 , g6928 , g6929 , g6930 , g6931 , g6932 , g6933 , g6934 , g6935 , g6936 , g6937 , g6938 , g6939 , g6940 , g6941 , g6942 , g6943 , g6944 , g6945 , g6946 , g6947 , g6948 , g6949 , g6950 , g6951 , g6952 , g6953 , g6954 , g6955 , g6956 , g6957 , g6958 , g6959 , g6960 , g6961 , g6962 , g6963 , g6964 , g6965 , g6966 , g6967 , g6968 , g6969 , g6970 , g6971 , g6972 , g6973 , g6974 , g6975 , g6976 , g6977 , g6978 , g6979 , g6980 , g6981 , g6982 , g6983 , g6984 , g6985 , g6986 , g6987 , g6988 , g6989 , g6990 , g6991 , g6992 , g6993 , g6994 , g6995 , g6996 , g6997 , g6998 , g6999 , g7000 , g7001 , g7002 , g7003 , g7004 , g7005 , g7006 , g7007 , g7008 , g7009 , g7010 , g7011 , g7012 , g7013 , g7014 , g7015 , g7016 , g7017 , g7018 , g7019 , g7020 , g7021 , g7022 , g7023 , g7024 , g7025 , g7026 , g7027 , g7028 , g7029 , g7030 , g7031 , g7032 , g7033 , g7034 , g7035 , g7036 , g7037 , g7038 , g7039 , g7040 , g7041 , g7042 , g7043 , g7044 , g7045 , g7046 , g7047 , g7048 , g7049 , g7050 , g7051 , g7052 , g7053 , g7054 , g7055 , g7056 , g7057 , g7058 , g7059 , g7060 , g7061 , g7062 , g7063 , g7064 , g7065 , g7066 , g7067 , g7068 , g7069 , g7070 , g7071 , g7072 , g7073 , g7074 , g7075 , g7076 , g7077 , g7078 , g7079 , g7080 , g7081 , g7082 , g7083 , g7084 , g7085 , g7086 , g7087 , g7088 , g7089 , g7090 , g7091 , g7092 , g7093 , g7094 , g7095 , g7096 , g7097 , g7098 , g7099 , g7100 , g7101 , g7102 , g7103 , g7104 , g7105 , g7106 , g7107 , g7108 , g7109 , g7110 , g7111 , g7112 , g7113 , g7114 , g7115 , g7116 , g7117 , g7118 , g7119 , g7120 , g7121 , g7122 , g7123 , g7124 , g7125 , g7126 , g7127 , g7128 , g7129 , g7130 , g7131 , g7132 , g7133 , g7134 , g7135 , g7136 , g7137 , g7138 , g7139 , g7140 , g7141 , g7142 , g7143 , g7144 , g7145 , g7146 , g7147 , g7148 , g7149 , g7150 , g7151 , g7152 , g7153 , g7154 , g7155 , g7156 , g7157 , g7158 , g7159 , g7160 , g7161 , g7162 , g7163 , g7164 , g7165 , g7166 , g7167 , g7168 , g7169 , g7170 , g7171 , g7172 , g7173 , g7174 , g7175 , g7176 , g7177 , g7178 , g7179 , g7180 , g7181 , g7182 , g7183 , g7184 , g7185 , g7186 , g7187 , g7188 , g7189 , g7190 , g7191 , g7192 , g7193 , g7194 , g7195 , g7196 , g7197 , g7198 , g7199 , g7200 , g7201 , g7202 , g7203 , g7204 , g7205 , g7206 , g7207 , g7208 , g7209 , g7210 , g7211 , g7212 , g7213 , g7214 , g7215 , g7216 , g7217 , g7218 , g7219 , g7220 , g7221 , g7222 , g7223 , g7224 , g7225 , g7226 , g7227 , g7228 , g7229 , g7230 , g7231 , g7232 , g7233 , g7234 , g7235 , g7236 , g7237 , g7238 , g7239 , g7240 , g7241 , g7242 , g7243 , g7244 , g7245 , g7246 , g7247 , g7248 , g7249 , g7250 , g7251 , g7252 , g7253 , g7254 , g7255 , g7256 , g7257 , g7258 , g7259 , g7260 , g7261 , g7262 , g7263 , g7264 , g7265 , g7266 , g7267 , g7268 , g7269 , g7270 , g7271 , g7272 , g7273 , g7274 , g7275 , g7276 , g7277 , g7278 , g7279 , g7280 , g7281 , g7282 , g7283 , g7284 , g7285 , g7286 , g7287 , g7288 , g7289 , g7290 , g7291 , g7292 , g7293 , g7294 , g7295 , g7296 , g7297 , g7298 , g7299 , g7300 , g7301 , g7302 , g7303 , g7304 , g7305 , g7306 , g7307 , g7308 , g7309 , g7310 , g7311 , g7312 , g7313 , g7314 , g7315 , g7316 , g7317 , g7318 , g7319 , g7320 , g7321 , g7322 , g7323 , g7324 , g7325 , g7326 , g7327 , g7328 , g7329 , g7330 , g7331 , g7332 , g7333 , g7334 , g7335 , g7336 , g7337 , g7338 , g7339 , g7340 , g7341 , g7342 , g7343 , g7344 , g7345 , g7346 , g7347 , g7348 , g7349 , g7350 , g7351 , g7352 , g7353 , g7354 , g7355 , g7356 , g7357 , g7358 , g7359 , g7360 , g7361 , g7362 , g7363 , g7364 , g7365 , g7366 , g7367 , g7368 , g7369 , g7370 , g7371 , g7372 , g7373 , g7374 , g7375 , g7376 , g7377 , g7378 , g7379 , g7380 , g7381 , g7382 , g7383 , g7384 , g7385 , g7386 , g7387 , g7388 , g7389 , g7390 , g7391 , g7392 , g7393 , g7394 , g7395 , g7396 , g7397 , g7398 , g7399 , g7400 , g7401 , g7402 , g7403 , g7404 , g7405 , g7406 , g7407 , g7408 , g7409 , g7410 , g7411 , g7412 , g7413 , g7414 , g7415 , g7416 , g7417 , g7418 , g7419 , g7420 , g7421 , g7422 , g7423 , g7424 , g7425 , g7426 , g7427 , g7428 , g7429 , g7430 , g7431 , g7432 , g7433 , g7434 , g7435 , g7436 , g7437 , g7438 , g7439 , g7440 , g7441 , g7442 , g7443 , g7444 , g7445 , g7446 , g7447 , g7448 , g7449 , g7450 , g7451 , g7452 , g7453 , g7454 , g7455 , g7456 , g7457 , g7458 , g7459 , g7460 , g7461 , g7462 , g7463 , g7464 , g7465 , g7466 , g7467 , g7468 , g7469 , g7470 , g7471 , g7472 , g7473 , g7474 , g7475 , g7476 , g7477 , g7478 , g7479 , g7480 , g7481 , g7482 , g7483 , g7484 , g7485 , g7486 , g7487 , g7488 , g7489 , g7490 , g7491 , g7492 , g7493 , g7494 , g7495 , g7496 , g7497 , g7498 , g7499 , g7500 , g7501 , g7502 , g7503 , g7504 , g7505 , g7506 , g7507 , g7508 , g7509 , g7510 , g7511 , g7512 , g7513 , g7514 , g7515 , g7516 , g7517 , g7518 , g7519 , g7520 , g7521 , g7522 , g7523 , g7524 , g7525 , g7526 , g7527 , g7528 , g7529 , g7530 , g7531 , g7532 , g7533 , g7534 , g7535 , g7536 , g7537 , g7538 , g7539 , g7540 , g7541 , g7542 , g7543 , g7544 , g7545 , g7546 , g7547 , g7548 , g7549 , g7550 , g7551 , g7552 , g7553 , g7554 , g7555 , g7556 , g7557 , g7558 , g7559 , g7560 , g7561 , g7562 , g7563 , g7564 , g7565 , g7566 , g7567 , g7568 , g7569 , g7570 , g7571 , g7572 , g7573 , g7574 , g7575 , g7576 , g7577 , g7578 , g7579 , g7580 , g7581 , g7582 , g7583 , g7584 , g7585 , g7586 , g7587 , g7588 , g7589 , g7590 , g7591 , g7592 , g7593 , g7594 , g7595 , g7596 , g7597 , g7598 , g7599 , g7600 , g7601 , g7602 , g7603 , g7604 , g7605 , g7606 , g7607 , g7608 , g7609 , g7610 , g7611 , g7612 , g7613 , g7614 , g7615 , g7616 , g7617 , g7618 , g7619 , g7620 , g7621 , g7622 , g7623 , g7624 , g7625 , g7626 , g7627 , g7628 , g7629 , g7630 , g7631 , g7632 , g7633 , g7634 , g7635 , g7636 , g7637 , g7638 , g7639 , g7640 , g7641 , g7642 , g7643 , g7644 , g7645 , g7646 , g7647 , g7648 , g7649 , g7650 , g7651 , g7652 , g7653 , g7654 , g7655 , g7656 , g7657 , g7658 , g7659 , g7660 , g7661 , g7662 , g7663 , g7664 , g7665 , g7666 , g7667 , g7668 , g7669 , g7670 , g7671 , g7672 , g7673 , g7674 , g7675 , g7676 , g7677 , g7678 , g7679 , g7680 , g7681 , g7682 , g7683 , g7684 , g7685 , g7686 , g7687 , g7688 , g7689 , g7690 , g7691 , g7692 , g7693 , g7694 , g7695 , g7696 , g7697 , g7698 , g7699 , g7700 , g7701 , g7702 , g7703 , g7704 , g7705 , g7706 , g7707 , g7708 , g7709 , g7710 , g7711 , g7712 , g7713 , g7714 , g7715 , g7716 , g7717 , g7718 , g7719 , g7720 , g7721 , g7722 , g7723 , g7724 , g7725 , g7726 , g7727 , g7728 , g7729 , g7730 , g7731 , g7732 , g7733 , g7734 , g7735 , g7736 , g7737 , g7738 , g7739 , g7740 , g7741 , g7742 , g7743 , g7744 , g7745 , g7746 , g7747 , g7748 , g7749 , g7750 , g7751 , g7752 , g7753 , g7754 , g7755 , g7756 , g7757 , g7758 , g7759 , g7760 , g7761 , g7762 , g7763 , g7764 , g7765 , g7766 , g7767 , g7768 , g7769 , g7770 , g7771 , g7772 , g7773 , g7774 , g7775 , g7776 , g7777 , g7778 , g7779 , g7780 , g7781 , g7782 , g7783 , g7784 , g7785 , g7786 , g7787 , g7788 , g7789 , g7790 , g7791 , g7792 , g7793 , g7794 , g7795 , g7796 , g7797 , g7798 , g7799 , g7800 , g7801 , g7802 , g7803 , g7804 , g7805 , g7806 , g7807 , g7808 , g7809 , g7810 , g7811 , g7812 , g7813 , g7814 , g7815 , g7816 , g7817 , g7818 , g7819 , g7820 , g7821 , g7822 , g7823 , g7824 , g7825 , g7826 , g7827 , g7828 , g7829 , g7830 , g7831 , g7832 , g7833 , g7834 , g7835 , g7836 , g7837 , g7838 , g7839 , g7840 , g7841 , g7842 , g7843 , g7844 , g7845 , g7846 , g7847 , g7848 , g7849 , g7850 , g7851 , g7852 , g7853 , g7854 , g7855 , g7856 , g7857 , g7858 , g7859 , g7860 , g7861 , g7862 , g7863 , g7864 , g7865 , g7866 , g7867 , g7868 , g7869 , g7870 , g7871 , g7872 , g7873 , g7874 , g7875 , g7876 , g7877 , g7878 , g7879 , g7880 , g7881 , g7882 , g7883 , g7884 , g7885 , g7886 , g7887 , g7888 , g7889 , g7890 , g7891 , g7892 , g7893 , g7894 , g7895 , g7896 , g7897 , g7898 , g7899 , g7900 , g7901 , g7902 , g7903 , g7904 , g7905 , g7906 , g7907 , g7908 , g7909 , g7910 , g7911 , g7912 , g7913 , g7914 , g7915 , g7916 , g7917 , g7918 , g7919 , g7920 , g7921 , g7922 , g7923 , g7924 , g7925 , g7926 , g7927 , g7928 , g7929 , g7930 , g7931 , g7932 , g7933 , g7934 , g7935 , g7936 , g7937 , g7938 , g7939 , g7940 , g7941 , g7942 , g7943 , g7944 , g7945 , g7946 , g7947 , g7948 , g7949 , g7950 , g7951 , g7952 , g7953 , g7954 , g7955 , g7956 , g7957 , g7958 , g7959 , g7960 , g7961 , g7962 , g7963 , g7964 , g7965 , g7966 , g7967 , g7968 , g7969 , g7970 , g7971 , g7972 , g7973 , g7974 , g7975 , g7976 , g7977 , g7978 , g7979 , g7980 , g7981 , g7982 , g7983 , g7984 , g7985 , g7986 , g7987 , g7988 , g7989 , g7990 , g7991 , g7992 , g7993 , g7994 , g7995 , g7996 , g7997 , g7998 , g7999 , g8000 , g8001 , g8002 , g8003 , g8004 , g8005 , g8006 , g8007 , g8008 , g8009 , g8010 , g8011 , g8012 , g8013 , g8014 , g8015 , g8016 , g8017 , g8018 , g8019 , g8020 , g8021 , g8022 , g8023 , g8024 , g8025 , g8026 , g8027 , g8028 , g8029 , g8030 , g8031 , g8032 , g8033 , g8034 , g8035 , g8036 , g8037 , g8038 , g8039 , g8040 , g8041 , g8042 , g8043 , g8044 , g8045 , g8046 , g8047 , g8048 , g8049 , g8050 , g8051 , g8052 , g8053 , g8054 , g8055 , g8056 , g8057 , g8058 , g8059 , g8060 , g8061 , g8062 , g8063 , g8064 , g8065 , g8066 , g8067 , g8068 , g8069 , g8070 , g8071 , g8072 , g8073 , g8074 , g8075 , g8076 , g8077 , g8078 , g8079 , g8080 , g8081 , g8082 , g8083 , g8084 , g8085 , g8086 , g8087 , g8088 , g8089 , g8090 , g8091 , g8092 , g8093 , g8094 , g8095 , g8096 , g8097 , g8098 , g8099 , g8100 , g8101 , g8102 , g8103 , g8104 , g8105 , g8106 , g8107 , g8108 , g8109 , g8110 , g8111 , g8112 , g8113 , g8114 , g8115 , g8116 , g8117 , g8118 , g8119 , g8120 , g8121 , g8122 , g8123 , g8124 , g8125 , g8126 , g8127 , g8128 , g8129 , g8130 , g8131 , g8132 , g8133 , g8134 , g8135 , g8136 , g8137 , g8138 , g8139 , g8140 , g8141 , g8142 , g8143 , g8144 , g8145 , g8146 , g8147 , g8148 , g8149 , g8150 , g8151 , g8152 , g8153 , g8154 , g8155 , g8156 , g8157 , g8158 , g8159 , g8160 , g8161 , g8162 , g8163 , g8164 , g8165 , g8166 , g8167 , g8168 , g8169 , g8170 , g8171 , g8172 , g8173 , g8174 , g8175 , g8176 , g8177 , g8178 , g8179 , g8180 , g8181 , g8182 , g8183 , g8184 , g8185 , g8186 , g8187 , g8188 , g8189 , g8190 , g8191 , g8192 , g8193 , g8194 , g8195 , g8196 , g8197 , g8198 , g8199 , g8200 , g8201 , g8202 , g8203 , g8204 , g8205 , g8206 , g8207 , g8208 , g8209 , g8210 , g8211 , g8212 , g8213 , g8214 , g8215 , g8216 , g8217 , g8218 , g8219 , g8220 , g8221 , g8222 , g8223 , g8224 , g8225 , g8226 , g8227 , g8228 , g8229 , g8230 , g8231 , g8232 , g8233 , g8234 , g8235 , g8236 , g8237 , g8238 , g8239 , g8240 , g8241 , g8242 , g8243 , g8244 , g8245 , g8246 , g8247 , g8248 , g8249 , g8250 , g8251 , g8252 , g8253 , g8254 , g8255 , g8256 , g8257 , g8258 , g8259 , g8260 , g8261 , g8262 , g8263 , g8264 , g8265 , g8266 , g8267 , g8268 , g8269 , g8270 , g8271 , g8272 , g8273 , g8274 , g8275 , g8276 , g8277 , g8278 , g8279 , g8280 , g8281 , g8282 , g8283 , g8284 , g8285 , g8286 , g8287 , g8288 , g8289 , g8290 , g8291 , g8292 , g8293 , g8294 , g8295 , g8296 , g8297 , g8298 , g8299 , g8300 , g8301 , g8302 , g8303 , g8304 , g8305 , g8306 , g8307 , g8308 , g8309 , g8310 , g8311 , g8312 , g8313 , g8314 , g8315 , g8316 , g8317 , g8318 , g8319 , g8320 , g8321 , g8322 , g8323 , g8324 , g8325 , g8326 , g8327 , g8328 , g8329 , g8330 , g8331 , g8332 , g8333 , g8334 , g8335 , g8336 , g8337 , g8338 , g8339 , g8340 , g8341 , g8342 , g8343 , g8344 , g8345 , g8346 , g8347 , g8348 , g8349 , g8350 , g8351 , g8352 , g8353 , g8354 , g8355 , g8356 , g8357 , g8358 , g8359 , g8360 , g8361 , g8362 , g8363 , g8364 , g8365 , g8366 , g8367 , g8368 , g8369 , g8370 , g8371 , g8372 , g8373 , g8374 , g8375 , g8376 , g8377 , g8378 , g8379 , g8380 , g8381 , g8382 , g8383 , g8384 , g8385 , g8386 , g8387 , g8388 , g8389 , g8390 , g8391 , g8392 , g8393 , g8394 , g8395 , g8396 , g8397 , g8398 , g8399 , g8400 , g8401 , g8402 , g8403 , g8404 , g8405 , g8406 , g8407 , g8408 , g8409 , g8410 , g8411 , g8412 , g8413 , g8414 , g8415 , g8416 , g8417 , g8418 , g8419 , g8420 , g8421 , g8422 , g8423 , g8424 , g8425 , g8426 , g8427 , g8428 , g8429 , g8430 , g8431 , g8432 , g8433 , g8434 , g8435 , g8436 , g8437 , g8438 , g8439 , g8440 , g8441 , g8442 , g8443 , g8444 , g8445 , g8446 , g8447 , g8448 , g8449 , g8450 , g8451 , g8452 , g8453 , g8454 , g8455 , g8456 , g8457 , g8458 , g8459 , g8460 , g8461 , g8462 , g8463 , g8464 , g8465 , g8466 , g8467 , g8468 , g8469 , g8470 , g8471 , g8472 , g8473 , g8474 , g8475 , g8476 , g8477 , g8478 , g8479 , g8480 , g8481 , g8482 , g8483 , g8484 , g8485 , g8486 , g8487 , g8488 , g8489 , g8490 , g8491 , g8492 , g8493 , g8494 , g8495 , g8496 , g8497 , g8498 , g8499 , g8500 , g8501 , g8502 , g8503 , g8504 , g8505 , g8506 , g8507 , g8508 , g8509 , g8510 , g8511 , g8512 , g8513 , g8514 , g8515 , g8516 , g8517 , g8518 , g8519 , g8520 , g8521 , g8522 , g8523 , g8524 , g8525 , g8526 , g8527 , g8528 , g8529 , g8530 , g8531 , g8532 , g8533 , g8534 , g8535 , g8536 , g8537 , g8538 , g8539 , g8540 , g8541 , g8542 , g8543 , g8544 , g8545 , g8546 , g8547 , g8548 , g8549 , g8550 , g8551 , g8552 , g8553 , g8554 , g8555 , g8556 , g8557 , g8558 , g8559 , g8560 , g8561 , g8562 , g8563 , g8564 , g8565 , g8566 , g8567 , g8568 , g8569 , g8570 , g8571 , g8572 , g8573 , g8574 , g8575 , g8576 , g8577 , g8578 , g8579 , g8580 , g8581 , g8582 , g8583 , g8584 , g8585 , g8586 , g8587 , g8588 , g8589 , g8590 , g8591 , g8592 , g8593 , g8594 , g8595 , g8596 , g8597 , g8598 , g8599 , g8600 , g8601 , g8602 , g8603 , g8604 , g8605 , g8606 , g8607 , g8608 , g8609 , g8610 , g8611 , g8612 , g8613 , g8614 , g8615 , g8616 , g8617 , g8618 , g8619 , g8620 , g8621 , g8622 , g8623 , g8624 , g8625 , g8626 , g8627 , g8628 , g8629 , g8630 , g8631 , g8632 , g8633 , g8634 , g8635 , g8636 , g8637 , g8638 , g8639 , g8640 , g8641 , g8642 , g8643 , g8644 , g8645 , g8646 , g8647 , g8648 , g8649 , g8650 , g8651 , g8652 , g8653 , g8654 , g8655 , g8656 , g8657 , g8658 , g8659 , g8660 , g8661 , g8662 , g8663 , g8664 , g8665 , g8666 , g8667 , g8668 , g8669 , g8670 , g8671 , g8672 , g8673 , g8674 , g8675 , g8676 , g8677 , g8678 , g8679 , g8680 , g8681 , g8682 , g8683 , g8684 , g8685 , g8686 , g8687 , g8688 , g8689 , g8690 , g8691 , g8692 , g8693 , g8694 , g8695 , g8696 , g8697 , g8698 , g8699 , g8700 , g8701 , g8702 , g8703 , g8704 , g8705 , g8706 , g8707 , g8708 , g8709 , g8710 , g8711 , g8712 , g8713 , g8714 , g8715 , g8716 , g8717 , g8718 , g8719 , g8720 , g8721 , g8722 , g8723 , g8724 , g8725 , g8726 , g8727 , g8728 , g8729 , g8730 , g8731 , g8732 , g8733 , g8734 , g8735 , g8736 , g8737 , g8738 , g8739 , g8740 , g8741 , g8742 , g8743 , g8744 , g8745 , g8746 , g8747 , g8748 , g8749 , g8750 , g8751 , g8752 , g8753 , g8754 , g8755 , g8756 , g8757 , g8758 , g8759 , g8760 , g8761 , g8762 , g8763 , g8764 , g8765 , g8766 , g8767 , g8768 , g8769 , g8770 , g8771 , g8772 , g8773 , g8774 , g8775 , g8776 , g8777 , g8778 , g8779 , g8780 , g8781 , g8782 , g8783 , g8784 , g8785 , g8786 , g8787 , g8788 , g8789 , g8790 , g8791 , g8792 , g8793 , g8794 , g8795 , g8796 , g8797 , g8798 , g8799 , g8800 , g8801 , g8802 , g8803 , g8804 , g8805 , g8806 , g8807 , g8808 , g8809 , g8810 , g8811 , g8812 , g8813 , g8814 , g8815 , g8816 , g8817 , g8818 , g8819 , g8820 , g8821 , g8822 , g8823 , g8824 , g8825 , g8826 , g8827 , g8828 , g8829 , g8830 , g8831 , g8832 , g8833 , g8834 , g8835 , g8836 , g8837 , g8838 , g8839 , g8840 , g8841 , g8842 , g8843 , g8844 , g8845 , g8846 , g8847 , g8848 , g8849 , g8850 , g8851 , g8852 , g8853 , g8854 , g8855 , g8856 , g8857 , g8858 , g8859 , g8860 , g8861 , g8862 , g8863 , g8864 , g8865 , g8866 , g8867 , g8868 , g8869 , g8870 , g8871 , g8872 , g8873 , g8874 , g8875 , g8876 , g8877 , g8878 , g8879 , g8880 , g8881 , g8882 , g8883 , g8884 , g8885 , g8886 , g8887 , g8888 , g8889 , g8890 , g8891 , g8892 , g8893 , g8894 , g8895 , g8896 , g8897 , g8898 , g8899 , g8900 , g8901 , g8902 , g8903 , g8904 , g8905 , g8906 , g8907 , g8908 , g8909 , g8910 , g8911 , g8912 , g8913 , g8914 , g8915 , g8916 , g8917 , g8918 , g8919 , g8920 , g8921 , g8922 , g8923 , g8924 , g8925 , g8926 , g8927 , g8928 , g8929 , g8930 , g8931 , g8932 , g8933 , g8934 , g8935 , g8936 , g8937 , g8938 , g8939 , g8940 , g8941 , g8942 , g8943 , g8944 , g8945 , g8946 , g8947 , g8948 , g8949 , g8950 , g8951 , g8952 , g8953 , g8954 , g8955 , g8956 , g8957 , g8958 , g8959 , g8960 , g8961 , g8962 , g8963 , g8964 , g8965 , g8966 , g8967 , g8968 , g8969 , g8970 , g8971 , g8972 , g8973 , g8974 , g8975 , g8976 , g8977 , g8978 );
input g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 , g98 , g99 , g100 , g101 , g102 , g103 , g104 , g105 , g106 , g107 , g108 , g109 , g110 , g111 , g112 , g113 , g114 , g115 , g116 , g117 , g118 , g119 , g120 , g121 , g122 , g123 , g124 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g136 , g137 , g138 , g139 , g140 , g141 , g142 , g143 , g144 , g145 , g146 , g147 , g148 , g149 , g150 , g151 , g152 , g153 , g154 , g155 , g156 , g157 , g158 , g159 , g160 , g161 , g162 , g163 , g164 , g165 , g166 , g167 , g168 , g169 , g170 , g171 , g172 , g173 , g174 , g175 , g176 , g177 , g178 , g179 , g180 , g181 , g182 , g183 , g184 , g185 , g186 , g187 , g188 , g189 , g190 , g191 , g192 , g193 , g194 , g195 , g196 , g197 , g198 , g199 , g200 , g201 , g202 , g203 , g204 , g205 , g206 , g207 , g208 , g209 , g210 , g211 , g212 , g213 , g214 , g215 , g216 , g217 , g218 , g219 , g220 , g221 , g222 , g223 , g224 , g225 , g226 , g227 , g228 , g229 , g230 , g231 , g232 , g233 , g234 , g235 , g236 , g237 , g238 , g239 , g240 , g241 , g242 , g243 , g244 , g245 , g246 , g247 , g248 , g249 , g250 , g251 , g252 , g253 , g254 , g255 , g256 , g257 , g258 , g259 , g260 , g261 , g262 , g263 , g264 , g265 , g266 , g267 , g268 , g269 , g270 , g271 , g272 , g273 , g274 , g275 , g276 , g277 , g278 , g279 , g280 , g281 , g282 , g283 , g284 , g285 , g286 , g287 , g288 , g289 , g290 , g291 , g292 , g293 , g294 , g295 , g296 , g297 , g298 , g299 , g300 , g301 , g302 , g303 , g304 , g305 , g306 , g307 , g308 , g309 , g310 , g311 , g312 , g313 , g314 , g315 , g316 , g317 , g318 , g319 , g320 , g321 , g322 , g323 , g324 , g325 , g326 , g327 , g328 , g329 , g330 , g331 , g332 , g333 , g334 , g335 , g336 , g337 , g338 , g339 , g340 , g341 , g342 , g343 , g344 , g345 , g346 , g347 , g348 , g349 , g350 , g351 , g352 , g353 , g354 , g355 , g356 , g357 , g358 , g359 , g360 , g361 , g362 , g363 , g364 , g365 , g366 , g367 , g368 , g369 , g370 , g371 , g372 , g373 , g374 , g375 , g376 , g377 , g378 , g379 , g380 , g381 , g382 , g383 , g384 , g385 , g386 , g387 , g388 , g389 , g390 , g391 , g392 , g393 , g394 , g395 , g396 , g397 , g398 , g399 , g400 , g401 , g402 , g403 , g404 , g405 , g406 , g407 , g408 , g409 , g410 , g411 , g412 , g413 , g414 , g415 , g416 , g417 , g418 , g419 , g420 , g421 , g422 , g423 , g424 , g425 , g426 , g427 , g428 , g429 , g430 , g431 , g432 , g433 , g434 , g435 , g436 , g437 , g438 , g439 , g440 , g441 , g442 , g443 , g444 , g445 , g446 , g447 , g448 , g449 , g450 , g451 , g452 , g453 , g454 , g455 , g456 , g457 , g458 , g459 , g460 , g461 , g462 , g463 , g464 , g465 , g466 , g467 , g468 , g469 , g470 , g471 , g472 , g473 , g474 , g475 , g476 , g477 , g478 , g479 , g480 , g481 , g482 , g483 , g484 , g485 , g486 , g487 , g488 , g489 , g490 , g491 , g492 , g493 , g494 , g495 , g496 , g497 , g498 , g499 , g500 , g501 , g502 , g503 , g504 , g505 , g506 , g507 , g508 , g509 , g510 , g511 , g512 , g513 , g514 , g515 , g516 , g517 , g518 , g519 , g520 , g521 , g522 , g523 , g524 , g525 , g526 , g527 , g528 , g529 , g530 , g531 , g532 , g533 , g534 , g535 , g536 , g537 , g538 , g539 , g540 , g541 , g542 , g543 , g544 , g545 , g546 , g547 , g548 , g549 , g550 , g551 , g552 , g553 , g554 , g555 , g556 , g557 , g558 , g559 , g560 , g561 , g562 , g563 , g564 , g565 , g566 , g567 , g568 , g569 , g570 , g571 , g572 , g573 , g574 , g575 , g576 , g577 , g578 , g579 , g580 , g581 , g582 , g583 , g584 , g585 , g586 , g587 , g588 , g589 , g590 , g591 , g592 , g593 , g594 , g595 , g596 , g597 , g598 , g599 , g600 , g601 , g602 , g603 , g604 , g605 , g606 , g607 , g608 , g609 , g610 , g611 , g612 , g613 , g614 , g615 , g616 , g617 , g618 , g619 , g620 , g621 , g622 , g623 , g624 , g625 , g626 , g627 , g628 , g629 , g630 , g631 , g632 , g633 , g634 , g635 , g636 , g637 , g638 , g639 , g640 , g641 , g642 , g643 , g644 , g645 , g646 , g647 , g648 , g649 , g650 , g651 , g652 , g653 , g654 , g655 , g656 , g657 , g658 , g659 , g660 , g661 , g662 , g663 , g664 , g665 , g666 , g667 , g668 , g669 , g670 , g671 , g672 , g673 , g674 , g675 , g676 , g677 , g678 , g679 , g680 , g681 , g682 , g683 , g684 , g685 , g686 , g687 , g688 , g689 , g690 , g691 , g692 , g693 , g694 , g695 , g696 , g697 , g698 , g699 , g700 , g701 , g702 , g703 , g704 , g705 , g706 , g707 , g708 , g709 , g710 , g711 , g712 , g713 , g714 , g715 , g716 , g717 , g718 , g719 , g720 , g721 , g722 , g723 , g724 , g725 , g726 , g727 , g728 , g729 , g730 , g731 , g732 , g733 , g734 , g735 , g736 , g737 , g738 , g739 , g740 , g741 , g742 , g743 , g744 , g745 , g746 , g747 , g748 , g749 , g750 , g751 , g752 , g753 , g754 , g755 , g756 , g757 , g758 , g759 , g760 , g761 , g762 , g763 , g764 , g765 , g766 , g767 , g768 , g769 , g770 , g771 , g772 , g773 , g774 , g775 , g776 , g777 , g778 , g779 , g780 , g781 , g782 , g783 , g784 , g785 , g786 , g787 , g788 , g789 , g790 , g791 , g792 , g793 , g794 , g795 , g796 , g797 , g798 , g799 , g800 , g801 , g802 , g803 , g804 , g805 , g806 , g807 , g808 , g809 , g810 , g811 , g812 , g813 , g814 , g815 , g816 , g817 , g818 , g819 , g820 , g821 , g822 , g823 , g824 , g825 , g826 , g827 , g828 , g829 , g830 , g831 , g832 , g833 , g834 , g835 , g836 , g837 , g838 , g839 , g840 , g841 , g842 , g843 , g844 , g845 , g846 , g847 , g848 , g849 , g850 , g851 , g852 , g853 , g854 , g855 , g856 , g857 , g858 , g859 , g860 , g861 , g862 , g863 , g864 , g865 , g866 , g867 , g868 , g869 , g870 , g871 , g872 , g873 , g874 , g875 , g876 , g877 , g878 , g879 , g880 , g881 , g882 , g883 , g884 , g885 , g886 , g887 , g888 , g889 , g890 , g891 , g892 , g893 , g894 , g895 , g896 , g897 , g898 , g899 , g900 , g901 , g902 , g903 , g904 , g905 , g906 , g907 , g908 , g909 , g910 , g911 , g912 , g913 , g914 , g915 , g916 , g917 , g918 , g919 , g920 , g921 , g922 , g923 , g924 , g925 , g926 , g927 , g928 , g929 , g930 , g931 , g932 , g933 , g934 , g935 , g936 , g937 , g938 , g939 , g940 , g941 , g942 , g943 , g944 , g945 , g946 , g947 , g948 , g949 , g950 , g951 , g952 , g953 , g954 , g955 , g956 , g957 , g958 , g959 , g960 , g961 , g962 , g963 , g964 , g965 , g966 , g967 , g968 , g969 , g970 , g971 , g972 , g973 , g974 , g975 , g976 , g977 , g978 , g979 , g980 , g981 , g982 , g983 , g984 , g985 , g986 , g987 , g988 , g989 , g990 , g991 , g992 , g993 , g994 , g995 , g996 , g997 , g998 , g999 , g1000 , g1001 , g1002 , g1003 , g1004 , g1005 , g1006 , g1007 , g1008 , g1009 , g1010 , g1011 , g1012 , g1013 , g1014 , g1015 , g1016 , g1017 , g1018 , g1019 , g1020 , g1021 , g1022 , g1023 , g1024 , g1025 , g1026 , g1027 , g1028 , g1029 , g1030 , g1031 , g1032 , g1033 , g1034 , g1035 , g1036 , g1037 , g1038 , g1039 , g1040 , g1041 , g1042 , g1043 , g1044 , g1045 , g1046 , g1047 , g1048 , g1049 , g1050 , g1051 , g1052 , g1053 , g1054 , g1055 , g1056 , g1057 , g1058 , g1059 , g1060 , g1061 , g1062 , g1063 , g1064 , g1065 , g1066 , g1067 , g1068 , g1069 , g1070 , g1071 , g1072 , g1073 , g1074 , g1075 , g1076 , g1077 , g1078 , g1079 , g1080 , g1081 , g1082 , g1083 , g1084 , g1085 , g1086 , g1087 , g1088 , g1089 , g1090 , g1091 , g1092 , g1093 , g1094 , g1095 , g1096 , g1097 , g1098 , g1099 , g1100 , g1101 , g1102 , g1103 , g1104 , g1105 , g1106 , g1107 , g1108 , g1109 , g1110 , g1111 , g1112 , g1113 , g1114 , g1115 , g1116 , g1117 , g1118 , g1119 , g1120 , g1121 , g1122 , g1123 , g1124 , g1125 , g1126 , g1127 , g1128 , g1129 , g1130 , g1131 , g1132 , g1133 , g1134 , g1135 , g1136 , g1137 , g1138 , g1139 , g1140 , g1141 , g1142 , g1143 , g1144 , g1145 , g1146 , g1147 , g1148 , g1149 , g1150 , g1151 , g1152 , g1153 , g1154 , g1155 , g1156 , g1157 , g1158 , g1159 , g1160 , g1161 , g1162 , g1163 , g1164 , g1165 , g1166 , g1167 , g1168 , g1169 , g1170 , g1171 , g1172 , g1173 , g1174 , g1175 , g1176 , g1177 , g1178 , g1179 , g1180 , g1181 , g1182 , g1183 , g1184 , g1185 , g1186 , g1187 , g1188 , g1189 , g1190 , g1191 , g1192 , g1193 , g1194 , g1195 , g1196 , g1197 , g1198 , g1199 , g1200 , g1201 , g1202 , g1203 , g1204 , g1205 , g1206 , g1207 , g1208 , g1209 , g1210 , g1211 , g1212 , g1213 , g1214 , g1215 , g1216 , g1217 , g1218 , g1219 , g1220 , g1221 , g1222 , g1223 , g1224 , g1225 , g1226 , g1227 , g1228 , g1229 , g1230 , g1231 , g1232 , g1233 , g1234 , g1235 , g1236 , g1237 , g1238 , g1239 , g1240 , g1241 , g1242 , g1243 , g1244 , g1245 , g1246 , g1247 , g1248 , g1249 , g1250 , g1251 , g1252 , g1253 , g1254 , g1255 , g1256 , g1257 , g1258 , g1259 , g1260 , g1261 , g1262 , g1263 , g1264 , g1265 , g1266 , g1267 , g1268 , g1269 , g1270 , g1271 , g1272 , g1273 , g1274 , g1275 , g1276 , g1277 , g1278 , g1279 , g1280 , g1281 , g1282 , g1283 , g1284 , g1285 , g1286 , g1287 , g1288 , g1289 , g1290 , g1291 , g1292 , g1293 , g1294 , g1295 , g1296 , g1297 , g1298 , g1299 , g1300 , g1301 , g1302 , g1303 , g1304 , g1305 , g1306 , g1307 , g1308 , g1309 , g1310 , g1311 , g1312 , g1313 , g1314 , g1315 , g1316 , g1317 , g1318 , g1319 , g1320 , g1321 , g1322 , g1323 , g1324 , g1325 , g1326 , g1327 , g1328 , g1329 , g1330 , g1331 , g1332 , g1333 , g1334 , g1335 , g1336 , g1337 , g1338 , g1339 , g1340 , g1341 , g1342 , g1343 , g1344 , g1345 , g1346 , g1347 , g1348 , g1349 , g1350 , g1351 , g1352 , g1353 , g1354 , g1355 , g1356 , g1357 , g1358 , g1359 , g1360 , g1361 , g1362 , g1363 , g1364 , g1365 , g1366 , g1367 , g1368 , g1369 , g1370 , g1371 , g1372 , g1373 , g1374 , g1375 , g1376 , g1377 , g1378 , g1379 , g1380 , g1381 , g1382 , g1383 , g1384 , g1385 , g1386 , g1387 , g1388 , g1389 , g1390 , g1391 , g1392 , g1393 , g1394 , g1395 , g1396 , g1397 , g1398 , g1399 , g1400 , g1401 , g1402 , g1403 , g1404 , g1405 , g1406 , g1407 , g1408 , g1409 , g1410 , g1411 , g1412 , g1413 , g1414 , g1415 , g1416 , g1417 , g1418 , g1419 , g1420 , g1421 , g1422 , g1423 , g1424 , g1425 , g1426 , g1427 , g1428 , g1429 , g1430 , g1431 , g1432 , g1433 , g1434 , g1435 , g1436 , g1437 , g1438 , g1439 , g1440 , g1441 , g1442 , g1443 , g1444 , g1445 , g1446 , g1447 , g1448 , g1449 , g1450 , g1451 , g1452 , g1453 , g1454 , g1455 , g1456 , g1457 , g1458 , g1459 , g1460 , g1461 , g1462 , g1463 , g1464 , g1465 , g1466 , g1467 , g1468 , g1469 , g1470 , g1471 , g1472 , g1473 , g1474 , g1475 , g1476 , g1477 , g1478 , g1479 , g1480 , g1481 , g1482 , g1483 , g1484 , g1485 , g1486 , g1487 , g1488 , g1489 , g1490 , g1491 , g1492 , g1493 , g1494 , g1495 , g1496 , g1497 , g1498 , g1499 , g1500 , g1501 , g1502 , g1503 , g1504 , g1505 , g1506 , g1507 , g1508 , g1509 , g1510 , g1511 , g1512 , g1513 , g1514 , g1515 , g1516 , g1517 , g1518 , g1519 , g1520 , g1521 , g1522 , g1523 , g1524 , g1525 , g1526 , g1527 , g1528 , g1529 , g1530 , g1531 , g1532 , g1533 , g1534 , g1535 , g1536 , g1537 , g1538 , g1539 , g1540 , g1541 , g1542 , g1543 , g1544 , g1545 , g1546 , g1547 , g1548 , g1549 , g1550 , g1551 , g1552 , g1553 , g1554 , g1555 , g1556 , g1557 , g1558 , g1559 , g1560 , g1561 , g1562 , g1563 , g1564 , g1565 , g1566 , g1567 , g1568 , g1569 , g1570 , g1571 , g1572 , g1573 , g1574 , g1575 , g1576 , g1577 , g1578 , g1579 , g1580 , g1581 , g1582 , g1583 , g1584 , g1585 , g1586 , g1587 , g1588 , g1589 , g1590 , g1591 , g1592 , g1593 , g1594 , g1595 , g1596 , g1597 , g1598 , g1599 , g1600 , g1601 , g1602 , g1603 , g1604 , g1605 , g1606 , g1607 , g1608 , g1609 , g1610 , g1611 , g1612 , g1613 , g1614 , g1615 , g1616 , g1617 , g1618 , g1619 , g1620 , g1621 , g1622 , g1623 , g1624 , g1625 , g1626 , g1627 , g1628 , g1629 , g1630 , g1631 , g1632 , g1633 , g1634 , g1635 , g1636 , g1637 , g1638 , g1639 , g1640 , g1641 , g1642 , g1643 , g1644 , g1645 , g1646 , g1647 , g1648 , g1649 , g1650 , g1651 , g1652 , g1653 , g1654 , g1655 , g1656 , g1657 , g1658 , g1659 , g1660 , g1661 , g1662 , g1663 , g1664 , g1665 , g1666 , g1667 , g1668 , g1669 , g1670 , g1671 , g1672 , g1673 , g1674 , g1675 , g1676 , g1677 , g1678 , g1679 , g1680 , g1681 , g1682 , g1683 , g1684 , g1685 , g1686 , g1687 , g1688 , g1689 , g1690 , g1691 , g1692 , g1693 , g1694 , g1695 , g1696 , g1697 , g1698 , g1699 , g1700 , g1701 , g1702 , g1703 , g1704 , g1705 , g1706 , g1707 , g1708 , g1709 , g1710 , g1711 , g1712 , g1713 , g1714 , g1715 , g1716 , g1717 , g1718 , g1719 , g1720 , g1721 , g1722 , g1723 , g1724 , g1725 , g1726 , g1727 , g1728 , g1729 , g1730 , g1731 , g1732 , g1733 , g1734 , g1735 , g1736 , g1737 , g1738 , g1739 , g1740 , g1741 , g1742 , g1743 , g1744 , g1745 , g1746 , g1747 , g1748 , g1749 , g1750 , g1751 , g1752 , g1753 , g1754 , g1755 , g1756 , g1757 , g1758 , g1759 , g1760 , g1761 , g1762 , g1763 , g1764 , g1765 , g1766 , g1767 , g1768 , g1769 , g1770 , g1771 , g1772 , g1773 , g1774 , g1775 , g1776 , g1777 , g1778 , g1779 , g1780 , g1781 , g1782 , g1783 , g1784 , g1785 , g1786 , g1787 , g1788 , g1789 , g1790 , g1791 , g1792 , g1793 , g1794 , g1795 , g1796 , g1797 , g1798 , g1799 , g1800 , g1801 , g1802 , g1803 , g1804 , g1805 , g1806 , g1807 , g1808 , g1809 , g1810 , g1811 , g1812 , g1813 , g1814 , g1815 , g1816 , g1817 , g1818 , g1819 , g1820 , g1821 , g1822 , g1823 , g1824 , g1825 , g1826 , g1827 , g1828 , g1829 , g1830 , g1831 , g1832 , g1833 , g1834 , g1835 , g1836 , g1837 , g1838 , g1839 , g1840 , g1841 , g1842 , g1843 , g1844 , g1845 , g1846 , g1847 , g1848 , g1849 , g1850 , g1851 , g1852 , g1853 , g1854 , g1855 , g1856 , g1857 , g1858 , g1859 , g1860 , g1861 , g1862 , g1863 , g1864 , g1865 , g1866 , g1867 , g1868 , g1869 , g1870 , g1871 , g1872 , g1873 ;
output g1874 , g1875 , g1876 , g1877 , g1878 , g1879 , g1880 , g1881 , g1882 , g1883 , g1884 , g1885 , g1886 , g1887 , g1888 , g1889 , g1890 , g1891 , g1892 , g1893 , g1894 , g1895 , g1896 , g1897 , g1898 , g1899 , g1900 , g1901 , g1902 , g1903 , g1904 , g1905 , g1906 , g1907 , g1908 , g1909 , g1910 , g1911 , g1912 , g1913 , g1914 , g1915 , g1916 , g1917 , g1918 , g1919 , g1920 , g1921 , g1922 , g1923 , g1924 , g1925 , g1926 , g1927 , g1928 , g1929 , g1930 , g1931 , g1932 , g1933 , g1934 , g1935 , g1936 , g1937 , g1938 , g1939 , g1940 , g1941 , g1942 , g1943 , g1944 , g1945 , g1946 , g1947 , g1948 , g1949 , g1950 , g1951 , g1952 , g1953 , g1954 , g1955 , g1956 , g1957 , g1958 , g1959 , g1960 , g1961 , g1962 , g1963 , g1964 , g1965 , g1966 , g1967 , g1968 , g1969 , g1970 , g1971 , g1972 , g1973 , g1974 , g1975 , g1976 , g1977 , g1978 , g1979 , g1980 , g1981 , g1982 , g1983 , g1984 , g1985 , g1986 , g1987 , g1988 , g1989 , g1990 , g1991 , g1992 , g1993 , g1994 , g1995 , g1996 , g1997 , g1998 , g1999 , g2000 , g2001 , g2002 , g2003 , g2004 , g2005 , g2006 , g2007 , g2008 , g2009 , g2010 , g2011 , g2012 , g2013 , g2014 , g2015 , g2016 , g2017 , g2018 , g2019 , g2020 , g2021 , g2022 , g2023 , g2024 , g2025 , g2026 , g2027 , g2028 , g2029 , g2030 , g2031 , g2032 , g2033 , g2034 , g2035 , g2036 , g2037 , g2038 , g2039 , g2040 , g2041 , g2042 , g2043 , g2044 , g2045 , g2046 , g2047 , g2048 , g2049 , g2050 , g2051 , g2052 , g2053 , g2054 , g2055 , g2056 , g2057 , g2058 , g2059 , g2060 , g2061 , g2062 , g2063 , g2064 , g2065 , g2066 , g2067 , g2068 , g2069 , g2070 , g2071 , g2072 , g2073 , g2074 , g2075 , g2076 , g2077 , g2078 , g2079 , g2080 , g2081 , g2082 , g2083 , g2084 , g2085 , g2086 , g2087 , g2088 , g2089 , g2090 , g2091 , g2092 , g2093 , g2094 , g2095 , g2096 , g2097 , g2098 , g2099 , g2100 , g2101 , g2102 , g2103 , g2104 , g2105 , g2106 , g2107 , g2108 , g2109 , g2110 , g2111 , g2112 , g2113 , g2114 , g2115 , g2116 , g2117 , g2118 , g2119 , g2120 , g2121 , g2122 , g2123 , g2124 , g2125 , g2126 , g2127 , g2128 , g2129 , g2130 , g2131 , g2132 , g2133 , g2134 , g2135 , g2136 , g2137 , g2138 , g2139 , g2140 , g2141 , g2142 , g2143 , g2144 , g2145 , g2146 , g2147 , g2148 , g2149 , g2150 , g2151 , g2152 , g2153 , g2154 , g2155 , g2156 , g2157 , g2158 , g2159 , g2160 , g2161 , g2162 , g2163 , g2164 , g2165 , g2166 , g2167 , g2168 , g2169 , g2170 , g2171 , g2172 , g2173 , g2174 , g2175 , g2176 , g2177 , g2178 , g2179 , g2180 , g2181 , g2182 , g2183 , g2184 , g2185 , g2186 , g2187 , g2188 , g2189 , g2190 , g2191 , g2192 , g2193 , g2194 , g2195 , g2196 , g2197 , g2198 , g2199 , g2200 , g2201 , g2202 , g2203 , g2204 , g2205 , g2206 , g2207 , g2208 , g2209 , g2210 , g2211 , g2212 , g2213 , g2214 , g2215 , g2216 , g2217 , g2218 , g2219 , g2220 , g2221 , g2222 , g2223 , g2224 , g2225 , g2226 , g2227 , g2228 , g2229 , g2230 , g2231 , g2232 , g2233 , g2234 , g2235 , g2236 , g2237 , g2238 , g2239 , g2240 , g2241 , g2242 , g2243 , g2244 , g2245 , g2246 , g2247 , g2248 , g2249 , g2250 , g2251 , g2252 , g2253 , g2254 , g2255 , g2256 , g2257 , g2258 , g2259 , g2260 , g2261 , g2262 , g2263 , g2264 , g2265 , g2266 , g2267 , g2268 , g2269 , g2270 , g2271 , g2272 , g2273 , g2274 , g2275 , g2276 , g2277 , g2278 , g2279 , g2280 , g2281 , g2282 , g2283 , g2284 , g2285 , g2286 , g2287 , g2288 , g2289 , g2290 , g2291 , g2292 , g2293 , g2294 , g2295 , g2296 , g2297 , g2298 , g2299 , g2300 , g2301 , g2302 , g2303 , g2304 , g2305 , g2306 , g2307 , g2308 , g2309 , g2310 , g2311 , g2312 , g2313 , g2314 , g2315 , g2316 , g2317 , g2318 , g2319 , g2320 , g2321 , g2322 , g2323 , g2324 , g2325 , g2326 , g2327 , g2328 , g2329 , g2330 , g2331 , g2332 , g2333 , g2334 , g2335 , g2336 , g2337 , g2338 , g2339 , g2340 , g2341 , g2342 , g2343 , g2344 , g2345 , g2346 , g2347 , g2348 , g2349 , g2350 , g2351 , g2352 , g2353 , g2354 , g2355 , g2356 , g2357 , g2358 , g2359 , g2360 , g2361 , g2362 , g2363 , g2364 , g2365 , g2366 , g2367 , g2368 , g2369 , g2370 , g2371 , g2372 , g2373 , g2374 , g2375 , g2376 , g2377 , g2378 , g2379 , g2380 , g2381 , g2382 , g2383 , g2384 , g2385 , g2386 , g2387 , g2388 , g2389 , g2390 , g2391 , g2392 , g2393 , g2394 , g2395 , g2396 , g2397 , g2398 , g2399 , g2400 , g2401 , g2402 , g2403 , g2404 , g2405 , g2406 , g2407 , g2408 , g2409 , g2410 , g2411 , g2412 , g2413 , g2414 , g2415 , g2416 , g2417 , g2418 , g2419 , g2420 , g2421 , g2422 , g2423 , g2424 , g2425 , g2426 , g2427 , g2428 , g2429 , g2430 , g2431 , g2432 , g2433 , g2434 , g2435 , g2436 , g2437 , g2438 , g2439 , g2440 , g2441 , g2442 , g2443 , g2444 , g2445 , g2446 , g2447 , g2448 , g2449 , g2450 , g2451 , g2452 , g2453 , g2454 , g2455 , g2456 , g2457 , g2458 , g2459 , g2460 , g2461 , g2462 , g2463 , g2464 , g2465 , g2466 , g2467 , g2468 , g2469 , g2470 , g2471 , g2472 , g2473 , g2474 , g2475 , g2476 , g2477 , g2478 , g2479 , g2480 , g2481 , g2482 , g2483 , g2484 , g2485 , g2486 , g2487 , g2488 , g2489 , g2490 , g2491 , g2492 , g2493 , g2494 , g2495 , g2496 , g2497 , g2498 , g2499 , g2500 , g2501 , g2502 , g2503 , g2504 , g2505 , g2506 , g2507 , g2508 , g2509 , g2510 , g2511 , g2512 , g2513 , g2514 , g2515 , g2516 , g2517 , g2518 , g2519 , g2520 , g2521 , g2522 , g2523 , g2524 , g2525 , g2526 , g2527 , g2528 , g2529 , g2530 , g2531 , g2532 , g2533 , g2534 , g2535 , g2536 , g2537 , g2538 , g2539 , g2540 , g2541 , g2542 , g2543 , g2544 , g2545 , g2546 , g2547 , g2548 , g2549 , g2550 , g2551 , g2552 , g2553 , g2554 , g2555 , g2556 , g2557 , g2558 , g2559 , g2560 , g2561 , g2562 , g2563 , g2564 , g2565 , g2566 , g2567 , g2568 , g2569 , g2570 , g2571 , g2572 , g2573 , g2574 , g2575 , g2576 , g2577 , g2578 , g2579 , g2580 , g2581 , g2582 , g2583 , g2584 , g2585 , g2586 , g2587 , g2588 , g2589 , g2590 , g2591 , g2592 , g2593 , g2594 , g2595 , g2596 , g2597 , g2598 , g2599 , g2600 , g2601 , g2602 , g2603 , g2604 , g2605 , g2606 , g2607 , g2608 , g2609 , g2610 , g2611 , g2612 , g2613 , g2614 , g2615 , g2616 , g2617 , g2618 , g2619 , g2620 , g2621 , g2622 , g2623 , g2624 , g2625 , g2626 , g2627 , g2628 , g2629 , g2630 , g2631 , g2632 , g2633 , g2634 , g2635 , g2636 , g2637 , g2638 , g2639 , g2640 , g2641 , g2642 , g2643 , g2644 , g2645 , g2646 , g2647 , g2648 , g2649 , g2650 , g2651 , g2652 , g2653 , g2654 , g2655 , g2656 , g2657 , g2658 , g2659 , g2660 , g2661 , g2662 , g2663 , g2664 , g2665 , g2666 , g2667 , g2668 , g2669 , g2670 , g2671 , g2672 , g2673 , g2674 , g2675 , g2676 , g2677 , g2678 , g2679 , g2680 , g2681 , g2682 , g2683 , g2684 , g2685 , g2686 , g2687 , g2688 , g2689 , g2690 , g2691 , g2692 , g2693 , g2694 , g2695 , g2696 , g2697 , g2698 , g2699 , g2700 , g2701 , g2702 , g2703 , g2704 , g2705 , g2706 , g2707 , g2708 , g2709 , g2710 , g2711 , g2712 , g2713 , g2714 , g2715 , g2716 , g2717 , g2718 , g2719 , g2720 , g2721 , g2722 , g2723 , g2724 , g2725 , g2726 , g2727 , g2728 , g2729 , g2730 , g2731 , g2732 , g2733 , g2734 , g2735 , g2736 , g2737 , g2738 , g2739 , g2740 , g2741 , g2742 , g2743 , g2744 , g2745 , g2746 , g2747 , g2748 , g2749 , g2750 , g2751 , g2752 , g2753 , g2754 , g2755 , g2756 , g2757 , g2758 , g2759 , g2760 , g2761 , g2762 , g2763 , g2764 , g2765 , g2766 , g2767 , g2768 , g2769 , g2770 , g2771 , g2772 , g2773 , g2774 , g2775 , g2776 , g2777 , g2778 , g2779 , g2780 , g2781 , g2782 , g2783 , g2784 , g2785 , g2786 , g2787 , g2788 , g2789 , g2790 , g2791 , g2792 , g2793 , g2794 , g2795 , g2796 , g2797 , g2798 , g2799 , g2800 , g2801 , g2802 , g2803 , g2804 , g2805 , g2806 , g2807 , g2808 , g2809 , g2810 , g2811 , g2812 , g2813 , g2814 , g2815 , g2816 , g2817 , g2818 , g2819 , g2820 , g2821 , g2822 , g2823 , g2824 , g2825 , g2826 , g2827 , g2828 , g2829 , g2830 , g2831 , g2832 , g2833 , g2834 , g2835 , g2836 , g2837 , g2838 , g2839 , g2840 , g2841 , g2842 , g2843 , g2844 , g2845 , g2846 , g2847 , g2848 , g2849 , g2850 , g2851 , g2852 , g2853 , g2854 , g2855 , g2856 , g2857 , g2858 , g2859 , g2860 , g2861 , g2862 , g2863 , g2864 , g2865 , g2866 , g2867 , g2868 , g2869 , g2870 , g2871 , g2872 , g2873 , g2874 , g2875 , g2876 , g2877 , g2878 , g2879 , g2880 , g2881 , g2882 , g2883 , g2884 , g2885 , g2886 , g2887 , g2888 , g2889 , g2890 , g2891 , g2892 , g2893 , g2894 , g2895 , g2896 , g2897 , g2898 , g2899 , g2900 , g2901 , g2902 , g2903 , g2904 , g2905 , g2906 , g2907 , g2908 , g2909 , g2910 , g2911 , g2912 , g2913 , g2914 , g2915 , g2916 , g2917 , g2918 , g2919 , g2920 , g2921 , g2922 , g2923 , g2924 , g2925 , g2926 , g2927 , g2928 , g2929 , g2930 , g2931 , g2932 , g2933 , g2934 , g2935 , g2936 , g2937 , g2938 , g2939 , g2940 , g2941 , g2942 , g2943 , g2944 , g2945 , g2946 , g2947 , g2948 , g2949 , g2950 , g2951 , g2952 , g2953 , g2954 , g2955 , g2956 , g2957 , g2958 , g2959 , g2960 , g2961 , g2962 , g2963 , g2964 , g2965 , g2966 , g2967 , g2968 , g2969 , g2970 , g2971 , g2972 , g2973 , g2974 , g2975 , g2976 , g2977 , g2978 , g2979 , g2980 , g2981 , g2982 , g2983 , g2984 , g2985 , g2986 , g2987 , g2988 , g2989 , g2990 , g2991 , g2992 , g2993 , g2994 , g2995 , g2996 , g2997 , g2998 , g2999 , g3000 , g3001 , g3002 , g3003 , g3004 , g3005 , g3006 , g3007 , g3008 , g3009 , g3010 , g3011 , g3012 , g3013 , g3014 , g3015 , g3016 , g3017 , g3018 , g3019 , g3020 , g3021 , g3022 , g3023 , g3024 , g3025 , g3026 , g3027 , g3028 , g3029 , g3030 , g3031 , g3032 , g3033 , g3034 , g3035 , g3036 , g3037 , g3038 , g3039 , g3040 , g3041 , g3042 , g3043 , g3044 , g3045 , g3046 , g3047 , g3048 , g3049 , g3050 , g3051 , g3052 , g3053 , g3054 , g3055 , g3056 , g3057 , g3058 , g3059 , g3060 , g3061 , g3062 , g3063 , g3064 , g3065 , g3066 , g3067 , g3068 , g3069 , g3070 , g3071 , g3072 , g3073 , g3074 , g3075 , g3076 , g3077 , g3078 , g3079 , g3080 , g3081 , g3082 , g3083 , g3084 , g3085 , g3086 , g3087 , g3088 , g3089 , g3090 , g3091 , g3092 , g3093 , g3094 , g3095 , g3096 , g3097 , g3098 , g3099 , g3100 , g3101 , g3102 , g3103 , g3104 , g3105 , g3106 , g3107 , g3108 , g3109 , g3110 , g3111 , g3112 , g3113 , g3114 , g3115 , g3116 , g3117 , g3118 , g3119 , g3120 , g3121 , g3122 , g3123 , g3124 , g3125 , g3126 , g3127 , g3128 , g3129 , g3130 , g3131 , g3132 , g3133 , g3134 , g3135 , g3136 , g3137 , g3138 , g3139 , g3140 , g3141 , g3142 , g3143 , g3144 , g3145 , g3146 , g3147 , g3148 , g3149 , g3150 , g3151 , g3152 , g3153 , g3154 , g3155 , g3156 , g3157 , g3158 , g3159 , g3160 , g3161 , g3162 , g3163 , g3164 , g3165 , g3166 , g3167 , g3168 , g3169 , g3170 , g3171 , g3172 , g3173 , g3174 , g3175 , g3176 , g3177 , g3178 , g3179 , g3180 , g3181 , g3182 , g3183 , g3184 , g3185 , g3186 , g3187 , g3188 , g3189 , g3190 , g3191 , g3192 , g3193 , g3194 , g3195 , g3196 , g3197 , g3198 , g3199 , g3200 , g3201 , g3202 , g3203 , g3204 , g3205 , g3206 , g3207 , g3208 , g3209 , g3210 , g3211 , g3212 , g3213 , g3214 , g3215 , g3216 , g3217 , g3218 , g3219 , g3220 , g3221 , g3222 , g3223 , g3224 , g3225 , g3226 , g3227 , g3228 , g3229 , g3230 , g3231 , g3232 , g3233 , g3234 , g3235 , g3236 , g3237 , g3238 , g3239 , g3240 , g3241 , g3242 , g3243 , g3244 , g3245 , g3246 , g3247 , g3248 , g3249 , g3250 , g3251 , g3252 , g3253 , g3254 , g3255 , g3256 , g3257 , g3258 , g3259 , g3260 , g3261 , g3262 , g3263 , g3264 , g3265 , g3266 , g3267 , g3268 , g3269 , g3270 , g3271 , g3272 , g3273 , g3274 , g3275 , g3276 , g3277 , g3278 , g3279 , g3280 , g3281 , g3282 , g3283 , g3284 , g3285 , g3286 , g3287 , g3288 , g3289 , g3290 , g3291 , g3292 , g3293 , g3294 , g3295 , g3296 , g3297 , g3298 , g3299 , g3300 , g3301 , g3302 , g3303 , g3304 , g3305 , g3306 , g3307 , g3308 , g3309 , g3310 , g3311 , g3312 , g3313 , g3314 , g3315 , g3316 , g3317 , g3318 , g3319 , g3320 , g3321 , g3322 , g3323 , g3324 , g3325 , g3326 , g3327 , g3328 , g3329 , g3330 , g3331 , g3332 , g3333 , g3334 , g3335 , g3336 , g3337 , g3338 , g3339 , g3340 , g3341 , g3342 , g3343 , g3344 , g3345 , g3346 , g3347 , g3348 , g3349 , g3350 , g3351 , g3352 , g3353 , g3354 , g3355 , g3356 , g3357 , g3358 , g3359 , g3360 , g3361 , g3362 , g3363 , g3364 , g3365 , g3366 , g3367 , g3368 , g3369 , g3370 , g3371 , g3372 , g3373 , g3374 , g3375 , g3376 , g3377 , g3378 , g3379 , g3380 , g3381 , g3382 , g3383 , g3384 , g3385 , g3386 , g3387 , g3388 , g3389 , g3390 , g3391 , g3392 , g3393 , g3394 , g3395 , g3396 , g3397 , g3398 , g3399 , g3400 , g3401 , g3402 , g3403 , g3404 , g3405 , g3406 , g3407 , g3408 , g3409 , g3410 , g3411 , g3412 , g3413 , g3414 , g3415 , g3416 , g3417 , g3418 , g3419 , g3420 , g3421 , g3422 , g3423 , g3424 , g3425 , g3426 , g3427 , g3428 , g3429 , g3430 , g3431 , g3432 , g3433 , g3434 , g3435 , g3436 , g3437 , g3438 , g3439 , g3440 , g3441 , g3442 , g3443 , g3444 , g3445 , g3446 , g3447 , g3448 , g3449 , g3450 , g3451 , g3452 , g3453 , g3454 , g3455 , g3456 , g3457 , g3458 , g3459 , g3460 , g3461 , g3462 , g3463 , g3464 , g3465 , g3466 , g3467 , g3468 , g3469 , g3470 , g3471 , g3472 , g3473 , g3474 , g3475 , g3476 , g3477 , g3478 , g3479 , g3480 , g3481 , g3482 , g3483 , g3484 , g3485 , g3486 , g3487 , g3488 , g3489 , g3490 , g3491 , g3492 , g3493 , g3494 , g3495 , g3496 , g3497 , g3498 , g3499 , g3500 , g3501 , g3502 , g3503 , g3504 , g3505 , g3506 , g3507 , g3508 , g3509 , g3510 , g3511 , g3512 , g3513 , g3514 , g3515 , g3516 , g3517 , g3518 , g3519 , g3520 , g3521 , g3522 , g3523 , g3524 , g3525 , g3526 , g3527 , g3528 , g3529 , g3530 , g3531 , g3532 , g3533 , g3534 , g3535 , g3536 , g3537 , g3538 , g3539 , g3540 , g3541 , g3542 , g3543 , g3544 , g3545 , g3546 , g3547 , g3548 , g3549 , g3550 , g3551 , g3552 , g3553 , g3554 , g3555 , g3556 , g3557 , g3558 , g3559 , g3560 , g3561 , g3562 , g3563 , g3564 , g3565 , g3566 , g3567 , g3568 , g3569 , g3570 , g3571 , g3572 , g3573 , g3574 , g3575 , g3576 , g3577 , g3578 , g3579 , g3580 , g3581 , g3582 , g3583 , g3584 , g3585 , g3586 , g3587 , g3588 , g3589 , g3590 , g3591 , g3592 , g3593 , g3594 , g3595 , g3596 , g3597 , g3598 , g3599 , g3600 , g3601 , g3602 , g3603 , g3604 , g3605 , g3606 , g3607 , g3608 , g3609 , g3610 , g3611 , g3612 , g3613 , g3614 , g3615 , g3616 , g3617 , g3618 , g3619 , g3620 , g3621 , g3622 , g3623 , g3624 , g3625 , g3626 , g3627 , g3628 , g3629 , g3630 , g3631 , g3632 , g3633 , g3634 , g3635 , g3636 , g3637 , g3638 , g3639 , g3640 , g3641 , g3642 , g3643 , g3644 , g3645 , g3646 , g3647 , g3648 , g3649 , g3650 , g3651 , g3652 , g3653 , g3654 , g3655 , g3656 , g3657 , g3658 , g3659 , g3660 , g3661 , g3662 , g3663 , g3664 , g3665 , g3666 , g3667 , g3668 , g3669 , g3670 , g3671 , g3672 , g3673 , g3674 , g3675 , g3676 , g3677 , g3678 , g3679 , g3680 , g3681 , g3682 , g3683 , g3684 , g3685 , g3686 , g3687 , g3688 , g3689 , g3690 , g3691 , g3692 , g3693 , g3694 , g3695 , g3696 , g3697 , g3698 , g3699 , g3700 , g3701 , g3702 , g3703 , g3704 , g3705 , g3706 , g3707 , g3708 , g3709 , g3710 , g3711 , g3712 , g3713 , g3714 , g3715 , g3716 , g3717 , g3718 , g3719 , g3720 , g3721 , g3722 , g3723 , g3724 , g3725 , g3726 , g3727 , g3728 , g3729 , g3730 , g3731 , g3732 , g3733 , g3734 , g3735 , g3736 , g3737 , g3738 , g3739 , g3740 , g3741 , g3742 , g3743 , g3744 , g3745 , g3746 , g3747 , g3748 , g3749 , g3750 , g3751 , g3752 , g3753 , g3754 , g3755 , g3756 , g3757 , g3758 , g3759 , g3760 , g3761 , g3762 , g3763 , g3764 , g3765 , g3766 , g3767 , g3768 , g3769 , g3770 , g3771 , g3772 , g3773 , g3774 , g3775 , g3776 , g3777 , g3778 , g3779 , g3780 , g3781 , g3782 , g3783 , g3784 , g3785 , g3786 , g3787 , g3788 , g3789 , g3790 , g3791 , g3792 , g3793 , g3794 , g3795 , g3796 , g3797 , g3798 , g3799 , g3800 , g3801 , g3802 , g3803 , g3804 , g3805 , g3806 , g3807 , g3808 , g3809 , g3810 , g3811 , g3812 , g3813 , g3814 , g3815 , g3816 , g3817 , g3818 , g3819 , g3820 , g3821 , g3822 , g3823 , g3824 , g3825 , g3826 , g3827 , g3828 , g3829 , g3830 , g3831 , g3832 , g3833 , g3834 , g3835 , g3836 , g3837 , g3838 , g3839 , g3840 , g3841 , g3842 , g3843 , g3844 , g3845 , g3846 , g3847 , g3848 , g3849 , g3850 , g3851 , g3852 , g3853 , g3854 , g3855 , g3856 , g3857 , g3858 , g3859 , g3860 , g3861 , g3862 , g3863 , g3864 , g3865 , g3866 , g3867 , g3868 , g3869 , g3870 , g3871 , g3872 , g3873 , g3874 , g3875 , g3876 , g3877 , g3878 , g3879 , g3880 , g3881 , g3882 , g3883 , g3884 , g3885 , g3886 , g3887 , g3888 , g3889 , g3890 , g3891 , g3892 , g3893 , g3894 , g3895 , g3896 , g3897 , g3898 , g3899 , g3900 , g3901 , g3902 , g3903 , g3904 , g3905 , g3906 , g3907 , g3908 , g3909 , g3910 , g3911 , g3912 , g3913 , g3914 , g3915 , g3916 , g3917 , g3918 , g3919 , g3920 , g3921 , g3922 , g3923 , g3924 , g3925 , g3926 , g3927 , g3928 , g3929 , g3930 , g3931 , g3932 , g3933 , g3934 , g3935 , g3936 , g3937 , g3938 , g3939 , g3940 , g3941 , g3942 , g3943 , g3944 , g3945 , g3946 , g3947 , g3948 , g3949 , g3950 , g3951 , g3952 , g3953 , g3954 , g3955 , g3956 , g3957 , g3958 , g3959 , g3960 , g3961 , g3962 , g3963 , g3964 , g3965 , g3966 , g3967 , g3968 , g3969 , g3970 , g3971 , g3972 , g3973 , g3974 , g3975 , g3976 , g3977 , g3978 , g3979 , g3980 , g3981 , g3982 , g3983 , g3984 , g3985 , g3986 , g3987 , g3988 , g3989 , g3990 , g3991 , g3992 , g3993 , g3994 , g3995 , g3996 , g3997 , g3998 , g3999 , g4000 , g4001 , g4002 , g4003 , g4004 , g4005 , g4006 , g4007 , g4008 , g4009 , g4010 , g4011 , g4012 , g4013 , g4014 , g4015 , g4016 , g4017 , g4018 , g4019 , g4020 , g4021 , g4022 , g4023 , g4024 , g4025 , g4026 , g4027 , g4028 , g4029 , g4030 , g4031 , g4032 , g4033 , g4034 , g4035 , g4036 , g4037 , g4038 , g4039 , g4040 , g4041 , g4042 , g4043 , g4044 , g4045 , g4046 , g4047 , g4048 , g4049 , g4050 , g4051 , g4052 , g4053 , g4054 , g4055 , g4056 , g4057 , g4058 , g4059 , g4060 , g4061 , g4062 , g4063 , g4064 , g4065 , g4066 , g4067 , g4068 , g4069 , g4070 , g4071 , g4072 , g4073 , g4074 , g4075 , g4076 , g4077 , g4078 , g4079 , g4080 , g4081 , g4082 , g4083 , g4084 , g4085 , g4086 , g4087 , g4088 , g4089 , g4090 , g4091 , g4092 , g4093 , g4094 , g4095 , g4096 , g4097 , g4098 , g4099 , g4100 , g4101 , g4102 , g4103 , g4104 , g4105 , g4106 , g4107 , g4108 , g4109 , g4110 , g4111 , g4112 , g4113 , g4114 , g4115 , g4116 , g4117 , g4118 , g4119 , g4120 , g4121 , g4122 , g4123 , g4124 , g4125 , g4126 , g4127 , g4128 , g4129 , g4130 , g4131 , g4132 , g4133 , g4134 , g4135 , g4136 , g4137 , g4138 , g4139 , g4140 , g4141 , g4142 , g4143 , g4144 , g4145 , g4146 , g4147 , g4148 , g4149 , g4150 , g4151 , g4152 , g4153 , g4154 , g4155 , g4156 , g4157 , g4158 , g4159 , g4160 , g4161 , g4162 , g4163 , g4164 , g4165 , g4166 , g4167 , g4168 , g4169 , g4170 , g4171 , g4172 , g4173 , g4174 , g4175 , g4176 , g4177 , g4178 , g4179 , g4180 , g4181 , g4182 , g4183 , g4184 , g4185 , g4186 , g4187 , g4188 , g4189 , g4190 , g4191 , g4192 , g4193 , g4194 , g4195 , g4196 , g4197 , g4198 , g4199 , g4200 , g4201 , g4202 , g4203 , g4204 , g4205 , g4206 , g4207 , g4208 , g4209 , g4210 , g4211 , g4212 , g4213 , g4214 , g4215 , g4216 , g4217 , g4218 , g4219 , g4220 , g4221 , g4222 , g4223 , g4224 , g4225 , g4226 , g4227 , g4228 , g4229 , g4230 , g4231 , g4232 , g4233 , g4234 , g4235 , g4236 , g4237 , g4238 , g4239 , g4240 , g4241 , g4242 , g4243 , g4244 , g4245 , g4246 , g4247 , g4248 , g4249 , g4250 , g4251 , g4252 , g4253 , g4254 , g4255 , g4256 , g4257 , g4258 , g4259 , g4260 , g4261 , g4262 , g4263 , g4264 , g4265 , g4266 , g4267 , g4268 , g4269 , g4270 , g4271 , g4272 , g4273 , g4274 , g4275 , g4276 , g4277 , g4278 , g4279 , g4280 , g4281 , g4282 , g4283 , g4284 , g4285 , g4286 , g4287 , g4288 , g4289 , g4290 , g4291 , g4292 , g4293 , g4294 , g4295 , g4296 , g4297 , g4298 , g4299 , g4300 , g4301 , g4302 , g4303 , g4304 , g4305 , g4306 , g4307 , g4308 , g4309 , g4310 , g4311 , g4312 , g4313 , g4314 , g4315 , g4316 , g4317 , g4318 , g4319 , g4320 , g4321 , g4322 , g4323 , g4324 , g4325 , g4326 , g4327 , g4328 , g4329 , g4330 , g4331 , g4332 , g4333 , g4334 , g4335 , g4336 , g4337 , g4338 , g4339 , g4340 , g4341 , g4342 , g4343 , g4344 , g4345 , g4346 , g4347 , g4348 , g4349 , g4350 , g4351 , g4352 , g4353 , g4354 , g4355 , g4356 , g4357 , g4358 , g4359 , g4360 , g4361 , g4362 , g4363 , g4364 , g4365 , g4366 , g4367 , g4368 , g4369 , g4370 , g4371 , g4372 , g4373 , g4374 , g4375 , g4376 , g4377 , g4378 , g4379 , g4380 , g4381 , g4382 , g4383 , g4384 , g4385 , g4386 , g4387 , g4388 , g4389 , g4390 , g4391 , g4392 , g4393 , g4394 , g4395 , g4396 , g4397 , g4398 , g4399 , g4400 , g4401 , g4402 , g4403 , g4404 , g4405 , g4406 , g4407 , g4408 , g4409 , g4410 , g4411 , g4412 , g4413 , g4414 , g4415 , g4416 , g4417 , g4418 , g4419 , g4420 , g4421 , g4422 , g4423 , g4424 , g4425 , g4426 , g4427 , g4428 , g4429 , g4430 , g4431 , g4432 , g4433 , g4434 , g4435 , g4436 , g4437 , g4438 , g4439 , g4440 , g4441 , g4442 , g4443 , g4444 , g4445 , g4446 , g4447 , g4448 , g4449 , g4450 , g4451 , g4452 , g4453 , g4454 , g4455 , g4456 , g4457 , g4458 , g4459 , g4460 , g4461 , g4462 , g4463 , g4464 , g4465 , g4466 , g4467 , g4468 , g4469 , g4470 , g4471 , g4472 , g4473 , g4474 , g4475 , g4476 , g4477 , g4478 , g4479 , g4480 , g4481 , g4482 , g4483 , g4484 , g4485 , g4486 , g4487 , g4488 , g4489 , g4490 , g4491 , g4492 , g4493 , g4494 , g4495 , g4496 , g4497 , g4498 , g4499 , g4500 , g4501 , g4502 , g4503 , g4504 , g4505 , g4506 , g4507 , g4508 , g4509 , g4510 , g4511 , g4512 , g4513 , g4514 , g4515 , g4516 , g4517 , g4518 , g4519 , g4520 , g4521 , g4522 , g4523 , g4524 , g4525 , g4526 , g4527 , g4528 , g4529 , g4530 , g4531 , g4532 , g4533 , g4534 , g4535 , g4536 , g4537 , g4538 , g4539 , g4540 , g4541 , g4542 , g4543 , g4544 , g4545 , g4546 , g4547 , g4548 , g4549 , g4550 , g4551 , g4552 , g4553 , g4554 , g4555 , g4556 , g4557 , g4558 , g4559 , g4560 , g4561 , g4562 , g4563 , g4564 , g4565 , g4566 , g4567 , g4568 , g4569 , g4570 , g4571 , g4572 , g4573 , g4574 , g4575 , g4576 , g4577 , g4578 , g4579 , g4580 , g4581 , g4582 , g4583 , g4584 , g4585 , g4586 , g4587 , g4588 , g4589 , g4590 , g4591 , g4592 , g4593 , g4594 , g4595 , g4596 , g4597 , g4598 , g4599 , g4600 , g4601 , g4602 , g4603 , g4604 , g4605 , g4606 , g4607 , g4608 , g4609 , g4610 , g4611 , g4612 , g4613 , g4614 , g4615 , g4616 , g4617 , g4618 , g4619 , g4620 , g4621 , g4622 , g4623 , g4624 , g4625 , g4626 , g4627 , g4628 , g4629 , g4630 , g4631 , g4632 , g4633 , g4634 , g4635 , g4636 , g4637 , g4638 , g4639 , g4640 , g4641 , g4642 , g4643 , g4644 , g4645 , g4646 , g4647 , g4648 , g4649 , g4650 , g4651 , g4652 , g4653 , g4654 , g4655 , g4656 , g4657 , g4658 , g4659 , g4660 , g4661 , g4662 , g4663 , g4664 , g4665 , g4666 , g4667 , g4668 , g4669 , g4670 , g4671 , g4672 , g4673 , g4674 , g4675 , g4676 , g4677 , g4678 , g4679 , g4680 , g4681 , g4682 , g4683 , g4684 , g4685 , g4686 , g4687 , g4688 , g4689 , g4690 , g4691 , g4692 , g4693 , g4694 , g4695 , g4696 , g4697 , g4698 , g4699 , g4700 , g4701 , g4702 , g4703 , g4704 , g4705 , g4706 , g4707 , g4708 , g4709 , g4710 , g4711 , g4712 , g4713 , g4714 , g4715 , g4716 , g4717 , g4718 , g4719 , g4720 , g4721 , g4722 , g4723 , g4724 , g4725 , g4726 , g4727 , g4728 , g4729 , g4730 , g4731 , g4732 , g4733 , g4734 , g4735 , g4736 , g4737 , g4738 , g4739 , g4740 , g4741 , g4742 , g4743 , g4744 , g4745 , g4746 , g4747 , g4748 , g4749 , g4750 , g4751 , g4752 , g4753 , g4754 , g4755 , g4756 , g4757 , g4758 , g4759 , g4760 , g4761 , g4762 , g4763 , g4764 , g4765 , g4766 , g4767 , g4768 , g4769 , g4770 , g4771 , g4772 , g4773 , g4774 , g4775 , g4776 , g4777 , g4778 , g4779 , g4780 , g4781 , g4782 , g4783 , g4784 , g4785 , g4786 , g4787 , g4788 , g4789 , g4790 , g4791 , g4792 , g4793 , g4794 , g4795 , g4796 , g4797 , g4798 , g4799 , g4800 , g4801 , g4802 , g4803 , g4804 , g4805 , g4806 , g4807 , g4808 , g4809 , g4810 , g4811 , g4812 , g4813 , g4814 , g4815 , g4816 , g4817 , g4818 , g4819 , g4820 , g4821 , g4822 , g4823 , g4824 , g4825 , g4826 , g4827 , g4828 , g4829 , g4830 , g4831 , g4832 , g4833 , g4834 , g4835 , g4836 , g4837 , g4838 , g4839 , g4840 , g4841 , g4842 , g4843 , g4844 , g4845 , g4846 , g4847 , g4848 , g4849 , g4850 , g4851 , g4852 , g4853 , g4854 , g4855 , g4856 , g4857 , g4858 , g4859 , g4860 , g4861 , g4862 , g4863 , g4864 , g4865 , g4866 , g4867 , g4868 , g4869 , g4870 , g4871 , g4872 , g4873 , g4874 , g4875 , g4876 , g4877 , g4878 , g4879 , g4880 , g4881 , g4882 , g4883 , g4884 , g4885 , g4886 , g4887 , g4888 , g4889 , g4890 , g4891 , g4892 , g4893 , g4894 , g4895 , g4896 , g4897 , g4898 , g4899 , g4900 , g4901 , g4902 , g4903 , g4904 , g4905 , g4906 , g4907 , g4908 , g4909 , g4910 , g4911 , g4912 , g4913 , g4914 , g4915 , g4916 , g4917 , g4918 , g4919 , g4920 , g4921 , g4922 , g4923 , g4924 , g4925 , g4926 , g4927 , g4928 , g4929 , g4930 , g4931 , g4932 , g4933 , g4934 , g4935 , g4936 , g4937 , g4938 , g4939 , g4940 , g4941 , g4942 , g4943 , g4944 , g4945 , g4946 , g4947 , g4948 , g4949 , g4950 , g4951 , g4952 , g4953 , g4954 , g4955 , g4956 , g4957 , g4958 , g4959 , g4960 , g4961 , g4962 , g4963 , g4964 , g4965 , g4966 , g4967 , g4968 , g4969 , g4970 , g4971 , g4972 , g4973 , g4974 , g4975 , g4976 , g4977 , g4978 , g4979 , g4980 , g4981 , g4982 , g4983 , g4984 , g4985 , g4986 , g4987 , g4988 , g4989 , g4990 , g4991 , g4992 , g4993 , g4994 , g4995 , g4996 , g4997 , g4998 , g4999 , g5000 , g5001 , g5002 , g5003 , g5004 , g5005 , g5006 , g5007 , g5008 , g5009 , g5010 , g5011 , g5012 , g5013 , g5014 , g5015 , g5016 , g5017 , g5018 , g5019 , g5020 , g5021 , g5022 , g5023 , g5024 , g5025 , g5026 , g5027 , g5028 , g5029 , g5030 , g5031 , g5032 , g5033 , g5034 , g5035 , g5036 , g5037 , g5038 , g5039 , g5040 , g5041 , g5042 , g5043 , g5044 , g5045 , g5046 , g5047 , g5048 , g5049 , g5050 , g5051 , g5052 , g5053 , g5054 , g5055 , g5056 , g5057 , g5058 , g5059 , g5060 , g5061 , g5062 , g5063 , g5064 , g5065 , g5066 , g5067 , g5068 , g5069 , g5070 , g5071 , g5072 , g5073 , g5074 , g5075 , g5076 , g5077 , g5078 , g5079 , g5080 , g5081 , g5082 , g5083 , g5084 , g5085 , g5086 , g5087 , g5088 , g5089 , g5090 , g5091 , g5092 , g5093 , g5094 , g5095 , g5096 , g5097 , g5098 , g5099 , g5100 , g5101 , g5102 , g5103 , g5104 , g5105 , g5106 , g5107 , g5108 , g5109 , g5110 , g5111 , g5112 , g5113 , g5114 , g5115 , g5116 , g5117 , g5118 , g5119 , g5120 , g5121 , g5122 , g5123 , g5124 , g5125 , g5126 , g5127 , g5128 , g5129 , g5130 , g5131 , g5132 , g5133 , g5134 , g5135 , g5136 , g5137 , g5138 , g5139 , g5140 , g5141 , g5142 , g5143 , g5144 , g5145 , g5146 , g5147 , g5148 , g5149 , g5150 , g5151 , g5152 , g5153 , g5154 , g5155 , g5156 , g5157 , g5158 , g5159 , g5160 , g5161 , g5162 , g5163 , g5164 , g5165 , g5166 , g5167 , g5168 , g5169 , g5170 , g5171 , g5172 , g5173 , g5174 , g5175 , g5176 , g5177 , g5178 , g5179 , g5180 , g5181 , g5182 , g5183 , g5184 , g5185 , g5186 , g5187 , g5188 , g5189 , g5190 , g5191 , g5192 , g5193 , g5194 , g5195 , g5196 , g5197 , g5198 , g5199 , g5200 , g5201 , g5202 , g5203 , g5204 , g5205 , g5206 , g5207 , g5208 , g5209 , g5210 , g5211 , g5212 , g5213 , g5214 , g5215 , g5216 , g5217 , g5218 , g5219 , g5220 , g5221 , g5222 , g5223 , g5224 , g5225 , g5226 , g5227 , g5228 , g5229 , g5230 , g5231 , g5232 , g5233 , g5234 , g5235 , g5236 , g5237 , g5238 , g5239 , g5240 , g5241 , g5242 , g5243 , g5244 , g5245 , g5246 , g5247 , g5248 , g5249 , g5250 , g5251 , g5252 , g5253 , g5254 , g5255 , g5256 , g5257 , g5258 , g5259 , g5260 , g5261 , g5262 , g5263 , g5264 , g5265 , g5266 , g5267 , g5268 , g5269 , g5270 , g5271 , g5272 , g5273 , g5274 , g5275 , g5276 , g5277 , g5278 , g5279 , g5280 , g5281 , g5282 , g5283 , g5284 , g5285 , g5286 , g5287 , g5288 , g5289 , g5290 , g5291 , g5292 , g5293 , g5294 , g5295 , g5296 , g5297 , g5298 , g5299 , g5300 , g5301 , g5302 , g5303 , g5304 , g5305 , g5306 , g5307 , g5308 , g5309 , g5310 , g5311 , g5312 , g5313 , g5314 , g5315 , g5316 , g5317 , g5318 , g5319 , g5320 , g5321 , g5322 , g5323 , g5324 , g5325 , g5326 , g5327 , g5328 , g5329 , g5330 , g5331 , g5332 , g5333 , g5334 , g5335 , g5336 , g5337 , g5338 , g5339 , g5340 , g5341 , g5342 , g5343 , g5344 , g5345 , g5346 , g5347 , g5348 , g5349 , g5350 , g5351 , g5352 , g5353 , g5354 , g5355 , g5356 , g5357 , g5358 , g5359 , g5360 , g5361 , g5362 , g5363 , g5364 , g5365 , g5366 , g5367 , g5368 , g5369 , g5370 , g5371 , g5372 , g5373 , g5374 , g5375 , g5376 , g5377 , g5378 , g5379 , g5380 , g5381 , g5382 , g5383 , g5384 , g5385 , g5386 , g5387 , g5388 , g5389 , g5390 , g5391 , g5392 , g5393 , g5394 , g5395 , g5396 , g5397 , g5398 , g5399 , g5400 , g5401 , g5402 , g5403 , g5404 , g5405 , g5406 , g5407 , g5408 , g5409 , g5410 , g5411 , g5412 , g5413 , g5414 , g5415 , g5416 , g5417 , g5418 , g5419 , g5420 , g5421 , g5422 , g5423 , g5424 , g5425 , g5426 , g5427 , g5428 , g5429 , g5430 , g5431 , g5432 , g5433 , g5434 , g5435 , g5436 , g5437 , g5438 , g5439 , g5440 , g5441 , g5442 , g5443 , g5444 , g5445 , g5446 , g5447 , g5448 , g5449 , g5450 , g5451 , g5452 , g5453 , g5454 , g5455 , g5456 , g5457 , g5458 , g5459 , g5460 , g5461 , g5462 , g5463 , g5464 , g5465 , g5466 , g5467 , g5468 , g5469 , g5470 , g5471 , g5472 , g5473 , g5474 , g5475 , g5476 , g5477 , g5478 , g5479 , g5480 , g5481 , g5482 , g5483 , g5484 , g5485 , g5486 , g5487 , g5488 , g5489 , g5490 , g5491 , g5492 , g5493 , g5494 , g5495 , g5496 , g5497 , g5498 , g5499 , g5500 , g5501 , g5502 , g5503 , g5504 , g5505 , g5506 , g5507 , g5508 , g5509 , g5510 , g5511 , g5512 , g5513 , g5514 , g5515 , g5516 , g5517 , g5518 , g5519 , g5520 , g5521 , g5522 , g5523 , g5524 , g5525 , g5526 , g5527 , g5528 , g5529 , g5530 , g5531 , g5532 , g5533 , g5534 , g5535 , g5536 , g5537 , g5538 , g5539 , g5540 , g5541 , g5542 , g5543 , g5544 , g5545 , g5546 , g5547 , g5548 , g5549 , g5550 , g5551 , g5552 , g5553 , g5554 , g5555 , g5556 , g5557 , g5558 , g5559 , g5560 , g5561 , g5562 , g5563 , g5564 , g5565 , g5566 , g5567 , g5568 , g5569 , g5570 , g5571 , g5572 , g5573 , g5574 , g5575 , g5576 , g5577 , g5578 , g5579 , g5580 , g5581 , g5582 , g5583 , g5584 , g5585 , g5586 , g5587 , g5588 , g5589 , g5590 , g5591 , g5592 , g5593 , g5594 , g5595 , g5596 , g5597 , g5598 , g5599 , g5600 , g5601 , g5602 , g5603 , g5604 , g5605 , g5606 , g5607 , g5608 , g5609 , g5610 , g5611 , g5612 , g5613 , g5614 , g5615 , g5616 , g5617 , g5618 , g5619 , g5620 , g5621 , g5622 , g5623 , g5624 , g5625 , g5626 , g5627 , g5628 , g5629 , g5630 , g5631 , g5632 , g5633 , g5634 , g5635 , g5636 , g5637 , g5638 , g5639 , g5640 , g5641 , g5642 , g5643 , g5644 , g5645 , g5646 , g5647 , g5648 , g5649 , g5650 , g5651 , g5652 , g5653 , g5654 , g5655 , g5656 , g5657 , g5658 , g5659 , g5660 , g5661 , g5662 , g5663 , g5664 , g5665 , g5666 , g5667 , g5668 , g5669 , g5670 , g5671 , g5672 , g5673 , g5674 , g5675 , g5676 , g5677 , g5678 , g5679 , g5680 , g5681 , g5682 , g5683 , g5684 , g5685 , g5686 , g5687 , g5688 , g5689 , g5690 , g5691 , g5692 , g5693 , g5694 , g5695 , g5696 , g5697 , g5698 , g5699 , g5700 , g5701 , g5702 , g5703 , g5704 , g5705 , g5706 , g5707 , g5708 , g5709 , g5710 , g5711 , g5712 , g5713 , g5714 , g5715 , g5716 , g5717 , g5718 , g5719 , g5720 , g5721 , g5722 , g5723 , g5724 , g5725 , g5726 , g5727 , g5728 , g5729 , g5730 , g5731 , g5732 , g5733 , g5734 , g5735 , g5736 , g5737 , g5738 , g5739 , g5740 , g5741 , g5742 , g5743 , g5744 , g5745 , g5746 , g5747 , g5748 , g5749 , g5750 , g5751 , g5752 , g5753 , g5754 , g5755 , g5756 , g5757 , g5758 , g5759 , g5760 , g5761 , g5762 , g5763 , g5764 , g5765 , g5766 , g5767 , g5768 , g5769 , g5770 , g5771 , g5772 , g5773 , g5774 , g5775 , g5776 , g5777 , g5778 , g5779 , g5780 , g5781 , g5782 , g5783 , g5784 , g5785 , g5786 , g5787 , g5788 , g5789 , g5790 , g5791 , g5792 , g5793 , g5794 , g5795 , g5796 , g5797 , g5798 , g5799 , g5800 , g5801 , g5802 , g5803 , g5804 , g5805 , g5806 , g5807 , g5808 , g5809 , g5810 , g5811 , g5812 , g5813 , g5814 , g5815 , g5816 , g5817 , g5818 , g5819 , g5820 , g5821 , g5822 , g5823 , g5824 , g5825 , g5826 , g5827 , g5828 , g5829 , g5830 , g5831 , g5832 , g5833 , g5834 , g5835 , g5836 , g5837 , g5838 , g5839 , g5840 , g5841 , g5842 , g5843 , g5844 , g5845 , g5846 , g5847 , g5848 , g5849 , g5850 , g5851 , g5852 , g5853 , g5854 , g5855 , g5856 , g5857 , g5858 , g5859 , g5860 , g5861 , g5862 , g5863 , g5864 , g5865 , g5866 , g5867 , g5868 , g5869 , g5870 , g5871 , g5872 , g5873 , g5874 , g5875 , g5876 , g5877 , g5878 , g5879 , g5880 , g5881 , g5882 , g5883 , g5884 , g5885 , g5886 , g5887 , g5888 , g5889 , g5890 , g5891 , g5892 , g5893 , g5894 , g5895 , g5896 , g5897 , g5898 , g5899 , g5900 , g5901 , g5902 , g5903 , g5904 , g5905 , g5906 , g5907 , g5908 , g5909 , g5910 , g5911 , g5912 , g5913 , g5914 , g5915 , g5916 , g5917 , g5918 , g5919 , g5920 , g5921 , g5922 , g5923 , g5924 , g5925 , g5926 , g5927 , g5928 , g5929 , g5930 , g5931 , g5932 , g5933 , g5934 , g5935 , g5936 , g5937 , g5938 , g5939 , g5940 , g5941 , g5942 , g5943 , g5944 , g5945 , g5946 , g5947 , g5948 , g5949 , g5950 , g5951 , g5952 , g5953 , g5954 , g5955 , g5956 , g5957 , g5958 , g5959 , g5960 , g5961 , g5962 , g5963 , g5964 , g5965 , g5966 , g5967 , g5968 , g5969 , g5970 , g5971 , g5972 , g5973 , g5974 , g5975 , g5976 , g5977 , g5978 , g5979 , g5980 , g5981 , g5982 , g5983 , g5984 , g5985 , g5986 , g5987 , g5988 , g5989 , g5990 , g5991 , g5992 , g5993 , g5994 , g5995 , g5996 , g5997 , g5998 , g5999 , g6000 , g6001 , g6002 , g6003 , g6004 , g6005 , g6006 , g6007 , g6008 , g6009 , g6010 , g6011 , g6012 , g6013 , g6014 , g6015 , g6016 , g6017 , g6018 , g6019 , g6020 , g6021 , g6022 , g6023 , g6024 , g6025 , g6026 , g6027 , g6028 , g6029 , g6030 , g6031 , g6032 , g6033 , g6034 , g6035 , g6036 , g6037 , g6038 , g6039 , g6040 , g6041 , g6042 , g6043 , g6044 , g6045 , g6046 , g6047 , g6048 , g6049 , g6050 , g6051 , g6052 , g6053 , g6054 , g6055 , g6056 , g6057 , g6058 , g6059 , g6060 , g6061 , g6062 , g6063 , g6064 , g6065 , g6066 , g6067 , g6068 , g6069 , g6070 , g6071 , g6072 , g6073 , g6074 , g6075 , g6076 , g6077 , g6078 , g6079 , g6080 , g6081 , g6082 , g6083 , g6084 , g6085 , g6086 , g6087 , g6088 , g6089 , g6090 , g6091 , g6092 , g6093 , g6094 , g6095 , g6096 , g6097 , g6098 , g6099 , g6100 , g6101 , g6102 , g6103 , g6104 , g6105 , g6106 , g6107 , g6108 , g6109 , g6110 , g6111 , g6112 , g6113 , g6114 , g6115 , g6116 , g6117 , g6118 , g6119 , g6120 , g6121 , g6122 , g6123 , g6124 , g6125 , g6126 , g6127 , g6128 , g6129 , g6130 , g6131 , g6132 , g6133 , g6134 , g6135 , g6136 , g6137 , g6138 , g6139 , g6140 , g6141 , g6142 , g6143 , g6144 , g6145 , g6146 , g6147 , g6148 , g6149 , g6150 , g6151 , g6152 , g6153 , g6154 , g6155 , g6156 , g6157 , g6158 , g6159 , g6160 , g6161 , g6162 , g6163 , g6164 , g6165 , g6166 , g6167 , g6168 , g6169 , g6170 , g6171 , g6172 , g6173 , g6174 , g6175 , g6176 , g6177 , g6178 , g6179 , g6180 , g6181 , g6182 , g6183 , g6184 , g6185 , g6186 , g6187 , g6188 , g6189 , g6190 , g6191 , g6192 , g6193 , g6194 , g6195 , g6196 , g6197 , g6198 , g6199 , g6200 , g6201 , g6202 , g6203 , g6204 , g6205 , g6206 , g6207 , g6208 , g6209 , g6210 , g6211 , g6212 , g6213 , g6214 , g6215 , g6216 , g6217 , g6218 , g6219 , g6220 , g6221 , g6222 , g6223 , g6224 , g6225 , g6226 , g6227 , g6228 , g6229 , g6230 , g6231 , g6232 , g6233 , g6234 , g6235 , g6236 , g6237 , g6238 , g6239 , g6240 , g6241 , g6242 , g6243 , g6244 , g6245 , g6246 , g6247 , g6248 , g6249 , g6250 , g6251 , g6252 , g6253 , g6254 , g6255 , g6256 , g6257 , g6258 , g6259 , g6260 , g6261 , g6262 , g6263 , g6264 , g6265 , g6266 , g6267 , g6268 , g6269 , g6270 , g6271 , g6272 , g6273 , g6274 , g6275 , g6276 , g6277 , g6278 , g6279 , g6280 , g6281 , g6282 , g6283 , g6284 , g6285 , g6286 , g6287 , g6288 , g6289 , g6290 , g6291 , g6292 , g6293 , g6294 , g6295 , g6296 , g6297 , g6298 , g6299 , g6300 , g6301 , g6302 , g6303 , g6304 , g6305 , g6306 , g6307 , g6308 , g6309 , g6310 , g6311 , g6312 , g6313 , g6314 , g6315 , g6316 , g6317 , g6318 , g6319 , g6320 , g6321 , g6322 , g6323 , g6324 , g6325 , g6326 , g6327 , g6328 , g6329 , g6330 , g6331 , g6332 , g6333 , g6334 , g6335 , g6336 , g6337 , g6338 , g6339 , g6340 , g6341 , g6342 , g6343 , g6344 , g6345 , g6346 , g6347 , g6348 , g6349 , g6350 , g6351 , g6352 , g6353 , g6354 , g6355 , g6356 , g6357 , g6358 , g6359 , g6360 , g6361 , g6362 , g6363 , g6364 , g6365 , g6366 , g6367 , g6368 , g6369 , g6370 , g6371 , g6372 , g6373 , g6374 , g6375 , g6376 , g6377 , g6378 , g6379 , g6380 , g6381 , g6382 , g6383 , g6384 , g6385 , g6386 , g6387 , g6388 , g6389 , g6390 , g6391 , g6392 , g6393 , g6394 , g6395 , g6396 , g6397 , g6398 , g6399 , g6400 , g6401 , g6402 , g6403 , g6404 , g6405 , g6406 , g6407 , g6408 , g6409 , g6410 , g6411 , g6412 , g6413 , g6414 , g6415 , g6416 , g6417 , g6418 , g6419 , g6420 , g6421 , g6422 , g6423 , g6424 , g6425 , g6426 , g6427 , g6428 , g6429 , g6430 , g6431 , g6432 , g6433 , g6434 , g6435 , g6436 , g6437 , g6438 , g6439 , g6440 , g6441 , g6442 , g6443 , g6444 , g6445 , g6446 , g6447 , g6448 , g6449 , g6450 , g6451 , g6452 , g6453 , g6454 , g6455 , g6456 , g6457 , g6458 , g6459 , g6460 , g6461 , g6462 , g6463 , g6464 , g6465 , g6466 , g6467 , g6468 , g6469 , g6470 , g6471 , g6472 , g6473 , g6474 , g6475 , g6476 , g6477 , g6478 , g6479 , g6480 , g6481 , g6482 , g6483 , g6484 , g6485 , g6486 , g6487 , g6488 , g6489 , g6490 , g6491 , g6492 , g6493 , g6494 , g6495 , g6496 , g6497 , g6498 , g6499 , g6500 , g6501 , g6502 , g6503 , g6504 , g6505 , g6506 , g6507 , g6508 , g6509 , g6510 , g6511 , g6512 , g6513 , g6514 , g6515 , g6516 , g6517 , g6518 , g6519 , g6520 , g6521 , g6522 , g6523 , g6524 , g6525 , g6526 , g6527 , g6528 , g6529 , g6530 , g6531 , g6532 , g6533 , g6534 , g6535 , g6536 , g6537 , g6538 , g6539 , g6540 , g6541 , g6542 , g6543 , g6544 , g6545 , g6546 , g6547 , g6548 , g6549 , g6550 , g6551 , g6552 , g6553 , g6554 , g6555 , g6556 , g6557 , g6558 , g6559 , g6560 , g6561 , g6562 , g6563 , g6564 , g6565 , g6566 , g6567 , g6568 , g6569 , g6570 , g6571 , g6572 , g6573 , g6574 , g6575 , g6576 , g6577 , g6578 , g6579 , g6580 , g6581 , g6582 , g6583 , g6584 , g6585 , g6586 , g6587 , g6588 , g6589 , g6590 , g6591 , g6592 , g6593 , g6594 , g6595 , g6596 , g6597 , g6598 , g6599 , g6600 , g6601 , g6602 , g6603 , g6604 , g6605 , g6606 , g6607 , g6608 , g6609 , g6610 , g6611 , g6612 , g6613 , g6614 , g6615 , g6616 , g6617 , g6618 , g6619 , g6620 , g6621 , g6622 , g6623 , g6624 , g6625 , g6626 , g6627 , g6628 , g6629 , g6630 , g6631 , g6632 , g6633 , g6634 , g6635 , g6636 , g6637 , g6638 , g6639 , g6640 , g6641 , g6642 , g6643 , g6644 , g6645 , g6646 , g6647 , g6648 , g6649 , g6650 , g6651 , g6652 , g6653 , g6654 , g6655 , g6656 , g6657 , g6658 , g6659 , g6660 , g6661 , g6662 , g6663 , g6664 , g6665 , g6666 , g6667 , g6668 , g6669 , g6670 , g6671 , g6672 , g6673 , g6674 , g6675 , g6676 , g6677 , g6678 , g6679 , g6680 , g6681 , g6682 , g6683 , g6684 , g6685 , g6686 , g6687 , g6688 , g6689 , g6690 , g6691 , g6692 , g6693 , g6694 , g6695 , g6696 , g6697 , g6698 , g6699 , g6700 , g6701 , g6702 , g6703 , g6704 , g6705 , g6706 , g6707 , g6708 , g6709 , g6710 , g6711 , g6712 , g6713 , g6714 , g6715 , g6716 , g6717 , g6718 , g6719 , g6720 , g6721 , g6722 , g6723 , g6724 , g6725 , g6726 , g6727 , g6728 , g6729 , g6730 , g6731 , g6732 , g6733 , g6734 , g6735 , g6736 , g6737 , g6738 , g6739 , g6740 , g6741 , g6742 , g6743 , g6744 , g6745 , g6746 , g6747 , g6748 , g6749 , g6750 , g6751 , g6752 , g6753 , g6754 , g6755 , g6756 , g6757 , g6758 , g6759 , g6760 , g6761 , g6762 , g6763 , g6764 , g6765 , g6766 , g6767 , g6768 , g6769 , g6770 , g6771 , g6772 , g6773 , g6774 , g6775 , g6776 , g6777 , g6778 , g6779 , g6780 , g6781 , g6782 , g6783 , g6784 , g6785 , g6786 , g6787 , g6788 , g6789 , g6790 , g6791 , g6792 , g6793 , g6794 , g6795 , g6796 , g6797 , g6798 , g6799 , g6800 , g6801 , g6802 , g6803 , g6804 , g6805 , g6806 , g6807 , g6808 , g6809 , g6810 , g6811 , g6812 , g6813 , g6814 , g6815 , g6816 , g6817 , g6818 , g6819 , g6820 , g6821 , g6822 , g6823 , g6824 , g6825 , g6826 , g6827 , g6828 , g6829 , g6830 , g6831 , g6832 , g6833 , g6834 , g6835 , g6836 , g6837 , g6838 , g6839 , g6840 , g6841 , g6842 , g6843 , g6844 , g6845 , g6846 , g6847 , g6848 , g6849 , g6850 , g6851 , g6852 , g6853 , g6854 , g6855 , g6856 , g6857 , g6858 , g6859 , g6860 , g6861 , g6862 , g6863 , g6864 , g6865 , g6866 , g6867 , g6868 , g6869 , g6870 , g6871 , g6872 , g6873 , g6874 , g6875 , g6876 , g6877 , g6878 , g6879 , g6880 , g6881 , g6882 , g6883 , g6884 , g6885 , g6886 , g6887 , g6888 , g6889 , g6890 , g6891 , g6892 , g6893 , g6894 , g6895 , g6896 , g6897 , g6898 , g6899 , g6900 , g6901 , g6902 , g6903 , g6904 , g6905 , g6906 , g6907 , g6908 , g6909 , g6910 , g6911 , g6912 , g6913 , g6914 , g6915 , g6916 , g6917 , g6918 , g6919 , g6920 , g6921 , g6922 , g6923 , g6924 , g6925 , g6926 , g6927 , g6928 , g6929 , g6930 , g6931 , g6932 , g6933 , g6934 , g6935 , g6936 , g6937 , g6938 , g6939 , g6940 , g6941 , g6942 , g6943 , g6944 , g6945 , g6946 , g6947 , g6948 , g6949 , g6950 , g6951 , g6952 , g6953 , g6954 , g6955 , g6956 , g6957 , g6958 , g6959 , g6960 , g6961 , g6962 , g6963 , g6964 , g6965 , g6966 , g6967 , g6968 , g6969 , g6970 , g6971 , g6972 , g6973 , g6974 , g6975 , g6976 , g6977 , g6978 , g6979 , g6980 , g6981 , g6982 , g6983 , g6984 , g6985 , g6986 , g6987 , g6988 , g6989 , g6990 , g6991 , g6992 , g6993 , g6994 , g6995 , g6996 , g6997 , g6998 , g6999 , g7000 , g7001 , g7002 , g7003 , g7004 , g7005 , g7006 , g7007 , g7008 , g7009 , g7010 , g7011 , g7012 , g7013 , g7014 , g7015 , g7016 , g7017 , g7018 , g7019 , g7020 , g7021 , g7022 , g7023 , g7024 , g7025 , g7026 , g7027 , g7028 , g7029 , g7030 , g7031 , g7032 , g7033 , g7034 , g7035 , g7036 , g7037 , g7038 , g7039 , g7040 , g7041 , g7042 , g7043 , g7044 , g7045 , g7046 , g7047 , g7048 , g7049 , g7050 , g7051 , g7052 , g7053 , g7054 , g7055 , g7056 , g7057 , g7058 , g7059 , g7060 , g7061 , g7062 , g7063 , g7064 , g7065 , g7066 , g7067 , g7068 , g7069 , g7070 , g7071 , g7072 , g7073 , g7074 , g7075 , g7076 , g7077 , g7078 , g7079 , g7080 , g7081 , g7082 , g7083 , g7084 , g7085 , g7086 , g7087 , g7088 , g7089 , g7090 , g7091 , g7092 , g7093 , g7094 , g7095 , g7096 , g7097 , g7098 , g7099 , g7100 , g7101 , g7102 , g7103 , g7104 , g7105 , g7106 , g7107 , g7108 , g7109 , g7110 , g7111 , g7112 , g7113 , g7114 , g7115 , g7116 , g7117 , g7118 , g7119 , g7120 , g7121 , g7122 , g7123 , g7124 , g7125 , g7126 , g7127 , g7128 , g7129 , g7130 , g7131 , g7132 , g7133 , g7134 , g7135 , g7136 , g7137 , g7138 , g7139 , g7140 , g7141 , g7142 , g7143 , g7144 , g7145 , g7146 , g7147 , g7148 , g7149 , g7150 , g7151 , g7152 , g7153 , g7154 , g7155 , g7156 , g7157 , g7158 , g7159 , g7160 , g7161 , g7162 , g7163 , g7164 , g7165 , g7166 , g7167 , g7168 , g7169 , g7170 , g7171 , g7172 , g7173 , g7174 , g7175 , g7176 , g7177 , g7178 , g7179 , g7180 , g7181 , g7182 , g7183 , g7184 , g7185 , g7186 , g7187 , g7188 , g7189 , g7190 , g7191 , g7192 , g7193 , g7194 , g7195 , g7196 , g7197 , g7198 , g7199 , g7200 , g7201 , g7202 , g7203 , g7204 , g7205 , g7206 , g7207 , g7208 , g7209 , g7210 , g7211 , g7212 , g7213 , g7214 , g7215 , g7216 , g7217 , g7218 , g7219 , g7220 , g7221 , g7222 , g7223 , g7224 , g7225 , g7226 , g7227 , g7228 , g7229 , g7230 , g7231 , g7232 , g7233 , g7234 , g7235 , g7236 , g7237 , g7238 , g7239 , g7240 , g7241 , g7242 , g7243 , g7244 , g7245 , g7246 , g7247 , g7248 , g7249 , g7250 , g7251 , g7252 , g7253 , g7254 , g7255 , g7256 , g7257 , g7258 , g7259 , g7260 , g7261 , g7262 , g7263 , g7264 , g7265 , g7266 , g7267 , g7268 , g7269 , g7270 , g7271 , g7272 , g7273 , g7274 , g7275 , g7276 , g7277 , g7278 , g7279 , g7280 , g7281 , g7282 , g7283 , g7284 , g7285 , g7286 , g7287 , g7288 , g7289 , g7290 , g7291 , g7292 , g7293 , g7294 , g7295 , g7296 , g7297 , g7298 , g7299 , g7300 , g7301 , g7302 , g7303 , g7304 , g7305 , g7306 , g7307 , g7308 , g7309 , g7310 , g7311 , g7312 , g7313 , g7314 , g7315 , g7316 , g7317 , g7318 , g7319 , g7320 , g7321 , g7322 , g7323 , g7324 , g7325 , g7326 , g7327 , g7328 , g7329 , g7330 , g7331 , g7332 , g7333 , g7334 , g7335 , g7336 , g7337 , g7338 , g7339 , g7340 , g7341 , g7342 , g7343 , g7344 , g7345 , g7346 , g7347 , g7348 , g7349 , g7350 , g7351 , g7352 , g7353 , g7354 , g7355 , g7356 , g7357 , g7358 , g7359 , g7360 , g7361 , g7362 , g7363 , g7364 , g7365 , g7366 , g7367 , g7368 , g7369 , g7370 , g7371 , g7372 , g7373 , g7374 , g7375 , g7376 , g7377 , g7378 , g7379 , g7380 , g7381 , g7382 , g7383 , g7384 , g7385 , g7386 , g7387 , g7388 , g7389 , g7390 , g7391 , g7392 , g7393 , g7394 , g7395 , g7396 , g7397 , g7398 , g7399 , g7400 , g7401 , g7402 , g7403 , g7404 , g7405 , g7406 , g7407 , g7408 , g7409 , g7410 , g7411 , g7412 , g7413 , g7414 , g7415 , g7416 , g7417 , g7418 , g7419 , g7420 , g7421 , g7422 , g7423 , g7424 , g7425 , g7426 , g7427 , g7428 , g7429 , g7430 , g7431 , g7432 , g7433 , g7434 , g7435 , g7436 , g7437 , g7438 , g7439 , g7440 , g7441 , g7442 , g7443 , g7444 , g7445 , g7446 , g7447 , g7448 , g7449 , g7450 , g7451 , g7452 , g7453 , g7454 , g7455 , g7456 , g7457 , g7458 , g7459 , g7460 , g7461 , g7462 , g7463 , g7464 , g7465 , g7466 , g7467 , g7468 , g7469 , g7470 , g7471 , g7472 , g7473 , g7474 , g7475 , g7476 , g7477 , g7478 , g7479 , g7480 , g7481 , g7482 , g7483 , g7484 , g7485 , g7486 , g7487 , g7488 , g7489 , g7490 , g7491 , g7492 , g7493 , g7494 , g7495 , g7496 , g7497 , g7498 , g7499 , g7500 , g7501 , g7502 , g7503 , g7504 , g7505 , g7506 , g7507 , g7508 , g7509 , g7510 , g7511 , g7512 , g7513 , g7514 , g7515 , g7516 , g7517 , g7518 , g7519 , g7520 , g7521 , g7522 , g7523 , g7524 , g7525 , g7526 , g7527 , g7528 , g7529 , g7530 , g7531 , g7532 , g7533 , g7534 , g7535 , g7536 , g7537 , g7538 , g7539 , g7540 , g7541 , g7542 , g7543 , g7544 , g7545 , g7546 , g7547 , g7548 , g7549 , g7550 , g7551 , g7552 , g7553 , g7554 , g7555 , g7556 , g7557 , g7558 , g7559 , g7560 , g7561 , g7562 , g7563 , g7564 , g7565 , g7566 , g7567 , g7568 , g7569 , g7570 , g7571 , g7572 , g7573 , g7574 , g7575 , g7576 , g7577 , g7578 , g7579 , g7580 , g7581 , g7582 , g7583 , g7584 , g7585 , g7586 , g7587 , g7588 , g7589 , g7590 , g7591 , g7592 , g7593 , g7594 , g7595 , g7596 , g7597 , g7598 , g7599 , g7600 , g7601 , g7602 , g7603 , g7604 , g7605 , g7606 , g7607 , g7608 , g7609 , g7610 , g7611 , g7612 , g7613 , g7614 , g7615 , g7616 , g7617 , g7618 , g7619 , g7620 , g7621 , g7622 , g7623 , g7624 , g7625 , g7626 , g7627 , g7628 , g7629 , g7630 , g7631 , g7632 , g7633 , g7634 , g7635 , g7636 , g7637 , g7638 , g7639 , g7640 , g7641 , g7642 , g7643 , g7644 , g7645 , g7646 , g7647 , g7648 , g7649 , g7650 , g7651 , g7652 , g7653 , g7654 , g7655 , g7656 , g7657 , g7658 , g7659 , g7660 , g7661 , g7662 , g7663 , g7664 , g7665 , g7666 , g7667 , g7668 , g7669 , g7670 , g7671 , g7672 , g7673 , g7674 , g7675 , g7676 , g7677 , g7678 , g7679 , g7680 , g7681 , g7682 , g7683 , g7684 , g7685 , g7686 , g7687 , g7688 , g7689 , g7690 , g7691 , g7692 , g7693 , g7694 , g7695 , g7696 , g7697 , g7698 , g7699 , g7700 , g7701 , g7702 , g7703 , g7704 , g7705 , g7706 , g7707 , g7708 , g7709 , g7710 , g7711 , g7712 , g7713 , g7714 , g7715 , g7716 , g7717 , g7718 , g7719 , g7720 , g7721 , g7722 , g7723 , g7724 , g7725 , g7726 , g7727 , g7728 , g7729 , g7730 , g7731 , g7732 , g7733 , g7734 , g7735 , g7736 , g7737 , g7738 , g7739 , g7740 , g7741 , g7742 , g7743 , g7744 , g7745 , g7746 , g7747 , g7748 , g7749 , g7750 , g7751 , g7752 , g7753 , g7754 , g7755 , g7756 , g7757 , g7758 , g7759 , g7760 , g7761 , g7762 , g7763 , g7764 , g7765 , g7766 , g7767 , g7768 , g7769 , g7770 , g7771 , g7772 , g7773 , g7774 , g7775 , g7776 , g7777 , g7778 , g7779 , g7780 , g7781 , g7782 , g7783 , g7784 , g7785 , g7786 , g7787 , g7788 , g7789 , g7790 , g7791 , g7792 , g7793 , g7794 , g7795 , g7796 , g7797 , g7798 , g7799 , g7800 , g7801 , g7802 , g7803 , g7804 , g7805 , g7806 , g7807 , g7808 , g7809 , g7810 , g7811 , g7812 , g7813 , g7814 , g7815 , g7816 , g7817 , g7818 , g7819 , g7820 , g7821 , g7822 , g7823 , g7824 , g7825 , g7826 , g7827 , g7828 , g7829 , g7830 , g7831 , g7832 , g7833 , g7834 , g7835 , g7836 , g7837 , g7838 , g7839 , g7840 , g7841 , g7842 , g7843 , g7844 , g7845 , g7846 , g7847 , g7848 , g7849 , g7850 , g7851 , g7852 , g7853 , g7854 , g7855 , g7856 , g7857 , g7858 , g7859 , g7860 , g7861 , g7862 , g7863 , g7864 , g7865 , g7866 , g7867 , g7868 , g7869 , g7870 , g7871 , g7872 , g7873 , g7874 , g7875 , g7876 , g7877 , g7878 , g7879 , g7880 , g7881 , g7882 , g7883 , g7884 , g7885 , g7886 , g7887 , g7888 , g7889 , g7890 , g7891 , g7892 , g7893 , g7894 , g7895 , g7896 , g7897 , g7898 , g7899 , g7900 , g7901 , g7902 , g7903 , g7904 , g7905 , g7906 , g7907 , g7908 , g7909 , g7910 , g7911 , g7912 , g7913 , g7914 , g7915 , g7916 , g7917 , g7918 , g7919 , g7920 , g7921 , g7922 , g7923 , g7924 , g7925 , g7926 , g7927 , g7928 , g7929 , g7930 , g7931 , g7932 , g7933 , g7934 , g7935 , g7936 , g7937 , g7938 , g7939 , g7940 , g7941 , g7942 , g7943 , g7944 , g7945 , g7946 , g7947 , g7948 , g7949 , g7950 , g7951 , g7952 , g7953 , g7954 , g7955 , g7956 , g7957 , g7958 , g7959 , g7960 , g7961 , g7962 , g7963 , g7964 , g7965 , g7966 , g7967 , g7968 , g7969 , g7970 , g7971 , g7972 , g7973 , g7974 , g7975 , g7976 , g7977 , g7978 , g7979 , g7980 , g7981 , g7982 , g7983 , g7984 , g7985 , g7986 , g7987 , g7988 , g7989 , g7990 , g7991 , g7992 , g7993 , g7994 , g7995 , g7996 , g7997 , g7998 , g7999 , g8000 , g8001 , g8002 , g8003 , g8004 , g8005 , g8006 , g8007 , g8008 , g8009 , g8010 , g8011 , g8012 , g8013 , g8014 , g8015 , g8016 , g8017 , g8018 , g8019 , g8020 , g8021 , g8022 , g8023 , g8024 , g8025 , g8026 , g8027 , g8028 , g8029 , g8030 , g8031 , g8032 , g8033 , g8034 , g8035 , g8036 , g8037 , g8038 , g8039 , g8040 , g8041 , g8042 , g8043 , g8044 , g8045 , g8046 , g8047 , g8048 , g8049 , g8050 , g8051 , g8052 , g8053 , g8054 , g8055 , g8056 , g8057 , g8058 , g8059 , g8060 , g8061 , g8062 , g8063 , g8064 , g8065 , g8066 , g8067 , g8068 , g8069 , g8070 , g8071 , g8072 , g8073 , g8074 , g8075 , g8076 , g8077 , g8078 , g8079 , g8080 , g8081 , g8082 , g8083 , g8084 , g8085 , g8086 , g8087 , g8088 , g8089 , g8090 , g8091 , g8092 , g8093 , g8094 , g8095 , g8096 , g8097 , g8098 , g8099 , g8100 , g8101 , g8102 , g8103 , g8104 , g8105 , g8106 , g8107 , g8108 , g8109 , g8110 , g8111 , g8112 , g8113 , g8114 , g8115 , g8116 , g8117 , g8118 , g8119 , g8120 , g8121 , g8122 , g8123 , g8124 , g8125 , g8126 , g8127 , g8128 , g8129 , g8130 , g8131 , g8132 , g8133 , g8134 , g8135 , g8136 , g8137 , g8138 , g8139 , g8140 , g8141 , g8142 , g8143 , g8144 , g8145 , g8146 , g8147 , g8148 , g8149 , g8150 , g8151 , g8152 , g8153 , g8154 , g8155 , g8156 , g8157 , g8158 , g8159 , g8160 , g8161 , g8162 , g8163 , g8164 , g8165 , g8166 , g8167 , g8168 , g8169 , g8170 , g8171 , g8172 , g8173 , g8174 , g8175 , g8176 , g8177 , g8178 , g8179 , g8180 , g8181 , g8182 , g8183 , g8184 , g8185 , g8186 , g8187 , g8188 , g8189 , g8190 , g8191 , g8192 , g8193 , g8194 , g8195 , g8196 , g8197 , g8198 , g8199 , g8200 , g8201 , g8202 , g8203 , g8204 , g8205 , g8206 , g8207 , g8208 , g8209 , g8210 , g8211 , g8212 , g8213 , g8214 , g8215 , g8216 , g8217 , g8218 , g8219 , g8220 , g8221 , g8222 , g8223 , g8224 , g8225 , g8226 , g8227 , g8228 , g8229 , g8230 , g8231 , g8232 , g8233 , g8234 , g8235 , g8236 , g8237 , g8238 , g8239 , g8240 , g8241 , g8242 , g8243 , g8244 , g8245 , g8246 , g8247 , g8248 , g8249 , g8250 , g8251 , g8252 , g8253 , g8254 , g8255 , g8256 , g8257 , g8258 , g8259 , g8260 , g8261 , g8262 , g8263 , g8264 , g8265 , g8266 , g8267 , g8268 , g8269 , g8270 , g8271 , g8272 , g8273 , g8274 , g8275 , g8276 , g8277 , g8278 , g8279 , g8280 , g8281 , g8282 , g8283 , g8284 , g8285 , g8286 , g8287 , g8288 , g8289 , g8290 , g8291 , g8292 , g8293 , g8294 , g8295 , g8296 , g8297 , g8298 , g8299 , g8300 , g8301 , g8302 , g8303 , g8304 , g8305 , g8306 , g8307 , g8308 , g8309 , g8310 , g8311 , g8312 , g8313 , g8314 , g8315 , g8316 , g8317 , g8318 , g8319 , g8320 , g8321 , g8322 , g8323 , g8324 , g8325 , g8326 , g8327 , g8328 , g8329 , g8330 , g8331 , g8332 , g8333 , g8334 , g8335 , g8336 , g8337 , g8338 , g8339 , g8340 , g8341 , g8342 , g8343 , g8344 , g8345 , g8346 , g8347 , g8348 , g8349 , g8350 , g8351 , g8352 , g8353 , g8354 , g8355 , g8356 , g8357 , g8358 , g8359 , g8360 , g8361 , g8362 , g8363 , g8364 , g8365 , g8366 , g8367 , g8368 , g8369 , g8370 , g8371 , g8372 , g8373 , g8374 , g8375 , g8376 , g8377 , g8378 , g8379 , g8380 , g8381 , g8382 , g8383 , g8384 , g8385 , g8386 , g8387 , g8388 , g8389 , g8390 , g8391 , g8392 , g8393 , g8394 , g8395 , g8396 , g8397 , g8398 , g8399 , g8400 , g8401 , g8402 , g8403 , g8404 , g8405 , g8406 , g8407 , g8408 , g8409 , g8410 , g8411 , g8412 , g8413 , g8414 , g8415 , g8416 , g8417 , g8418 , g8419 , g8420 , g8421 , g8422 , g8423 , g8424 , g8425 , g8426 , g8427 , g8428 , g8429 , g8430 , g8431 , g8432 , g8433 , g8434 , g8435 , g8436 , g8437 , g8438 , g8439 , g8440 , g8441 , g8442 , g8443 , g8444 , g8445 , g8446 , g8447 , g8448 , g8449 , g8450 , g8451 , g8452 , g8453 , g8454 , g8455 , g8456 , g8457 , g8458 , g8459 , g8460 , g8461 , g8462 , g8463 , g8464 , g8465 , g8466 , g8467 , g8468 , g8469 , g8470 , g8471 , g8472 , g8473 , g8474 , g8475 , g8476 , g8477 , g8478 , g8479 , g8480 , g8481 , g8482 , g8483 , g8484 , g8485 , g8486 , g8487 , g8488 , g8489 , g8490 , g8491 , g8492 , g8493 , g8494 , g8495 , g8496 , g8497 , g8498 , g8499 , g8500 , g8501 , g8502 , g8503 , g8504 , g8505 , g8506 , g8507 , g8508 , g8509 , g8510 , g8511 , g8512 , g8513 , g8514 , g8515 , g8516 , g8517 , g8518 , g8519 , g8520 , g8521 , g8522 , g8523 , g8524 , g8525 , g8526 , g8527 , g8528 , g8529 , g8530 , g8531 , g8532 , g8533 , g8534 , g8535 , g8536 , g8537 , g8538 , g8539 , g8540 , g8541 , g8542 , g8543 , g8544 , g8545 , g8546 , g8547 , g8548 , g8549 , g8550 , g8551 , g8552 , g8553 , g8554 , g8555 , g8556 , g8557 , g8558 , g8559 , g8560 , g8561 , g8562 , g8563 , g8564 , g8565 , g8566 , g8567 , g8568 , g8569 , g8570 , g8571 , g8572 , g8573 , g8574 , g8575 , g8576 , g8577 , g8578 , g8579 , g8580 , g8581 , g8582 , g8583 , g8584 , g8585 , g8586 , g8587 , g8588 , g8589 , g8590 , g8591 , g8592 , g8593 , g8594 , g8595 , g8596 , g8597 , g8598 , g8599 , g8600 , g8601 , g8602 , g8603 , g8604 , g8605 , g8606 , g8607 , g8608 , g8609 , g8610 , g8611 , g8612 , g8613 , g8614 , g8615 , g8616 , g8617 , g8618 , g8619 , g8620 , g8621 , g8622 , g8623 , g8624 , g8625 , g8626 , g8627 , g8628 , g8629 , g8630 , g8631 , g8632 , g8633 , g8634 , g8635 , g8636 , g8637 , g8638 , g8639 , g8640 , g8641 , g8642 , g8643 , g8644 , g8645 , g8646 , g8647 , g8648 , g8649 , g8650 , g8651 , g8652 , g8653 , g8654 , g8655 , g8656 , g8657 , g8658 , g8659 , g8660 , g8661 , g8662 , g8663 , g8664 , g8665 , g8666 , g8667 , g8668 , g8669 , g8670 , g8671 , g8672 , g8673 , g8674 , g8675 , g8676 , g8677 , g8678 , g8679 , g8680 , g8681 , g8682 , g8683 , g8684 , g8685 , g8686 , g8687 , g8688 , g8689 , g8690 , g8691 , g8692 , g8693 , g8694 , g8695 , g8696 , g8697 , g8698 , g8699 , g8700 , g8701 , g8702 , g8703 , g8704 , g8705 , g8706 , g8707 , g8708 , g8709 , g8710 , g8711 , g8712 , g8713 , g8714 , g8715 , g8716 , g8717 , g8718 , g8719 , g8720 , g8721 , g8722 , g8723 , g8724 , g8725 , g8726 , g8727 , g8728 , g8729 , g8730 , g8731 , g8732 , g8733 , g8734 , g8735 , g8736 , g8737 , g8738 , g8739 , g8740 , g8741 , g8742 , g8743 , g8744 , g8745 , g8746 , g8747 , g8748 , g8749 , g8750 , g8751 , g8752 , g8753 , g8754 , g8755 , g8756 , g8757 , g8758 , g8759 , g8760 , g8761 , g8762 , g8763 , g8764 , g8765 , g8766 , g8767 , g8768 , g8769 , g8770 , g8771 , g8772 , g8773 , g8774 , g8775 , g8776 , g8777 , g8778 , g8779 , g8780 , g8781 , g8782 , g8783 , g8784 , g8785 , g8786 , g8787 , g8788 , g8789 , g8790 , g8791 , g8792 , g8793 , g8794 , g8795 , g8796 , g8797 , g8798 , g8799 , g8800 , g8801 , g8802 , g8803 , g8804 , g8805 , g8806 , g8807 , g8808 , g8809 , g8810 , g8811 , g8812 , g8813 , g8814 , g8815 , g8816 , g8817 , g8818 , g8819 , g8820 , g8821 , g8822 , g8823 , g8824 , g8825 , g8826 , g8827 , g8828 , g8829 , g8830 , g8831 , g8832 , g8833 , g8834 , g8835 , g8836 , g8837 , g8838 , g8839 , g8840 , g8841 , g8842 , g8843 , g8844 , g8845 , g8846 , g8847 , g8848 , g8849 , g8850 , g8851 , g8852 , g8853 , g8854 , g8855 , g8856 , g8857 , g8858 , g8859 , g8860 , g8861 , g8862 , g8863 , g8864 , g8865 , g8866 , g8867 , g8868 , g8869 , g8870 , g8871 , g8872 , g8873 , g8874 , g8875 , g8876 , g8877 , g8878 , g8879 , g8880 , g8881 , g8882 , g8883 , g8884 , g8885 , g8886 , g8887 , g8888 , g8889 , g8890 , g8891 , g8892 , g8893 , g8894 , g8895 , g8896 , g8897 , g8898 , g8899 , g8900 , g8901 , g8902 , g8903 , g8904 , g8905 , g8906 , g8907 , g8908 , g8909 , g8910 , g8911 , g8912 , g8913 , g8914 , g8915 , g8916 , g8917 , g8918 , g8919 , g8920 , g8921 , g8922 , g8923 , g8924 , g8925 , g8926 , g8927 , g8928 , g8929 , g8930 , g8931 , g8932 , g8933 , g8934 , g8935 , g8936 , g8937 , g8938 , g8939 , g8940 , g8941 , g8942 , g8943 , g8944 , g8945 , g8946 , g8947 , g8948 , g8949 , g8950 , g8951 , g8952 , g8953 , g8954 , g8955 , g8956 , g8957 , g8958 , g8959 , g8960 , g8961 , g8962 , g8963 , g8964 , g8965 , g8966 , g8967 , g8968 , g8969 , g8970 , g8971 , g8972 , g8973 , g8974 , g8975 , g8976 , g8977 , g8978 ;

wire n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , 
     n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , 
     n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , 
     n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , 
     n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , 
     n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , 
     n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , 
     n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , 
     n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , 
     n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , 
     n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , 
     n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , 
     n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , 
     n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , 
     n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , 
     n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , 
     n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , 
     n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , 
     n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , 
     n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , 
     n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , 
     n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , 
     n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , 
     n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , 
     n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , 
     n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , 
     n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , 
     n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , 
     n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , 
     n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , 
     n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , 
     n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , 
     n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , 
     n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , 
     n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , 
     n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , 
     n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , 
     n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , 
     n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , 
     n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , 
     n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , 
     n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , 
     n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , 
     n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , 
     n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , 
     n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , 
     n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , 
     n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , 
     n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , 
     n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , 
     n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , 
     n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , 
     n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , 
     n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , 
     n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , 
     n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , 
     n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , 
     n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , 
     n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , 
     n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , 
     n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , 
     n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , 
     n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , 
     n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , 
     n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , 
     n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , 
     n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , 
     n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , 
     n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , 
     n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , 
     n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , 
     n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , 
     n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , 
     n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , 
     n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , 
     n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , 
     n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , 
     n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , 
     n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , 
     n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , 
     n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , 
     n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , 
     n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , 
     n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , 
     n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , 
     n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , 
     n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , 
     n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , 
     n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , 
     n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , 
     n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , 
     n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , 
     n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , 
     n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , 
     n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , 
     n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , 
     n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , 
     n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , 
     n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , 
     n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , 
     n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , 
     n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , 
     n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , 
     n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , 
     n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , 
     n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , 
     n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , 
     n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , 
     n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , 
     n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , 
     n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , 
     n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , 
     n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , 
     n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , 
     n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , 
     n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , 
     n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , 
     n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , 
     n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , 
     n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , 
     n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , 
     n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , 
     n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , 
     n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , 
     n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , 
     n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , 
     n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , 
     n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , 
     n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , 
     n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , 
     n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , 
     n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , 
     n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , 
     n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , 
     n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , 
     n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , 
     n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , 
     n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , 
     n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , 
     n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , 
     n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , 
     n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , 
     n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , 
     n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , 
     n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , 
     n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , 
     n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , 
     n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , 
     n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , 
     n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , 
     n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , 
     n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , 
     n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , 
     n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , 
     n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , 
     n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , 
     n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , 
     n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , 
     n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , 
     n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , 
     n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , 
     n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , 
     n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , 
     n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , 
     n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , 
     n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , 
     n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , 
     n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , 
     n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , 
     n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , 
     n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , 
     n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , 
     n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , 
     n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , 
     n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , 
     n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , 
     n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , 
     n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , 
     n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , 
     n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , 
     n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , 
     n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , 
     n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , 
     n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , 
     n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , 
     n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , 
     n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , 
     n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , 
     n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , 
     n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , 
     n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , 
     n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , 
     n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , 
     n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , 
     n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , 
     n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , 
     n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , 
     n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , 
     n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , 
     n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , 
     n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , 
     n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , 
     n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , 
     n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , 
     n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , 
     n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , 
     n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , 
     n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , 
     n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , 
     n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , 
     n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , 
     n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , 
     n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , 
     n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , 
     n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , 
     n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , 
     n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , 
     n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , 
     n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , 
     n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , 
     n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , 
     n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , 
     n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , 
     n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , 
     n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , 
     n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , 
     n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , 
     n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , 
     n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , 
     n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , 
     n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , 
     n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , 
     n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , 
     n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , 
     n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , 
     n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , 
     n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , 
     n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , 
     n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , 
     n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , 
     n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , 
     n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , 
     n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , 
     n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , 
     n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , 
     n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , 
     n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , 
     n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , 
     n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , 
     n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , 
     n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , 
     n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , 
     n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , 
     n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , 
     n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , 
     n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , 
     n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , 
     n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , 
     n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , 
     n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , 
     n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , 
     n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , 
     n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , 
     n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , 
     n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , 
     n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , 
     n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , 
     n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , 
     n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , 
     n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , 
     n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , 
     n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , 
     n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , 
     n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , 
     n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , 
     n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , 
     n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , 
     n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , 
     n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , 
     n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , 
     n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , 
     n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , 
     n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , 
     n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , 
     n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , 
     n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , 
     n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , 
     n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , 
     n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , 
     n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , 
     n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , 
     n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , 
     n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , 
     n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , 
     n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , 
     n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , 
     n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , 
     n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , 
     n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , 
     n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , 
     n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , 
     n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , 
     n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , 
     n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , 
     n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , 
     n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , 
     n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , 
     n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , 
     n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , 
     n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , 
     n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , 
     n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , 
     n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , 
     n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , 
     n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , 
     n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , 
     n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , 
     n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , 
     n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , 
     n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , 
     n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , 
     n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , 
     n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , 
     n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , 
     n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , 
     n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , 
     n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , 
     n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , 
     n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , 
     n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , 
     n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , 
     n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , 
     n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , 
     n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , 
     n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , 
     n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , 
     n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , 
     n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , 
     n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , 
     n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , 
     n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , 
     n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , 
     n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , 
     n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , 
     n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , 
     n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , 
     n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , 
     n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , 
     n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , 
     n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , 
     n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , 
     n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , 
     n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , 
     n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , 
     n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , 
     n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , 
     n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , 
     n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , 
     n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , 
     n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , 
     n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , 
     n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , 
     n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , 
     n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , 
     n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , 
     n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , 
     n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , 
     n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , 
     n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , 
     n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , 
     n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , 
     n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , 
     n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , 
     n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , 
     n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , 
     n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , 
     n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , 
     n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , 
     n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , 
     n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , 
     n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , 
     n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , 
     n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , 
     n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , 
     n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , 
     n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , 
     n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , 
     n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , 
     n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , 
     n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , 
     n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , 
     n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , 
     n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , 
     n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , 
     n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , 
     n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , 
     n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , 
     n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , 
     n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , 
     n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , 
     n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , 
     n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , 
     n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , 
     n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , 
     n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , 
     n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , 
     n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , 
     n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , 
     n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , 
     n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , 
     n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , 
     n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , 
     n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , 
     n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , 
     n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , 
     n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , 
     n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , 
     n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , 
     n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , 
     n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , 
     n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , 
     n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , 
     n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , 
     n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , 
     n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , 
     n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , 
     n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , 
     n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , 
     n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , 
     n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , 
     n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , 
     n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , 
     n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , 
     n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , 
     n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , 
     n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , 
     n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , 
     n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , 
     n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , 
     n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , 
     n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , 
     n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , 
     n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , 
     n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , 
     n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , 
     n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , 
     n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , 
     n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , 
     n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , 
     n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , 
     n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , 
     n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , 
     n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , 
     n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , 
     n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , 
     n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , 
     n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , 
     n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , 
     n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , 
     n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , 
     n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , 
     n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , 
     n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , 
     n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , 
     n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , 
     n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , 
     n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , 
     n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , 
     n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , 
     n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , 
     n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , 
     n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , 
     n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , 
     n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , 
     n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , 
     n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , 
     n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , 
     n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , 
     n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , 
     n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , 
     n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , 
     n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , 
     n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , 
     n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , 
     n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , 
     n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , 
     n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , 
     n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , 
     n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , 
     n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , 
     n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , 
     n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , 
     n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , 
     n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , 
     n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , 
     n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , 
     n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , 
     n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , 
     n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , 
     n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , 
     n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , 
     n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , 
     n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , 
     n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , 
     n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , 
     n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , 
     n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , 
     n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , 
     n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , 
     n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , 
     n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , 
     n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , 
     n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , 
     n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , 
     n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , 
     n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , 
     n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , 
     n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , 
     n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , 
     n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , 
     n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , 
     n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , 
     n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , 
     n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , 
     n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , 
     n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , 
     n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , 
     n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , 
     n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , 
     n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , 
     n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , 
     n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , 
     n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , 
     n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , 
     n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , 
     n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , 
     n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , 
     n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , 
     n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , 
     n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , 
     n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , 
     n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , 
     n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , 
     n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , 
     n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , 
     n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , 
     n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , 
     n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , 
     n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , 
     n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , 
     n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , 
     n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , 
     n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , 
     n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , 
     n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , 
     n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , 
     n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , 
     n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , 
     n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , 
     n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , 
     n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , 
     n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , 
     n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , 
     n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , 
     n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , 
     n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , 
     n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , 
     n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , 
     n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , 
     n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , 
     n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , 
     n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , 
     n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , 
     n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , 
     n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , 
     n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , 
     n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , 
     n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , 
     n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , 
     n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , 
     n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , 
     n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , 
     n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , 
     n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , 
     n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , 
     n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , 
     n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , 
     n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , 
     n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , 
     n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , 
     n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , 
     n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , 
     n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , 
     n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , 
     n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , 
     n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , 
     n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , 
     n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , 
     n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , 
     n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , 
     n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , 
     n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , 
     n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , 
     n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , 
     n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , 
     n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , 
     n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , 
     n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , 
     n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , 
     n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , 
     n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , 
     n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , 
     n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , 
     n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , 
     n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , 
     n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , 
     n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , 
     n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , 
     n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , 
     n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , 
     n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , 
     n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , 
     n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , 
     n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , 
     n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , 
     n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , 
     n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , 
     n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , 
     n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , 
     n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , 
     n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , 
     n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , 
     n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , 
     n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , 
     n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , 
     n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , 
     n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , 
     n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , 
     n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , 
     n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , 
     n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , 
     n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , 
     n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , 
     n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , 
     n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , 
     n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , 
     n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , 
     n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , 
     n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , 
     n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , 
     n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , 
     n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , 
     n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , 
     n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , 
     n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , 
     n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , 
     n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , 
     n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , 
     n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , 
     n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , 
     n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , 
     n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , 
     n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , 
     n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , 
     n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , 
     n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , 
     n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , 
     n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , 
     n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , 
     n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , 
     n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , 
     n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , 
     n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , 
     n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , 
     n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , 
     n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , 
     n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , 
     n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , 
     n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , 
     n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , 
     n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , 
     n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , 
     n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , 
     n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , 
     n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , 
     n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , 
     n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , 
     n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , 
     n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , 
     n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , 
     n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , 
     n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , 
     n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , 
     n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , 
     n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , 
     n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , 
     n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , 
     n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , 
     n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , 
     n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , 
     n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , 
     n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , 
     n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , 
     n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , 
     n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , 
     n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , 
     n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , 
     n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , 
     n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , 
     n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , 
     n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , 
     n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , 
     n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , 
     n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , 
     n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , 
     n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , 
     n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , 
     n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , 
     n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , 
     n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , 
     n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , 
     n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , 
     n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , 
     n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , 
     n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , 
     n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , 
     n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , 
     n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , 
     n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , 
     n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , 
     n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , 
     n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , 
     n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , 
     n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , 
     n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , 
     n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , 
     n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , 
     n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , 
     n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , 
     n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , 
     n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , 
     n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , 
     n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , 
     n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , 
     n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , 
     n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , 
     n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , 
     n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , 
     n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , 
     n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , 
     n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , 
     n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , 
     n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , 
     n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , 
     n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , 
     n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , 
     n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , 
     n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , 
     n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , 
     n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , 
     n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , 
     n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , 
     n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , 
     n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , 
     n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , 
     n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , 
     n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , 
     n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , 
     n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , 
     n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , 
     n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , 
     n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , 
     n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , 
     n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , 
     n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , 
     n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , 
     n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , 
     n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , 
     n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , 
     n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , 
     n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , 
     n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , 
     n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , 
     n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , 
     n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , 
     n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , 
     n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , 
     n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , 
     n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , 
     n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , 
     n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , 
     n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , 
     n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , 
     n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , 
     n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , 
     n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , 
     n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , 
     n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , 
     n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , 
     n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , 
     n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , 
     n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , 
     n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , 
     n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , 
     n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , 
     n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , 
     n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , 
     n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , 
     n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , 
     n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , 
     n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , 
     n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , 
     n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , 
     n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , 
     n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , 
     n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , 
     n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , 
     n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , 
     n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , 
     n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , 
     n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , 
     n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , 
     n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , 
     n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , 
     n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , 
     n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , 
     n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , 
     n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , 
     n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , 
     n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , 
     n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , 
     n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , 
     n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , 
     n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , 
     n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , 
     n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , 
     n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , 
     n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , 
     n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , 
     n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , 
     n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , 
     n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , 
     n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , 
     n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , 
     n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , 
     n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , 
     n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , 
     n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , 
     n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , 
     n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , 
     n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , 
     n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , 
     n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , 
     n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , 
     n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , 
     n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , 
     n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , 
     n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , 
     n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , 
     n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , 
     n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , 
     n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , 
     n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , 
     n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , 
     n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , 
     n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , 
     n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , 
     n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , 
     n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , 
     n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , 
     n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , 
     n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , 
     n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , 
     n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , 
     n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , 
     n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , 
     n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , 
     n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , 
     n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , 
     n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , 
     n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , 
     n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , 
     n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , 
     n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , 
     n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , 
     n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , 
     n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , 
     n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , 
     n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , 
     n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , 
     n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , 
     n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , 
     n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , 
     n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , 
     n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , 
     n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , 
     n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , 
     n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , 
     n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , 
     n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , 
     n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , 
     n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , 
     n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , 
     n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , 
     n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , 
     n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , 
     n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , 
     n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , 
     n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , 
     n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , 
     n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , 
     n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , 
     n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , 
     n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , 
     n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , 
     n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , 
     n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , 
     n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , 
     n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , 
     n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , 
     n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , 
     n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , 
     n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , 
     n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , 
     n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , 
     n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , 
     n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , 
     n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , 
     n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , 
     n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , 
     n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , 
     n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , 
     n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , 
     n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , 
     n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , 
     n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , 
     n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , 
     n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , 
     n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , 
     n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , 
     n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , 
     n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , 
     n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , 
     n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , 
     n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , 
     n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , 
     n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , 
     n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , 
     n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , 
     n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , 
     n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , 
     n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , 
     n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , 
     n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , 
     n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , 
     n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , 
     n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , 
     n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , 
     n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , 
     n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , 
     n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , 
     n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , 
     n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , 
     n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , 
     n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , 
     n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , 
     n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , 
     n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , 
     n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , 
     n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , 
     n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , 
     n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , 
     n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , 
     n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , 
     n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , 
     n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , 
     n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , 
     n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , 
     n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , 
     n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , 
     n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , 
     n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , 
     n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , 
     n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , 
     n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , 
     n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , 
     n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , 
     n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , 
     n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , 
     n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , 
     n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , 
     n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , 
     n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , 
     n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , 
     n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , 
     n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , 
     n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , 
     n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , 
     n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , 
     n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , 
     n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , 
     n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , 
     n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , 
     n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , 
     n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , 
     n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , 
     n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , 
     n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , 
     n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , 
     n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , 
     n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , 
     n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , 
     n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , 
     n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , 
     n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , 
     n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , 
     n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , 
     n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , 
     n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , 
     n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , 
     n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , 
     n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , 
     n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , 
     n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , 
     n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , 
     n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , 
     n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , 
     n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , 
     n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , 
     n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , 
     n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , 
     n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , 
     n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , 
     n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , 
     n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , 
     n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , 
     n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , 
     n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , 
     n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , 
     n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , 
     n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , 
     n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , 
     n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , 
     n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , 
     n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , 
     n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , 
     n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , 
     n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , 
     n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , 
     n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , 
     n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , 
     n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , 
     n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , 
     n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , 
     n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , 
     n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , 
     n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , 
     n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , 
     n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , 
     n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , 
     n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , 
     n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , 
     n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , 
     n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , 
     n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , 
     n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , 
     n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , 
     n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , 
     n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , 
     n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , 
     n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , 
     n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , 
     n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , 
     n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , 
     n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , 
     n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , 
     n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , 
     n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , 
     n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , 
     n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , 
     n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , 
     n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , 
     n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , 
     n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , 
     n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , 
     n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , 
     n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , 
     n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , 
     n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , 
     n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , 
     n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , 
     n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , 
     n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , 
     n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , 
     n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , 
     n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , 
     n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , 
     n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , 
     n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , 
     n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , 
     n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , 
     n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , 
     n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , 
     n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , 
     n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , 
     n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , 
     n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , 
     n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , 
     n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , 
     n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , 
     n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , 
     n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , 
     n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , 
     n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , 
     n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , 
     n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , 
     n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , 
     n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , 
     n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , 
     n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , 
     n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , 
     n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , 
     n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , 
     n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , 
     n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , 
     n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , 
     n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , 
     n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , 
     n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , 
     n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , 
     n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , 
     n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , 
     n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , 
     n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , 
     n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , 
     n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , 
     n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , 
     n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , 
     n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , 
     n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , 
     n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , 
     n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , 
     n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , 
     n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , 
     n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , 
     n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , 
     n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , 
     n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , 
     n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , 
     n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , 
     n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , 
     n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , 
     n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , 
     n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , 
     n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , 
     n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , 
     n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , 
     n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , 
     n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , 
     n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , 
     n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , 
     n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , 
     n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , 
     n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , 
     n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , 
     n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , 
     n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , 
     n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , 
     n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , 
     n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , 
     n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , 
     n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , 
     n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , 
     n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , 
     n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , 
     n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , 
     n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , 
     n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , 
     n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , 
     n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , 
     n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , 
     n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , 
     n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , 
     n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , 
     n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , 
     n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , 
     n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , 
     n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , 
     n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , 
     n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , 
     n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , 
     n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , 
     n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , 
     n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , 
     n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , 
     n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , 
     n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , 
     n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , 
     n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , 
     n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , 
     n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , 
     n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , 
     n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , 
     n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , 
     n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , 
     n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , 
     n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , 
     n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , 
     n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , 
     n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , 
     n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , 
     n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , 
     n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , 
     n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , 
     n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , 
     n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , 
     n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , 
     n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , 
     n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , 
     n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , 
     n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , 
     n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , 
     n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , 
     n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , 
     n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , 
     n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , 
     n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , 
     n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , 
     n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , 
     n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , 
     n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , 
     n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , 
     n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , 
     n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , 
     n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , 
     n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , 
     n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , 
     n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , 
     n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , 
     n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , 
     n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , 
     n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , 
     n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , 
     n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , 
     n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , 
     n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , 
     n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , 
     n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , 
     n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , 
     n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , 
     n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , 
     n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , 
     n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , 
     n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , 
     n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , 
     n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , 
     n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , 
     n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , 
     n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , 
     n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , 
     n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , 
     n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , 
     n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , 
     n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , 
     n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , 
     n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , 
     n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , 
     n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , 
     n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , 
     n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , 
     n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , 
     n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , 
     n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , 
     n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , 
     n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , 
     n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , 
     n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , 
     n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , 
     n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , 
     n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , 
     n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , 
     n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , 
     n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , 
     n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , 
     n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , 
     n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , 
     n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , 
     n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , 
     n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , 
     n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , 
     n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , 
     n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , 
     n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , 
     n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , 
     n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , 
     n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , 
     n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , 
     n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , 
     n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , 
     n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , 
     n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , 
     n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , 
     n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , 
     n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , 
     n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , 
     n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , 
     n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , 
     n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , 
     n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , 
     n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , 
     n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , 
     n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , 
     n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , 
     n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , 
     n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , 
     n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , 
     n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , 
     n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , 
     n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , 
     n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , 
     n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , 
     n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , 
     n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , 
     n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , 
     n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , 
     n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , 
     n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , 
     n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , 
     n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , 
     n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , 
     n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , 
     n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , 
     n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , 
     n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , 
     n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , 
     n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , 
     n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , 
     n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , 
     n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , 
     n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , 
     n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , 
     n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , 
     n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , 
     n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , 
     n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , 
     n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , 
     n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , 
     n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , 
     n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , 
     n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , 
     n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , 
     n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , 
     n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , 
     n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , 
     n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , 
     n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , 
     n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , 
     n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , 
     n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , 
     n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , 
     n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , 
     n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , 
     n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , 
     n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , 
     n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , 
     n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , 
     n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , 
     n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , 
     n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , 
     n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , 
     n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , 
     n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , 
     n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , 
     n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , 
     n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , 
     n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , 
     n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , 
     n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , 
     n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , 
     n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , 
     n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , 
     n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , 
     n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , 
     n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , 
     n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , 
     n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , 
     n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , 
     n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , 
     n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , 
     n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , 
     n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , 
     n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , 
     n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , 
     n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , 
     n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , 
     n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , 
     n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , 
     n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , 
     n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , 
     n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , 
     n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , 
     n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , 
     n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , 
     n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , 
     n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , 
     n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , 
     n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , 
     n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , 
     n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , 
     n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , 
     n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , 
     n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , 
     n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , 
     n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , 
     n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , 
     n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , 
     n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , 
     n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , 
     n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , 
     n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , 
     n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , 
     n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , 
     n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , 
     n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , 
     n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , 
     n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , 
     n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , 
     n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , 
     n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , 
     n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , 
     n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , 
     n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , 
     n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , 
     n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , 
     n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , 
     n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , 
     n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , 
     n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , 
     n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , 
     n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , 
     n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , 
     n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , 
     n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , 
     n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , 
     n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , 
     n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , 
     n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , 
     n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , 
     n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , 
     n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , 
     n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , 
     n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , 
     n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , 
     n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , 
     n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , 
     n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , 
     n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , 
     n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , 
     n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , 
     n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , 
     n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , 
     n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , 
     n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , 
     n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , 
     n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , 
     n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , 
     n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , 
     n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , 
     n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , 
     n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , 
     n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , 
     n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , 
     n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , 
     n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , 
     n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , 
     n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , 
     n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , 
     n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , 
     n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , 
     n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , 
     n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , 
     n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , 
     n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , 
     n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , 
     n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , 
     n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , 
     n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , 
     n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , 
     n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , 
     n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , 
     n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , 
     n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , 
     n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , 
     n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , 
     n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , 
     n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , 
     n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , 
     n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , 
     n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , 
     n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , 
     n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , 
     n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , 
     n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , 
     n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , 
     n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , 
     n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , 
     n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , 
     n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , 
     n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , 
     n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , 
     n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , 
     n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , 
     n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , 
     n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , 
     n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , 
     n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , 
     n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , 
     n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , 
     n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , 
     n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , 
     n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , 
     n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , 
     n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , 
     n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , 
     n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , 
     n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , 
     n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , 
     n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , 
     n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , 
     n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , 
     n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , 
     n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , 
     n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , 
     n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , 
     n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , 
     n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , 
     n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , 
     n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , 
     n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , 
     n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , 
     n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , 
     n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , 
     n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , 
     n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , 
     n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , 
     n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , 
     n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , 
     n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , 
     n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , 
     n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , 
     n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , 
     n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , 
     n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , 
     n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , 
     n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , 
     n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , 
     n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , 
     n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , 
     n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , 
     n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , 
     n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , 
     n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , 
     n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , 
     n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , 
     n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , 
     n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , 
     n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , 
     n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , 
     n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , 
     n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , 
     n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , 
     n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , 
     n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , 
     n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , 
     n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , 
     n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , 
     n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , 
     n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , 
     n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , 
     n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , 
     n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , 
     n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , 
     n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , 
     n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , 
     n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , 
     n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , 
     n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , 
     n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , 
     n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , 
     n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , 
     n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , 
     n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , 
     n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , 
     n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , 
     n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , 
     n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , 
     n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , 
     n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , 
     n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , 
     n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , 
     n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , 
     n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , 
     n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , 
     n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , 
     n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , 
     n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , 
     n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , 
     n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , 
     n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , 
     n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , 
     n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , 
     n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , 
     n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , 
     n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , 
     n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , 
     n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , 
     n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , 
     n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , 
     n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , 
     n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , 
     n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , 
     n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , 
     n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , 
     n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , 
     n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , 
     n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , 
     n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , 
     n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , 
     n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , 
     n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , 
     n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , 
     n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , 
     n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , 
     n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , 
     n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , 
     n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , 
     n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , 
     n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , 
     n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , 
     n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , 
     n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , 
     n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , 
     n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , 
     n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , 
     n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , 
     n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , 
     n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , 
     n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , 
     n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , 
     n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , 
     n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , 
     n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , 
     n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , 
     n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , 
     n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , 
     n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , 
     n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , 
     n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , 
     n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , 
     n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , 
     n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , 
     n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , 
     n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , 
     n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , 
     n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , 
     n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , 
     n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , 
     n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , 
     n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , 
     n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , 
     n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , 
     n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , 
     n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , 
     n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , 
     n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , 
     n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , 
     n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , 
     n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , 
     n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , 
     n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , 
     n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , 
     n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , 
     n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , 
     n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , 
     n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , 
     n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , 
     n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , 
     n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , 
     n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , 
     n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , 
     n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , 
     n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , 
     n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , 
     n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , 
     n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , 
     n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , 
     n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , 
     n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , 
     n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , 
     n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , 
     n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , 
     n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , 
     n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , 
     n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , 
     n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , 
     n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , 
     n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , 
     n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , 
     n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , 
     n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , 
     n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , 
     n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , 
     n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , 
     n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , 
     n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , 
     n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , 
     n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , 
     n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , 
     n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , 
     n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , 
     n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , 
     n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , 
     n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , 
     n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , 
     n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , 
     n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , 
     n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , 
     n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , 
     n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , 
     n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , 
     n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , 
     n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , 
     n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , 
     n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , 
     n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , 
     n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , 
     n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , 
     n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , 
     n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , 
     n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , 
     n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , 
     n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , 
     n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , 
     n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , 
     n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , 
     n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , 
     n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , 
     n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , 
     n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , 
     n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , 
     n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , 
     n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , 
     n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , 
     n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , 
     n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , 
     n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , 
     n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , 
     n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , 
     n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , 
     n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , 
     n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , 
     n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , 
     n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , 
     n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , 
     n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , 
     n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , 
     n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , 
     n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , 
     n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , 
     n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , 
     n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , 
     n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , 
     n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , 
     n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , 
     n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , 
     n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , 
     n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , 
     n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , 
     n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , 
     n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , 
     n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , 
     n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , 
     n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , 
     n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , 
     n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , 
     n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , 
     n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , 
     n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , 
     n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , 
     n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , 
     n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , 
     n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , 
     n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , 
     n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , 
     n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , 
     n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , 
     n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , 
     n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , 
     n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , 
     n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , 
     n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , 
     n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , 
     n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , 
     n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , 
     n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , 
     n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , 
     n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , 
     n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , 
     n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , 
     n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , 
     n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , 
     n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , 
     n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , 
     n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , 
     n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , 
     n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , 
     n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , 
     n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , 
     n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , 
     n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , 
     n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , 
     n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , 
     n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , 
     n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , 
     n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , 
     n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , 
     n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , 
     n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , 
     n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , 
     n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , 
     n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , 
     n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , 
     n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , 
     n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , 
     n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , 
     n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , 
     n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , 
     n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , 
     n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , 
     n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , 
     n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , 
     n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , 
     n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , 
     n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , 
     n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , 
     n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , 
     n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , 
     n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , 
     n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , 
     n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , 
     n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , 
     n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , 
     n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , 
     n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , 
     n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , 
     n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , 
     n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , 
     n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , 
     n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , 
     n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , 
     n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , 
     n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , 
     n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , 
     n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , 
     n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , 
     n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , 
     n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , 
     n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , 
     n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , 
     n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , 
     n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , 
     n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , 
     n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , 
     n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , 
     n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , 
     n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , 
     n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , 
     n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , 
     n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , 
     n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , 
     n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , 
     n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , 
     n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , 
     n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , 
     n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , 
     n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , 
     n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , 
     n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , 
     n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , 
     n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , 
     n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , 
     n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , 
     n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , 
     n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , 
     n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , 
     n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , 
     n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , 
     n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , 
     n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , 
     n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , 
     n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , 
     n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , 
     n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , 
     n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , 
     n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , 
     n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , 
     n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , 
     n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , 
     n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , 
     n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , 
     n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , 
     n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , 
     n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , 
     n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , 
     n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , 
     n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , 
     n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , 
     n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , 
     n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , 
     n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , 
     n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , 
     n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , 
     n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , 
     n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , 
     n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , 
     n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , 
     n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , 
     n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , 
     n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , 
     n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , 
     n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , 
     n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , 
     n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , 
     n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , 
     n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , 
     n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , 
     n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , 
     n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , 
     n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , 
     n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , 
     n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , 
     n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , 
     n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , 
     n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , 
     n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , 
     n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , 
     n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , 
     n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , 
     n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , 
     n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , 
     n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , 
     n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , 
     n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , 
     n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , 
     n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , 
     n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , 
     n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , 
     n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , 
     n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , 
     n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , 
     n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , 
     n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , 
     n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , 
     n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , 
     n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , 
     n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , 
     n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , 
     n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , 
     n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , 
     n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , 
     n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , 
     n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , 
     n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , 
     n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , 
     n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , 
     n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , 
     n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , 
     n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , 
     n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , 
     n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , 
     n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , 
     n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , 
     n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , 
     n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , 
     n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , 
     n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , 
     n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , 
     n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , 
     n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , 
     n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , 
     n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , 
     n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , 
     n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , 
     n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , 
     n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , 
     n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , 
     n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , 
     n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , 
     n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , 
     n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , 
     n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , 
     n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , 
     n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , 
     n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , 
     n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , 
     n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , 
     n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , 
     n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , 
     n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , 
     n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , 
     n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , 
     n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , 
     n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , 
     n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , 
     n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , 
     n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , 
     n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , 
     n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , 
     n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , 
     n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , 
     n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , 
     n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , 
     n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , 
     n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , 
     n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , 
     n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , 
     n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , 
     n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , 
     n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , 
     n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , 
     n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , 
     n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , 
     n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , 
     n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , 
     n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , 
     n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , 
     n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , 
     n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , 
     n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , 
     n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , 
     n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , 
     n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , 
     n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , 
     n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , 
     n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , 
     n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , 
     n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , 
     n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , 
     n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , 
     n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , 
     n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , 
     n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , 
     n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , 
     n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , 
     n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , 
     n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , 
     n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , 
     n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , 
     n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , 
     n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , 
     n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , 
     n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , 
     n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , 
     n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , 
     n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , 
     n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , 
     n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , 
     n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , 
     n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , 
     n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , 
     n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , 
     n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , 
     n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , 
     n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , 
     n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , 
     n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , 
     n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , 
     n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , 
     n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , 
     n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , 
     n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , 
     n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , 
     n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , 
     n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , 
     n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , 
     n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , 
     n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , 
     n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , 
     n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , 
     n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , 
     n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , 
     n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , 
     n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , 
     n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , 
     n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , 
     n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , 
     n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , 
     n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , 
     n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , 
     n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , 
     n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , 
     n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , 
     n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , 
     n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , 
     n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , 
     n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , 
     n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , 
     n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , 
     n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , 
     n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , 
     n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , 
     n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , 
     n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , 
     n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , 
     n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , 
     n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , 
     n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , 
     n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , 
     n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , 
     n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , 
     n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , 
     n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , 
     n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , 
     n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , 
     n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , 
     n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , 
     n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , 
     n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , 
     n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , 
     n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , 
     n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , 
     n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , 
     n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , 
     n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , 
     n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , 
     n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , 
     n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , 
     n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , 
     n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , 
     n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , 
     n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , 
     n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , 
     n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , 
     n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , 
     n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , 
     n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , 
     n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , 
     n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , 
     n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , 
     n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , 
     n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , 
     n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , 
     n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , 
     n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , 
     n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , 
     n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , 
     n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , 
     n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , 
     n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , 
     n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , 
     n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , 
     n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , 
     n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , 
     n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , 
     n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , 
     n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , 
     n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , 
     n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , 
     n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , 
     n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , 
     n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , 
     n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , 
     n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , 
     n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , 
     n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , 
     n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , 
     n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , 
     n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , 
     n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , 
     n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , 
     n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , 
     n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , 
     n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , 
     n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , 
     n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , 
     n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , 
     n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , 
     n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , 
     n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , 
     n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , 
     n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , 
     n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , 
     n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , 
     n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , 
     n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , 
     n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , 
     n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , 
     n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , 
     n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , 
     n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , 
     n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , 
     n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , 
     n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , 
     n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , 
     n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , 
     n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , 
     n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , 
     n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , 
     n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , 
     n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , 
     n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , 
     n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , 
     n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , 
     n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , 
     n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , 
     n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , 
     n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , 
     n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , 
     n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , 
     n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , 
     n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , 
     n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , 
     n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , 
     n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , 
     n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , 
     n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , 
     n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , 
     n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , 
     n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , 
     n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , 
     n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , 
     n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , 
     n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , 
     n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , 
     n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , 
     n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , 
     n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , 
     n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , 
     n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , 
     n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , 
     n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , 
     n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , 
     n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , 
     n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , 
     n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , 
     n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , 
     n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , 
     n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , 
     n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , 
     n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , 
     n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , 
     n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , 
     n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , 
     n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , 
     n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , 
     n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , 
     n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , 
     n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , 
     n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , 
     n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , 
     n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , 
     n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , 
     n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , 
     n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , 
     n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , 
     n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , 
     n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , 
     n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , 
     n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , 
     n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , 
     n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , 
     n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , 
     n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , 
     n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , 
     n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , 
     n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , 
     n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , 
     n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , 
     n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , 
     n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , 
     n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , 
     n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , 
     n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , 
     n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , 
     n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , 
     n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , 
     n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , 
     n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , 
     n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , 
     n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , 
     n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , 
     n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , 
     n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , 
     n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , 
     n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , 
     n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , 
     n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , 
     n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , 
     n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , 
     n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , 
     n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , 
     n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , 
     n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , 
     n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , 
     n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , 
     n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , 
     n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , 
     n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , 
     n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , 
     n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , 
     n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , 
     n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , 
     n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , 
     n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , 
     n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , 
     n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , 
     n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , 
     n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , 
     n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , 
     n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , 
     n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , 
     n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , 
     n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , 
     n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , 
     n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , 
     n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , 
     n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , 
     n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , 
     n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , 
     n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , 
     n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , 
     n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , 
     n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , 
     n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , 
     n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , 
     n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , 
     n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , 
     n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , 
     n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , 
     n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , 
     n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , 
     n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , 
     n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , 
     n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , 
     n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , 
     n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , 
     n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , 
     n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , 
     n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , 
     n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , 
     n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , 
     n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , 
     n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , 
     n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , 
     n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , 
     n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , 
     n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , 
     n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , 
     n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , 
     n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , 
     n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , 
     n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , 
     n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , 
     n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , 
     n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , 
     n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , 
     n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , 
     n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , 
     n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , 
     n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , 
     n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , 
     n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , 
     n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , 
     n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , 
     n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , 
     n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , 
     n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , 
     n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , 
     n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , 
     n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , 
     n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , 
     n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , 
     n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , 
     n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , 
     n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , 
     n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , 
     n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , 
     n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , 
     n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , 
     n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , 
     n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , 
     n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , 
     n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , 
     n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , 
     n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , 
     n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , 
     n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , 
     n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , 
     n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , 
     n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , 
     n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , 
     n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , 
     n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , 
     n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , 
     n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , 
     n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , 
     n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , 
     n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , 
     n24080 , n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , 
     n24090 , n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , 
     n24100 , n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , 
     n24110 , n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , 
     n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , 
     n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , 
     n24140 , n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , 
     n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , 
     n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , 
     n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , 
     n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , 
     n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , 
     n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , 
     n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , 
     n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , 
     n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , 
     n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , 
     n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , 
     n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , 
     n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , 
     n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , 
     n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , 
     n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , 
     n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , 
     n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , 
     n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , 
     n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , 
     n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , 
     n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , 
     n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , 
     n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , 
     n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , 
     n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , 
     n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , 
     n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , 
     n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , 
     n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , n24449 , 
     n24450 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , 
     n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , 
     n24470 , n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , n24479 , 
     n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , 
     n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , 
     n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , 
     n24510 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , 
     n24520 , n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , 
     n24530 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , 
     n24540 , n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , 
     n24550 , n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , 
     n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , 
     n24570 , n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , 
     n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , 
     n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , 
     n24600 , n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , 
     n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , 
     n24620 , n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , n24629 , 
     n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , n24639 , 
     n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , 
     n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , 
     n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , 
     n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , 
     n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , 
     n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , 
     n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , 
     n24710 , n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , 
     n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , 
     n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , 
     n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , 
     n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , 
     n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , n24767 , n24768 , n24769 , 
     n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , 
     n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , 
     n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , 
     n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , 
     n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , 
     n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , n24829 , 
     n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , 
     n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , 
     n24850 , n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , 
     n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , 
     n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , 
     n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , 
     n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , 
     n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , 
     n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , 
     n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , 
     n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , 
     n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , 
     n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , 
     n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , 
     n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , 
     n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , 
     n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , n24999 , 
     n25000 , n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , n25009 , 
     n25010 , n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , 
     n25020 , n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , n25029 , 
     n25030 , n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , n25039 , 
     n25040 , n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , n25049 , 
     n25050 , n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , n25059 , 
     n25060 , n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , n25069 , 
     n25070 , n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , n25079 , 
     n25080 , n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , n25089 , 
     n25090 , n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , n25099 , 
     n25100 , n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , n25109 , 
     n25110 , n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , n25119 , 
     n25120 , n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , n25127 , n25128 , n25129 , 
     n25130 , n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , n25139 , 
     n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , n25149 , 
     n25150 , n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , n25159 , 
     n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , n25169 , 
     n25170 , n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , n25179 , 
     n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , n25189 , 
     n25190 , n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , n25199 , 
     n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , n25209 , 
     n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , n25219 , 
     n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , n25229 , 
     n25230 , n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , n25239 , 
     n25240 , n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , n25249 , 
     n25250 , n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , n25259 , 
     n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , 
     n25270 , n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , n25279 , 
     n25280 , n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , n25289 , 
     n25290 , n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , n25299 , 
     n25300 , n25301 , n25302 , n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , n25309 , 
     n25310 , n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , n25319 , 
     n25320 , n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , n25329 , 
     n25330 , n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , n25337 , n25338 , n25339 , 
     n25340 , n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , n25347 , n25348 , n25349 , 
     n25350 , n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , n25357 , n25358 , n25359 , 
     n25360 , n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , n25369 , 
     n25370 , n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , n25379 , 
     n25380 , n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , n25389 , 
     n25390 , n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , n25399 , 
     n25400 , n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , n25409 , 
     n25410 , n25411 , n25412 , n25413 , n25414 , n25415 , n25416 , n25417 , n25418 , n25419 , 
     n25420 , n25421 , n25422 , n25423 , n25424 , n25425 , n25426 , n25427 , n25428 , n25429 , 
     n25430 , n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , n25439 , 
     n25440 , n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , n25449 , 
     n25450 , n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , n25459 , 
     n25460 , n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , n25469 , 
     n25470 , n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , n25479 , 
     n25480 , n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , n25489 , 
     n25490 , n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , n25499 , 
     n25500 , n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , n25509 , 
     n25510 , n25511 , n25512 , n25513 , n25514 , n25515 , n25516 , n25517 , n25518 , n25519 , 
     n25520 , n25521 , n25522 , n25523 , n25524 , n25525 , n25526 , n25527 , n25528 , n25529 , 
     n25530 , n25531 , n25532 , n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , n25539 , 
     n25540 , n25541 , n25542 , n25543 , n25544 , n25545 , n25546 , n25547 , n25548 , n25549 , 
     n25550 , n25551 , n25552 , n25553 , n25554 , n25555 , n25556 , n25557 , n25558 , n25559 , 
     n25560 , n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , n25567 , n25568 , n25569 , 
     n25570 , n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , n25577 , n25578 , n25579 , 
     n25580 , n25581 , n25582 , n25583 , n25584 , n25585 , n25586 , n25587 , n25588 , n25589 , 
     n25590 , n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , n25597 , n25598 , n25599 , 
     n25600 , n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , n25607 , n25608 , n25609 , 
     n25610 , n25611 , n25612 , n25613 , n25614 , n25615 , n25616 , n25617 , n25618 , n25619 , 
     n25620 , n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , n25627 , n25628 , n25629 , 
     n25630 , n25631 , n25632 , n25633 , n25634 , n25635 , n25636 , n25637 , n25638 , n25639 , 
     n25640 , n25641 , n25642 , n25643 , n25644 , n25645 , n25646 , n25647 , n25648 , n25649 , 
     n25650 , n25651 , n25652 , n25653 , n25654 , n25655 , n25656 , n25657 , n25658 , n25659 , 
     n25660 , n25661 , n25662 , n25663 , n25664 , n25665 , n25666 , n25667 , n25668 , n25669 , 
     n25670 , n25671 , n25672 , n25673 , n25674 , n25675 , n25676 , n25677 , n25678 , n25679 , 
     n25680 , n25681 , n25682 , n25683 , n25684 , n25685 , n25686 , n25687 , n25688 , n25689 , 
     n25690 , n25691 , n25692 , n25693 , n25694 , n25695 , n25696 , n25697 , n25698 , n25699 , 
     n25700 , n25701 , n25702 , n25703 , n25704 , n25705 , n25706 , n25707 , n25708 , n25709 , 
     n25710 , n25711 , n25712 , n25713 , n25714 , n25715 , n25716 , n25717 , n25718 , n25719 , 
     n25720 , n25721 , n25722 , n25723 , n25724 , n25725 , n25726 , n25727 , n25728 , n25729 , 
     n25730 , n25731 , n25732 , n25733 , n25734 , n25735 , n25736 , n25737 , n25738 , n25739 , 
     n25740 , n25741 , n25742 , n25743 , n25744 , n25745 , n25746 , n25747 , n25748 , n25749 , 
     n25750 , n25751 , n25752 , n25753 , n25754 , n25755 , n25756 , n25757 , n25758 , n25759 , 
     n25760 , n25761 , n25762 , n25763 , n25764 , n25765 , n25766 , n25767 , n25768 , n25769 , 
     n25770 , n25771 , n25772 , n25773 , n25774 , n25775 , n25776 , n25777 , n25778 , n25779 , 
     n25780 , n25781 , n25782 , n25783 , n25784 , n25785 , n25786 , n25787 , n25788 , n25789 , 
     n25790 , n25791 , n25792 , n25793 , n25794 , n25795 , n25796 , n25797 , n25798 , n25799 , 
     n25800 , n25801 , n25802 , n25803 , n25804 , n25805 , n25806 , n25807 , n25808 , n25809 , 
     n25810 , n25811 , n25812 , n25813 , n25814 , n25815 , n25816 , n25817 , n25818 , n25819 , 
     n25820 , n25821 , n25822 , n25823 , n25824 , n25825 , n25826 , n25827 , n25828 , n25829 , 
     n25830 , n25831 , n25832 , n25833 , n25834 , n25835 , n25836 , n25837 , n25838 , n25839 , 
     n25840 , n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , n25847 , n25848 , n25849 , 
     n25850 , n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , n25857 , n25858 , n25859 , 
     n25860 , n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , n25867 , n25868 , n25869 , 
     n25870 , n25871 , n25872 , n25873 , n25874 , n25875 , n25876 , n25877 , n25878 , n25879 , 
     n25880 , n25881 , n25882 , n25883 , n25884 , n25885 , n25886 , n25887 , n25888 , n25889 , 
     n25890 , n25891 , n25892 , n25893 , n25894 , n25895 , n25896 , n25897 , n25898 , n25899 , 
     n25900 , n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , n25907 , n25908 , n25909 , 
     n25910 , n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , n25917 , n25918 , n25919 , 
     n25920 , n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , n25927 , n25928 , n25929 , 
     n25930 , n25931 , n25932 , n25933 , n25934 , n25935 , n25936 , n25937 , n25938 , n25939 , 
     n25940 , n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , n25947 , n25948 , n25949 , 
     n25950 , n25951 , n25952 , n25953 , n25954 , n25955 , n25956 , n25957 , n25958 , n25959 , 
     n25960 , n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , n25967 , n25968 , n25969 , 
     n25970 , n25971 , n25972 , n25973 , n25974 , n25975 , n25976 , n25977 , n25978 , n25979 , 
     n25980 , n25981 , n25982 , n25983 , n25984 , n25985 , n25986 , n25987 , n25988 , n25989 , 
     n25990 , n25991 , n25992 , n25993 , n25994 , n25995 , n25996 , n25997 , n25998 , n25999 , 
     n26000 , n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , n26007 , n26008 , n26009 , 
     n26010 , n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , n26017 , n26018 , n26019 , 
     n26020 , n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , n26027 , n26028 , n26029 , 
     n26030 , n26031 , n26032 , n26033 , n26034 , n26035 , n26036 , n26037 , n26038 , n26039 , 
     n26040 , n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , n26047 , n26048 , n26049 , 
     n26050 , n26051 , n26052 , n26053 , n26054 , n26055 , n26056 , n26057 , n26058 , n26059 , 
     n26060 , n26061 , n26062 , n26063 , n26064 , n26065 , n26066 , n26067 , n26068 , n26069 , 
     n26070 , n26071 , n26072 , n26073 , n26074 , n26075 , n26076 , n26077 , n26078 , n26079 , 
     n26080 , n26081 , n26082 , n26083 , n26084 , n26085 , n26086 , n26087 , n26088 , n26089 , 
     n26090 , n26091 , n26092 , n26093 , n26094 , n26095 , n26096 , n26097 , n26098 , n26099 , 
     n26100 , n26101 , n26102 , n26103 , n26104 , n26105 , n26106 , n26107 , n26108 , n26109 , 
     n26110 , n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , n26117 , n26118 , n26119 , 
     n26120 , n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , n26127 , n26128 , n26129 , 
     n26130 , n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , n26137 , n26138 , n26139 , 
     n26140 , n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , n26147 , n26148 , n26149 , 
     n26150 , n26151 , n26152 , n26153 , n26154 , n26155 , n26156 , n26157 , n26158 , n26159 , 
     n26160 , n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , n26167 , n26168 , n26169 , 
     n26170 , n26171 , n26172 , n26173 , n26174 , n26175 , n26176 , n26177 , n26178 , n26179 , 
     n26180 , n26181 , n26182 , n26183 , n26184 , n26185 , n26186 , n26187 , n26188 , n26189 , 
     n26190 , n26191 , n26192 , n26193 , n26194 , n26195 , n26196 , n26197 , n26198 , n26199 , 
     n26200 , n26201 , n26202 , n26203 , n26204 , n26205 , n26206 , n26207 , n26208 , n26209 , 
     n26210 , n26211 , n26212 , n26213 , n26214 , n26215 , n26216 , n26217 , n26218 , n26219 , 
     n26220 , n26221 , n26222 , n26223 , n26224 , n26225 , n26226 , n26227 , n26228 , n26229 , 
     n26230 , n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , n26237 , n26238 , n26239 , 
     n26240 , n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , n26247 , n26248 , n26249 , 
     n26250 , n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , n26257 , n26258 , n26259 , 
     n26260 , n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , n26267 , n26268 , n26269 , 
     n26270 , n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , n26277 , n26278 , n26279 , 
     n26280 , n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , n26287 , n26288 , n26289 , 
     n26290 , n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , n26297 , n26298 , n26299 , 
     n26300 , n26301 , n26302 , n26303 , n26304 , n26305 , n26306 , n26307 , n26308 , n26309 , 
     n26310 , n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , n26317 , n26318 , n26319 , 
     n26320 , n26321 , n26322 , n26323 , n26324 , n26325 , n26326 , n26327 , n26328 , n26329 , 
     n26330 , n26331 , n26332 , n26333 , n26334 , n26335 , n26336 , n26337 , n26338 , n26339 , 
     n26340 , n26341 , n26342 , n26343 , n26344 , n26345 , n26346 , n26347 , n26348 , n26349 , 
     n26350 , n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , n26357 , n26358 , n26359 , 
     n26360 , n26361 , n26362 , n26363 , n26364 , n26365 , n26366 , n26367 , n26368 , n26369 , 
     n26370 , n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , n26377 , n26378 , n26379 , 
     n26380 , n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , n26387 , n26388 , n26389 , 
     n26390 , n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , n26397 , n26398 , n26399 , 
     n26400 , n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , n26407 , n26408 , n26409 , 
     n26410 , n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , n26417 , n26418 , n26419 , 
     n26420 , n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , n26427 , n26428 , n26429 , 
     n26430 , n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , n26437 , n26438 , n26439 , 
     n26440 , n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , n26447 , n26448 , n26449 , 
     n26450 , n26451 , n26452 , n26453 , n26454 , n26455 , n26456 , n26457 , n26458 , n26459 , 
     n26460 , n26461 , n26462 , n26463 , n26464 , n26465 , n26466 , n26467 , n26468 , n26469 , 
     n26470 , n26471 , n26472 , n26473 , n26474 , n26475 , n26476 , n26477 , n26478 , n26479 , 
     n26480 , n26481 , n26482 , n26483 , n26484 , n26485 , n26486 , n26487 , n26488 , n26489 , 
     n26490 , n26491 , n26492 , n26493 , n26494 , n26495 , n26496 , n26497 , n26498 , n26499 , 
     n26500 , n26501 , n26502 , n26503 , n26504 , n26505 , n26506 , n26507 , n26508 , n26509 , 
     n26510 , n26511 , n26512 , n26513 , n26514 , n26515 , n26516 , n26517 , n26518 , n26519 , 
     n26520 , n26521 , n26522 , n26523 , n26524 , n26525 , n26526 , n26527 , n26528 , n26529 , 
     n26530 , n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , n26537 , n26538 , n26539 , 
     n26540 , n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , n26547 , n26548 , n26549 , 
     n26550 , n26551 , n26552 , n26553 , n26554 , n26555 , n26556 , n26557 , n26558 , n26559 , 
     n26560 , n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , n26567 , n26568 , n26569 , 
     n26570 , n26571 , n26572 , n26573 , n26574 , n26575 , n26576 , n26577 , n26578 , n26579 , 
     n26580 , n26581 , n26582 , n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , n26589 , 
     n26590 , n26591 , n26592 , n26593 , n26594 , n26595 , n26596 , n26597 , n26598 , n26599 , 
     n26600 , n26601 , n26602 , n26603 , n26604 , n26605 , n26606 , n26607 , n26608 , n26609 , 
     n26610 , n26611 , n26612 , n26613 , n26614 , n26615 , n26616 , n26617 , n26618 , n26619 , 
     n26620 , n26621 , n26622 , n26623 , n26624 , n26625 , n26626 , n26627 , n26628 , n26629 , 
     n26630 , n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , n26637 , n26638 , n26639 , 
     n26640 , n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , n26647 , n26648 , n26649 , 
     n26650 , n26651 , n26652 , n26653 , n26654 , n26655 , n26656 , n26657 , n26658 , n26659 , 
     n26660 , n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , n26667 , n26668 , n26669 , 
     n26670 , n26671 , n26672 , n26673 , n26674 , n26675 , n26676 , n26677 , n26678 , n26679 , 
     n26680 , n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , n26687 , n26688 , n26689 , 
     n26690 , n26691 , n26692 , n26693 , n26694 , n26695 , n26696 , n26697 , n26698 , n26699 , 
     n26700 , n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , n26707 , n26708 , n26709 , 
     n26710 , n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , n26717 , n26718 , n26719 , 
     n26720 , n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , n26727 , n26728 , n26729 , 
     n26730 , n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , n26737 , n26738 , n26739 , 
     n26740 , n26741 , n26742 , n26743 , n26744 , n26745 , n26746 , n26747 , n26748 , n26749 , 
     n26750 , n26751 , n26752 , n26753 , n26754 , n26755 , n26756 , n26757 , n26758 , n26759 , 
     n26760 , n26761 , n26762 , n26763 , n26764 , n26765 , n26766 , n26767 , n26768 , n26769 , 
     n26770 , n26771 , n26772 , n26773 , n26774 , n26775 , n26776 , n26777 , n26778 , n26779 , 
     n26780 , n26781 , n26782 , n26783 , n26784 , n26785 , n26786 , n26787 , n26788 , n26789 , 
     n26790 , n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , n26797 , n26798 , n26799 , 
     n26800 , n26801 , n26802 , n26803 , n26804 , n26805 , n26806 , n26807 , n26808 , n26809 , 
     n26810 , n26811 , n26812 , n26813 , n26814 , n26815 , n26816 , n26817 , n26818 , n26819 , 
     n26820 , n26821 , n26822 , n26823 , n26824 , n26825 , n26826 , n26827 , n26828 , n26829 , 
     n26830 , n26831 , n26832 , n26833 , n26834 , n26835 , n26836 , n26837 , n26838 , n26839 , 
     n26840 , n26841 , n26842 , n26843 , n26844 , n26845 , n26846 , n26847 , n26848 , n26849 , 
     n26850 , n26851 , n26852 , n26853 , n26854 , n26855 , n26856 , n26857 , n26858 , n26859 , 
     n26860 , n26861 , n26862 , n26863 , n26864 , n26865 , n26866 , n26867 , n26868 , n26869 , 
     n26870 , n26871 , n26872 , n26873 , n26874 , n26875 , n26876 , n26877 , n26878 , n26879 , 
     n26880 , n26881 , n26882 , n26883 , n26884 , n26885 , n26886 , n26887 , n26888 , n26889 , 
     n26890 , n26891 , n26892 , n26893 , n26894 , n26895 , n26896 , n26897 , n26898 , n26899 , 
     n26900 , n26901 , n26902 , n26903 , n26904 , n26905 , n26906 , n26907 , n26908 , n26909 , 
     n26910 , n26911 , n26912 , n26913 , n26914 , n26915 , n26916 , n26917 , n26918 , n26919 , 
     n26920 , n26921 , n26922 , n26923 , n26924 , n26925 , n26926 , n26927 , n26928 , n26929 , 
     n26930 , n26931 , n26932 , n26933 , n26934 , n26935 , n26936 , n26937 , n26938 , n26939 , 
     n26940 , n26941 , n26942 , n26943 , n26944 , n26945 , n26946 , n26947 , n26948 , n26949 , 
     n26950 , n26951 , n26952 , n26953 , n26954 , n26955 , n26956 , n26957 , n26958 , n26959 , 
     n26960 , n26961 , n26962 , n26963 , n26964 , n26965 , n26966 , n26967 , n26968 , n26969 , 
     n26970 , n26971 , n26972 , n26973 , n26974 , n26975 , n26976 , n26977 , n26978 , n26979 , 
     n26980 , n26981 , n26982 , n26983 , n26984 , n26985 , n26986 , n26987 , n26988 , n26989 , 
     n26990 , n26991 , n26992 , n26993 , n26994 , n26995 , n26996 , n26997 , n26998 , n26999 , 
     n27000 , n27001 , n27002 , n27003 , n27004 , n27005 , n27006 , n27007 , n27008 , n27009 , 
     n27010 , n27011 , n27012 , n27013 , n27014 , n27015 , n27016 , n27017 , n27018 , n27019 , 
     n27020 , n27021 , n27022 , n27023 , n27024 , n27025 , n27026 , n27027 , n27028 , n27029 , 
     n27030 , n27031 , n27032 , n27033 , n27034 , n27035 , n27036 , n27037 , n27038 , n27039 , 
     n27040 , n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , n27047 , n27048 , n27049 , 
     n27050 , n27051 , n27052 , n27053 , n27054 , n27055 , n27056 , n27057 , n27058 , n27059 , 
     n27060 , n27061 , n27062 , n27063 , n27064 , n27065 , n27066 , n27067 , n27068 , n27069 , 
     n27070 , n27071 , n27072 , n27073 , n27074 , n27075 , n27076 , n27077 , n27078 , n27079 , 
     n27080 , n27081 , n27082 , n27083 , n27084 , n27085 , n27086 , n27087 , n27088 , n27089 , 
     n27090 , n27091 , n27092 , n27093 , n27094 , n27095 , n27096 , n27097 , n27098 , n27099 , 
     n27100 , n27101 , n27102 , n27103 , n27104 , n27105 , n27106 , n27107 , n27108 , n27109 , 
     n27110 , n27111 , n27112 , n27113 , n27114 , n27115 , n27116 , n27117 , n27118 , n27119 , 
     n27120 , n27121 , n27122 , n27123 , n27124 , n27125 , n27126 , n27127 , n27128 , n27129 , 
     n27130 , n27131 , n27132 , n27133 , n27134 , n27135 , n27136 , n27137 , n27138 , n27139 , 
     n27140 , n27141 , n27142 , n27143 , n27144 , n27145 , n27146 , n27147 , n27148 , n27149 , 
     n27150 , n27151 , n27152 , n27153 , n27154 , n27155 , n27156 , n27157 , n27158 , n27159 , 
     n27160 , n27161 , n27162 , n27163 , n27164 , n27165 , n27166 , n27167 , n27168 , n27169 , 
     n27170 , n27171 , n27172 , n27173 , n27174 , n27175 , n27176 , n27177 , n27178 , n27179 , 
     n27180 , n27181 , n27182 , n27183 , n27184 , n27185 , n27186 , n27187 , n27188 , n27189 , 
     n27190 , n27191 , n27192 , n27193 , n27194 , n27195 , n27196 , n27197 , n27198 , n27199 , 
     n27200 , n27201 , n27202 , n27203 , n27204 , n27205 , n27206 , n27207 , n27208 , n27209 , 
     n27210 , n27211 , n27212 , n27213 , n27214 , n27215 , n27216 , n27217 , n27218 , n27219 , 
     n27220 , n27221 , n27222 , n27223 , n27224 , n27225 , n27226 , n27227 , n27228 , n27229 , 
     n27230 , n27231 , n27232 , n27233 , n27234 , n27235 , n27236 , n27237 , n27238 , n27239 , 
     n27240 , n27241 , n27242 , n27243 , n27244 , n27245 , n27246 , n27247 , n27248 , n27249 , 
     n27250 , n27251 , n27252 , n27253 , n27254 , n27255 , n27256 , n27257 , n27258 , n27259 , 
     n27260 , n27261 , n27262 , n27263 , n27264 , n27265 , n27266 , n27267 , n27268 , n27269 , 
     n27270 , n27271 , n27272 , n27273 , n27274 , n27275 , n27276 , n27277 , n27278 , n27279 , 
     n27280 , n27281 , n27282 , n27283 , n27284 , n27285 , n27286 , n27287 , n27288 , n27289 , 
     n27290 , n27291 , n27292 , n27293 , n27294 , n27295 , n27296 , n27297 , n27298 , n27299 , 
     n27300 , n27301 , n27302 , n27303 , n27304 , n27305 , n27306 , n27307 , n27308 , n27309 , 
     n27310 , n27311 , n27312 , n27313 , n27314 , n27315 , n27316 , n27317 , n27318 , n27319 , 
     n27320 , n27321 , n27322 , n27323 , n27324 , n27325 , n27326 , n27327 , n27328 , n27329 , 
     n27330 , n27331 , n27332 , n27333 , n27334 , n27335 , n27336 , n27337 , n27338 , n27339 , 
     n27340 , n27341 , n27342 , n27343 , n27344 , n27345 , n27346 , n27347 , n27348 , n27349 , 
     n27350 , n27351 , n27352 , n27353 , n27354 , n27355 , n27356 , n27357 , n27358 , n27359 , 
     n27360 , n27361 , n27362 , n27363 , n27364 , n27365 , n27366 , n27367 , n27368 , n27369 , 
     n27370 , n27371 , n27372 , n27373 , n27374 , n27375 , n27376 , n27377 , n27378 , n27379 , 
     n27380 , n27381 , n27382 , n27383 , n27384 , n27385 , n27386 , n27387 , n27388 , n27389 , 
     n27390 , n27391 , n27392 , n27393 , n27394 , n27395 , n27396 , n27397 , n27398 , n27399 , 
     n27400 , n27401 , n27402 , n27403 , n27404 , n27405 , n27406 , n27407 , n27408 , n27409 , 
     n27410 , n27411 , n27412 , n27413 , n27414 , n27415 , n27416 , n27417 , n27418 , n27419 , 
     n27420 , n27421 , n27422 , n27423 , n27424 , n27425 , n27426 , n27427 , n27428 , n27429 , 
     n27430 , n27431 , n27432 , n27433 , n27434 , n27435 , n27436 , n27437 , n27438 , n27439 , 
     n27440 , n27441 , n27442 , n27443 , n27444 , n27445 , n27446 , n27447 , n27448 , n27449 , 
     n27450 , n27451 , n27452 , n27453 , n27454 , n27455 , n27456 , n27457 , n27458 , n27459 , 
     n27460 , n27461 , n27462 , n27463 , n27464 , n27465 , n27466 , n27467 , n27468 , n27469 , 
     n27470 , n27471 , n27472 , n27473 , n27474 , n27475 , n27476 , n27477 , n27478 , n27479 , 
     n27480 , n27481 , n27482 , n27483 , n27484 , n27485 , n27486 , n27487 , n27488 , n27489 , 
     n27490 , n27491 , n27492 , n27493 , n27494 , n27495 , n27496 , n27497 , n27498 , n27499 , 
     n27500 , n27501 , n27502 , n27503 , n27504 , n27505 , n27506 , n27507 , n27508 , n27509 , 
     n27510 , n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , n27517 , n27518 , n27519 , 
     n27520 , n27521 , n27522 , n27523 , n27524 , n27525 , n27526 , n27527 , n27528 , n27529 , 
     n27530 , n27531 , n27532 , n27533 , n27534 , n27535 , n27536 , n27537 , n27538 , n27539 , 
     n27540 , n27541 , n27542 , n27543 , n27544 , n27545 , n27546 , n27547 , n27548 , n27549 , 
     n27550 , n27551 , n27552 , n27553 , n27554 , n27555 , n27556 , n27557 , n27558 , n27559 , 
     n27560 , n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , n27567 , n27568 , n27569 , 
     n27570 , n27571 , n27572 , n27573 , n27574 , n27575 , n27576 , n27577 , n27578 , n27579 , 
     n27580 , n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , n27587 , n27588 , n27589 , 
     n27590 , n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , n27597 , n27598 , n27599 , 
     n27600 , n27601 , n27602 , n27603 , n27604 , n27605 , n27606 , n27607 , n27608 , n27609 , 
     n27610 , n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , n27617 , n27618 , n27619 , 
     n27620 , n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , n27627 , n27628 , n27629 , 
     n27630 , n27631 , n27632 , n27633 , n27634 , n27635 , n27636 , n27637 , n27638 , n27639 , 
     n27640 , n27641 , n27642 , n27643 , n27644 , n27645 , n27646 , n27647 , n27648 , n27649 , 
     n27650 , n27651 , n27652 , n27653 , n27654 , n27655 , n27656 , n27657 , n27658 , n27659 , 
     n27660 , n27661 , n27662 , n27663 , n27664 , n27665 , n27666 , n27667 , n27668 , n27669 , 
     n27670 , n27671 , n27672 , n27673 , n27674 , n27675 , n27676 , n27677 , n27678 , n27679 , 
     n27680 , n27681 , n27682 , n27683 , n27684 , n27685 , n27686 , n27687 , n27688 , n27689 , 
     n27690 , n27691 , n27692 , n27693 , n27694 , n27695 , n27696 , n27697 , n27698 , n27699 , 
     n27700 , n27701 , n27702 , n27703 , n27704 , n27705 , n27706 , n27707 , n27708 , n27709 , 
     n27710 , n27711 , n27712 , n27713 , n27714 , n27715 , n27716 , n27717 , n27718 , n27719 , 
     n27720 , n27721 , n27722 , n27723 , n27724 , n27725 , n27726 , n27727 , n27728 , n27729 , 
     n27730 , n27731 , n27732 , n27733 , n27734 , n27735 , n27736 , n27737 , n27738 , n27739 , 
     n27740 , n27741 , n27742 , n27743 , n27744 , n27745 , n27746 , n27747 , n27748 , n27749 , 
     n27750 , n27751 , n27752 , n27753 , n27754 , n27755 , n27756 , n27757 , n27758 , n27759 , 
     n27760 , n27761 , n27762 , n27763 , n27764 , n27765 , n27766 , n27767 , n27768 , n27769 , 
     n27770 , n27771 , n27772 , n27773 , n27774 , n27775 , n27776 , n27777 , n27778 , n27779 , 
     n27780 , n27781 , n27782 , n27783 , n27784 , n27785 , n27786 , n27787 , n27788 , n27789 , 
     n27790 , n27791 , n27792 , n27793 , n27794 , n27795 , n27796 , n27797 , n27798 , n27799 , 
     n27800 , n27801 , n27802 , n27803 , n27804 , n27805 , n27806 , n27807 , n27808 , n27809 , 
     n27810 , n27811 , n27812 , n27813 , n27814 , n27815 , n27816 , n27817 , n27818 , n27819 , 
     n27820 , n27821 , n27822 , n27823 , n27824 , n27825 , n27826 , n27827 , n27828 , n27829 , 
     n27830 , n27831 , n27832 , n27833 , n27834 , n27835 , n27836 , n27837 , n27838 , n27839 , 
     n27840 , n27841 , n27842 , n27843 , n27844 , n27845 , n27846 , n27847 , n27848 , n27849 , 
     n27850 , n27851 , n27852 , n27853 , n27854 , n27855 , n27856 , n27857 , n27858 , n27859 , 
     n27860 , n27861 , n27862 , n27863 , n27864 , n27865 , n27866 , n27867 , n27868 , n27869 , 
     n27870 , n27871 , n27872 , n27873 , n27874 , n27875 , n27876 , n27877 , n27878 , n27879 , 
     n27880 , n27881 , n27882 , n27883 , n27884 , n27885 , n27886 , n27887 , n27888 , n27889 , 
     n27890 , n27891 , n27892 , n27893 , n27894 , n27895 , n27896 , n27897 , n27898 , n27899 , 
     n27900 , n27901 , n27902 , n27903 , n27904 , n27905 , n27906 , n27907 , n27908 , n27909 , 
     n27910 , n27911 , n27912 , n27913 , n27914 , n27915 , n27916 , n27917 , n27918 , n27919 , 
     n27920 , n27921 , n27922 , n27923 , n27924 , n27925 , n27926 , n27927 , n27928 , n27929 , 
     n27930 , n27931 , n27932 , n27933 , n27934 , n27935 , n27936 , n27937 , n27938 , n27939 , 
     n27940 , n27941 , n27942 , n27943 , n27944 , n27945 , n27946 , n27947 , n27948 , n27949 , 
     n27950 , n27951 , n27952 , n27953 , n27954 , n27955 , n27956 , n27957 , n27958 , n27959 , 
     n27960 , n27961 , n27962 , n27963 , n27964 , n27965 , n27966 , n27967 , n27968 , n27969 , 
     n27970 , n27971 , n27972 , n27973 , n27974 , n27975 , n27976 , n27977 , n27978 , n27979 , 
     n27980 , n27981 , n27982 , n27983 , n27984 , n27985 , n27986 , n27987 , n27988 , n27989 , 
     n27990 , n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , n27997 , n27998 , n27999 , 
     n28000 , n28001 , n28002 , n28003 , n28004 , n28005 , n28006 , n28007 , n28008 , n28009 , 
     n28010 , n28011 , n28012 , n28013 , n28014 , n28015 , n28016 , n28017 , n28018 , n28019 , 
     n28020 , n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , n28027 , n28028 , n28029 , 
     n28030 , n28031 , n28032 , n28033 , n28034 , n28035 , n28036 , n28037 , n28038 , n28039 , 
     n28040 , n28041 , n28042 , n28043 , n28044 , n28045 , n28046 , n28047 , n28048 , n28049 , 
     n28050 , n28051 , n28052 , n28053 , n28054 , n28055 , n28056 , n28057 , n28058 , n28059 , 
     n28060 , n28061 , n28062 , n28063 , n28064 , n28065 , n28066 , n28067 , n28068 , n28069 , 
     n28070 , n28071 , n28072 , n28073 , n28074 , n28075 , n28076 , n28077 , n28078 , n28079 , 
     n28080 , n28081 , n28082 , n28083 , n28084 , n28085 , n28086 , n28087 , n28088 , n28089 , 
     n28090 , n28091 , n28092 , n28093 , n28094 , n28095 , n28096 , n28097 , n28098 , n28099 , 
     n28100 , n28101 , n28102 , n28103 , n28104 , n28105 , n28106 , n28107 , n28108 , n28109 , 
     n28110 , n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , n28117 , n28118 , n28119 , 
     n28120 , n28121 , n28122 , n28123 , n28124 , n28125 , n28126 , n28127 , n28128 , n28129 , 
     n28130 , n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , n28137 , n28138 , n28139 , 
     n28140 , n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , n28147 , n28148 , n28149 , 
     n28150 , n28151 , n28152 , n28153 , n28154 , n28155 , n28156 , n28157 , n28158 , n28159 , 
     n28160 , n28161 , n28162 , n28163 , n28164 , n28165 , n28166 , n28167 , n28168 , n28169 , 
     n28170 , n28171 , n28172 , n28173 , n28174 , n28175 , n28176 , n28177 , n28178 , n28179 , 
     n28180 , n28181 , n28182 , n28183 , n28184 , n28185 , n28186 , n28187 , n28188 , n28189 , 
     n28190 , n28191 , n28192 , n28193 , n28194 , n28195 , n28196 , n28197 , n28198 , n28199 , 
     n28200 , n28201 , n28202 , n28203 , n28204 , n28205 , n28206 , n28207 , n28208 , n28209 , 
     n28210 , n28211 , n28212 , n28213 , n28214 , n28215 , n28216 , n28217 , n28218 , n28219 , 
     n28220 , n28221 , n28222 , n28223 , n28224 , n28225 , n28226 , n28227 , n28228 , n28229 , 
     n28230 , n28231 , n28232 , n28233 , n28234 , n28235 , n28236 , n28237 , n28238 , n28239 , 
     n28240 , n28241 , n28242 , n28243 , n28244 , n28245 , n28246 , n28247 , n28248 , n28249 , 
     n28250 , n28251 , n28252 , n28253 , n28254 , n28255 , n28256 , n28257 , n28258 , n28259 , 
     n28260 , n28261 , n28262 , n28263 , n28264 , n28265 , n28266 , n28267 , n28268 , n28269 , 
     n28270 , n28271 , n28272 , n28273 , n28274 , n28275 , n28276 , n28277 , n28278 , n28279 , 
     n28280 , n28281 , n28282 , n28283 , n28284 , n28285 , n28286 , n28287 , n28288 , n28289 , 
     n28290 , n28291 , n28292 , n28293 , n28294 , n28295 , n28296 , n28297 , n28298 , n28299 , 
     n28300 , n28301 , n28302 , n28303 , n28304 , n28305 , n28306 , n28307 , n28308 , n28309 , 
     n28310 , n28311 , n28312 , n28313 , n28314 , n28315 , n28316 , n28317 , n28318 , n28319 , 
     n28320 , n28321 , n28322 , n28323 , n28324 , n28325 , n28326 , n28327 , n28328 , n28329 , 
     n28330 , n28331 , n28332 , n28333 , n28334 , n28335 , n28336 , n28337 , n28338 , n28339 , 
     n28340 , n28341 , n28342 , n28343 , n28344 , n28345 , n28346 , n28347 , n28348 , n28349 , 
     n28350 , n28351 , n28352 , n28353 , n28354 , n28355 , n28356 , n28357 , n28358 , n28359 , 
     n28360 , n28361 , n28362 , n28363 , n28364 , n28365 , n28366 , n28367 , n28368 , n28369 , 
     n28370 , n28371 , n28372 , n28373 , n28374 , n28375 , n28376 , n28377 , n28378 , n28379 , 
     n28380 , n28381 , n28382 , n28383 , n28384 , n28385 , n28386 , n28387 , n28388 , n28389 , 
     n28390 , n28391 , n28392 , n28393 , n28394 , n28395 , n28396 , n28397 , n28398 , n28399 , 
     n28400 , n28401 , n28402 , n28403 , n28404 , n28405 , n28406 , n28407 , n28408 , n28409 , 
     n28410 , n28411 , n28412 , n28413 , n28414 , n28415 , n28416 , n28417 , n28418 , n28419 , 
     n28420 , n28421 , n28422 , n28423 , n28424 , n28425 , n28426 , n28427 , n28428 , n28429 , 
     n28430 , n28431 , n28432 , n28433 , n28434 , n28435 , n28436 , n28437 , n28438 , n28439 , 
     n28440 , n28441 , n28442 , n28443 , n28444 , n28445 , n28446 , n28447 , n28448 , n28449 , 
     n28450 , n28451 , n28452 , n28453 , n28454 , n28455 , n28456 , n28457 , n28458 , n28459 , 
     n28460 , n28461 , n28462 , n28463 , n28464 , n28465 , n28466 , n28467 , n28468 , n28469 , 
     n28470 , n28471 , n28472 , n28473 , n28474 , n28475 , n28476 , n28477 , n28478 , n28479 , 
     n28480 , n28481 , n28482 , n28483 , n28484 , n28485 , n28486 , n28487 , n28488 , n28489 , 
     n28490 , n28491 , n28492 , n28493 , n28494 , n28495 , n28496 , n28497 , n28498 , n28499 , 
     n28500 , n28501 , n28502 , n28503 , n28504 , n28505 , n28506 , n28507 , n28508 , n28509 , 
     n28510 , n28511 , n28512 , n28513 , n28514 , n28515 , n28516 , n28517 , n28518 , n28519 , 
     n28520 , n28521 , n28522 , n28523 , n28524 , n28525 , n28526 , n28527 , n28528 , n28529 , 
     n28530 , n28531 , n28532 , n28533 , n28534 , n28535 , n28536 , n28537 , n28538 , n28539 , 
     n28540 , n28541 , n28542 , n28543 , n28544 , n28545 , n28546 , n28547 , n28548 , n28549 , 
     n28550 , n28551 , n28552 , n28553 , n28554 , n28555 , n28556 , n28557 , n28558 , n28559 , 
     n28560 , n28561 , n28562 , n28563 , n28564 , n28565 , n28566 , n28567 , n28568 , n28569 , 
     n28570 , n28571 , n28572 , n28573 , n28574 , n28575 , n28576 , n28577 , n28578 , n28579 , 
     n28580 , n28581 , n28582 , n28583 , n28584 , n28585 , n28586 , n28587 , n28588 , n28589 , 
     n28590 , n28591 , n28592 , n28593 , n28594 , n28595 , n28596 , n28597 , n28598 , n28599 , 
     n28600 , n28601 , n28602 , n28603 , n28604 , n28605 , n28606 , n28607 , n28608 , n28609 , 
     n28610 , n28611 , n28612 , n28613 , n28614 , n28615 , n28616 , n28617 , n28618 , n28619 , 
     n28620 , n28621 , n28622 , n28623 , n28624 , n28625 , n28626 , n28627 , n28628 , n28629 , 
     n28630 , n28631 , n28632 , n28633 , n28634 , n28635 , n28636 , n28637 , n28638 , n28639 , 
     n28640 , n28641 , n28642 , n28643 , n28644 , n28645 , n28646 , n28647 , n28648 , n28649 , 
     n28650 , n28651 , n28652 , n28653 , n28654 , n28655 , n28656 , n28657 , n28658 , n28659 , 
     n28660 , n28661 , n28662 , n28663 , n28664 , n28665 , n28666 , n28667 , n28668 , n28669 , 
     n28670 , n28671 , n28672 , n28673 , n28674 , n28675 , n28676 , n28677 , n28678 , n28679 , 
     n28680 , n28681 , n28682 , n28683 , n28684 , n28685 , n28686 , n28687 , n28688 , n28689 , 
     n28690 , n28691 , n28692 , n28693 , n28694 , n28695 , n28696 , n28697 , n28698 , n28699 , 
     n28700 , n28701 , n28702 , n28703 , n28704 , n28705 , n28706 , n28707 , n28708 , n28709 , 
     n28710 , n28711 , n28712 , n28713 , n28714 , n28715 , n28716 , n28717 , n28718 , n28719 , 
     n28720 , n28721 , n28722 , n28723 , n28724 , n28725 , n28726 , n28727 , n28728 , n28729 , 
     n28730 , n28731 , n28732 , n28733 , n28734 , n28735 , n28736 , n28737 , n28738 , n28739 , 
     n28740 , n28741 , n28742 , n28743 , n28744 , n28745 , n28746 , n28747 , n28748 , n28749 , 
     n28750 , n28751 , n28752 , n28753 , n28754 , n28755 , n28756 , n28757 , n28758 , n28759 , 
     n28760 , n28761 , n28762 , n28763 , n28764 , n28765 , n28766 , n28767 , n28768 , n28769 , 
     n28770 , n28771 , n28772 , n28773 , n28774 , n28775 , n28776 , n28777 , n28778 , n28779 , 
     n28780 , n28781 , n28782 , n28783 , n28784 , n28785 , n28786 , n28787 , n28788 , n28789 , 
     n28790 , n28791 , n28792 , n28793 , n28794 , n28795 , n28796 , n28797 , n28798 , n28799 , 
     n28800 , n28801 , n28802 , n28803 , n28804 , n28805 , n28806 , n28807 , n28808 , n28809 , 
     n28810 , n28811 , n28812 , n28813 , n28814 , n28815 , n28816 , n28817 , n28818 , n28819 , 
     n28820 , n28821 , n28822 , n28823 , n28824 , n28825 , n28826 , n28827 , n28828 , n28829 , 
     n28830 , n28831 , n28832 , n28833 , n28834 , n28835 , n28836 , n28837 , n28838 , n28839 , 
     n28840 , n28841 , n28842 , n28843 , n28844 , n28845 , n28846 , n28847 , n28848 , n28849 , 
     n28850 , n28851 , n28852 , n28853 , n28854 , n28855 , n28856 , n28857 , n28858 , n28859 , 
     n28860 , n28861 , n28862 , n28863 , n28864 , n28865 , n28866 , n28867 , n28868 , n28869 , 
     n28870 , n28871 , n28872 , n28873 , n28874 , n28875 , n28876 , n28877 , n28878 , n28879 , 
     n28880 , n28881 , n28882 , n28883 , n28884 , n28885 , n28886 , n28887 , n28888 , n28889 , 
     n28890 , n28891 , n28892 , n28893 , n28894 , n28895 , n28896 , n28897 , n28898 , n28899 , 
     n28900 , n28901 , n28902 , n28903 , n28904 , n28905 , n28906 , n28907 , n28908 , n28909 , 
     n28910 , n28911 , n28912 , n28913 , n28914 , n28915 , n28916 , n28917 , n28918 , n28919 , 
     n28920 , n28921 , n28922 , n28923 , n28924 , n28925 , n28926 , n28927 , n28928 , n28929 , 
     n28930 , n28931 , n28932 , n28933 , n28934 , n28935 , n28936 , n28937 , n28938 , n28939 , 
     n28940 , n28941 , n28942 , n28943 , n28944 , n28945 , n28946 , n28947 , n28948 , n28949 , 
     n28950 , n28951 , n28952 , n28953 , n28954 , n28955 , n28956 , n28957 , n28958 , n28959 , 
     n28960 , n28961 , n28962 , n28963 , n28964 , n28965 , n28966 , n28967 , n28968 , n28969 , 
     n28970 , n28971 , n28972 , n28973 , n28974 , n28975 , n28976 , n28977 , n28978 , n28979 , 
     n28980 , n28981 , n28982 , n28983 , n28984 , n28985 , n28986 , n28987 , n28988 , n28989 , 
     n28990 , n28991 , n28992 , n28993 , n28994 , n28995 , n28996 , n28997 , n28998 , n28999 , 
     n29000 , n29001 , n29002 , n29003 , n29004 , n29005 , n29006 , n29007 , n29008 , n29009 , 
     n29010 , n29011 , n29012 , n29013 , n29014 , n29015 , n29016 , n29017 , n29018 , n29019 , 
     n29020 , n29021 , n29022 , n29023 , n29024 , n29025 , n29026 , n29027 , n29028 , n29029 , 
     n29030 , n29031 , n29032 , n29033 , n29034 , n29035 , n29036 , n29037 , n29038 , n29039 , 
     n29040 , n29041 , n29042 , n29043 , n29044 , n29045 , n29046 , n29047 , n29048 , n29049 , 
     n29050 , n29051 , n29052 , n29053 , n29054 , n29055 , n29056 , n29057 , n29058 , n29059 , 
     n29060 , n29061 , n29062 , n29063 , n29064 , n29065 , n29066 , n29067 , n29068 , n29069 , 
     n29070 , n29071 , n29072 , n29073 , n29074 , n29075 , n29076 , n29077 , n29078 , n29079 , 
     n29080 , n29081 , n29082 , n29083 , n29084 , n29085 , n29086 , n29087 , n29088 , n29089 , 
     n29090 , n29091 , n29092 , n29093 , n29094 , n29095 , n29096 , n29097 , n29098 , n29099 , 
     n29100 , n29101 , n29102 , n29103 , n29104 , n29105 , n29106 , n29107 , n29108 , n29109 , 
     n29110 , n29111 , n29112 , n29113 , n29114 , n29115 , n29116 , n29117 , n29118 , n29119 , 
     n29120 , n29121 , n29122 , n29123 , n29124 , n29125 , n29126 , n29127 , n29128 , n29129 , 
     n29130 , n29131 , n29132 , n29133 , n29134 , n29135 , n29136 , n29137 , n29138 , n29139 , 
     n29140 , n29141 , n29142 , n29143 , n29144 , n29145 , n29146 , n29147 , n29148 , n29149 , 
     n29150 , n29151 , n29152 , n29153 , n29154 , n29155 , n29156 , n29157 , n29158 , n29159 , 
     n29160 , n29161 , n29162 , n29163 , n29164 , n29165 , n29166 , n29167 , n29168 , n29169 , 
     n29170 , n29171 , n29172 , n29173 , n29174 , n29175 , n29176 , n29177 , n29178 , n29179 , 
     n29180 , n29181 , n29182 , n29183 , n29184 , n29185 , n29186 , n29187 , n29188 , n29189 , 
     n29190 , n29191 , n29192 , n29193 , n29194 , n29195 , n29196 , n29197 , n29198 , n29199 , 
     n29200 , n29201 , n29202 , n29203 , n29204 , n29205 , n29206 , n29207 , n29208 , n29209 , 
     n29210 , n29211 , n29212 , n29213 , n29214 , n29215 , n29216 , n29217 , n29218 , n29219 , 
     n29220 , n29221 , n29222 , n29223 , n29224 , n29225 , n29226 , n29227 , n29228 , n29229 , 
     n29230 , n29231 , n29232 , n29233 , n29234 , n29235 , n29236 , n29237 , n29238 , n29239 , 
     n29240 , n29241 , n29242 , n29243 , n29244 , n29245 , n29246 , n29247 , n29248 , n29249 , 
     n29250 , n29251 , n29252 , n29253 , n29254 , n29255 , n29256 , n29257 , n29258 , n29259 , 
     n29260 , n29261 , n29262 , n29263 , n29264 , n29265 , n29266 , n29267 , n29268 , n29269 , 
     n29270 , n29271 , n29272 , n29273 , n29274 , n29275 , n29276 , n29277 , n29278 , n29279 , 
     n29280 , n29281 , n29282 , n29283 , n29284 , n29285 , n29286 , n29287 , n29288 , n29289 , 
     n29290 , n29291 , n29292 , n29293 , n29294 , n29295 , n29296 , n29297 , n29298 , n29299 , 
     n29300 , n29301 , n29302 , n29303 , n29304 , n29305 , n29306 , n29307 , n29308 , n29309 , 
     n29310 , n29311 , n29312 , n29313 , n29314 , n29315 , n29316 , n29317 , n29318 , n29319 , 
     n29320 , n29321 , n29322 , n29323 , n29324 , n29325 , n29326 , n29327 , n29328 , n29329 , 
     n29330 , n29331 , n29332 , n29333 , n29334 , n29335 , n29336 , n29337 , n29338 , n29339 , 
     n29340 , n29341 , n29342 , n29343 , n29344 , n29345 , n29346 , n29347 , n29348 , n29349 , 
     n29350 , n29351 , n29352 , n29353 , n29354 , n29355 , n29356 , n29357 , n29358 , n29359 , 
     n29360 , n29361 , n29362 , n29363 , n29364 , n29365 , n29366 , n29367 , n29368 , n29369 , 
     n29370 , n29371 , n29372 , n29373 , n29374 , n29375 , n29376 , n29377 , n29378 , n29379 , 
     n29380 , n29381 , n29382 , n29383 , n29384 , n29385 , n29386 , n29387 , n29388 , n29389 , 
     n29390 , n29391 , n29392 , n29393 , n29394 , n29395 , n29396 , n29397 , n29398 , n29399 , 
     n29400 , n29401 , n29402 , n29403 , n29404 , n29405 , n29406 , n29407 , n29408 , n29409 , 
     n29410 , n29411 , n29412 , n29413 , n29414 , n29415 , n29416 , n29417 , n29418 , n29419 , 
     n29420 , n29421 , n29422 , n29423 , n29424 , n29425 , n29426 , n29427 , n29428 , n29429 , 
     n29430 , n29431 , n29432 , n29433 , n29434 , n29435 , n29436 , n29437 , n29438 , n29439 , 
     n29440 , n29441 , n29442 , n29443 , n29444 , n29445 , n29446 , n29447 , n29448 , n29449 , 
     n29450 , n29451 , n29452 , n29453 , n29454 , n29455 , n29456 , n29457 , n29458 , n29459 , 
     n29460 , n29461 , n29462 , n29463 , n29464 , n29465 , n29466 , n29467 , n29468 , n29469 , 
     n29470 , n29471 , n29472 , n29473 , n29474 , n29475 , n29476 , n29477 , n29478 , n29479 , 
     n29480 , n29481 , n29482 , n29483 , n29484 , n29485 , n29486 , n29487 , n29488 , n29489 , 
     n29490 , n29491 , n29492 , n29493 , n29494 , n29495 , n29496 , n29497 , n29498 , n29499 , 
     n29500 , n29501 , n29502 , n29503 , n29504 , n29505 , n29506 , n29507 , n29508 , n29509 , 
     n29510 , n29511 , n29512 , n29513 , n29514 , n29515 , n29516 , n29517 , n29518 , n29519 , 
     n29520 , n29521 , n29522 , n29523 , n29524 , n29525 , n29526 , n29527 , n29528 , n29529 , 
     n29530 , n29531 , n29532 , n29533 , n29534 , n29535 , n29536 , n29537 , n29538 , n29539 , 
     n29540 , n29541 , n29542 , n29543 , n29544 , n29545 , n29546 , n29547 , n29548 , n29549 , 
     n29550 , n29551 , n29552 , n29553 , n29554 , n29555 , n29556 , n29557 , n29558 , n29559 , 
     n29560 , n29561 , n29562 , n29563 , n29564 , n29565 , n29566 , n29567 , n29568 , n29569 , 
     n29570 , n29571 , n29572 , n29573 , n29574 , n29575 , n29576 , n29577 , n29578 , n29579 , 
     n29580 , n29581 , n29582 , n29583 , n29584 , n29585 , n29586 , n29587 , n29588 , n29589 , 
     n29590 , n29591 , n29592 , n29593 , n29594 , n29595 , n29596 , n29597 , n29598 , n29599 , 
     n29600 , n29601 , n29602 , n29603 , n29604 , n29605 , n29606 , n29607 , n29608 , n29609 , 
     n29610 , n29611 , n29612 , n29613 , n29614 , n29615 , n29616 , n29617 , n29618 , n29619 , 
     n29620 , n29621 , n29622 , n29623 , n29624 , n29625 , n29626 , n29627 , n29628 , n29629 , 
     n29630 , n29631 , n29632 , n29633 , n29634 , n29635 , n29636 , n29637 , n29638 , n29639 , 
     n29640 , n29641 , n29642 , n29643 , n29644 , n29645 , n29646 , n29647 , n29648 , n29649 , 
     n29650 , n29651 , n29652 , n29653 , n29654 , n29655 , n29656 , n29657 , n29658 , n29659 , 
     n29660 , n29661 , n29662 , n29663 , n29664 , n29665 , n29666 , n29667 , n29668 , n29669 , 
     n29670 , n29671 , n29672 , n29673 , n29674 , n29675 , n29676 , n29677 , n29678 , n29679 , 
     n29680 , n29681 , n29682 , n29683 , n29684 , n29685 , n29686 , n29687 , n29688 , n29689 , 
     n29690 , n29691 , n29692 , n29693 , n29694 , n29695 , n29696 , n29697 , n29698 , n29699 , 
     n29700 , n29701 , n29702 , n29703 , n29704 , n29705 , n29706 , n29707 , n29708 , n29709 , 
     n29710 , n29711 , n29712 , n29713 , n29714 , n29715 , n29716 , n29717 , n29718 , n29719 , 
     n29720 , n29721 , n29722 , n29723 , n29724 , n29725 , n29726 , n29727 , n29728 , n29729 , 
     n29730 , n29731 , n29732 , n29733 , n29734 , n29735 , n29736 , n29737 , n29738 , n29739 , 
     n29740 , n29741 , n29742 , n29743 , n29744 , n29745 , n29746 , n29747 , n29748 , n29749 , 
     n29750 , n29751 , n29752 , n29753 , n29754 , n29755 , n29756 , n29757 , n29758 , n29759 , 
     n29760 , n29761 , n29762 , n29763 , n29764 , n29765 , n29766 , n29767 , n29768 , n29769 , 
     n29770 , n29771 , n29772 , n29773 , n29774 , n29775 , n29776 , n29777 , n29778 , n29779 , 
     n29780 , n29781 , n29782 , n29783 , n29784 , n29785 , n29786 , n29787 , n29788 , n29789 , 
     n29790 , n29791 , n29792 , n29793 , n29794 , n29795 , n29796 , n29797 , n29798 , n29799 , 
     n29800 , n29801 , n29802 , n29803 , n29804 , n29805 , n29806 , n29807 , n29808 , n29809 , 
     n29810 , n29811 , n29812 , n29813 , n29814 , n29815 , n29816 , n29817 , n29818 , n29819 , 
     n29820 , n29821 , n29822 , n29823 , n29824 , n29825 , n29826 , n29827 , n29828 , n29829 , 
     n29830 , n29831 , n29832 , n29833 , n29834 , n29835 , n29836 , n29837 , n29838 , n29839 , 
     n29840 , n29841 , n29842 , n29843 , n29844 , n29845 , n29846 , n29847 , n29848 , n29849 , 
     n29850 , n29851 , n29852 , n29853 , n29854 , n29855 , n29856 , n29857 , n29858 , n29859 , 
     n29860 , n29861 , n29862 , n29863 , n29864 , n29865 , n29866 , n29867 , n29868 , n29869 , 
     n29870 , n29871 , n29872 , n29873 , n29874 , n29875 , n29876 , n29877 , n29878 , n29879 , 
     n29880 , n29881 , n29882 , n29883 , n29884 , n29885 , n29886 , n29887 , n29888 , n29889 , 
     n29890 , n29891 , n29892 , n29893 , n29894 , n29895 , n29896 , n29897 , n29898 , n29899 , 
     n29900 , n29901 , n29902 , n29903 , n29904 , n29905 , n29906 , n29907 , n29908 , n29909 , 
     n29910 , n29911 , n29912 , n29913 , n29914 , n29915 , n29916 , n29917 , n29918 , n29919 , 
     n29920 , n29921 , n29922 , n29923 , n29924 , n29925 , n29926 , n29927 , n29928 , n29929 , 
     n29930 , n29931 , n29932 , n29933 , n29934 , n29935 , n29936 , n29937 , n29938 , n29939 , 
     n29940 , n29941 , n29942 , n29943 , n29944 , n29945 , n29946 , n29947 , n29948 , n29949 , 
     n29950 , n29951 , n29952 , n29953 , n29954 , n29955 , n29956 , n29957 , n29958 , n29959 , 
     n29960 , n29961 , n29962 , n29963 , n29964 , n29965 , n29966 , n29967 , n29968 , n29969 , 
     n29970 , n29971 , n29972 , n29973 , n29974 , n29975 , n29976 , n29977 , n29978 , n29979 , 
     n29980 , n29981 , n29982 , n29983 , n29984 , n29985 , n29986 , n29987 , n29988 , n29989 , 
     n29990 , n29991 , n29992 , n29993 , n29994 , n29995 , n29996 , n29997 , n29998 , n29999 , 
     n30000 , n30001 , n30002 , n30003 , n30004 , n30005 , n30006 , n30007 , n30008 , n30009 , 
     n30010 , n30011 , n30012 , n30013 , n30014 , n30015 , n30016 , n30017 , n30018 , n30019 , 
     n30020 , n30021 , n30022 , n30023 , n30024 , n30025 , n30026 , n30027 , n30028 , n30029 , 
     n30030 , n30031 , n30032 , n30033 , n30034 , n30035 , n30036 , n30037 , n30038 , n30039 , 
     n30040 , n30041 , n30042 , n30043 , n30044 , n30045 , n30046 , n30047 , n30048 , n30049 , 
     n30050 , n30051 , n30052 , n30053 , n30054 , n30055 , n30056 , n30057 , n30058 , n30059 , 
     n30060 , n30061 , n30062 , n30063 , n30064 , n30065 , n30066 , n30067 , n30068 , n30069 , 
     n30070 , n30071 , n30072 , n30073 , n30074 , n30075 , n30076 , n30077 , n30078 , n30079 , 
     n30080 , n30081 , n30082 , n30083 , n30084 , n30085 , n30086 , n30087 , n30088 , n30089 , 
     n30090 , n30091 , n30092 , n30093 , n30094 , n30095 , n30096 , n30097 , n30098 , n30099 , 
     n30100 , n30101 , n30102 , n30103 , n30104 , n30105 , n30106 , n30107 , n30108 , n30109 , 
     n30110 , n30111 , n30112 , n30113 , n30114 , n30115 , n30116 , n30117 , n30118 , n30119 , 
     n30120 , n30121 , n30122 , n30123 , n30124 , n30125 , n30126 , n30127 , n30128 , n30129 , 
     n30130 , n30131 , n30132 , n30133 , n30134 , n30135 , n30136 , n30137 , n30138 , n30139 , 
     n30140 , n30141 , n30142 , n30143 , n30144 , n30145 , n30146 , n30147 , n30148 , n30149 , 
     n30150 , n30151 , n30152 , n30153 , n30154 , n30155 , n30156 , n30157 , n30158 , n30159 , 
     n30160 , n30161 , n30162 , n30163 , n30164 , n30165 , n30166 , n30167 , n30168 , n30169 , 
     n30170 , n30171 , n30172 , n30173 , n30174 , n30175 , n30176 , n30177 , n30178 , n30179 , 
     n30180 , n30181 , n30182 , n30183 , n30184 , n30185 , n30186 , n30187 , n30188 , n30189 , 
     n30190 , n30191 , n30192 , n30193 , n30194 , n30195 , n30196 , n30197 , n30198 , n30199 , 
     n30200 , n30201 , n30202 , n30203 , n30204 , n30205 , n30206 , n30207 , n30208 , n30209 , 
     n30210 , n30211 , n30212 , n30213 , n30214 , n30215 , n30216 , n30217 , n30218 , n30219 , 
     n30220 , n30221 , n30222 , n30223 , n30224 , n30225 , n30226 , n30227 , n30228 , n30229 , 
     n30230 , n30231 , n30232 , n30233 , n30234 , n30235 , n30236 , n30237 , n30238 , n30239 , 
     n30240 , n30241 , n30242 , n30243 , n30244 , n30245 , n30246 , n30247 , n30248 , n30249 , 
     n30250 , n30251 , n30252 , n30253 , n30254 , n30255 , n30256 , n30257 , n30258 , n30259 , 
     n30260 , n30261 , n30262 , n30263 , n30264 , n30265 , n30266 , n30267 , n30268 , n30269 , 
     n30270 , n30271 , n30272 , n30273 , n30274 , n30275 , n30276 , n30277 , n30278 , n30279 , 
     n30280 , n30281 , n30282 , n30283 , n30284 , n30285 , n30286 , n30287 , n30288 , n30289 , 
     n30290 , n30291 , n30292 , n30293 , n30294 , n30295 , n30296 , n30297 , n30298 , n30299 , 
     n30300 , n30301 , n30302 , n30303 , n30304 , n30305 , n30306 , n30307 , n30308 , n30309 , 
     n30310 , n30311 , n30312 , n30313 , n30314 , n30315 , n30316 , n30317 , n30318 , n30319 , 
     n30320 , n30321 , n30322 , n30323 , n30324 , n30325 , n30326 , n30327 , n30328 , n30329 , 
     n30330 , n30331 , n30332 , n30333 , n30334 , n30335 , n30336 , n30337 , n30338 , n30339 , 
     n30340 , n30341 , n30342 , n30343 , n30344 , n30345 , n30346 , n30347 , n30348 , n30349 , 
     n30350 , n30351 , n30352 , n30353 , n30354 , n30355 , n30356 , n30357 , n30358 , n30359 , 
     n30360 , n30361 , n30362 , n30363 , n30364 , n30365 , n30366 , n30367 , n30368 , n30369 , 
     n30370 , n30371 , n30372 , n30373 , n30374 , n30375 , n30376 , n30377 , n30378 , n30379 , 
     n30380 , n30381 , n30382 , n30383 , n30384 , n30385 , n30386 , n30387 , n30388 , n30389 , 
     n30390 , n30391 , n30392 , n30393 , n30394 , n30395 , n30396 , n30397 , n30398 , n30399 , 
     n30400 , n30401 , n30402 ;
buf ( n1 , g0 );
buf ( n2 , g1 );
buf ( n3  , g2 );
buf ( n4  , g3 );
buf ( n5  , g4 );
buf ( n6  , g5 );
buf ( n7  , g6 );
buf ( n8  , g7 );
buf ( n9  , g8 );
buf ( n10  , g9 );
buf ( n11  , g10 );
buf ( n12  , g11 );
buf ( n13  , g12 );
buf ( n14  , g13 );
buf ( n15  , g14 );
buf ( n16  , g15 );
buf ( n17  , g16 );
buf ( n18  , g17 );
buf ( n19  , g18 );
buf ( n20  , g19 );
buf ( n21  , g20 );
buf ( n22  , g21 );
buf ( n23  , g22 );
buf ( n24  , g23 );
buf ( n25  , g24 );
buf ( n26  , g25 );
buf ( n27  , g26 );
buf ( n28  , g27 );
buf ( n29  , g28 );
buf ( n30  , g29 );
buf ( n31  , g30 );
buf ( n32  , g31 );
buf ( n33  , g32 );
buf ( n34  , g33 );
buf ( n35  , g34 );
buf ( n36  , g35 );
buf ( n37  , g36 );
buf ( n38  , g37 );
buf ( n39  , g38 );
buf ( n40  , g39 );
buf ( n41  , g40 );
buf ( n42  , g41 );
buf ( n43  , g42 );
buf ( n44  , g43 );
buf ( n45  , g44 );
buf ( n46  , g45 );
buf ( n47  , g46 );
buf ( n48  , g47 );
buf ( n49  , g48 );
buf ( n50  , g49 );
buf ( n51  , g50 );
buf ( n52  , g51 );
buf ( n53 , g52 );
buf ( n54 , g53 );
buf ( n55 , g54 );
buf ( n56  , g55 );
buf ( n57  , g56 );
buf ( n58  , g57 );
buf ( n59  , g58 );
buf ( n60  , g59 );
buf ( n61  , g60 );
buf ( n62  , g61 );
buf ( n63  , g62 );
buf ( n64  , g63 );
buf ( n65  , g64 );
buf ( n66  , g65 );
buf ( n67  , g66 );
buf ( n68  , g67 );
buf ( n69  , g68 );
buf ( n70  , g69 );
buf ( n71  , g70 );
buf ( n72 , g71 );
buf ( n73 , g72 );
buf ( n74 , g73 );
buf ( n75 , g74 );
buf ( n76 , g75 );
buf ( n77 , g76 );
buf ( n78  , g77 );
buf ( n79  , g78 );
buf ( n80  , g79 );
buf ( n81  , g80 );
buf ( n82  , g81 );
buf ( n83  , g82 );
buf ( n84  , g83 );
buf ( n85  , g84 );
buf ( n86  , g85 );
buf ( n87  , g86 );
buf ( n88 , g87 );
buf ( n89  , g88 );
buf ( n90  , g89 );
buf ( n91  , g90 );
buf ( n92  , g91 );
buf ( n93  , g92 );
buf ( n94  , g93 );
buf ( n95  , g94 );
buf ( n96  , g95 );
buf ( n97  , g96 );
buf ( n98  , g97 );
buf ( n99  , g98 );
buf ( n100  , g99 );
buf ( n101  , g100 );
buf ( n102  , g101 );
buf ( n103  , g102 );
buf ( n104  , g103 );
buf ( n105  , g104 );
buf ( n106  , g105 );
buf ( n107  , g106 );
buf ( n108  , g107 );
buf ( n109  , g108 );
buf ( n110  , g109 );
buf ( n111  , g110 );
buf ( n112  , g111 );
buf ( n113  , g112 );
buf ( n114  , g113 );
buf ( n115  , g114 );
buf ( n116  , g115 );
buf ( n117  , g116 );
buf ( n118  , g117 );
buf ( n119  , g118 );
buf ( n120  , g119 );
buf ( n121  , g120 );
buf ( n122  , g121 );
buf ( n123  , g122 );
buf ( n124  , g123 );
buf ( n125  , g124 );
buf ( n126  , g125 );
buf ( n127  , g126 );
buf ( n128  , g127 );
buf ( n129  , g128 );
buf ( n130  , g129 );
buf ( n131  , g130 );
buf ( n132  , g131 );
buf ( n133  , g132 );
buf ( n134  , g133 );
buf ( n135  , g134 );
buf ( n136  , g135 );
buf ( n137  , g136 );
buf ( n138  , g137 );
buf ( n139  , g138 );
buf ( n140  , g139 );
buf ( n141  , g140 );
buf ( n142  , g141 );
buf ( n143  , g142 );
buf ( n144  , g143 );
buf ( n145  , g144 );
buf ( n146  , g145 );
buf ( n147  , g146 );
buf ( n148  , g147 );
buf ( n149  , g148 );
buf ( n150  , g149 );
buf ( n151  , g150 );
buf ( n152  , g151 );
buf ( n153  , g152 );
buf ( n154  , g153 );
buf ( n155  , g154 );
buf ( n156  , g155 );
buf ( n157  , g156 );
buf ( n158  , g157 );
buf ( n159  , g158 );
buf ( n160  , g159 );
buf ( n161  , g160 );
buf ( n162  , g161 );
buf ( n163  , g162 );
buf ( n164  , g163 );
buf ( n165  , g164 );
buf ( n166  , g165 );
buf ( n167  , g166 );
buf ( n168  , g167 );
buf ( n169  , g168 );
buf ( n170  , g169 );
buf ( n171  , g170 );
buf ( n172  , g171 );
buf ( n173  , g172 );
buf ( n174  , g173 );
buf ( n175  , g174 );
buf ( n176  , g175 );
buf ( n177  , g176 );
buf ( n178  , g177 );
buf ( n179  , g178 );
buf ( n180  , g179 );
buf ( n181  , g180 );
buf ( n182  , g181 );
buf ( n183  , g182 );
buf ( n184  , g183 );
buf ( n185  , g184 );
buf ( n186  , g185 );
buf ( n187  , g186 );
buf ( n188  , g187 );
buf ( n189  , g188 );
buf ( n190  , g189 );
buf ( n191  , g190 );
buf ( n192  , g191 );
buf ( n193  , g192 );
buf ( n194  , g193 );
buf ( n195  , g194 );
buf ( n196  , g195 );
buf ( n197  , g196 );
buf ( n198  , g197 );
buf ( n199  , g198 );
buf ( n200  , g199 );
buf ( n201  , g200 );
buf ( n202  , g201 );
buf ( n203  , g202 );
buf ( n204  , g203 );
buf ( n205  , g204 );
buf ( n206  , g205 );
buf ( n207  , g206 );
buf ( n208  , g207 );
buf ( n209  , g208 );
buf ( n210  , g209 );
buf ( n211  , g210 );
buf ( n212  , g211 );
buf ( n213  , g212 );
buf ( n214  , g213 );
buf ( n215  , g214 );
buf ( n216  , g215 );
buf ( n217  , g216 );
buf ( n218  , g217 );
buf ( n219  , g218 );
buf ( n220  , g219 );
buf ( n221  , g220 );
buf ( n222  , g221 );
buf ( n223  , g222 );
buf ( n224  , g223 );
buf ( n225  , g224 );
buf ( n226  , g225 );
buf ( n227  , g226 );
buf ( n228  , g227 );
buf ( n229  , g228 );
buf ( n230  , g229 );
buf ( n231  , g230 );
buf ( n232  , g231 );
buf ( n233  , g232 );
buf ( n234  , g233 );
buf ( n235  , g234 );
buf ( n236  , g235 );
buf ( n237  , g236 );
buf ( n238  , g237 );
buf ( n239  , g238 );
buf ( n240  , g239 );
buf ( n241  , g240 );
buf ( n242  , g241 );
buf ( n243  , g242 );
buf ( n244  , g243 );
buf ( n245  , g244 );
buf ( n246  , g245 );
buf ( n247  , g246 );
buf ( n248  , g247 );
buf ( n249  , g248 );
buf ( n250  , g249 );
buf ( n251  , g250 );
buf ( n252  , g251 );
buf ( n253  , g252 );
buf ( n254  , g253 );
buf ( n255  , g254 );
buf ( n256  , g255 );
buf ( n257  , g256 );
buf ( n258  , g257 );
buf ( n259  , g258 );
buf ( n260  , g259 );
buf ( n261  , g260 );
buf ( n262  , g261 );
buf ( n263  , g262 );
buf ( n264  , g263 );
buf ( n265  , g264 );
buf ( n266  , g265 );
buf ( n267  , g266 );
buf ( n268  , g267 );
buf ( n269  , g268 );
buf ( n270  , g269 );
buf ( n271  , g270 );
buf ( n272  , g271 );
buf ( n273  , g272 );
buf ( n274  , g273 );
buf ( n275  , g274 );
buf ( n276  , g275 );
buf ( n277  , g276 );
buf ( n278  , g277 );
buf ( n279  , g278 );
buf ( n280  , g279 );
buf ( n281  , g280 );
buf ( n282  , g281 );
buf ( n283  , g282 );
buf ( n284  , g283 );
buf ( n285  , g284 );
buf ( n286  , g285 );
buf ( n287  , g286 );
buf ( n288  , g287 );
buf ( n289  , g288 );
buf ( n290  , g289 );
buf ( n291  , g290 );
buf ( n292  , g291 );
buf ( n293  , g292 );
buf ( n294  , g293 );
buf ( n295  , g294 );
buf ( n296  , g295 );
buf ( n297  , g296 );
buf ( n298  , g297 );
buf ( n299  , g298 );
buf ( n300  , g299 );
buf ( n301  , g300 );
buf ( n302  , g301 );
buf ( n303  , g302 );
buf ( n304  , g303 );
buf ( n305  , g304 );
buf ( n306  , g305 );
buf ( n307  , g306 );
buf ( n308  , g307 );
buf ( n309  , g308 );
buf ( n310  , g309 );
buf ( n311  , g310 );
buf ( n312  , g311 );
buf ( n313  , g312 );
buf ( n314  , g313 );
buf ( n315  , g314 );
buf ( n316  , g315 );
buf ( n317  , g316 );
buf ( n318  , g317 );
buf ( n319  , g318 );
buf ( n320  , g319 );
buf ( n321  , g320 );
buf ( n322  , g321 );
buf ( n323  , g322 );
buf ( n324  , g323 );
buf ( n325  , g324 );
buf ( n326  , g325 );
buf ( n327  , g326 );
buf ( n328  , g327 );
buf ( n329  , g328 );
buf ( n330  , g329 );
buf ( n331  , g330 );
buf ( n332  , g331 );
buf ( n333  , g332 );
buf ( n334  , g333 );
buf ( n335  , g334 );
buf ( n336  , g335 );
buf ( n337  , g336 );
buf ( n338  , g337 );
buf ( n339  , g338 );
buf ( n340  , g339 );
buf ( n341  , g340 );
buf ( n342  , g341 );
buf ( n343  , g342 );
buf ( n344  , g343 );
buf ( n345  , g344 );
buf ( n346  , g345 );
buf ( n347  , g346 );
buf ( n348  , g347 );
buf ( n349  , g348 );
buf ( n350  , g349 );
buf ( n351  , g350 );
buf ( n352  , g351 );
buf ( n353  , g352 );
buf ( n354  , g353 );
buf ( n355  , g354 );
buf ( n356  , g355 );
buf ( n357  , g356 );
buf ( n358  , g357 );
buf ( n359  , g358 );
buf ( n360  , g359 );
buf ( n361  , g360 );
buf ( n362  , g361 );
buf ( n363  , g362 );
buf ( n364  , g363 );
buf ( n365  , g364 );
buf ( n366  , g365 );
buf ( n367  , g366 );
buf ( n368  , g367 );
buf ( n369  , g368 );
buf ( n370  , g369 );
buf ( n371  , g370 );
buf ( n372  , g371 );
buf ( n373  , g372 );
buf ( n374  , g373 );
buf ( n375  , g374 );
buf ( n376  , g375 );
buf ( n377  , g376 );
buf ( n378  , g377 );
buf ( n379  , g378 );
buf ( n380  , g379 );
buf ( n381  , g380 );
buf ( n382  , g381 );
buf ( n383  , g382 );
buf ( n384  , g383 );
buf ( n385  , g384 );
buf ( n386  , g385 );
buf ( n387  , g386 );
buf ( n388  , g387 );
buf ( n389  , g388 );
buf ( n390  , g389 );
buf ( n391  , g390 );
buf ( n392  , g391 );
buf ( n393  , g392 );
buf ( n394  , g393 );
buf ( n395  , g394 );
buf ( n396  , g395 );
buf ( n397  , g396 );
buf ( n398  , g397 );
buf ( n399  , g398 );
buf ( n400  , g399 );
buf ( n401  , g400 );
buf ( n402  , g401 );
buf ( n403  , g402 );
buf ( n404  , g403 );
buf ( n405  , g404 );
buf ( n406  , g405 );
buf ( n407  , g406 );
buf ( n408  , g407 );
buf ( n409  , g408 );
buf ( n410  , g409 );
buf ( n411  , g410 );
buf ( n412  , g411 );
buf ( n413  , g412 );
buf ( n414  , g413 );
buf ( n415  , g414 );
buf ( n416  , g415 );
buf ( n417  , g416 );
buf ( n418  , g417 );
buf ( n419  , g418 );
buf ( n420  , g419 );
buf ( n421  , g420 );
buf ( n422  , g421 );
buf ( n423  , g422 );
buf ( n424  , g423 );
buf ( n425  , g424 );
buf ( n426  , g425 );
buf ( n427  , g426 );
buf ( n428  , g427 );
buf ( n429  , g428 );
buf ( n430  , g429 );
buf ( n431  , g430 );
buf ( n432  , g431 );
buf ( n433  , g432 );
buf ( n434  , g433 );
buf ( n435  , g434 );
buf ( n436  , g435 );
buf ( n437  , g436 );
buf ( n438  , g437 );
buf ( n439  , g438 );
buf ( n440  , g439 );
buf ( n441  , g440 );
buf ( n442  , g441 );
buf ( n443  , g442 );
buf ( n444  , g443 );
buf ( n445  , g444 );
buf ( n446  , g445 );
buf ( n447  , g446 );
buf ( n448  , g447 );
buf ( n449  , g448 );
buf ( n450  , g449 );
buf ( n451  , g450 );
buf ( n452  , g451 );
buf ( n453  , g452 );
buf ( n454  , g453 );
buf ( n455  , g454 );
buf ( n456  , g455 );
buf ( n457  , g456 );
buf ( n458  , g457 );
buf ( n459  , g458 );
buf ( n460  , g459 );
buf ( n461  , g460 );
buf ( n462  , g461 );
buf ( n463  , g462 );
buf ( n464  , g463 );
buf ( n465  , g464 );
buf ( n466  , g465 );
buf ( n467  , g466 );
buf ( n468  , g467 );
buf ( n469  , g468 );
buf ( n470  , g469 );
buf ( n471  , g470 );
buf ( n472  , g471 );
buf ( n473  , g472 );
buf ( n474  , g473 );
buf ( n475  , g474 );
buf ( n476  , g475 );
buf ( n477  , g476 );
buf ( n478  , g477 );
buf ( n479  , g478 );
buf ( n480  , g479 );
buf ( n481  , g480 );
buf ( n482  , g481 );
buf ( n483  , g482 );
buf ( n484  , g483 );
buf ( n485  , g484 );
buf ( n486  , g485 );
buf ( n487  , g486 );
buf ( n488  , g487 );
buf ( n489  , g488 );
buf ( n490  , g489 );
buf ( n491  , g490 );
buf ( n492  , g491 );
buf ( n493  , g492 );
buf ( n494  , g493 );
buf ( n495  , g494 );
buf ( n496  , g495 );
buf ( n497  , g496 );
buf ( n498  , g497 );
buf ( n499  , g498 );
buf ( n500  , g499 );
buf ( n501  , g500 );
buf ( n502  , g501 );
buf ( n503  , g502 );
buf ( n504  , g503 );
buf ( n505  , g504 );
buf ( n506  , g505 );
buf ( n507  , g506 );
buf ( n508  , g507 );
buf ( n509  , g508 );
buf ( n510  , g509 );
buf ( n511  , g510 );
buf ( n512  , g511 );
buf ( n513  , g512 );
buf ( n514  , g513 );
buf ( n515  , g514 );
buf ( n516  , g515 );
buf ( n517  , g516 );
buf ( n518  , g517 );
buf ( n519  , g518 );
buf ( n520  , g519 );
buf ( n521  , g520 );
buf ( n522  , g521 );
buf ( n523  , g522 );
buf ( n524  , g523 );
buf ( n525  , g524 );
buf ( n526  , g525 );
buf ( n527  , g526 );
buf ( n528  , g527 );
buf ( n529  , g528 );
buf ( n530  , g529 );
buf ( n531  , g530 );
buf ( n532  , g531 );
buf ( n533  , g532 );
buf ( n534  , g533 );
buf ( n535  , g534 );
buf ( n536  , g535 );
buf ( n537  , g536 );
buf ( n538  , g537 );
buf ( n539  , g538 );
buf ( n540  , g539 );
buf ( n541  , g540 );
buf ( n542  , g541 );
buf ( n543  , g542 );
buf ( n544  , g543 );
buf ( n545  , g544 );
buf ( n546  , g545 );
buf ( n547  , g546 );
buf ( n548  , g547 );
buf ( n549  , g548 );
buf ( n550  , g549 );
buf ( n551  , g550 );
buf ( n552  , g551 );
buf ( n553  , g552 );
buf ( n554  , g553 );
buf ( n555  , g554 );
buf ( n556  , g555 );
buf ( n557  , g556 );
buf ( n558  , g557 );
buf ( n559  , g558 );
buf ( n560  , g559 );
buf ( n561  , g560 );
buf ( n562  , g561 );
buf ( n563  , g562 );
buf ( n564  , g563 );
buf ( n565  , g564 );
buf ( n566  , g565 );
buf ( n567  , g566 );
buf ( n568  , g567 );
buf ( n569  , g568 );
buf ( n570  , g569 );
buf ( n571  , g570 );
buf ( n572  , g571 );
buf ( n573  , g572 );
buf ( n574  , g573 );
buf ( n575  , g574 );
buf ( n576  , g575 );
buf ( n577  , g576 );
buf ( n578  , g577 );
buf ( n579  , g578 );
buf ( n580  , g579 );
buf ( n581  , g580 );
buf ( n582  , g581 );
buf ( n583  , g582 );
buf ( n584  , g583 );
buf ( n585  , g584 );
buf ( n586  , g585 );
buf ( n587  , g586 );
buf ( n588  , g587 );
buf ( n589  , g588 );
buf ( n590  , g589 );
buf ( n591  , g590 );
buf ( n592  , g591 );
buf ( n593  , g592 );
buf ( n594  , g593 );
buf ( n595  , g594 );
buf ( n596  , g595 );
buf ( n597  , g596 );
buf ( n598  , g597 );
buf ( n599  , g598 );
buf ( n600  , g599 );
buf ( n601  , g600 );
buf ( n602  , g601 );
buf ( n603  , g602 );
buf ( n604  , g603 );
buf ( n605  , g604 );
buf ( n606  , g605 );
buf ( n607  , g606 );
buf ( n608  , g607 );
buf ( n609  , g608 );
buf ( n610  , g609 );
buf ( n611  , g610 );
buf ( n612  , g611 );
buf ( n613  , g612 );
buf ( n614  , g613 );
buf ( n615  , g614 );
buf ( n616  , g615 );
buf ( n617  , g616 );
buf ( n618  , g617 );
buf ( n619  , g618 );
buf ( n620  , g619 );
buf ( n621  , g620 );
buf ( n622  , g621 );
buf ( n623  , g622 );
buf ( n624  , g623 );
buf ( n625  , g624 );
buf ( n626  , g625 );
buf ( n627  , g626 );
buf ( n628  , g627 );
buf ( n629  , g628 );
buf ( n630  , g629 );
buf ( n631  , g630 );
buf ( n632  , g631 );
buf ( n633  , g632 );
buf ( n634  , g633 );
buf ( n635  , g634 );
buf ( n636  , g635 );
buf ( n637  , g636 );
buf ( n638  , g637 );
buf ( n639  , g638 );
buf ( n640  , g639 );
buf ( n641  , g640 );
buf ( n642  , g641 );
buf ( n643  , g642 );
buf ( n644  , g643 );
buf ( n645  , g644 );
buf ( n646  , g645 );
buf ( n647  , g646 );
buf ( n648  , g647 );
buf ( n649  , g648 );
buf ( n650  , g649 );
buf ( n651  , g650 );
buf ( n652  , g651 );
buf ( n653  , g652 );
buf ( n654  , g653 );
buf ( n655  , g654 );
buf ( n656  , g655 );
buf ( n657  , g656 );
buf ( n658  , g657 );
buf ( n659  , g658 );
buf ( n660  , g659 );
buf ( n661  , g660 );
buf ( n662  , g661 );
buf ( n663  , g662 );
buf ( n664  , g663 );
buf ( n665  , g664 );
buf ( n666  , g665 );
buf ( n667  , g666 );
buf ( n668  , g667 );
buf ( n669  , g668 );
buf ( n670  , g669 );
buf ( n671  , g670 );
buf ( n672  , g671 );
buf ( n673  , g672 );
buf ( n674  , g673 );
buf ( n675  , g674 );
buf ( n676  , g675 );
buf ( n677  , g676 );
buf ( n678  , g677 );
buf ( n679  , g678 );
buf ( n680  , g679 );
buf ( n681  , g680 );
buf ( n682  , g681 );
buf ( n683  , g682 );
buf ( n684  , g683 );
buf ( n685  , g684 );
buf ( n686  , g685 );
buf ( n687  , g686 );
buf ( n688  , g687 );
buf ( n689  , g688 );
buf ( n690  , g689 );
buf ( n691  , g690 );
buf ( n692  , g691 );
buf ( n693  , g692 );
buf ( n694  , g693 );
buf ( n695  , g694 );
buf ( n696  , g695 );
buf ( n697  , g696 );
buf ( n698  , g697 );
buf ( n699  , g698 );
buf ( n700  , g699 );
buf ( n701  , g700 );
buf ( n702  , g701 );
buf ( n703  , g702 );
buf ( n704  , g703 );
buf ( n705  , g704 );
buf ( n706  , g705 );
buf ( n707  , g706 );
buf ( n708  , g707 );
buf ( n709  , g708 );
buf ( n710  , g709 );
buf ( n711  , g710 );
buf ( n712  , g711 );
buf ( n713  , g712 );
buf ( n714  , g713 );
buf ( n715  , g714 );
buf ( n716  , g715 );
buf ( n717  , g716 );
buf ( n718  , g717 );
buf ( n719  , g718 );
buf ( n720  , g719 );
buf ( n721  , g720 );
buf ( n722  , g721 );
buf ( n723  , g722 );
buf ( n724  , g723 );
buf ( n725  , g724 );
buf ( n726  , g725 );
buf ( n727  , g726 );
buf ( n728  , g727 );
buf ( n729  , g728 );
buf ( n730  , g729 );
buf ( n731  , g730 );
buf ( n732  , g731 );
buf ( n733  , g732 );
buf ( n734  , g733 );
buf ( n735  , g734 );
buf ( n736  , g735 );
buf ( n737  , g736 );
buf ( n738  , g737 );
buf ( n739  , g738 );
buf ( n740  , g739 );
buf ( n741  , g740 );
buf ( n742  , g741 );
buf ( n743  , g742 );
buf ( n744  , g743 );
buf ( n745  , g744 );
buf ( n746  , g745 );
buf ( n747  , g746 );
buf ( n748  , g747 );
buf ( n749  , g748 );
buf ( n750  , g749 );
buf ( n751  , g750 );
buf ( n752  , g751 );
buf ( n753  , g752 );
buf ( n754  , g753 );
buf ( n755  , g754 );
buf ( n756  , g755 );
buf ( n757  , g756 );
buf ( n758  , g757 );
buf ( n759  , g758 );
buf ( n760  , g759 );
buf ( n761  , g760 );
buf ( n762  , g761 );
buf ( n763  , g762 );
buf ( n764  , g763 );
buf ( n765  , g764 );
buf ( n766  , g765 );
buf ( n767  , g766 );
buf ( n768  , g767 );
buf ( n769  , g768 );
buf ( n770  , g769 );
buf ( n771  , g770 );
buf ( n772  , g771 );
buf ( n773  , g772 );
buf ( n774  , g773 );
buf ( n775  , g774 );
buf ( n776  , g775 );
buf ( n777  , g776 );
buf ( n778  , g777 );
buf ( n779  , g778 );
buf ( n780  , g779 );
buf ( n781  , g780 );
buf ( n782  , g781 );
buf ( n783  , g782 );
buf ( n784  , g783 );
buf ( n785  , g784 );
buf ( n786  , g785 );
buf ( n787  , g786 );
buf ( n788  , g787 );
buf ( n789  , g788 );
buf ( n790  , g789 );
buf ( n791  , g790 );
buf ( n792  , g791 );
buf ( n793  , g792 );
buf ( n794  , g793 );
buf ( n795  , g794 );
buf ( n796  , g795 );
buf ( n797  , g796 );
buf ( n798  , g797 );
buf ( n799  , g798 );
buf ( n800  , g799 );
buf ( n801  , g800 );
buf ( n802  , g801 );
buf ( n803  , g802 );
buf ( n804  , g803 );
buf ( n805  , g804 );
buf ( n806  , g805 );
buf ( n807  , g806 );
buf ( n808  , g807 );
buf ( n809  , g808 );
buf ( n810  , g809 );
buf ( n811  , g810 );
buf ( n812  , g811 );
buf ( n813  , g812 );
buf ( n814  , g813 );
buf ( n815  , g814 );
buf ( n816  , g815 );
buf ( n817  , g816 );
buf ( n818  , g817 );
buf ( n819  , g818 );
buf ( n820  , g819 );
buf ( n821  , g820 );
buf ( n822  , g821 );
buf ( n823  , g822 );
buf ( n824  , g823 );
buf ( n825  , g824 );
buf ( n826  , g825 );
buf ( n827  , g826 );
buf ( n828  , g827 );
buf ( n829  , g828 );
buf ( n830  , g829 );
buf ( n831  , g830 );
buf ( n832  , g831 );
buf ( n833  , g832 );
buf ( n834  , g833 );
buf ( n835  , g834 );
buf ( n836  , g835 );
buf ( n837  , g836 );
buf ( n838  , g837 );
buf ( n839  , g838 );
buf ( n840  , g839 );
buf ( n841  , g840 );
buf ( n842  , g841 );
buf ( n843  , g842 );
buf ( n844  , g843 );
buf ( n845  , g844 );
buf ( n846  , g845 );
buf ( n847  , g846 );
buf ( n848  , g847 );
buf ( n849  , g848 );
buf ( n850  , g849 );
buf ( n851  , g850 );
buf ( n852  , g851 );
buf ( n853  , g852 );
buf ( n854  , g853 );
buf ( n855  , g854 );
buf ( n856  , g855 );
buf ( n857  , g856 );
buf ( n858  , g857 );
buf ( n859  , g858 );
buf ( n860  , g859 );
buf ( n861  , g860 );
buf ( n862  , g861 );
buf ( n863  , g862 );
buf ( n864  , g863 );
buf ( n865  , g864 );
buf ( n866  , g865 );
buf ( n867  , g866 );
buf ( n868  , g867 );
buf ( n869  , g868 );
buf ( n870  , g869 );
buf ( n871  , g870 );
buf ( n872  , g871 );
buf ( n873  , g872 );
buf ( n874  , g873 );
buf ( n875  , g874 );
buf ( n876  , g875 );
buf ( n877  , g876 );
buf ( n878  , g877 );
buf ( n879  , g878 );
buf ( n880  , g879 );
buf ( n881  , g880 );
buf ( n882  , g881 );
buf ( n883  , g882 );
buf ( n884  , g883 );
buf ( n885  , g884 );
buf ( n886  , g885 );
buf ( n887  , g886 );
buf ( n888  , g887 );
buf ( n889  , g888 );
buf ( n890  , g889 );
buf ( n891  , g890 );
buf ( n892  , g891 );
buf ( n893  , g892 );
buf ( n894  , g893 );
buf ( n895  , g894 );
buf ( n896  , g895 );
buf ( n897  , g896 );
buf ( n898  , g897 );
buf ( n899  , g898 );
buf ( n900  , g899 );
buf ( n901  , g900 );
buf ( n902  , g901 );
buf ( n903  , g902 );
buf ( n904  , g903 );
buf ( n905  , g904 );
buf ( n906  , g905 );
buf ( n907  , g906 );
buf ( n908  , g907 );
buf ( n909  , g908 );
buf ( n910  , g909 );
buf ( n911  , g910 );
buf ( n912  , g911 );
buf ( n913  , g912 );
buf ( n914  , g913 );
buf ( n915  , g914 );
buf ( n916  , g915 );
buf ( n917  , g916 );
buf ( n918  , g917 );
buf ( n919  , g918 );
buf ( n920  , g919 );
buf ( n921  , g920 );
buf ( n922  , g921 );
buf ( n923  , g922 );
buf ( n924  , g923 );
buf ( n925  , g924 );
buf ( n926  , g925 );
buf ( n927  , g926 );
buf ( n928  , g927 );
buf ( n929  , g928 );
buf ( n930  , g929 );
buf ( n931  , g930 );
buf ( n932  , g931 );
buf ( n933  , g932 );
buf ( n934  , g933 );
buf ( n935  , g934 );
buf ( n936  , g935 );
buf ( n937  , g936 );
buf ( n938  , g937 );
buf ( n939  , g938 );
buf ( n940  , g939 );
buf ( n941  , g940 );
buf ( n942  , g941 );
buf ( n943  , g942 );
buf ( n944  , g943 );
buf ( n945  , g944 );
buf ( n946  , g945 );
buf ( n947  , g946 );
buf ( n948  , g947 );
buf ( n949  , g948 );
buf ( n950  , g949 );
buf ( n951  , g950 );
buf ( n952  , g951 );
buf ( n953  , g952 );
buf ( n954  , g953 );
buf ( n955  , g954 );
buf ( n956  , g955 );
buf ( n957  , g956 );
buf ( n958  , g957 );
buf ( n959  , g958 );
buf ( n960  , g959 );
buf ( n961  , g960 );
buf ( n962  , g961 );
buf ( n963  , g962 );
buf ( n964  , g963 );
buf ( n965  , g964 );
buf ( n966  , g965 );
buf ( n967  , g966 );
buf ( n968  , g967 );
buf ( n969  , g968 );
buf ( n970  , g969 );
buf ( n971  , g970 );
buf ( n972  , g971 );
buf ( n973  , g972 );
buf ( n974  , g973 );
buf ( n975  , g974 );
buf ( n976  , g975 );
buf ( n977  , g976 );
buf ( n978  , g977 );
buf ( n979  , g978 );
buf ( n980  , g979 );
buf ( n981  , g980 );
buf ( n982  , g981 );
buf ( n983  , g982 );
buf ( n984  , g983 );
buf ( n985  , g984 );
buf ( n986  , g985 );
buf ( n987  , g986 );
buf ( n988  , g987 );
buf ( n989  , g988 );
buf ( n990  , g989 );
buf ( n991  , g990 );
buf ( n992  , g991 );
buf ( n993  , g992 );
buf ( n994  , g993 );
buf ( n995  , g994 );
buf ( n996  , g995 );
buf ( n997  , g996 );
buf ( n998  , g997 );
buf ( n999  , g998 );
buf ( n1000  , g999 );
buf ( n1001  , g1000 );
buf ( n1002  , g1001 );
buf ( n1003  , g1002 );
buf ( n1004  , g1003 );
buf ( n1005  , g1004 );
buf ( n1006  , g1005 );
buf ( n1007  , g1006 );
buf ( n1008  , g1007 );
buf ( n1009  , g1008 );
buf ( n1010  , g1009 );
buf ( n1011  , g1010 );
buf ( n1012  , g1011 );
buf ( n1013  , g1012 );
buf ( n1014  , g1013 );
buf ( n1015  , g1014 );
buf ( n1016  , g1015 );
buf ( n1017  , g1016 );
buf ( n1018  , g1017 );
buf ( n1019  , g1018 );
buf ( n1020  , g1019 );
buf ( n1021  , g1020 );
buf ( n1022  , g1021 );
buf ( n1023  , g1022 );
buf ( n1024  , g1023 );
buf ( n1025  , g1024 );
buf ( n1026  , g1025 );
buf ( n1027  , g1026 );
buf ( n1028  , g1027 );
buf ( n1029  , g1028 );
buf ( n1030  , g1029 );
buf ( n1031  , g1030 );
buf ( n1032  , g1031 );
buf ( n1033  , g1032 );
buf ( n1034  , g1033 );
buf ( n1035  , g1034 );
buf ( n1036  , g1035 );
buf ( n1037  , g1036 );
buf ( n1038  , g1037 );
buf ( n1039  , g1038 );
buf ( n1040  , g1039 );
buf ( n1041  , g1040 );
buf ( n1042  , g1041 );
buf ( n1043  , g1042 );
buf ( n1044  , g1043 );
buf ( n1045  , g1044 );
buf ( n1046  , g1045 );
buf ( n1047  , g1046 );
buf ( n1048  , g1047 );
buf ( n1049  , g1048 );
buf ( n1050  , g1049 );
buf ( n1051  , g1050 );
buf ( n1052  , g1051 );
buf ( n1053  , g1052 );
buf ( n1054  , g1053 );
buf ( n1055  , g1054 );
buf ( n1056  , g1055 );
buf ( n1057  , g1056 );
buf ( n1058  , g1057 );
buf ( n1059  , g1058 );
buf ( n1060  , g1059 );
buf ( n1061  , g1060 );
buf ( n1062  , g1061 );
buf ( n1063  , g1062 );
buf ( n1064  , g1063 );
buf ( n1065  , g1064 );
buf ( n1066  , g1065 );
buf ( n1067  , g1066 );
buf ( n1068  , g1067 );
buf ( n1069  , g1068 );
buf ( n1070  , g1069 );
buf ( n1071  , g1070 );
buf ( n1072  , g1071 );
buf ( n1073  , g1072 );
buf ( n1074  , g1073 );
buf ( n1075  , g1074 );
buf ( n1076  , g1075 );
buf ( n1077  , g1076 );
buf ( n1078  , g1077 );
buf ( n1079  , g1078 );
buf ( n1080  , g1079 );
buf ( n1081  , g1080 );
buf ( n1082  , g1081 );
buf ( n1083  , g1082 );
buf ( n1084  , g1083 );
buf ( n1085  , g1084 );
buf ( n1086  , g1085 );
buf ( n1087  , g1086 );
buf ( n1088  , g1087 );
buf ( n1089  , g1088 );
buf ( n1090  , g1089 );
buf ( n1091  , g1090 );
buf ( n1092  , g1091 );
buf ( n1093  , g1092 );
buf ( n1094  , g1093 );
buf ( n1095  , g1094 );
buf ( n1096  , g1095 );
buf ( n1097  , g1096 );
buf ( n1098  , g1097 );
buf ( n1099  , g1098 );
buf ( n1100  , g1099 );
buf ( n1101  , g1100 );
buf ( n1102  , g1101 );
buf ( n1103  , g1102 );
buf ( n1104  , g1103 );
buf ( n1105  , g1104 );
buf ( n1106  , g1105 );
buf ( n1107  , g1106 );
buf ( n1108  , g1107 );
buf ( n1109  , g1108 );
buf ( n1110  , g1109 );
buf ( n1111  , g1110 );
buf ( n1112  , g1111 );
buf ( n1113  , g1112 );
buf ( n1114  , g1113 );
buf ( n1115  , g1114 );
buf ( n1116  , g1115 );
buf ( n1117  , g1116 );
buf ( n1118  , g1117 );
buf ( n1119  , g1118 );
buf ( n1120  , g1119 );
buf ( n1121  , g1120 );
buf ( n1122  , g1121 );
buf ( n1123  , g1122 );
buf ( n1124  , g1123 );
buf ( n1125  , g1124 );
buf ( n1126  , g1125 );
buf ( n1127  , g1126 );
buf ( n1128  , g1127 );
buf ( n1129  , g1128 );
buf ( n1130  , g1129 );
buf ( n1131  , g1130 );
buf ( n1132  , g1131 );
buf ( n1133  , g1132 );
buf ( n1134  , g1133 );
buf ( n1135  , g1134 );
buf ( n1136  , g1135 );
buf ( n1137  , g1136 );
buf ( n1138  , g1137 );
buf ( n1139  , g1138 );
buf ( n1140  , g1139 );
buf ( n1141  , g1140 );
buf ( n1142  , g1141 );
buf ( n1143  , g1142 );
buf ( n1144  , g1143 );
buf ( n1145  , g1144 );
buf ( n1146  , g1145 );
buf ( n1147  , g1146 );
buf ( n1148  , g1147 );
buf ( n1149  , g1148 );
buf ( n1150  , g1149 );
buf ( n1151  , g1150 );
buf ( n1152  , g1151 );
buf ( n1153  , g1152 );
buf ( n1154  , g1153 );
buf ( n1155  , g1154 );
buf ( n1156  , g1155 );
buf ( n1157  , g1156 );
buf ( n1158  , g1157 );
buf ( n1159  , g1158 );
buf ( n1160  , g1159 );
buf ( n1161  , g1160 );
buf ( n1162  , g1161 );
buf ( n1163  , g1162 );
buf ( n1164  , g1163 );
buf ( n1165  , g1164 );
buf ( n1166  , g1165 );
buf ( n1167  , g1166 );
buf ( n1168  , g1167 );
buf ( n1169  , g1168 );
buf ( n1170  , g1169 );
buf ( n1171  , g1170 );
buf ( n1172  , g1171 );
buf ( n1173  , g1172 );
buf ( n1174  , g1173 );
buf ( n1175  , g1174 );
buf ( n1176  , g1175 );
buf ( n1177  , g1176 );
buf ( n1178  , g1177 );
buf ( n1179  , g1178 );
buf ( n1180  , g1179 );
buf ( n1181  , g1180 );
buf ( n1182  , g1181 );
buf ( n1183  , g1182 );
buf ( n1184  , g1183 );
buf ( n1185  , g1184 );
buf ( n1186  , g1185 );
buf ( n1187  , g1186 );
buf ( n1188  , g1187 );
buf ( n1189  , g1188 );
buf ( n1190  , g1189 );
buf ( n1191  , g1190 );
buf ( n1192  , g1191 );
buf ( n1193  , g1192 );
buf ( n1194  , g1193 );
buf ( n1195  , g1194 );
buf ( n1196  , g1195 );
buf ( n1197  , g1196 );
buf ( n1198  , g1197 );
buf ( n1199  , g1198 );
buf ( n1200  , g1199 );
buf ( n1201  , g1200 );
buf ( n1202  , g1201 );
buf ( n1203  , g1202 );
buf ( n1204  , g1203 );
buf ( n1205  , g1204 );
buf ( n1206  , g1205 );
buf ( n1207  , g1206 );
buf ( n1208  , g1207 );
buf ( n1209  , g1208 );
buf ( n1210  , g1209 );
buf ( n1211  , g1210 );
buf ( n1212  , g1211 );
buf ( n1213  , g1212 );
buf ( n1214  , g1213 );
buf ( n1215  , g1214 );
buf ( n1216  , g1215 );
buf ( n1217  , g1216 );
buf ( n1218  , g1217 );
buf ( n1219  , g1218 );
buf ( n1220  , g1219 );
buf ( n1221  , g1220 );
buf ( n1222  , g1221 );
buf ( n1223  , g1222 );
buf ( n1224  , g1223 );
buf ( n1225  , g1224 );
buf ( n1226  , g1225 );
buf ( n1227  , g1226 );
buf ( n1228  , g1227 );
buf ( n1229  , g1228 );
buf ( n1230  , g1229 );
buf ( n1231  , g1230 );
buf ( n1232  , g1231 );
buf ( n1233  , g1232 );
buf ( n1234  , g1233 );
buf ( n1235  , g1234 );
buf ( n1236  , g1235 );
buf ( n1237  , g1236 );
buf ( n1238  , g1237 );
buf ( n1239  , g1238 );
buf ( n1240  , g1239 );
buf ( n1241  , g1240 );
buf ( n1242  , g1241 );
buf ( n1243  , g1242 );
buf ( n1244  , g1243 );
buf ( n1245  , g1244 );
buf ( n1246  , g1245 );
buf ( n1247  , g1246 );
buf ( n1248  , g1247 );
buf ( n1249  , g1248 );
buf ( n1250  , g1249 );
buf ( n1251  , g1250 );
buf ( n1252  , g1251 );
buf ( n1253  , g1252 );
buf ( n1254  , g1253 );
buf ( n1255  , g1254 );
buf ( n1256  , g1255 );
buf ( n1257  , g1256 );
buf ( n1258  , g1257 );
buf ( n1259  , g1258 );
buf ( n1260  , g1259 );
buf ( n1261  , g1260 );
buf ( n1262  , g1261 );
buf ( n1263  , g1262 );
buf ( n1264  , g1263 );
buf ( n1265  , g1264 );
buf ( n1266  , g1265 );
buf ( n1267  , g1266 );
buf ( n1268  , g1267 );
buf ( n1269  , g1268 );
buf ( n1270  , g1269 );
buf ( n1271  , g1270 );
buf ( n1272  , g1271 );
buf ( n1273  , g1272 );
buf ( n1274  , g1273 );
buf ( n1275  , g1274 );
buf ( n1276  , g1275 );
buf ( n1277  , g1276 );
buf ( n1278  , g1277 );
buf ( n1279  , g1278 );
buf ( n1280  , g1279 );
buf ( n1281  , g1280 );
buf ( n1282  , g1281 );
buf ( n1283  , g1282 );
buf ( n1284  , g1283 );
buf ( n1285  , g1284 );
buf ( n1286  , g1285 );
buf ( n1287  , g1286 );
buf ( n1288  , g1287 );
buf ( n1289  , g1288 );
buf ( n1290  , g1289 );
buf ( n1291  , g1290 );
buf ( n1292  , g1291 );
buf ( n1293  , g1292 );
buf ( n1294  , g1293 );
buf ( n1295  , g1294 );
buf ( n1296  , g1295 );
buf ( n1297  , g1296 );
buf ( n1298  , g1297 );
buf ( n1299  , g1298 );
buf ( n1300  , g1299 );
buf ( n1301  , g1300 );
buf ( n1302  , g1301 );
buf ( n1303  , g1302 );
buf ( n1304  , g1303 );
buf ( n1305  , g1304 );
buf ( n1306  , g1305 );
buf ( n1307  , g1306 );
buf ( n1308  , g1307 );
buf ( n1309  , g1308 );
buf ( n1310  , g1309 );
buf ( n1311  , g1310 );
buf ( n1312  , g1311 );
buf ( n1313  , g1312 );
buf ( n1314  , g1313 );
buf ( n1315  , g1314 );
buf ( n1316  , g1315 );
buf ( n1317  , g1316 );
buf ( n1318  , g1317 );
buf ( n1319  , g1318 );
buf ( n1320  , g1319 );
buf ( n1321  , g1320 );
buf ( n1322  , g1321 );
buf ( n1323  , g1322 );
buf ( n1324  , g1323 );
buf ( n1325  , g1324 );
buf ( n1326  , g1325 );
buf ( n1327  , g1326 );
buf ( n1328  , g1327 );
buf ( n1329  , g1328 );
buf ( n1330  , g1329 );
buf ( n1331  , g1330 );
buf ( n1332  , g1331 );
buf ( n1333  , g1332 );
buf ( n1334  , g1333 );
buf ( n1335  , g1334 );
buf ( n1336  , g1335 );
buf ( n1337  , g1336 );
buf ( n1338  , g1337 );
buf ( n1339  , g1338 );
buf ( n1340  , g1339 );
buf ( n1341  , g1340 );
buf ( n1342  , g1341 );
buf ( n1343  , g1342 );
buf ( n1344  , g1343 );
buf ( n1345  , g1344 );
buf ( n1346  , g1345 );
buf ( n1347  , g1346 );
buf ( n1348  , g1347 );
buf ( n1349  , g1348 );
buf ( n1350  , g1349 );
buf ( n1351  , g1350 );
buf ( n1352  , g1351 );
buf ( n1353  , g1352 );
buf ( n1354  , g1353 );
buf ( n1355  , g1354 );
buf ( n1356  , g1355 );
buf ( n1357  , g1356 );
buf ( n1358  , g1357 );
buf ( n1359  , g1358 );
buf ( n1360  , g1359 );
buf ( n1361  , g1360 );
buf ( n1362  , g1361 );
buf ( n1363  , g1362 );
buf ( n1364  , g1363 );
buf ( n1365  , g1364 );
buf ( n1366  , g1365 );
buf ( n1367  , g1366 );
buf ( n1368  , g1367 );
buf ( n1369  , g1368 );
buf ( n1370  , g1369 );
buf ( n1371  , g1370 );
buf ( n1372  , g1371 );
buf ( n1373  , g1372 );
buf ( n1374  , g1373 );
buf ( n1375  , g1374 );
buf ( n1376  , g1375 );
buf ( n1377  , g1376 );
buf ( n1378  , g1377 );
buf ( n1379  , g1378 );
buf ( n1380  , g1379 );
buf ( n1381  , g1380 );
buf ( n1382  , g1381 );
buf ( n1383  , g1382 );
buf ( n1384  , g1383 );
buf ( n1385  , g1384 );
buf ( n1386  , g1385 );
buf ( n1387  , g1386 );
buf ( n1388  , g1387 );
buf ( n1389  , g1388 );
buf ( n1390  , g1389 );
buf ( n1391  , g1390 );
buf ( n1392  , g1391 );
buf ( n1393  , g1392 );
buf ( n1394  , g1393 );
buf ( n1395  , g1394 );
buf ( n1396  , g1395 );
buf ( n1397  , g1396 );
buf ( n1398  , g1397 );
buf ( n1399  , g1398 );
buf ( n1400  , g1399 );
buf ( n1401  , g1400 );
buf ( n1402  , g1401 );
buf ( n1403  , g1402 );
buf ( n1404  , g1403 );
buf ( n1405  , g1404 );
buf ( n1406  , g1405 );
buf ( n1407  , g1406 );
buf ( n1408  , g1407 );
buf ( n1409  , g1408 );
buf ( n1410  , g1409 );
buf ( n1411  , g1410 );
buf ( n1412  , g1411 );
buf ( n1413  , g1412 );
buf ( n1414  , g1413 );
buf ( n1415  , g1414 );
buf ( n1416  , g1415 );
buf ( n1417  , g1416 );
buf ( n1418  , g1417 );
buf ( n1419  , g1418 );
buf ( n1420  , g1419 );
buf ( n1421  , g1420 );
buf ( n1422  , g1421 );
buf ( n1423  , g1422 );
buf ( n1424  , g1423 );
buf ( n1425  , g1424 );
buf ( n1426  , g1425 );
buf ( n1427  , g1426 );
buf ( n1428  , g1427 );
buf ( n1429  , g1428 );
buf ( n1430  , g1429 );
buf ( n1431  , g1430 );
buf ( n1432  , g1431 );
buf ( n1433  , g1432 );
buf ( n1434  , g1433 );
buf ( n1435  , g1434 );
buf ( n1436  , g1435 );
buf ( n1437  , g1436 );
buf ( n1438  , g1437 );
buf ( n1439  , g1438 );
buf ( n1440  , g1439 );
buf ( n1441  , g1440 );
buf ( n1442  , g1441 );
buf ( n1443  , g1442 );
buf ( n1444  , g1443 );
buf ( n1445  , g1444 );
buf ( n1446  , g1445 );
buf ( n1447  , g1446 );
buf ( n1448  , g1447 );
buf ( n1449  , g1448 );
buf ( n1450  , g1449 );
buf ( n1451  , g1450 );
buf ( n1452  , g1451 );
buf ( n1453  , g1452 );
buf ( n1454  , g1453 );
buf ( n1455  , g1454 );
buf ( n1456  , g1455 );
buf ( n1457  , g1456 );
buf ( n1458  , g1457 );
buf ( n1459  , g1458 );
buf ( n1460  , g1459 );
buf ( n1461  , g1460 );
buf ( n1462  , g1461 );
buf ( n1463  , g1462 );
buf ( n1464  , g1463 );
buf ( n1465  , g1464 );
buf ( n1466  , g1465 );
buf ( n1467  , g1466 );
buf ( n1468  , g1467 );
buf ( n1469  , g1468 );
buf ( n1470  , g1469 );
buf ( n1471  , g1470 );
buf ( n1472  , g1471 );
buf ( n1473  , g1472 );
buf ( n1474  , g1473 );
buf ( n1475  , g1474 );
buf ( n1476  , g1475 );
buf ( n1477  , g1476 );
buf ( n1478  , g1477 );
buf ( n1479  , g1478 );
buf ( n1480  , g1479 );
buf ( n1481  , g1480 );
buf ( n1482  , g1481 );
buf ( n1483  , g1482 );
buf ( n1484  , g1483 );
buf ( n1485  , g1484 );
buf ( n1486  , g1485 );
buf ( n1487  , g1486 );
buf ( n1488  , g1487 );
buf ( n1489  , g1488 );
buf ( n1490  , g1489 );
buf ( n1491  , g1490 );
buf ( n1492  , g1491 );
buf ( n1493  , g1492 );
buf ( n1494  , g1493 );
buf ( n1495  , g1494 );
buf ( n1496  , g1495 );
buf ( n1497  , g1496 );
buf ( n1498  , g1497 );
buf ( n1499  , g1498 );
buf ( n1500  , g1499 );
buf ( n1501  , g1500 );
buf ( n1502  , g1501 );
buf ( n1503  , g1502 );
buf ( n1504  , g1503 );
buf ( n1505  , g1504 );
buf ( n1506  , g1505 );
buf ( n1507  , g1506 );
buf ( n1508  , g1507 );
buf ( n1509  , g1508 );
buf ( n1510  , g1509 );
buf ( n1511  , g1510 );
buf ( n1512  , g1511 );
buf ( n1513  , g1512 );
buf ( n1514  , g1513 );
buf ( n1515  , g1514 );
buf ( n1516  , g1515 );
buf ( n1517  , g1516 );
buf ( n1518  , g1517 );
buf ( n1519  , g1518 );
buf ( n1520  , g1519 );
buf ( n1521  , g1520 );
buf ( n1522  , g1521 );
buf ( n1523  , g1522 );
buf ( n1524  , g1523 );
buf ( n1525  , g1524 );
buf ( n1526  , g1525 );
buf ( n1527  , g1526 );
buf ( n1528  , g1527 );
buf ( n1529  , g1528 );
buf ( n1530  , g1529 );
buf ( n1531  , g1530 );
buf ( n1532  , g1531 );
buf ( n1533  , g1532 );
buf ( n1534  , g1533 );
buf ( n1535  , g1534 );
buf ( n1536  , g1535 );
buf ( n1537  , g1536 );
buf ( n1538  , g1537 );
buf ( n1539  , g1538 );
buf ( n1540  , g1539 );
buf ( n1541  , g1540 );
buf ( n1542  , g1541 );
buf ( n1543  , g1542 );
buf ( n1544  , g1543 );
buf ( n1545  , g1544 );
buf ( n1546  , g1545 );
buf ( n1547  , g1546 );
buf ( n1548  , g1547 );
buf ( n1549  , g1548 );
buf ( n1550  , g1549 );
buf ( n1551  , g1550 );
buf ( n1552  , g1551 );
buf ( n1553  , g1552 );
buf ( n1554  , g1553 );
buf ( n1555  , g1554 );
buf ( n1556  , g1555 );
buf ( n1557  , g1556 );
buf ( n1558  , g1557 );
buf ( n1559  , g1558 );
buf ( n1560  , g1559 );
buf ( n1561  , g1560 );
buf ( n1562  , g1561 );
buf ( n1563  , g1562 );
buf ( n1564  , g1563 );
buf ( n1565  , g1564 );
buf ( n1566  , g1565 );
buf ( n1567  , g1566 );
buf ( n1568  , g1567 );
buf ( n1569  , g1568 );
buf ( n1570  , g1569 );
buf ( n1571  , g1570 );
buf ( n1572  , g1571 );
buf ( n1573  , g1572 );
buf ( n1574  , g1573 );
buf ( n1575  , g1574 );
buf ( n1576  , g1575 );
buf ( n1577  , g1576 );
buf ( n1578  , g1577 );
buf ( n1579  , g1578 );
buf ( n1580  , g1579 );
buf ( n1581  , g1580 );
buf ( n1582  , g1581 );
buf ( n1583  , g1582 );
buf ( n1584  , g1583 );
buf ( n1585  , g1584 );
buf ( n1586  , g1585 );
buf ( n1587  , g1586 );
buf ( n1588  , g1587 );
buf ( n1589  , g1588 );
buf ( n1590  , g1589 );
buf ( n1591  , g1590 );
buf ( n1592  , g1591 );
buf ( n1593  , g1592 );
buf ( n1594  , g1593 );
buf ( n1595  , g1594 );
buf ( n1596  , g1595 );
buf ( n1597  , g1596 );
buf ( n1598  , g1597 );
buf ( n1599  , g1598 );
buf ( n1600  , g1599 );
buf ( n1601  , g1600 );
buf ( n1602  , g1601 );
buf ( n1603  , g1602 );
buf ( n1604  , g1603 );
buf ( n1605  , g1604 );
buf ( n1606  , g1605 );
buf ( n1607  , g1606 );
buf ( n1608  , g1607 );
buf ( n1609  , g1608 );
buf ( n1610  , g1609 );
buf ( n1611  , g1610 );
buf ( n1612  , g1611 );
buf ( n1613  , g1612 );
buf ( n1614  , g1613 );
buf ( n1615  , g1614 );
buf ( n1616  , g1615 );
buf ( n1617  , g1616 );
buf ( n1618  , g1617 );
buf ( n1619  , g1618 );
buf ( n1620  , g1619 );
buf ( n1621  , g1620 );
buf ( n1622  , g1621 );
buf ( n1623  , g1622 );
buf ( n1624  , g1623 );
buf ( n1625  , g1624 );
buf ( n1626  , g1625 );
buf ( n1627  , g1626 );
buf ( n1628  , g1627 );
buf ( n1629  , g1628 );
buf ( n1630  , g1629 );
buf ( n1631  , g1630 );
buf ( n1632  , g1631 );
buf ( n1633  , g1632 );
buf ( n1634  , g1633 );
buf ( n1635  , g1634 );
buf ( n1636  , g1635 );
buf ( n1637  , g1636 );
buf ( n1638  , g1637 );
buf ( n1639  , g1638 );
buf ( n1640  , g1639 );
buf ( n1641  , g1640 );
buf ( n1642  , g1641 );
buf ( n1643  , g1642 );
buf ( n1644  , g1643 );
buf ( n1645  , g1644 );
buf ( n1646  , g1645 );
buf ( n1647  , g1646 );
buf ( n1648  , g1647 );
buf ( n1649  , g1648 );
buf ( n1650  , g1649 );
buf ( n1651  , g1650 );
buf ( n1652  , g1651 );
buf ( n1653  , g1652 );
buf ( n1654  , g1653 );
buf ( n1655  , g1654 );
buf ( n1656  , g1655 );
buf ( n1657  , g1656 );
buf ( n1658  , g1657 );
buf ( n1659  , g1658 );
buf ( n1660  , g1659 );
buf ( n1661  , g1660 );
buf ( n1662  , g1661 );
buf ( n1663  , g1662 );
buf ( n1664  , g1663 );
buf ( n1665  , g1664 );
buf ( n1666  , g1665 );
buf ( n1667  , g1666 );
buf ( n1668  , g1667 );
buf ( n1669  , g1668 );
buf ( n1670  , g1669 );
buf ( n1671  , g1670 );
buf ( n1672  , g1671 );
buf ( n1673  , g1672 );
buf ( n1674  , g1673 );
buf ( n1675  , g1674 );
buf ( n1676  , g1675 );
buf ( n1677  , g1676 );
buf ( n1678  , g1677 );
buf ( n1679  , g1678 );
buf ( n1680  , g1679 );
buf ( n1681  , g1680 );
buf ( n1682  , g1681 );
buf ( n1683  , g1682 );
buf ( n1684  , g1683 );
buf ( n1685  , g1684 );
buf ( n1686  , g1685 );
buf ( n1687  , g1686 );
buf ( n1688  , g1687 );
buf ( n1689  , g1688 );
buf ( n1690  , g1689 );
buf ( n1691  , g1690 );
buf ( n1692  , g1691 );
buf ( n1693  , g1692 );
buf ( n1694  , g1693 );
buf ( n1695  , g1694 );
buf ( n1696  , g1695 );
buf ( n1697  , g1696 );
buf ( n1698  , g1697 );
buf ( n1699  , g1698 );
buf ( n1700  , g1699 );
buf ( n1701  , g1700 );
buf ( n1702  , g1701 );
buf ( n1703  , g1702 );
buf ( n1704  , g1703 );
buf ( n1705  , g1704 );
buf ( n1706  , g1705 );
buf ( n1707  , g1706 );
buf ( n1708  , g1707 );
buf ( n1709  , g1708 );
buf ( n1710  , g1709 );
buf ( n1711  , g1710 );
buf ( n1712  , g1711 );
buf ( n1713  , g1712 );
buf ( n1714  , g1713 );
buf ( n1715  , g1714 );
buf ( n1716  , g1715 );
buf ( n1717  , g1716 );
buf ( n1718  , g1717 );
buf ( n1719  , g1718 );
buf ( n1720  , g1719 );
buf ( n1721  , g1720 );
buf ( n1722  , g1721 );
buf ( n1723  , g1722 );
buf ( n1724  , g1723 );
buf ( n1725  , g1724 );
buf ( n1726  , g1725 );
buf ( n1727  , g1726 );
buf ( n1728  , g1727 );
buf ( n1729  , g1728 );
buf ( n1730  , g1729 );
buf ( n1731  , g1730 );
buf ( n1732  , g1731 );
buf ( n1733  , g1732 );
buf ( n1734  , g1733 );
buf ( n1735  , g1734 );
buf ( n1736  , g1735 );
buf ( n1737  , g1736 );
buf ( n1738  , g1737 );
buf ( n1739  , g1738 );
buf ( n1740  , g1739 );
buf ( n1741  , g1740 );
buf ( n1742  , g1741 );
buf ( n1743  , g1742 );
buf ( n1744  , g1743 );
buf ( n1745  , g1744 );
buf ( n1746  , g1745 );
buf ( n1747  , g1746 );
buf ( n1748  , g1747 );
buf ( n1749  , g1748 );
buf ( n1750  , g1749 );
buf ( n1751  , g1750 );
buf ( n1752  , g1751 );
buf ( n1753  , g1752 );
buf ( n1754  , g1753 );
buf ( n1755  , g1754 );
buf ( n1756  , g1755 );
buf ( n1757  , g1756 );
buf ( n1758  , g1757 );
buf ( n1759  , g1758 );
buf ( n1760  , g1759 );
buf ( n1761  , g1760 );
buf ( n1762  , g1761 );
buf ( n1763  , g1762 );
buf ( n1764  , g1763 );
buf ( n1765  , g1764 );
buf ( n1766  , g1765 );
buf ( n1767  , g1766 );
buf ( n1768  , g1767 );
buf ( n1769  , g1768 );
buf ( n1770  , g1769 );
buf ( n1771  , g1770 );
buf ( n1772  , g1771 );
buf ( n1773  , g1772 );
buf ( n1774  , g1773 );
buf ( n1775  , g1774 );
buf ( n1776  , g1775 );
buf ( n1777  , g1776 );
buf ( n1778  , g1777 );
buf ( n1779  , g1778 );
buf ( n1780  , g1779 );
buf ( n1781  , g1780 );
buf ( n1782  , g1781 );
buf ( n1783  , g1782 );
buf ( n1784  , g1783 );
buf ( n1785  , g1784 );
buf ( n1786  , g1785 );
buf ( n1787  , g1786 );
buf ( n1788  , g1787 );
buf ( n1789  , g1788 );
buf ( n1790  , g1789 );
buf ( n1791  , g1790 );
buf ( n1792  , g1791 );
buf ( n1793  , g1792 );
buf ( n1794  , g1793 );
buf ( n1795  , g1794 );
buf ( n1796  , g1795 );
buf ( n1797  , g1796 );
buf ( n1798  , g1797 );
buf ( n1799  , g1798 );
buf ( n1800  , g1799 );
buf ( n1801  , g1800 );
buf ( n1802  , g1801 );
buf ( n1803  , g1802 );
buf ( n1804  , g1803 );
buf ( n1805  , g1804 );
buf ( n1806  , g1805 );
buf ( n1807  , g1806 );
buf ( n1808  , g1807 );
buf ( n1809  , g1808 );
buf ( n1810  , g1809 );
buf ( n1811  , g1810 );
buf ( n1812  , g1811 );
buf ( n1813  , g1812 );
buf ( n1814  , g1813 );
buf ( n1815  , g1814 );
buf ( n1816  , g1815 );
buf ( n1817  , g1816 );
buf ( n1818  , g1817 );
buf ( n1819  , g1818 );
buf ( n1820  , g1819 );
buf ( n1821  , g1820 );
buf ( n1822  , g1821 );
buf ( n1823  , g1822 );
buf ( n1824  , g1823 );
buf ( n1825  , g1824 );
buf ( n1826  , g1825 );
buf ( n1827  , g1826 );
buf ( n1828  , g1827 );
buf ( n1829  , g1828 );
buf ( n1830  , g1829 );
buf ( n1831  , g1830 );
buf ( n1832  , g1831 );
buf ( n1833  , g1832 );
buf ( n1834  , g1833 );
buf ( n1835  , g1834 );
buf ( n1836  , g1835 );
buf ( n1837  , g1836 );
buf ( n1838  , g1837 );
buf ( n1839  , g1838 );
buf ( n1840  , g1839 );
buf ( n1841  , g1840 );
buf ( n1842  , g1841 );
buf ( n1843  , g1842 );
buf ( n1844  , g1843 );
buf ( n1845  , g1844 );
buf ( n1846  , g1845 );
buf ( n1847  , g1846 );
buf ( n1848  , g1847 );
buf ( n1849  , g1848 );
buf ( n1850  , g1849 );
buf ( n1851  , g1850 );
buf ( n1852  , g1851 );
buf ( n1853  , g1852 );
buf ( n1854  , g1853 );
buf ( n1855  , g1854 );
buf ( n1856  , g1855 );
buf ( n1857  , g1856 );
buf ( n1858  , g1857 );
buf ( n1859  , g1858 );
buf ( n1860  , g1859 );
buf ( n1861  , g1860 );
buf ( n1862  , g1861 );
buf ( n1863  , g1862 );
buf ( n1864  , g1863 );
buf ( n1865  , g1864 );
buf ( n1866  , g1865 );
buf ( n1867  , g1866 );
buf ( n1868  , g1867 );
buf ( n1869  , g1868 );
buf ( n1870  , g1869 );
buf ( n1871  , g1870 );
buf ( n1872  , g1871 );
buf ( n1873  , g1872 );
buf ( n1874  , g1873 );
buf ( g1874 , n1875  );
buf ( g1875 , n1876  );
buf ( g1876 , n1877  );
buf ( g1877 , n1878  );
buf ( g1878 , n1879  );
buf ( g1879 , n1880  );
buf ( g1880 , n1881  );
buf ( g1881 , n1882  );
buf ( g1882 , n1883  );
buf ( g1883 , n1884  );
buf ( g1884 , n1885  );
buf ( g1885 , n1886  );
buf ( g1886 , n1887  );
buf ( g1887 , n1888  );
buf ( g1888 , n1889  );
buf ( g1889 , n1890  );
buf ( g1890 , n1891  );
buf ( g1891 , n1892  );
buf ( g1892 , n1893  );
buf ( g1893 , n1894  );
buf ( g1894 , n1895  );
buf ( g1895 , n1896  );
buf ( g1896 , n1897  );
buf ( g1897 , n1898  );
buf ( g1898 , n1899  );
buf ( g1899 , n1900  );
buf ( g1900 , n1901  );
buf ( g1901 , n1902  );
buf ( g1902 , n1903  );
buf ( g1903 , n1904  );
buf ( g1904 , n1905  );
buf ( g1905 , n1906  );
buf ( g1906 , n1907 );
buf ( g1907 , n1908 );
buf ( g1908 , n1909 );
buf ( g1909 , n1910  );
buf ( g1910 , n1911  );
buf ( g1911 , n1912  );
buf ( g1912 , n1913  );
buf ( g1913 , n1914  );
buf ( g1914 , n1915  );
buf ( g1915 , n1916  );
buf ( g1916 , n1917  );
buf ( g1917 , n1918  );
buf ( g1918 , n1919  );
buf ( g1919 , n1920  );
buf ( g1920 , n1921  );
buf ( g1921 , n1922  );
buf ( g1922 , n1923  );
buf ( g1923 , n1924  );
buf ( g1924 , n1925  );
buf ( g1925 , n1926 );
buf ( g1926 , n1927 );
buf ( g1927 , n1928  );
buf ( g1928 , n1929  );
buf ( g1929 , n1930  );
buf ( g1930 , n1931  );
buf ( g1931 , n1932  );
buf ( g1932 , n1933  );
buf ( g1933 , n1934  );
buf ( g1934 , n1935  );
buf ( g1935 , n1936 );
buf ( g1936 , n1937 );
buf ( g1937 , n1938 );
buf ( g1938 , n1939 );
buf ( g1939 , n1940  );
buf ( g1940 , n1941  );
buf ( g1941 , n1942 );
buf ( g1942 , n1943  );
buf ( g1943 , n1944  );
buf ( g1944 , n1945  );
buf ( g1945 , n1946  );
buf ( g1946 , n1947  );
buf ( g1947 , n1948  );
buf ( g1948 , n1949  );
buf ( g1949 , n1950  );
buf ( g1950 , n1951  );
buf ( g1951 , n1952  );
buf ( g1952 , n1953  );
buf ( g1953 , n1954  );
buf ( g1954 , n1955  );
buf ( g1955 , n1956  );
buf ( g1956 , n1957  );
buf ( g1957 , n1958  );
buf ( g1958 , n1959  );
buf ( g1959 , n1960  );
buf ( g1960 , n1961  );
buf ( g1961 , n1962  );
buf ( g1962 , n1963  );
buf ( g1963 , n1964  );
buf ( g1964 , n1965  );
buf ( g1965 , n1966  );
buf ( g1966 , n1967  );
buf ( g1967 , n1968  );
buf ( g1968 , n1969  );
buf ( g1969 , n1970  );
buf ( g1970 , n1971  );
buf ( g1971 , n1972  );
buf ( g1972 , n1973  );
buf ( g1973 , n1974  );
buf ( g1974 , n1975  );
buf ( g1975 , n1976  );
buf ( g1976 , n1977  );
buf ( g1977 , n1978  );
buf ( g1978 , n1979  );
buf ( g1979 , n1980  );
buf ( g1980 , n1981  );
buf ( g1981 , n1982  );
buf ( g1982 , n1983  );
buf ( g1983 , n1984  );
buf ( g1984 , n1985  );
buf ( g1985 , n1986  );
buf ( g1986 , n1987  );
buf ( g1987 , n1988  );
buf ( g1988 , n1989  );
buf ( g1989 , n1990  );
buf ( g1990 , n1991  );
buf ( g1991 , n1992  );
buf ( g1992 , n1993  );
buf ( g1993 , n1994 );
buf ( g1994 , n1995 );
buf ( g1995 , n1996  );
buf ( g1996 , n1997  );
buf ( g1997 , n1998  );
buf ( g1998 , n1999  );
buf ( g1999 , n2000  );
buf ( g2000 , n2001  );
buf ( g2001 , n2002  );
buf ( g2002 , n2003  );
buf ( g2003 , n2004  );
buf ( g2004 , n2005  );
buf ( g2005 , n2006  );
buf ( g2006 , n2007  );
buf ( g2007 , n2008  );
buf ( g2008 , n2009  );
buf ( g2009 , n2010  );
buf ( g2010 , n2011  );
buf ( g2011 , n2012  );
buf ( g2012 , n2013  );
buf ( g2013 , n2014  );
buf ( g2014 , n2015  );
buf ( g2015 , n2016  );
buf ( g2016 , n2017  );
buf ( g2017 , n2018  );
buf ( g2018 , n2019  );
buf ( g2019 , n2020  );
buf ( g2020 , n2021  );
buf ( g2021 , n2022  );
buf ( g2022 , n2023  );
buf ( g2023 , n2024  );
buf ( g2024 , n2025  );
buf ( g2025 , n2026  );
buf ( g2026 , n2027  );
buf ( g2027 , n2028  );
buf ( g2028 , n2029  );
buf ( g2029 , n2030  );
buf ( g2030 , n2031  );
buf ( g2031 , n2032  );
buf ( g2032 , n2033  );
buf ( g2033 , n2034  );
buf ( g2034 , n2035  );
buf ( g2035 , n2036  );
buf ( g2036 , n2037  );
buf ( g2037 , n2038  );
buf ( g2038 , n2039  );
buf ( g2039 , n2040  );
buf ( g2040 , n2041  );
buf ( g2041 , n2042  );
buf ( g2042 , n2043  );
buf ( g2043 , n2044  );
buf ( g2044 , n2045  );
buf ( g2045 , n2046  );
buf ( g2046 , n2047  );
buf ( g2047 , n2048  );
buf ( g2048 , n2049  );
buf ( g2049 , n2050  );
buf ( g2050 , n2051  );
buf ( g2051 , n2052  );
buf ( g2052 , n2053  );
buf ( g2053 , n2054  );
buf ( g2054 , n2055  );
buf ( g2055 , n2056  );
buf ( g2056 , n2057  );
buf ( g2057 , n2058  );
buf ( g2058 , n2059  );
buf ( g2059 , n2060  );
buf ( g2060 , n2061  );
buf ( g2061 , n2062  );
buf ( g2062 , n2063  );
buf ( g2063 , n2064  );
buf ( g2064 , n2065  );
buf ( g2065 , n2066  );
buf ( g2066 , n2067  );
buf ( g2067 , n2068  );
buf ( g2068 , n2069  );
buf ( g2069 , n2070  );
buf ( g2070 , n2071  );
buf ( g2071 , n2072  );
buf ( g2072 , n2073  );
buf ( g2073 , n2074  );
buf ( g2074 , n2075  );
buf ( g2075 , n2076  );
buf ( g2076 , n2077  );
buf ( g2077 , n2078  );
buf ( g2078 , n2079  );
buf ( g2079 , n2080  );
buf ( g2080 , n2081  );
buf ( g2081 , n2082  );
buf ( g2082 , n2083  );
buf ( g2083 , n2084  );
buf ( g2084 , n2085  );
buf ( g2085 , n2086  );
buf ( g2086 , n2087  );
buf ( g2087 , n2088  );
buf ( g2088 , n2089  );
buf ( g2089 , n2090  );
buf ( g2090 , n2091  );
buf ( g2091 , n2092  );
buf ( g2092 , n2093  );
buf ( g2093 , n2094  );
buf ( g2094 , n2095  );
buf ( g2095 , n2096  );
buf ( g2096 , n2097  );
buf ( g2097 , n2098  );
buf ( g2098 , n2099  );
buf ( g2099 , n2100  );
buf ( g2100 , n2101  );
buf ( g2101 , n2102  );
buf ( g2102 , n2103  );
buf ( g2103 , n2104  );
buf ( g2104 , n2105  );
buf ( g2105 , n2106  );
buf ( g2106 , n2107  );
buf ( g2107 , n2108  );
buf ( g2108 , n2109  );
buf ( g2109 , n2110  );
buf ( g2110 , n2111  );
buf ( g2111 , n2112  );
buf ( g2112 , n2113  );
buf ( g2113 , n2114  );
buf ( g2114 , n2115  );
buf ( g2115 , n2116  );
buf ( g2116 , n2117  );
buf ( g2117 , n2118  );
buf ( g2118 , n2119  );
buf ( g2119 , n2120  );
buf ( g2120 , n2121  );
buf ( g2121 , n2122  );
buf ( g2122 , n2123  );
buf ( g2123 , n2124  );
buf ( g2124 , n2125  );
buf ( g2125 , n2126  );
buf ( g2126 , n2127  );
buf ( g2127 , n2128  );
buf ( g2128 , n2129  );
buf ( g2129 , n2130  );
buf ( g2130 , n2131  );
buf ( g2131 , n2132  );
buf ( g2132 , n2133  );
buf ( g2133 , n2134  );
buf ( g2134 , n2135  );
buf ( g2135 , n2136  );
buf ( g2136 , n2137  );
buf ( g2137 , n2138  );
buf ( g2138 , n2139  );
buf ( g2139 , n2140  );
buf ( g2140 , n2141  );
buf ( g2141 , n2142  );
buf ( g2142 , n2143  );
buf ( g2143 , n2144  );
buf ( g2144 , n2145  );
buf ( g2145 , n2146  );
buf ( g2146 , n2147  );
buf ( g2147 , n2148  );
buf ( g2148 , n2149  );
buf ( g2149 , n2150  );
buf ( g2150 , n2151  );
buf ( g2151 , n2152  );
buf ( g2152 , n2153  );
buf ( g2153 , n2154  );
buf ( g2154 , n2155  );
buf ( g2155 , n2156  );
buf ( g2156 , n2157  );
buf ( g2157 , n2158  );
buf ( g2158 , n2159  );
buf ( g2159 , n2160  );
buf ( g2160 , n2161  );
buf ( g2161 , n2162  );
buf ( g2162 , n2163  );
buf ( g2163 , n2164  );
buf ( g2164 , n2165  );
buf ( g2165 , n2166  );
buf ( g2166 , n2167  );
buf ( g2167 , n2168  );
buf ( g2168 , n2169  );
buf ( g2169 , n2170  );
buf ( g2170 , n2171  );
buf ( g2171 , n2172  );
buf ( g2172 , n2173  );
buf ( g2173 , n2174  );
buf ( g2174 , n2175  );
buf ( g2175 , n2176  );
buf ( g2176 , n2177  );
buf ( g2177 , n2178  );
buf ( g2178 , n2179  );
buf ( g2179 , n2180  );
buf ( g2180 , n2181  );
buf ( g2181 , n2182  );
buf ( g2182 , n2183  );
buf ( g2183 , n2184  );
buf ( g2184 , n2185  );
buf ( g2185 , n2186  );
buf ( g2186 , n2187  );
buf ( g2187 , n2188  );
buf ( g2188 , n2189  );
buf ( g2189 , n2190  );
buf ( g2190 , n2191  );
buf ( g2191 , n2192  );
buf ( g2192 , n2193  );
buf ( g2193 , n2194  );
buf ( g2194 , n2195  );
buf ( g2195 , n2196  );
buf ( g2196 , n2197  );
buf ( g2197 , n2198  );
buf ( g2198 , n2199  );
buf ( g2199 , n2200  );
buf ( g2200 , n2201  );
buf ( g2201 , n2202  );
buf ( g2202 , n2203  );
buf ( g2203 , n2204  );
buf ( g2204 , n2205  );
buf ( g2205 , n2206  );
buf ( g2206 , n2207  );
buf ( g2207 , n2208  );
buf ( g2208 , n2209  );
buf ( g2209 , n2210  );
buf ( g2210 , n2211  );
buf ( g2211 , n2212  );
buf ( g2212 , n2213  );
buf ( g2213 , n2214  );
buf ( g2214 , n2215  );
buf ( g2215 , n2216  );
buf ( g2216 , n2217  );
buf ( g2217 , n2218  );
buf ( g2218 , n2219  );
buf ( g2219 , n2220  );
buf ( g2220 , n2221  );
buf ( g2221 , n2222  );
buf ( g2222 , n2223  );
buf ( g2223 , n2224  );
buf ( g2224 , n2225  );
buf ( g2225 , n2226  );
buf ( g2226 , n2227  );
buf ( g2227 , n2228  );
buf ( g2228 , n2229  );
buf ( g2229 , n2230  );
buf ( g2230 , n2231  );
buf ( g2231 , n2232  );
buf ( g2232 , n2233  );
buf ( g2233 , n2234  );
buf ( g2234 , n2235  );
buf ( g2235 , n2236  );
buf ( g2236 , n2237  );
buf ( g2237 , n2238  );
buf ( g2238 , n2239  );
buf ( g2239 , n2240  );
buf ( g2240 , n2241  );
buf ( g2241 , n2242  );
buf ( g2242 , n2243  );
buf ( g2243 , n2244  );
buf ( g2244 , n2245  );
buf ( g2245 , n2246  );
buf ( g2246 , n2247  );
buf ( g2247 , n2248  );
buf ( g2248 , n2249  );
buf ( g2249 , n2250  );
buf ( g2250 , n2251  );
buf ( g2251 , n2252  );
buf ( g2252 , n2253  );
buf ( g2253 , n2254  );
buf ( g2254 , n2255  );
buf ( g2255 , n2256  );
buf ( g2256 , n2257  );
buf ( g2257 , n2258  );
buf ( g2258 , n2259  );
buf ( g2259 , n2260  );
buf ( g2260 , n2261  );
buf ( g2261 , n2262  );
buf ( g2262 , n2263  );
buf ( g2263 , n2264  );
buf ( g2264 , n2265  );
buf ( g2265 , n2266  );
buf ( g2266 , n2267  );
buf ( g2267 , n2268  );
buf ( g2268 , n2269  );
buf ( g2269 , n2270  );
buf ( g2270 , n2271  );
buf ( g2271 , n2272  );
buf ( g2272 , n2273  );
buf ( g2273 , n2274  );
buf ( g2274 , n2275  );
buf ( g2275 , n2276  );
buf ( g2276 , n2277  );
buf ( g2277 , n2278  );
buf ( g2278 , n2279  );
buf ( g2279 , n2280  );
buf ( g2280 , n2281  );
buf ( g2281 , n2282  );
buf ( g2282 , n2283  );
buf ( g2283 , n2284  );
buf ( g2284 , n2285  );
buf ( g2285 , n2286  );
buf ( g2286 , n2287  );
buf ( g2287 , n2288  );
buf ( g2288 , n2289  );
buf ( g2289 , n2290  );
buf ( g2290 , n2291  );
buf ( g2291 , n2292  );
buf ( g2292 , n2293  );
buf ( g2293 , n2294  );
buf ( g2294 , n2295  );
buf ( g2295 , n2296  );
buf ( g2296 , n2297  );
buf ( g2297 , n2298  );
buf ( g2298 , n2299  );
buf ( g2299 , n2300  );
buf ( g2300 , n2301  );
buf ( g2301 , n2302  );
buf ( g2302 , n2303  );
buf ( g2303 , n2304  );
buf ( g2304 , n2305  );
buf ( g2305 , n2306  );
buf ( g2306 , n2307  );
buf ( g2307 , n2308  );
buf ( g2308 , n2309  );
buf ( g2309 , n2310  );
buf ( g2310 , n2311  );
buf ( g2311 , n2312  );
buf ( g2312 , n2313  );
buf ( g2313 , n2314  );
buf ( g2314 , n2315  );
buf ( g2315 , n2316  );
buf ( g2316 , n2317  );
buf ( g2317 , n2318  );
buf ( g2318 , n2319  );
buf ( g2319 , n2320  );
buf ( g2320 , n2321  );
buf ( g2321 , n2322  );
buf ( g2322 , n2323  );
buf ( g2323 , n2324  );
buf ( g2324 , n2325  );
buf ( g2325 , n2326  );
buf ( g2326 , n2327  );
buf ( g2327 , n2328  );
buf ( g2328 , n2329  );
buf ( g2329 , n2330  );
buf ( g2330 , n2331  );
buf ( g2331 , n2332  );
buf ( g2332 , n2333  );
buf ( g2333 , n2334  );
buf ( g2334 , n2335  );
buf ( g2335 , n2336  );
buf ( g2336 , n2337  );
buf ( g2337 , n2338  );
buf ( g2338 , n2339  );
buf ( g2339 , n2340  );
buf ( g2340 , n2341  );
buf ( g2341 , n2342  );
buf ( g2342 , n2343  );
buf ( g2343 , n2344  );
buf ( g2344 , n2345  );
buf ( g2345 , n2346  );
buf ( g2346 , n2347  );
buf ( g2347 , n2348  );
buf ( g2348 , n2349  );
buf ( g2349 , n2350  );
buf ( g2350 , n2351  );
buf ( g2351 , n2352  );
buf ( g2352 , n2353  );
buf ( g2353 , n2354  );
buf ( g2354 , n2355  );
buf ( g2355 , n2356  );
buf ( g2356 , n2357  );
buf ( g2357 , n2358  );
buf ( g2358 , n2359  );
buf ( g2359 , n2360  );
buf ( g2360 , n2361  );
buf ( g2361 , n2362  );
buf ( g2362 , n2363  );
buf ( g2363 , n2364  );
buf ( g2364 , n2365  );
buf ( g2365 , n2366  );
buf ( g2366 , n2367  );
buf ( g2367 , n2368  );
buf ( g2368 , n2369  );
buf ( g2369 , n2370  );
buf ( g2370 , n2371  );
buf ( g2371 , n2372  );
buf ( g2372 , n2373  );
buf ( g2373 , n2374  );
buf ( g2374 , n2375  );
buf ( g2375 , n2376  );
buf ( g2376 , n2377  );
buf ( g2377 , n2378  );
buf ( g2378 , n2379  );
buf ( g2379 , n2380  );
buf ( g2380 , n2381  );
buf ( g2381 , n2382  );
buf ( g2382 , n2383  );
buf ( g2383 , n2384  );
buf ( g2384 , n2385  );
buf ( g2385 , n2386  );
buf ( g2386 , n2387  );
buf ( g2387 , n2388  );
buf ( g2388 , n2389  );
buf ( g2389 , n2390  );
buf ( g2390 , n2391  );
buf ( g2391 , n2392  );
buf ( g2392 , n2393  );
buf ( g2393 , n2394  );
buf ( g2394 , n2395  );
buf ( g2395 , n2396  );
buf ( g2396 , n2397  );
buf ( g2397 , n2398  );
buf ( g2398 , n2399  );
buf ( g2399 , n2400  );
buf ( g2400 , n2401  );
buf ( g2401 , n2402  );
buf ( g2402 , n2403  );
buf ( g2403 , n2404  );
buf ( g2404 , n2405  );
buf ( g2405 , n2406  );
buf ( g2406 , n2407  );
buf ( g2407 , n2408  );
buf ( g2408 , n2409  );
buf ( g2409 , n2410  );
buf ( g2410 , n2411  );
buf ( g2411 , n2412  );
buf ( g2412 , n2413  );
buf ( g2413 , n2414  );
buf ( g2414 , n2415  );
buf ( g2415 , n2416  );
buf ( g2416 , n2417  );
buf ( g2417 , n2418  );
buf ( g2418 , n2419  );
buf ( g2419 , n2420  );
buf ( g2420 , n2421  );
buf ( g2421 , n2422  );
buf ( g2422 , n2423  );
buf ( g2423 , n2424  );
buf ( g2424 , n2425  );
buf ( g2425 , n2426  );
buf ( g2426 , n2427  );
buf ( g2427 , n2428  );
buf ( g2428 , n2429  );
buf ( g2429 , n2430  );
buf ( g2430 , n2431  );
buf ( g2431 , n2432  );
buf ( g2432 , n2433  );
buf ( g2433 , n2434  );
buf ( g2434 , n2435  );
buf ( g2435 , n2436  );
buf ( g2436 , n2437  );
buf ( g2437 , n2438  );
buf ( g2438 , n2439  );
buf ( g2439 , n2440  );
buf ( g2440 , n2441  );
buf ( g2441 , n2442  );
buf ( g2442 , n2443  );
buf ( g2443 , n2444  );
buf ( g2444 , n2445  );
buf ( g2445 , n2446  );
buf ( g2446 , n2447  );
buf ( g2447 , n2448  );
buf ( g2448 , n2449  );
buf ( g2449 , n2450  );
buf ( g2450 , n2451  );
buf ( g2451 , n2452  );
buf ( g2452 , n2453  );
buf ( g2453 , n2454  );
buf ( g2454 , n2455  );
buf ( g2455 , n2456  );
buf ( g2456 , n2457  );
buf ( g2457 , n2458  );
buf ( g2458 , n2459  );
buf ( g2459 , n2460  );
buf ( g2460 , n2461  );
buf ( g2461 , n2462  );
buf ( g2462 , n2463  );
buf ( g2463 , n2464  );
buf ( g2464 , n2465  );
buf ( g2465 , n2466  );
buf ( g2466 , n2467  );
buf ( g2467 , n2468  );
buf ( g2468 , n2469  );
buf ( g2469 , n2470  );
buf ( g2470 , n2471  );
buf ( g2471 , n2472  );
buf ( g2472 , n2473  );
buf ( g2473 , n2474  );
buf ( g2474 , n2475  );
buf ( g2475 , n2476  );
buf ( g2476 , n2477  );
buf ( g2477 , n2478  );
buf ( g2478 , n2479  );
buf ( g2479 , n2480  );
buf ( g2480 , n2481  );
buf ( g2481 , n2482  );
buf ( g2482 , n2483  );
buf ( g2483 , n2484  );
buf ( g2484 , n2485  );
buf ( g2485 , n2486  );
buf ( g2486 , n2487  );
buf ( g2487 , n2488  );
buf ( g2488 , n2489  );
buf ( g2489 , n2490  );
buf ( g2490 , n2491  );
buf ( g2491 , n2492  );
buf ( g2492 , n2493  );
buf ( g2493 , n2494  );
buf ( g2494 , n2495  );
buf ( g2495 , n2496  );
buf ( g2496 , n2497  );
buf ( g2497 , n2498  );
buf ( g2498 , n2499  );
buf ( g2499 , n2500  );
buf ( g2500 , n2501  );
buf ( g2501 , n2502  );
buf ( g2502 , n2503  );
buf ( g2503 , n2504  );
buf ( g2504 , n2505  );
buf ( g2505 , n2506  );
buf ( g2506 , n2507  );
buf ( g2507 , n2508  );
buf ( g2508 , n2509  );
buf ( g2509 , n2510  );
buf ( g2510 , n2511  );
buf ( g2511 , n2512  );
buf ( g2512 , n2513  );
buf ( g2513 , n2514  );
buf ( g2514 , n2515  );
buf ( g2515 , n2516  );
buf ( g2516 , n2517  );
buf ( g2517 , n2518  );
buf ( g2518 , n2519  );
buf ( g2519 , n2520  );
buf ( g2520 , n2521  );
buf ( g2521 , n2522  );
buf ( g2522 , n2523  );
buf ( g2523 , n2524  );
buf ( g2524 , n2525  );
buf ( g2525 , n2526  );
buf ( g2526 , n2527  );
buf ( g2527 , n2528  );
buf ( g2528 , n2529  );
buf ( g2529 , n2530  );
buf ( g2530 , n2531  );
buf ( g2531 , n2532  );
buf ( g2532 , n2533  );
buf ( g2533 , n2534  );
buf ( g2534 , n2535  );
buf ( g2535 , n2536  );
buf ( g2536 , n2537  );
buf ( g2537 , n2538  );
buf ( g2538 , n2539  );
buf ( g2539 , n2540  );
buf ( g2540 , n2541  );
buf ( g2541 , n2542  );
buf ( g2542 , n2543  );
buf ( g2543 , n2544  );
buf ( g2544 , n2545  );
buf ( g2545 , n2546  );
buf ( g2546 , n2547  );
buf ( g2547 , n2548  );
buf ( g2548 , n2549  );
buf ( g2549 , n2550  );
buf ( g2550 , n2551  );
buf ( g2551 , n2552  );
buf ( g2552 , n2553  );
buf ( g2553 , n2554  );
buf ( g2554 , n2555  );
buf ( g2555 , n2556  );
buf ( g2556 , n2557  );
buf ( g2557 , n2558  );
buf ( g2558 , n2559  );
buf ( g2559 , n2560  );
buf ( g2560 , n2561  );
buf ( g2561 , n2562  );
buf ( g2562 , n2563  );
buf ( g2563 , n2564  );
buf ( g2564 , n2565  );
buf ( g2565 , n2566  );
buf ( g2566 , n2567  );
buf ( g2567 , n2568  );
buf ( g2568 , n2569  );
buf ( g2569 , n2570  );
buf ( g2570 , n2571  );
buf ( g2571 , n2572  );
buf ( g2572 , n2573  );
buf ( g2573 , n2574  );
buf ( g2574 , n2575  );
buf ( g2575 , n2576  );
buf ( g2576 , n2577  );
buf ( g2577 , n2578  );
buf ( g2578 , n2579  );
buf ( g2579 , n2580  );
buf ( g2580 , n2581  );
buf ( g2581 , n2582  );
buf ( g2582 , n2583  );
buf ( g2583 , n2584  );
buf ( g2584 , n2585  );
buf ( g2585 , n2586  );
buf ( g2586 , n2587  );
buf ( g2587 , n2588  );
buf ( g2588 , n2589  );
buf ( g2589 , n2590  );
buf ( g2590 , n2591  );
buf ( g2591 , n2592  );
buf ( g2592 , n2593  );
buf ( g2593 , n2594  );
buf ( g2594 , n2595  );
buf ( g2595 , n2596  );
buf ( g2596 , n2597  );
buf ( g2597 , n2598  );
buf ( g2598 , n2599  );
buf ( g2599 , n2600  );
buf ( g2600 , n2601  );
buf ( g2601 , n2602  );
buf ( g2602 , n2603  );
buf ( g2603 , n2604  );
buf ( g2604 , n2605  );
buf ( g2605 , n2606  );
buf ( g2606 , n2607  );
buf ( g2607 , n2608  );
buf ( g2608 , n2609  );
buf ( g2609 , n2610  );
buf ( g2610 , n2611  );
buf ( g2611 , n2612  );
buf ( g2612 , n2613  );
buf ( g2613 , n2614  );
buf ( g2614 , n2615  );
buf ( g2615 , n2616  );
buf ( g2616 , n2617  );
buf ( g2617 , n2618  );
buf ( g2618 , n2619  );
buf ( g2619 , n2620  );
buf ( g2620 , n2621  );
buf ( g2621 , n2622  );
buf ( g2622 , n2623  );
buf ( g2623 , n2624  );
buf ( g2624 , n2625  );
buf ( g2625 , n2626  );
buf ( g2626 , n2627  );
buf ( g2627 , n2628  );
buf ( g2628 , n2629  );
buf ( g2629 , n2630  );
buf ( g2630 , n2631  );
buf ( g2631 , n2632  );
buf ( g2632 , n2633  );
buf ( g2633 , n2634  );
buf ( g2634 , n2635  );
buf ( g2635 , n2636  );
buf ( g2636 , n2637  );
buf ( g2637 , n2638  );
buf ( g2638 , n2639  );
buf ( g2639 , n2640  );
buf ( g2640 , n2641  );
buf ( g2641 , n2642  );
buf ( g2642 , n2643  );
buf ( g2643 , n2644  );
buf ( g2644 , n2645  );
buf ( g2645 , n2646  );
buf ( g2646 , n2647  );
buf ( g2647 , n2648  );
buf ( g2648 , n2649  );
buf ( g2649 , n2650  );
buf ( g2650 , n2651  );
buf ( g2651 , n2652  );
buf ( g2652 , n2653  );
buf ( g2653 , n2654  );
buf ( g2654 , n2655  );
buf ( g2655 , n2656  );
buf ( g2656 , n2657  );
buf ( g2657 , n2658  );
buf ( g2658 , n2659  );
buf ( g2659 , n2660  );
buf ( g2660 , n2661  );
buf ( g2661 , n2662  );
buf ( g2662 , n2663  );
buf ( g2663 , n2664  );
buf ( g2664 , n2665  );
buf ( g2665 , n2666  );
buf ( g2666 , n2667  );
buf ( g2667 , n2668  );
buf ( g2668 , n2669  );
buf ( g2669 , n2670  );
buf ( g2670 , n2671  );
buf ( g2671 , n2672  );
buf ( g2672 , n2673  );
buf ( g2673 , n2674  );
buf ( g2674 , n2675  );
buf ( g2675 , n2676  );
buf ( g2676 , n2677  );
buf ( g2677 , n2678  );
buf ( g2678 , n2679  );
buf ( g2679 , n2680  );
buf ( g2680 , n2681  );
buf ( g2681 , n2682  );
buf ( g2682 , n2683  );
buf ( g2683 , n2684  );
buf ( g2684 , n2685  );
buf ( g2685 , n2686  );
buf ( g2686 , n2687  );
buf ( g2687 , n2688  );
buf ( g2688 , n2689  );
buf ( g2689 , n2690  );
buf ( g2690 , n2691  );
buf ( g2691 , n2692  );
buf ( g2692 , n2693  );
buf ( g2693 , n2694  );
buf ( g2694 , n2695  );
buf ( g2695 , n2696  );
buf ( g2696 , n2697  );
buf ( g2697 , n2698  );
buf ( g2698 , n2699  );
buf ( g2699 , n2700  );
buf ( g2700 , n2701  );
buf ( g2701 , n2702  );
buf ( g2702 , n2703  );
buf ( g2703 , n2704  );
buf ( g2704 , n2705  );
buf ( g2705 , n2706  );
buf ( g2706 , n2707  );
buf ( g2707 , n2708  );
buf ( g2708 , n2709  );
buf ( g2709 , n2710  );
buf ( g2710 , n2711  );
buf ( g2711 , n2712  );
buf ( g2712 , n2713  );
buf ( g2713 , n2714  );
buf ( g2714 , n2715  );
buf ( g2715 , n2716  );
buf ( g2716 , n2717  );
buf ( g2717 , n2718  );
buf ( g2718 , n2719  );
buf ( g2719 , n2720  );
buf ( g2720 , n2721  );
buf ( g2721 , n2722  );
buf ( g2722 , n2723  );
buf ( g2723 , n2724  );
buf ( g2724 , n2725  );
buf ( g2725 , n2726  );
buf ( g2726 , n2727  );
buf ( g2727 , n2728  );
buf ( g2728 , n2729  );
buf ( g2729 , n2730  );
buf ( g2730 , n2731  );
buf ( g2731 , n2732  );
buf ( g2732 , n2733  );
buf ( g2733 , n2734  );
buf ( g2734 , n2735  );
buf ( g2735 , n2736  );
buf ( g2736 , n2737  );
buf ( g2737 , n2738  );
buf ( g2738 , n2739  );
buf ( g2739 , n2740  );
buf ( g2740 , n2741  );
buf ( g2741 , n2742  );
buf ( g2742 , n2743  );
buf ( g2743 , n2744  );
buf ( g2744 , n2745  );
buf ( g2745 , n2746  );
buf ( g2746 , n2747  );
buf ( g2747 , n2748  );
buf ( g2748 , n2749  );
buf ( g2749 , n2750  );
buf ( g2750 , n2751  );
buf ( g2751 , n2752  );
buf ( g2752 , n2753  );
buf ( g2753 , n2754  );
buf ( g2754 , n2755  );
buf ( g2755 , n2756  );
buf ( g2756 , n2757  );
buf ( g2757 , n2758  );
buf ( g2758 , n2759  );
buf ( g2759 , n2760  );
buf ( g2760 , n2761  );
buf ( g2761 , n2762  );
buf ( g2762 , n2763  );
buf ( g2763 , n2764  );
buf ( g2764 , n2765  );
buf ( g2765 , n2766  );
buf ( g2766 , n2767  );
buf ( g2767 , n2768  );
buf ( g2768 , n2769  );
buf ( g2769 , n2770  );
buf ( g2770 , n2771  );
buf ( g2771 , n2772  );
buf ( g2772 , n2773  );
buf ( g2773 , n2774  );
buf ( g2774 , n2775  );
buf ( g2775 , n2776  );
buf ( g2776 , n2777  );
buf ( g2777 , n2778  );
buf ( g2778 , n2779  );
buf ( g2779 , n2780  );
buf ( g2780 , n2781  );
buf ( g2781 , n2782  );
buf ( g2782 , n2783  );
buf ( g2783 , n2784  );
buf ( g2784 , n2785  );
buf ( g2785 , n2786  );
buf ( g2786 , n2787  );
buf ( g2787 , n2788  );
buf ( g2788 , n2789  );
buf ( g2789 , n2790  );
buf ( g2790 , n2791  );
buf ( g2791 , n2792  );
buf ( g2792 , n2793  );
buf ( g2793 , n2794  );
buf ( g2794 , n2795  );
buf ( g2795 , n2796  );
buf ( g2796 , n2797  );
buf ( g2797 , n2798  );
buf ( g2798 , n2799  );
buf ( g2799 , n2800  );
buf ( g2800 , n2801  );
buf ( g2801 , n2802  );
buf ( g2802 , n2803  );
buf ( g2803 , n2804  );
buf ( g2804 , n2805  );
buf ( g2805 , n2806  );
buf ( g2806 , n2807  );
buf ( g2807 , n2808  );
buf ( g2808 , n2809  );
buf ( g2809 , n2810  );
buf ( g2810 , n2811  );
buf ( g2811 , n2812  );
buf ( g2812 , n2813  );
buf ( g2813 , n2814  );
buf ( g2814 , n2815  );
buf ( g2815 , n2816  );
buf ( g2816 , n2817  );
buf ( g2817 , n2818  );
buf ( g2818 , n2819  );
buf ( g2819 , n2820  );
buf ( g2820 , n2821  );
buf ( g2821 , n2822  );
buf ( g2822 , n2823  );
buf ( g2823 , n2824  );
buf ( g2824 , n2825  );
buf ( g2825 , n2826  );
buf ( g2826 , n2827  );
buf ( g2827 , n2828  );
buf ( g2828 , n2829  );
buf ( g2829 , n2830  );
buf ( g2830 , n2831  );
buf ( g2831 , n2832  );
buf ( g2832 , n2833  );
buf ( g2833 , n2834  );
buf ( g2834 , n2835  );
buf ( g2835 , n2836  );
buf ( g2836 , n2837  );
buf ( g2837 , n2838  );
buf ( g2838 , n2839  );
buf ( g2839 , n2840  );
buf ( g2840 , n2841  );
buf ( g2841 , n2842  );
buf ( g2842 , n2843  );
buf ( g2843 , n2844  );
buf ( g2844 , n2845  );
buf ( g2845 , n2846  );
buf ( g2846 , n2847  );
buf ( g2847 , n2848  );
buf ( g2848 , n2849  );
buf ( g2849 , n2850  );
buf ( g2850 , n2851  );
buf ( g2851 , n2852  );
buf ( g2852 , n2853  );
buf ( g2853 , n2854  );
buf ( g2854 , n2855  );
buf ( g2855 , n2856  );
buf ( g2856 , n2857  );
buf ( g2857 , n2858  );
buf ( g2858 , n2859  );
buf ( g2859 , n2860  );
buf ( g2860 , n2861  );
buf ( g2861 , n2862  );
buf ( g2862 , n2863  );
buf ( g2863 , n2864  );
buf ( g2864 , n2865  );
buf ( g2865 , n2866  );
buf ( g2866 , n2867  );
buf ( g2867 , n2868  );
buf ( g2868 , n2869  );
buf ( g2869 , n2870  );
buf ( g2870 , n2871  );
buf ( g2871 , n2872  );
buf ( g2872 , n2873  );
buf ( g2873 , n2874  );
buf ( g2874 , n2875  );
buf ( g2875 , n2876  );
buf ( g2876 , n2877  );
buf ( g2877 , n2878  );
buf ( g2878 , n2879  );
buf ( g2879 , n2880  );
buf ( g2880 , n2881  );
buf ( g2881 , n2882  );
buf ( g2882 , n2883  );
buf ( g2883 , n2884  );
buf ( g2884 , n2885  );
buf ( g2885 , n2886  );
buf ( g2886 , n2887  );
buf ( g2887 , n2888  );
buf ( g2888 , n2889  );
buf ( g2889 , n2890  );
buf ( g2890 , n2891  );
buf ( g2891 , n2892  );
buf ( g2892 , n2893  );
buf ( g2893 , n2894  );
buf ( g2894 , n2895  );
buf ( g2895 , n2896  );
buf ( g2896 , n2897  );
buf ( g2897 , n2898  );
buf ( g2898 , n2899  );
buf ( g2899 , n2900  );
buf ( g2900 , n2901  );
buf ( g2901 , n2902  );
buf ( g2902 , n2903  );
buf ( g2903 , n2904  );
buf ( g2904 , n2905  );
buf ( g2905 , n2906  );
buf ( g2906 , n2907  );
buf ( g2907 , n2908  );
buf ( g2908 , n2909  );
buf ( g2909 , n2910  );
buf ( g2910 , n2911  );
buf ( g2911 , n2912  );
buf ( g2912 , n2913  );
buf ( g2913 , n2914  );
buf ( g2914 , n2915  );
buf ( g2915 , n2916  );
buf ( g2916 , n2917  );
buf ( g2917 , n2918  );
buf ( g2918 , n2919  );
buf ( g2919 , n2920  );
buf ( g2920 , n2921  );
buf ( g2921 , n2922  );
buf ( g2922 , n2923  );
buf ( g2923 , n2924  );
buf ( g2924 , n2925  );
buf ( g2925 , n2926  );
buf ( g2926 , n2927  );
buf ( g2927 , n2928  );
buf ( g2928 , n2929  );
buf ( g2929 , n2930  );
buf ( g2930 , n2931  );
buf ( g2931 , n2932  );
buf ( g2932 , n2933  );
buf ( g2933 , n2934  );
buf ( g2934 , n2935  );
buf ( g2935 , n2936  );
buf ( g2936 , n2937  );
buf ( g2937 , n2938  );
buf ( g2938 , n2939  );
buf ( g2939 , n2940  );
buf ( g2940 , n2941  );
buf ( g2941 , n2942  );
buf ( g2942 , n2943  );
buf ( g2943 , n2944  );
buf ( g2944 , n2945  );
buf ( g2945 , n2946  );
buf ( g2946 , n2947  );
buf ( g2947 , n2948  );
buf ( g2948 , n2949  );
buf ( g2949 , n2950  );
buf ( g2950 , n2951  );
buf ( g2951 , n2952  );
buf ( g2952 , n2953  );
buf ( g2953 , n2954  );
buf ( g2954 , n2955  );
buf ( g2955 , n2956  );
buf ( g2956 , n2957  );
buf ( g2957 , n2958  );
buf ( g2958 , n2959  );
buf ( g2959 , n2960  );
buf ( g2960 , n2961  );
buf ( g2961 , n2962  );
buf ( g2962 , n2963  );
buf ( g2963 , n2964  );
buf ( g2964 , n2965  );
buf ( g2965 , n2966  );
buf ( g2966 , n2967  );
buf ( g2967 , n2968  );
buf ( g2968 , n2969  );
buf ( g2969 , n2970  );
buf ( g2970 , n2971  );
buf ( g2971 , n2972  );
buf ( g2972 , n2973  );
buf ( g2973 , n2974  );
buf ( g2974 , n2975  );
buf ( g2975 , n2976  );
buf ( g2976 , n2977  );
buf ( g2977 , n2978  );
buf ( g2978 , n2979  );
buf ( g2979 , n2980  );
buf ( g2980 , n2981  );
buf ( g2981 , n2982  );
buf ( g2982 , n2983  );
buf ( g2983 , n2984  );
buf ( g2984 , n2985  );
buf ( g2985 , n2986  );
buf ( g2986 , n2987  );
buf ( g2987 , n2988  );
buf ( g2988 , n2989  );
buf ( g2989 , n2990  );
buf ( g2990 , n2991  );
buf ( g2991 , n2992  );
buf ( g2992 , n2993  );
buf ( g2993 , n2994  );
buf ( g2994 , n2995  );
buf ( g2995 , n2996  );
buf ( g2996 , n2997  );
buf ( g2997 , n2998  );
buf ( g2998 , n2999  );
buf ( g2999 , n3000  );
buf ( g3000 , n3001  );
buf ( g3001 , n3002  );
buf ( g3002 , n3003  );
buf ( g3003 , n3004  );
buf ( g3004 , n3005  );
buf ( g3005 , n3006  );
buf ( g3006 , n3007  );
buf ( g3007 , n3008  );
buf ( g3008 , n3009  );
buf ( g3009 , n3010  );
buf ( g3010 , n3011  );
buf ( g3011 , n3012  );
buf ( g3012 , n3013  );
buf ( g3013 , n3014  );
buf ( g3014 , n3015  );
buf ( g3015 , n3016  );
buf ( g3016 , n3017  );
buf ( g3017 , n3018  );
buf ( g3018 , n3019  );
buf ( g3019 , n3020  );
buf ( g3020 , n3021  );
buf ( g3021 , n3022  );
buf ( g3022 , n3023  );
buf ( g3023 , n3024  );
buf ( g3024 , n3025  );
buf ( g3025 , n3026  );
buf ( g3026 , n3027  );
buf ( g3027 , n3028  );
buf ( g3028 , n3029  );
buf ( g3029 , n3030  );
buf ( g3030 , n3031  );
buf ( g3031 , n3032  );
buf ( g3032 , n3033  );
buf ( g3033 , n3034  );
buf ( g3034 , n3035  );
buf ( g3035 , n3036  );
buf ( g3036 , n3037  );
buf ( g3037 , n3038  );
buf ( g3038 , n3039  );
buf ( g3039 , n3040  );
buf ( g3040 , n3041  );
buf ( g3041 , n3042  );
buf ( g3042 , n3043  );
buf ( g3043 , n3044  );
buf ( g3044 , n3045  );
buf ( g3045 , n3046  );
buf ( g3046 , n3047  );
buf ( g3047 , n3048  );
buf ( g3048 , n3049  );
buf ( g3049 , n3050  );
buf ( g3050 , n3051  );
buf ( g3051 , n3052  );
buf ( g3052 , n3053  );
buf ( g3053 , n3054  );
buf ( g3054 , n3055  );
buf ( g3055 , n3056  );
buf ( g3056 , n3057  );
buf ( g3057 , n3058  );
buf ( g3058 , n3059  );
buf ( g3059 , n3060  );
buf ( g3060 , n3061  );
buf ( g3061 , n3062  );
buf ( g3062 , n3063  );
buf ( g3063 , n3064  );
buf ( g3064 , n3065  );
buf ( g3065 , n3066  );
buf ( g3066 , n3067  );
buf ( g3067 , n3068  );
buf ( g3068 , n3069  );
buf ( g3069 , n3070  );
buf ( g3070 , n3071  );
buf ( g3071 , n3072  );
buf ( g3072 , n3073  );
buf ( g3073 , n3074  );
buf ( g3074 , n3075  );
buf ( g3075 , n3076  );
buf ( g3076 , n3077  );
buf ( g3077 , n3078  );
buf ( g3078 , n3079  );
buf ( g3079 , n3080  );
buf ( g3080 , n3081  );
buf ( g3081 , n3082  );
buf ( g3082 , n3083  );
buf ( g3083 , n3084  );
buf ( g3084 , n3085  );
buf ( g3085 , n3086  );
buf ( g3086 , n3087  );
buf ( g3087 , n3088  );
buf ( g3088 , n3089  );
buf ( g3089 , n3090  );
buf ( g3090 , n3091  );
buf ( g3091 , n3092  );
buf ( g3092 , n3093  );
buf ( g3093 , n3094  );
buf ( g3094 , n3095  );
buf ( g3095 , n3096  );
buf ( g3096 , n3097  );
buf ( g3097 , n3098  );
buf ( g3098 , n3099  );
buf ( g3099 , n3100  );
buf ( g3100 , n3101  );
buf ( g3101 , n3102  );
buf ( g3102 , n3103  );
buf ( g3103 , n3104  );
buf ( g3104 , n3105  );
buf ( g3105 , n3106  );
buf ( g3106 , n3107  );
buf ( g3107 , n3108  );
buf ( g3108 , n3109  );
buf ( g3109 , n3110  );
buf ( g3110 , n3111  );
buf ( g3111 , n3112  );
buf ( g3112 , n3113  );
buf ( g3113 , n3114  );
buf ( g3114 , n3115  );
buf ( g3115 , n3116  );
buf ( g3116 , n3117  );
buf ( g3117 , n3118  );
buf ( g3118 , n3119  );
buf ( g3119 , n3120  );
buf ( g3120 , n3121  );
buf ( g3121 , n3122  );
buf ( g3122 , n3123  );
buf ( g3123 , n3124  );
buf ( g3124 , n3125  );
buf ( g3125 , n3126  );
buf ( g3126 , n3127  );
buf ( g3127 , n3128  );
buf ( g3128 , n3129  );
buf ( g3129 , n3130  );
buf ( g3130 , n3131  );
buf ( g3131 , n3132  );
buf ( g3132 , n3133  );
buf ( g3133 , n3134  );
buf ( g3134 , n3135  );
buf ( g3135 , n3136  );
buf ( g3136 , n3137  );
buf ( g3137 , n3138  );
buf ( g3138 , n3139  );
buf ( g3139 , n3140  );
buf ( g3140 , n3141  );
buf ( g3141 , n3142  );
buf ( g3142 , n3143  );
buf ( g3143 , n3144  );
buf ( g3144 , n3145  );
buf ( g3145 , n3146  );
buf ( g3146 , n3147  );
buf ( g3147 , n3148  );
buf ( g3148 , n3149  );
buf ( g3149 , n3150  );
buf ( g3150 , n3151  );
buf ( g3151 , n3152  );
buf ( g3152 , n3153  );
buf ( g3153 , n3154  );
buf ( g3154 , n3155  );
buf ( g3155 , n3156  );
buf ( g3156 , n3157  );
buf ( g3157 , n3158  );
buf ( g3158 , n3159  );
buf ( g3159 , n3160  );
buf ( g3160 , n3161  );
buf ( g3161 , n3162  );
buf ( g3162 , n3163  );
buf ( g3163 , n3164  );
buf ( g3164 , n3165  );
buf ( g3165 , n3166  );
buf ( g3166 , n3167  );
buf ( g3167 , n3168  );
buf ( g3168 , n3169  );
buf ( g3169 , n3170  );
buf ( g3170 , n3171  );
buf ( g3171 , n3172  );
buf ( g3172 , n3173  );
buf ( g3173 , n3174  );
buf ( g3174 , n3175  );
buf ( g3175 , n3176  );
buf ( g3176 , n3177  );
buf ( g3177 , n3178  );
buf ( g3178 , n3179  );
buf ( g3179 , n3180  );
buf ( g3180 , n3181  );
buf ( g3181 , n3182  );
buf ( g3182 , n3183  );
buf ( g3183 , n3184  );
buf ( g3184 , n3185  );
buf ( g3185 , n3186  );
buf ( g3186 , n3187  );
buf ( g3187 , n3188  );
buf ( g3188 , n3189  );
buf ( g3189 , n3190  );
buf ( g3190 , n3191  );
buf ( g3191 , n3192  );
buf ( g3192 , n3193  );
buf ( g3193 , n3194  );
buf ( g3194 , n3195  );
buf ( g3195 , n3196  );
buf ( g3196 , n3197  );
buf ( g3197 , n3198  );
buf ( g3198 , n3199  );
buf ( g3199 , n3200  );
buf ( g3200 , n3201  );
buf ( g3201 , n3202  );
buf ( g3202 , n3203  );
buf ( g3203 , n3204  );
buf ( g3204 , n3205  );
buf ( g3205 , n3206  );
buf ( g3206 , n3207  );
buf ( g3207 , n3208  );
buf ( g3208 , n3209  );
buf ( g3209 , n3210  );
buf ( g3210 , n3211  );
buf ( g3211 , n3212  );
buf ( g3212 , n3213  );
buf ( g3213 , n3214  );
buf ( g3214 , n3215  );
buf ( g3215 , n3216  );
buf ( g3216 , n3217  );
buf ( g3217 , n3218  );
buf ( g3218 , n3219  );
buf ( g3219 , n3220  );
buf ( g3220 , n3221  );
buf ( g3221 , n3222  );
buf ( g3222 , n3223  );
buf ( g3223 , n3224  );
buf ( g3224 , n3225  );
buf ( g3225 , n3226  );
buf ( g3226 , n3227  );
buf ( g3227 , n3228  );
buf ( g3228 , n3229  );
buf ( g3229 , n3230  );
buf ( g3230 , n3231  );
buf ( g3231 , n3232  );
buf ( g3232 , n3233  );
buf ( g3233 , n3234  );
buf ( g3234 , n3235  );
buf ( g3235 , n3236  );
buf ( g3236 , n3237  );
buf ( g3237 , n3238  );
buf ( g3238 , n3239  );
buf ( g3239 , n3240  );
buf ( g3240 , n3241  );
buf ( g3241 , n3242  );
buf ( g3242 , n3243  );
buf ( g3243 , n3244  );
buf ( g3244 , n3245  );
buf ( g3245 , n3246  );
buf ( g3246 , n3247  );
buf ( g3247 , n3248  );
buf ( g3248 , n3249  );
buf ( g3249 , n3250  );
buf ( g3250 , n3251  );
buf ( g3251 , n3252  );
buf ( g3252 , n3253  );
buf ( g3253 , n3254  );
buf ( g3254 , n3255  );
buf ( g3255 , n3256  );
buf ( g3256 , n3257  );
buf ( g3257 , n3258  );
buf ( g3258 , n3259  );
buf ( g3259 , n3260  );
buf ( g3260 , n3261  );
buf ( g3261 , n3262  );
buf ( g3262 , n3263  );
buf ( g3263 , n3264  );
buf ( g3264 , n3265  );
buf ( g3265 , n3266  );
buf ( g3266 , n3267  );
buf ( g3267 , n3268  );
buf ( g3268 , n3269  );
buf ( g3269 , n3270  );
buf ( g3270 , n3271  );
buf ( g3271 , n3272  );
buf ( g3272 , n3273  );
buf ( g3273 , n3274  );
buf ( g3274 , n3275  );
buf ( g3275 , n3276  );
buf ( g3276 , n3277  );
buf ( g3277 , n3278  );
buf ( g3278 , n3279  );
buf ( g3279 , n3280  );
buf ( g3280 , n3281  );
buf ( g3281 , n3282  );
buf ( g3282 , n3283  );
buf ( g3283 , n3284  );
buf ( g3284 , n3285  );
buf ( g3285 , n3286  );
buf ( g3286 , n3287  );
buf ( g3287 , n3288  );
buf ( g3288 , n3289  );
buf ( g3289 , n3290  );
buf ( g3290 , n3291  );
buf ( g3291 , n3292  );
buf ( g3292 , n3293  );
buf ( g3293 , n3294  );
buf ( g3294 , n3295  );
buf ( g3295 , n3296  );
buf ( g3296 , n3297  );
buf ( g3297 , n3298  );
buf ( g3298 , n3299  );
buf ( g3299 , n3300  );
buf ( g3300 , n3301  );
buf ( g3301 , n3302  );
buf ( g3302 , n3303  );
buf ( g3303 , n3304  );
buf ( g3304 , n3305  );
buf ( g3305 , n3306  );
buf ( g3306 , n3307  );
buf ( g3307 , n3308  );
buf ( g3308 , n3309  );
buf ( g3309 , n3310  );
buf ( g3310 , n3311  );
buf ( g3311 , n3312  );
buf ( g3312 , n3313  );
buf ( g3313 , n3314  );
buf ( g3314 , n3315  );
buf ( g3315 , n3316  );
buf ( g3316 , n3317  );
buf ( g3317 , n3318  );
buf ( g3318 , n3319  );
buf ( g3319 , n3320  );
buf ( g3320 , n3321  );
buf ( g3321 , n3322  );
buf ( g3322 , n3323  );
buf ( g3323 , n3324  );
buf ( g3324 , n3325  );
buf ( g3325 , n3326  );
buf ( g3326 , n3327  );
buf ( g3327 , n3328  );
buf ( g3328 , n3329  );
buf ( g3329 , n3330  );
buf ( g3330 , n3331  );
buf ( g3331 , n3332  );
buf ( g3332 , n3333  );
buf ( g3333 , n3334  );
buf ( g3334 , n3335  );
buf ( g3335 , n3336  );
buf ( g3336 , n3337  );
buf ( g3337 , n3338  );
buf ( g3338 , n3339  );
buf ( g3339 , n3340  );
buf ( g3340 , n3341  );
buf ( g3341 , n3342  );
buf ( g3342 , n3343  );
buf ( g3343 , n3344  );
buf ( g3344 , n3345  );
buf ( g3345 , n3346  );
buf ( g3346 , n3347  );
buf ( g3347 , n3348  );
buf ( g3348 , n3349  );
buf ( g3349 , n3350  );
buf ( g3350 , n3351  );
buf ( g3351 , n3352  );
buf ( g3352 , n3353  );
buf ( g3353 , n3354  );
buf ( g3354 , n3355  );
buf ( g3355 , n3356  );
buf ( g3356 , n3357  );
buf ( g3357 , n3358  );
buf ( g3358 , n3359  );
buf ( g3359 , n3360  );
buf ( g3360 , n3361  );
buf ( g3361 , n3362  );
buf ( g3362 , n3363  );
buf ( g3363 , n3364  );
buf ( g3364 , n3365  );
buf ( g3365 , n3366  );
buf ( g3366 , n3367  );
buf ( g3367 , n3368  );
buf ( g3368 , n3369  );
buf ( g3369 , n3370  );
buf ( g3370 , n3371  );
buf ( g3371 , n3372  );
buf ( g3372 , n3373  );
buf ( g3373 , n3374  );
buf ( g3374 , n3375  );
buf ( g3375 , n3376  );
buf ( g3376 , n3377  );
buf ( g3377 , n3378  );
buf ( g3378 , n3379  );
buf ( g3379 , n3380  );
buf ( g3380 , n3381  );
buf ( g3381 , n3382  );
buf ( g3382 , n3383  );
buf ( g3383 , n3384  );
buf ( g3384 , n3385  );
buf ( g3385 , n3386  );
buf ( g3386 , n3387  );
buf ( g3387 , n3388  );
buf ( g3388 , n3389  );
buf ( g3389 , n3390  );
buf ( g3390 , n3391  );
buf ( g3391 , n3392  );
buf ( g3392 , n3393  );
buf ( g3393 , n3394  );
buf ( g3394 , n3395  );
buf ( g3395 , n3396  );
buf ( g3396 , n3397  );
buf ( g3397 , n3398  );
buf ( g3398 , n3399  );
buf ( g3399 , n3400  );
buf ( g3400 , n3401  );
buf ( g3401 , n3402  );
buf ( g3402 , n3403  );
buf ( g3403 , n3404  );
buf ( g3404 , n3405  );
buf ( g3405 , n3406  );
buf ( g3406 , n3407  );
buf ( g3407 , n3408  );
buf ( g3408 , n3409  );
buf ( g3409 , n3410  );
buf ( g3410 , n3411  );
buf ( g3411 , n3412  );
buf ( g3412 , n3413  );
buf ( g3413 , n3414  );
buf ( g3414 , n3415  );
buf ( g3415 , n3416  );
buf ( g3416 , n3417  );
buf ( g3417 , n3418  );
buf ( g3418 , n3419  );
buf ( g3419 , n3420  );
buf ( g3420 , n3421  );
buf ( g3421 , n3422  );
buf ( g3422 , n3423  );
buf ( g3423 , n3424  );
buf ( g3424 , n3425  );
buf ( g3425 , n3426  );
buf ( g3426 , n3427  );
buf ( g3427 , n3428  );
buf ( g3428 , n3429  );
buf ( g3429 , n3430  );
buf ( g3430 , n3431  );
buf ( g3431 , n3432  );
buf ( g3432 , n3433  );
buf ( g3433 , n3434  );
buf ( g3434 , n3435  );
buf ( g3435 , n3436  );
buf ( g3436 , n3437  );
buf ( g3437 , n3438  );
buf ( g3438 , n3439  );
buf ( g3439 , n3440  );
buf ( g3440 , n3441  );
buf ( g3441 , n3442  );
buf ( g3442 , n3443  );
buf ( g3443 , n3444  );
buf ( g3444 , n3445  );
buf ( g3445 , n3446  );
buf ( g3446 , n3447  );
buf ( g3447 , n3448  );
buf ( g3448 , n3449  );
buf ( g3449 , n3450  );
buf ( g3450 , n3451  );
buf ( g3451 , n3452  );
buf ( g3452 , n3453  );
buf ( g3453 , n3454  );
buf ( g3454 , n3455  );
buf ( g3455 , n3456  );
buf ( g3456 , n3457  );
buf ( g3457 , n3458  );
buf ( g3458 , n3459  );
buf ( g3459 , n3460  );
buf ( g3460 , n3461  );
buf ( g3461 , n3462  );
buf ( g3462 , n3463  );
buf ( g3463 , n3464  );
buf ( g3464 , n3465  );
buf ( g3465 , n3466  );
buf ( g3466 , n3467  );
buf ( g3467 , n3468  );
buf ( g3468 , n3469  );
buf ( g3469 , n3470  );
buf ( g3470 , n3471  );
buf ( g3471 , n3472  );
buf ( g3472 , n3473  );
buf ( g3473 , n3474  );
buf ( g3474 , n3475  );
buf ( g3475 , n3476  );
buf ( g3476 , n3477  );
buf ( g3477 , n3478  );
buf ( g3478 , n3479  );
buf ( g3479 , n3480  );
buf ( g3480 , n3481  );
buf ( g3481 , n3482  );
buf ( g3482 , n3483  );
buf ( g3483 , n3484  );
buf ( g3484 , n3485  );
buf ( g3485 , n3486  );
buf ( g3486 , n3487  );
buf ( g3487 , n3488  );
buf ( g3488 , n3489  );
buf ( g3489 , n3490  );
buf ( g3490 , n3491  );
buf ( g3491 , n3492  );
buf ( g3492 , n3493  );
buf ( g3493 , n3494  );
buf ( g3494 , n3495  );
buf ( g3495 , n3496  );
buf ( g3496 , n3497  );
buf ( g3497 , n3498  );
buf ( g3498 , n3499  );
buf ( g3499 , n3500  );
buf ( g3500 , n3501  );
buf ( g3501 , n3502  );
buf ( g3502 , n3503  );
buf ( g3503 , n3504  );
buf ( g3504 , n3505  );
buf ( g3505 , n3506  );
buf ( g3506 , n3507  );
buf ( g3507 , n3508  );
buf ( g3508 , n3509  );
buf ( g3509 , n3510  );
buf ( g3510 , n3511  );
buf ( g3511 , n3512  );
buf ( g3512 , n3513  );
buf ( g3513 , n3514  );
buf ( g3514 , n3515  );
buf ( g3515 , n3516  );
buf ( g3516 , n3517  );
buf ( g3517 , n3518  );
buf ( g3518 , n3519  );
buf ( g3519 , n3520  );
buf ( g3520 , n3521  );
buf ( g3521 , n3522  );
buf ( g3522 , n3523  );
buf ( g3523 , n3524  );
buf ( g3524 , n3525  );
buf ( g3525 , n3526  );
buf ( g3526 , n3527  );
buf ( g3527 , n3528  );
buf ( g3528 , n3529  );
buf ( g3529 , n3530  );
buf ( g3530 , n3531  );
buf ( g3531 , n3532  );
buf ( g3532 , n3533  );
buf ( g3533 , n3534  );
buf ( g3534 , n3535  );
buf ( g3535 , n3536  );
buf ( g3536 , n3537  );
buf ( g3537 , n3538  );
buf ( g3538 , n3539  );
buf ( g3539 , n3540  );
buf ( g3540 , n3541  );
buf ( g3541 , n3542  );
buf ( g3542 , n3543  );
buf ( g3543 , n3544  );
buf ( g3544 , n3545  );
buf ( g3545 , n3546  );
buf ( g3546 , n3547  );
buf ( g3547 , n3548  );
buf ( g3548 , n3549  );
buf ( g3549 , n3550  );
buf ( g3550 , n3551  );
buf ( g3551 , n3552  );
buf ( g3552 , n3553  );
buf ( g3553 , n3554  );
buf ( g3554 , n3555  );
buf ( g3555 , n3556  );
buf ( g3556 , n3557  );
buf ( g3557 , n3558  );
buf ( g3558 , n3559  );
buf ( g3559 , n3560  );
buf ( g3560 , n3561  );
buf ( g3561 , n3562  );
buf ( g3562 , n3563  );
buf ( g3563 , n3564  );
buf ( g3564 , n3565  );
buf ( g3565 , n3566  );
buf ( g3566 , n3567  );
buf ( g3567 , n3568  );
buf ( g3568 , n3569  );
buf ( g3569 , n3570  );
buf ( g3570 , n3571  );
buf ( g3571 , n3572  );
buf ( g3572 , n3573  );
buf ( g3573 , n3574  );
buf ( g3574 , n3575  );
buf ( g3575 , n3576  );
buf ( g3576 , n3577  );
buf ( g3577 , n3578  );
buf ( g3578 , n3579  );
buf ( g3579 , n3580  );
buf ( g3580 , n3581  );
buf ( g3581 , n3582  );
buf ( g3582 , n3583  );
buf ( g3583 , n3584  );
buf ( g3584 , n3585  );
buf ( g3585 , n3586  );
buf ( g3586 , n3587  );
buf ( g3587 , n3588  );
buf ( g3588 , n3589  );
buf ( g3589 , n3590  );
buf ( g3590 , n3591  );
buf ( g3591 , n3592  );
buf ( g3592 , n3593  );
buf ( g3593 , n3594  );
buf ( g3594 , n3595  );
buf ( g3595 , n3596  );
buf ( g3596 , n3597  );
buf ( g3597 , n3598  );
buf ( g3598 , n3599  );
buf ( g3599 , n3600  );
buf ( g3600 , n3601  );
buf ( g3601 , n3602  );
buf ( g3602 , n3603  );
buf ( g3603 , n3604  );
buf ( g3604 , n3605  );
buf ( g3605 , n3606  );
buf ( g3606 , n3607  );
buf ( g3607 , n3608  );
buf ( g3608 , n3609  );
buf ( g3609 , n3610  );
buf ( g3610 , n3611  );
buf ( g3611 , n3612  );
buf ( g3612 , n3613  );
buf ( g3613 , n3614  );
buf ( g3614 , n3615  );
buf ( g3615 , n3616  );
buf ( g3616 , n3617  );
buf ( g3617 , n3618  );
buf ( g3618 , n3619  );
buf ( g3619 , n3620  );
buf ( g3620 , n3621  );
buf ( g3621 , n3622  );
buf ( g3622 , n3623  );
buf ( g3623 , n3624  );
buf ( g3624 , n3625  );
buf ( g3625 , n3626  );
buf ( g3626 , n3627  );
buf ( g3627 , n3628  );
buf ( g3628 , n3629  );
buf ( g3629 , n3630  );
buf ( g3630 , n3631  );
buf ( g3631 , n3632  );
buf ( g3632 , n3633  );
buf ( g3633 , n3634  );
buf ( g3634 , n3635  );
buf ( g3635 , n3636  );
buf ( g3636 , n3637  );
buf ( g3637 , n3638  );
buf ( g3638 , n3639  );
buf ( g3639 , n3640  );
buf ( g3640 , n3641  );
buf ( g3641 , n3642  );
buf ( g3642 , n3643  );
buf ( g3643 , n3644  );
buf ( g3644 , n3645  );
buf ( g3645 , n3646  );
buf ( g3646 , n3647  );
buf ( g3647 , n3648  );
buf ( g3648 , n3649  );
buf ( g3649 , n3650  );
buf ( g3650 , n3651  );
buf ( g3651 , n3652  );
buf ( g3652 , n3653  );
buf ( g3653 , n3654  );
buf ( g3654 , n3655  );
buf ( g3655 , n3656  );
buf ( g3656 , n3657  );
buf ( g3657 , n3658  );
buf ( g3658 , n3659  );
buf ( g3659 , n3660  );
buf ( g3660 , n3661  );
buf ( g3661 , n3662  );
buf ( g3662 , n3663  );
buf ( g3663 , n3664  );
buf ( g3664 , n3665  );
buf ( g3665 , n3666  );
buf ( g3666 , n3667  );
buf ( g3667 , n3668  );
buf ( g3668 , n3669  );
buf ( g3669 , n3670  );
buf ( g3670 , n3671  );
buf ( g3671 , n3672  );
buf ( g3672 , n3673  );
buf ( g3673 , n3674  );
buf ( g3674 , n3675  );
buf ( g3675 , n3676  );
buf ( g3676 , n3677  );
buf ( g3677 , n3678  );
buf ( g3678 , n3679  );
buf ( g3679 , n3680  );
buf ( g3680 , n3681  );
buf ( g3681 , n3682  );
buf ( g3682 , n3683  );
buf ( g3683 , n3684  );
buf ( g3684 , n3685  );
buf ( g3685 , n3686  );
buf ( g3686 , n3687  );
buf ( g3687 , n3688  );
buf ( g3688 , n3689  );
buf ( g3689 , n3690  );
buf ( g3690 , n3691  );
buf ( g3691 , n3692  );
buf ( g3692 , n3693  );
buf ( g3693 , n3694  );
buf ( g3694 , n3695  );
buf ( g3695 , n3696  );
buf ( g3696 , n3697  );
buf ( g3697 , n3698  );
buf ( g3698 , n3699  );
buf ( g3699 , n3700  );
buf ( g3700 , n3701  );
buf ( g3701 , n3702  );
buf ( g3702 , n3703  );
buf ( g3703 , n3704  );
buf ( g3704 , n3705  );
buf ( g3705 , n3706  );
buf ( g3706 , n3707  );
buf ( g3707 , n3708  );
buf ( g3708 , n3709  );
buf ( g3709 , n3710  );
buf ( g3710 , n3711  );
buf ( g3711 , n3712  );
buf ( g3712 , n3713  );
buf ( g3713 , n3714  );
buf ( g3714 , n3715  );
buf ( g3715 , n3716  );
buf ( g3716 , n3717  );
buf ( g3717 , n3718  );
buf ( g3718 , n3719  );
buf ( g3719 , n3720  );
buf ( g3720 , n3721  );
buf ( g3721 , n3722  );
buf ( g3722 , n3723  );
buf ( g3723 , n3724  );
buf ( g3724 , n3725  );
buf ( g3725 , n3726  );
buf ( g3726 , n3727  );
buf ( g3727 , n3728  );
buf ( g3728 , n3729  );
buf ( g3729 , n3730  );
buf ( g3730 , n3731  );
buf ( g3731 , n3732  );
buf ( g3732 , n3733  );
buf ( g3733 , n3734  );
buf ( g3734 , n3735  );
buf ( g3735 , n3736  );
buf ( g3736 , n3737  );
buf ( g3737 , n3738  );
buf ( g3738 , n3739  );
buf ( g3739 , n3740  );
buf ( g3740 , n3741  );
buf ( g3741 , n3742  );
buf ( g3742 , n3743  );
buf ( g3743 , n3744  );
buf ( g3744 , n3745  );
buf ( g3745 , n3746  );
buf ( g3746 , n3747  );
buf ( g3747 , n3748  );
buf ( g3748 , n3749  );
buf ( g3749 , n3750  );
buf ( g3750 , n3751  );
buf ( g3751 , n3752  );
buf ( g3752 , n3753  );
buf ( g3753 , n3754  );
buf ( g3754 , n3755  );
buf ( g3755 , n3756  );
buf ( g3756 , n3757  );
buf ( g3757 , n3758  );
buf ( g3758 , n3759  );
buf ( g3759 , n3760  );
buf ( g3760 , n3761  );
buf ( g3761 , n3762  );
buf ( g3762 , n3763  );
buf ( g3763 , n3764  );
buf ( g3764 , n3765  );
buf ( g3765 , n3766  );
buf ( g3766 , n3767  );
buf ( g3767 , n3768  );
buf ( g3768 , n3769  );
buf ( g3769 , n3770  );
buf ( g3770 , n3771  );
buf ( g3771 , n3772  );
buf ( g3772 , n3773  );
buf ( g3773 , n3774  );
buf ( g3774 , n3775  );
buf ( g3775 , n3776  );
buf ( g3776 , n3777  );
buf ( g3777 , n3778  );
buf ( g3778 , n3779  );
buf ( g3779 , n3780  );
buf ( g3780 , n3781  );
buf ( g3781 , n3782  );
buf ( g3782 , n3783  );
buf ( g3783 , n3784  );
buf ( g3784 , n3785  );
buf ( g3785 , n3786  );
buf ( g3786 , n3787  );
buf ( g3787 , n3788  );
buf ( g3788 , n3789  );
buf ( g3789 , n3790  );
buf ( g3790 , n3791  );
buf ( g3791 , n3792  );
buf ( g3792 , n3793  );
buf ( g3793 , n3794  );
buf ( g3794 , n3795  );
buf ( g3795 , n3796  );
buf ( g3796 , n3797  );
buf ( g3797 , n3798  );
buf ( g3798 , n3799  );
buf ( g3799 , n3800  );
buf ( g3800 , n3801  );
buf ( g3801 , n3802  );
buf ( g3802 , n3803  );
buf ( g3803 , n3804  );
buf ( g3804 , n3805  );
buf ( g3805 , n3806  );
buf ( g3806 , n3807  );
buf ( g3807 , n3808  );
buf ( g3808 , n3809  );
buf ( g3809 , n3810  );
buf ( g3810 , n3811  );
buf ( g3811 , n3812  );
buf ( g3812 , n3813  );
buf ( g3813 , n3814  );
buf ( g3814 , n3815  );
buf ( g3815 , n3816  );
buf ( g3816 , n3817  );
buf ( g3817 , n3818  );
buf ( g3818 , n3819  );
buf ( g3819 , n3820  );
buf ( g3820 , n3821  );
buf ( g3821 , n3822  );
buf ( g3822 , n3823  );
buf ( g3823 , n3824  );
buf ( g3824 , n3825  );
buf ( g3825 , n3826  );
buf ( g3826 , n3827  );
buf ( g3827 , n3828  );
buf ( g3828 , n3829  );
buf ( g3829 , n3830  );
buf ( g3830 , n3831  );
buf ( g3831 , n3832  );
buf ( g3832 , n3833  );
buf ( g3833 , n3834  );
buf ( g3834 , n3835  );
buf ( g3835 , n3836  );
buf ( g3836 , n3837  );
buf ( g3837 , n3838  );
buf ( g3838 , n3839  );
buf ( g3839 , n3840  );
buf ( g3840 , n3841  );
buf ( g3841 , n3842  );
buf ( g3842 , n3843  );
buf ( g3843 , n3844  );
buf ( g3844 , n3845  );
buf ( g3845 , n3846  );
buf ( g3846 , n3847  );
buf ( g3847 , n3848  );
buf ( g3848 , n3849  );
buf ( g3849 , n3850  );
buf ( g3850 , n3851  );
buf ( g3851 , n3852  );
buf ( g3852 , n3853  );
buf ( g3853 , n3854  );
buf ( g3854 , n3855  );
buf ( g3855 , n3856  );
buf ( g3856 , n3857  );
buf ( g3857 , n3858  );
buf ( g3858 , n3859  );
buf ( g3859 , n3860  );
buf ( g3860 , n3861  );
buf ( g3861 , n3862  );
buf ( g3862 , n3863  );
buf ( g3863 , n3864  );
buf ( g3864 , n3865  );
buf ( g3865 , n3866  );
buf ( g3866 , n3867  );
buf ( g3867 , n3868  );
buf ( g3868 , n3869  );
buf ( g3869 , n3870  );
buf ( g3870 , n3871  );
buf ( g3871 , n3872  );
buf ( g3872 , n3873  );
buf ( g3873 , n3874  );
buf ( g3874 , n3875  );
buf ( g3875 , n3876  );
buf ( g3876 , n3877  );
buf ( g3877 , n3878  );
buf ( g3878 , n3879  );
buf ( g3879 , n3880  );
buf ( g3880 , n3881  );
buf ( g3881 , n3882  );
buf ( g3882 , n3883  );
buf ( g3883 , n3884  );
buf ( g3884 , n3885  );
buf ( g3885 , n3886  );
buf ( g3886 , n3887  );
buf ( g3887 , n3888  );
buf ( g3888 , n3889  );
buf ( g3889 , n3890  );
buf ( g3890 , n3891  );
buf ( g3891 , n3892  );
buf ( g3892 , n3893  );
buf ( g3893 , n3894  );
buf ( g3894 , n3895  );
buf ( g3895 , n3896  );
buf ( g3896 , n3897  );
buf ( g3897 , n3898  );
buf ( g3898 , n3899  );
buf ( g3899 , n3900  );
buf ( g3900 , n3901  );
buf ( g3901 , n3902  );
buf ( g3902 , n3903  );
buf ( g3903 , n3904  );
buf ( g3904 , n3905  );
buf ( g3905 , n3906  );
buf ( g3906 , n3907  );
buf ( g3907 , n3908  );
buf ( g3908 , n3909  );
buf ( g3909 , n3910  );
buf ( g3910 , n3911  );
buf ( g3911 , n3912  );
buf ( g3912 , n3913  );
buf ( g3913 , n3914  );
buf ( g3914 , n3915  );
buf ( g3915 , n3916  );
buf ( g3916 , n3917  );
buf ( g3917 , n3918  );
buf ( g3918 , n3919  );
buf ( g3919 , n3920  );
buf ( g3920 , n3921  );
buf ( g3921 , n3922  );
buf ( g3922 , n3923  );
buf ( g3923 , n3924  );
buf ( g3924 , n3925  );
buf ( g3925 , n3926  );
buf ( g3926 , n3927  );
buf ( g3927 , n3928  );
buf ( g3928 , n3929  );
buf ( g3929 , n3930  );
buf ( g3930 , n3931  );
buf ( g3931 , n3932  );
buf ( g3932 , n3933  );
buf ( g3933 , n3934  );
buf ( g3934 , n3935  );
buf ( g3935 , n3936  );
buf ( g3936 , n3937  );
buf ( g3937 , n3938  );
buf ( g3938 , n3939  );
buf ( g3939 , n3940  );
buf ( g3940 , n3941  );
buf ( g3941 , n3942  );
buf ( g3942 , n3943  );
buf ( g3943 , n3944  );
buf ( g3944 , n3945  );
buf ( g3945 , n3946  );
buf ( g3946 , n3947  );
buf ( g3947 , n3948  );
buf ( g3948 , n3949  );
buf ( g3949 , n3950  );
buf ( g3950 , n3951  );
buf ( g3951 , n3952  );
buf ( g3952 , n3953  );
buf ( g3953 , n3954  );
buf ( g3954 , n3955  );
buf ( g3955 , n3956  );
buf ( g3956 , n3957  );
buf ( g3957 , n3958  );
buf ( g3958 , n3959  );
buf ( g3959 , n3960  );
buf ( g3960 , n3961  );
buf ( g3961 , n3962  );
buf ( g3962 , n3963  );
buf ( g3963 , n3964  );
buf ( g3964 , n3965  );
buf ( g3965 , n3966  );
buf ( g3966 , n3967  );
buf ( g3967 , n3968  );
buf ( g3968 , n3969  );
buf ( g3969 , n3970  );
buf ( g3970 , n3971  );
buf ( g3971 , n3972  );
buf ( g3972 , n3973  );
buf ( g3973 , n3974  );
buf ( g3974 , n3975  );
buf ( g3975 , n3976  );
buf ( g3976 , n3977  );
buf ( g3977 , n3978  );
buf ( g3978 , n3979  );
buf ( g3979 , n3980  );
buf ( g3980 , n3981  );
buf ( g3981 , n3982  );
buf ( g3982 , n3983  );
buf ( g3983 , n3984  );
buf ( g3984 , n3985  );
buf ( g3985 , n3986  );
buf ( g3986 , n3987  );
buf ( g3987 , n3988  );
buf ( g3988 , n3989  );
buf ( g3989 , n3990  );
buf ( g3990 , n3991  );
buf ( g3991 , n3992  );
buf ( g3992 , n3993  );
buf ( g3993 , n3994  );
buf ( g3994 , n3995  );
buf ( g3995 , n3996  );
buf ( g3996 , n3997  );
buf ( g3997 , n3998  );
buf ( g3998 , n3999  );
buf ( g3999 , n4000  );
buf ( g4000 , n4001  );
buf ( g4001 , n4002  );
buf ( g4002 , n4003  );
buf ( g4003 , n4004  );
buf ( g4004 , n4005  );
buf ( g4005 , n4006  );
buf ( g4006 , n4007  );
buf ( g4007 , n4008  );
buf ( g4008 , n4009  );
buf ( g4009 , n4010  );
buf ( g4010 , n4011  );
buf ( g4011 , n4012  );
buf ( g4012 , n4013  );
buf ( g4013 , n4014  );
buf ( g4014 , n4015  );
buf ( g4015 , n4016  );
buf ( g4016 , n4017  );
buf ( g4017 , n4018  );
buf ( g4018 , n4019  );
buf ( g4019 , n4020  );
buf ( g4020 , n4021  );
buf ( g4021 , n4022  );
buf ( g4022 , n4023  );
buf ( g4023 , n4024  );
buf ( g4024 , n4025  );
buf ( g4025 , n4026  );
buf ( g4026 , n4027  );
buf ( g4027 , n4028  );
buf ( g4028 , n4029  );
buf ( g4029 , n4030  );
buf ( g4030 , n4031  );
buf ( g4031 , n4032  );
buf ( g4032 , n4033  );
buf ( g4033 , n4034  );
buf ( g4034 , n4035  );
buf ( g4035 , n4036  );
buf ( g4036 , n4037  );
buf ( g4037 , n4038  );
buf ( g4038 , n4039  );
buf ( g4039 , n4040  );
buf ( g4040 , n4041  );
buf ( g4041 , n4042  );
buf ( g4042 , n4043  );
buf ( g4043 , n4044  );
buf ( g4044 , n4045  );
buf ( g4045 , n4046  );
buf ( g4046 , n4047  );
buf ( g4047 , n4048  );
buf ( g4048 , n4049  );
buf ( g4049 , n4050  );
buf ( g4050 , n4051  );
buf ( g4051 , n4052  );
buf ( g4052 , n4053  );
buf ( g4053 , n4054  );
buf ( g4054 , n4055  );
buf ( g4055 , n4056  );
buf ( g4056 , n4057  );
buf ( g4057 , n4058  );
buf ( g4058 , n4059  );
buf ( g4059 , n4060  );
buf ( g4060 , n4061  );
buf ( g4061 , n4062  );
buf ( g4062 , n4063  );
buf ( g4063 , n4064  );
buf ( g4064 , n4065  );
buf ( g4065 , n4066  );
buf ( g4066 , n4067  );
buf ( g4067 , n4068  );
buf ( g4068 , n4069  );
buf ( g4069 , n4070  );
buf ( g4070 , n4071  );
buf ( g4071 , n4072  );
buf ( g4072 , n4073  );
buf ( g4073 , n4074  );
buf ( g4074 , n4075  );
buf ( g4075 , n4076  );
buf ( g4076 , n4077  );
buf ( g4077 , n4078  );
buf ( g4078 , n4079  );
buf ( g4079 , n4080  );
buf ( g4080 , n4081  );
buf ( g4081 , n4082  );
buf ( g4082 , n4083  );
buf ( g4083 , n4084  );
buf ( g4084 , n4085  );
buf ( g4085 , n4086  );
buf ( g4086 , n4087  );
buf ( g4087 , n4088  );
buf ( g4088 , n4089  );
buf ( g4089 , n4090  );
buf ( g4090 , n4091  );
buf ( g4091 , n4092  );
buf ( g4092 , n4093  );
buf ( g4093 , n4094  );
buf ( g4094 , n4095  );
buf ( g4095 , n4096  );
buf ( g4096 , n4097  );
buf ( g4097 , n4098  );
buf ( g4098 , n4099  );
buf ( g4099 , n4100  );
buf ( g4100 , n4101  );
buf ( g4101 , n4102  );
buf ( g4102 , n4103  );
buf ( g4103 , n4104  );
buf ( g4104 , n4105  );
buf ( g4105 , n4106  );
buf ( g4106 , n4107  );
buf ( g4107 , n4108  );
buf ( g4108 , n4109  );
buf ( g4109 , n4110  );
buf ( g4110 , n4111  );
buf ( g4111 , n4112  );
buf ( g4112 , n4113  );
buf ( g4113 , n4114  );
buf ( g4114 , n4115  );
buf ( g4115 , n4116  );
buf ( g4116 , n4117  );
buf ( g4117 , n4118  );
buf ( g4118 , n4119  );
buf ( g4119 , n4120  );
buf ( g4120 , n4121  );
buf ( g4121 , n4122  );
buf ( g4122 , n4123  );
buf ( g4123 , n4124  );
buf ( g4124 , n4125  );
buf ( g4125 , n4126  );
buf ( g4126 , n4127  );
buf ( g4127 , n4128  );
buf ( g4128 , n4129  );
buf ( g4129 , n4130  );
buf ( g4130 , n4131  );
buf ( g4131 , n4132  );
buf ( g4132 , n4133  );
buf ( g4133 , n4134  );
buf ( g4134 , n4135  );
buf ( g4135 , n4136  );
buf ( g4136 , n4137  );
buf ( g4137 , n4138  );
buf ( g4138 , n4139  );
buf ( g4139 , n4140  );
buf ( g4140 , n4141  );
buf ( g4141 , n4142  );
buf ( g4142 , n4143  );
buf ( g4143 , n4144  );
buf ( g4144 , n4145  );
buf ( g4145 , n4146  );
buf ( g4146 , n4147  );
buf ( g4147 , n4148  );
buf ( g4148 , n4149  );
buf ( g4149 , n4150  );
buf ( g4150 , n4151  );
buf ( g4151 , n4152  );
buf ( g4152 , n4153  );
buf ( g4153 , n4154  );
buf ( g4154 , n4155  );
buf ( g4155 , n4156  );
buf ( g4156 , n4157  );
buf ( g4157 , n4158  );
buf ( g4158 , n4159  );
buf ( g4159 , n4160  );
buf ( g4160 , n4161  );
buf ( g4161 , n4162  );
buf ( g4162 , n4163  );
buf ( g4163 , n4164  );
buf ( g4164 , n4165  );
buf ( g4165 , n4166  );
buf ( g4166 , n4167  );
buf ( g4167 , n4168  );
buf ( g4168 , n4169  );
buf ( g4169 , n4170  );
buf ( g4170 , n4171  );
buf ( g4171 , n4172  );
buf ( g4172 , n4173  );
buf ( g4173 , n4174  );
buf ( g4174 , n4175  );
buf ( g4175 , n4176  );
buf ( g4176 , n4177  );
buf ( g4177 , n4178  );
buf ( g4178 , n4179  );
buf ( g4179 , n4180  );
buf ( g4180 , n4181  );
buf ( g4181 , n4182  );
buf ( g4182 , n4183  );
buf ( g4183 , n4184  );
buf ( g4184 , n4185  );
buf ( g4185 , n4186  );
buf ( g4186 , n4187  );
buf ( g4187 , n4188  );
buf ( g4188 , n4189  );
buf ( g4189 , n4190  );
buf ( g4190 , n4191  );
buf ( g4191 , n4192  );
buf ( g4192 , n4193  );
buf ( g4193 , n4194  );
buf ( g4194 , n4195  );
buf ( g4195 , n4196  );
buf ( g4196 , n4197  );
buf ( g4197 , n4198  );
buf ( g4198 , n4199  );
buf ( g4199 , n4200  );
buf ( g4200 , n4201  );
buf ( g4201 , n4202  );
buf ( g4202 , n4203  );
buf ( g4203 , n4204  );
buf ( g4204 , n4205  );
buf ( g4205 , n4206  );
buf ( g4206 , n4207  );
buf ( g4207 , n4208  );
buf ( g4208 , n4209  );
buf ( g4209 , n4210  );
buf ( g4210 , n4211  );
buf ( g4211 , n4212  );
buf ( g4212 , n4213  );
buf ( g4213 , n4214  );
buf ( g4214 , n4215  );
buf ( g4215 , n4216  );
buf ( g4216 , n4217  );
buf ( g4217 , n4218  );
buf ( g4218 , n4219  );
buf ( g4219 , n4220  );
buf ( g4220 , n4221  );
buf ( g4221 , n4222  );
buf ( g4222 , n4223  );
buf ( g4223 , n4224  );
buf ( g4224 , n4225  );
buf ( g4225 , n4226  );
buf ( g4226 , n4227  );
buf ( g4227 , n4228  );
buf ( g4228 , n4229  );
buf ( g4229 , n4230  );
buf ( g4230 , n4231  );
buf ( g4231 , n4232  );
buf ( g4232 , n4233  );
buf ( g4233 , n4234  );
buf ( g4234 , n4235  );
buf ( g4235 , n4236  );
buf ( g4236 , n4237  );
buf ( g4237 , n4238  );
buf ( g4238 , n4239  );
buf ( g4239 , n4240  );
buf ( g4240 , n4241  );
buf ( g4241 , n4242  );
buf ( g4242 , n4243  );
buf ( g4243 , n4244  );
buf ( g4244 , n4245  );
buf ( g4245 , n4246  );
buf ( g4246 , n4247  );
buf ( g4247 , n4248  );
buf ( g4248 , n4249  );
buf ( g4249 , n4250  );
buf ( g4250 , n4251  );
buf ( g4251 , n4252  );
buf ( g4252 , n4253  );
buf ( g4253 , n4254  );
buf ( g4254 , n4255  );
buf ( g4255 , n4256  );
buf ( g4256 , n4257  );
buf ( g4257 , n4258  );
buf ( g4258 , n4259  );
buf ( g4259 , n4260  );
buf ( g4260 , n4261  );
buf ( g4261 , n4262  );
buf ( g4262 , n4263  );
buf ( g4263 , n4264  );
buf ( g4264 , n4265  );
buf ( g4265 , n4266  );
buf ( g4266 , n4267  );
buf ( g4267 , n4268  );
buf ( g4268 , n4269  );
buf ( g4269 , n4270  );
buf ( g4270 , n4271  );
buf ( g4271 , n4272  );
buf ( g4272 , n4273  );
buf ( g4273 , n4274  );
buf ( g4274 , n4275  );
buf ( g4275 , n4276  );
buf ( g4276 , n4277  );
buf ( g4277 , n4278  );
buf ( g4278 , n4279  );
buf ( g4279 , n4280  );
buf ( g4280 , n4281  );
buf ( g4281 , n4282  );
buf ( g4282 , n4283  );
buf ( g4283 , n4284  );
buf ( g4284 , n4285  );
buf ( g4285 , n4286  );
buf ( g4286 , n4287  );
buf ( g4287 , n4288  );
buf ( g4288 , n4289  );
buf ( g4289 , n4290  );
buf ( g4290 , n4291  );
buf ( g4291 , n4292  );
buf ( g4292 , n4293  );
buf ( g4293 , n4294  );
buf ( g4294 , n4295  );
buf ( g4295 , n4296  );
buf ( g4296 , n4297  );
buf ( g4297 , n4298  );
buf ( g4298 , n4299  );
buf ( g4299 , n4300  );
buf ( g4300 , n4301  );
buf ( g4301 , n4302  );
buf ( g4302 , n4303  );
buf ( g4303 , n4304  );
buf ( g4304 , n4305  );
buf ( g4305 , n4306  );
buf ( g4306 , n4307  );
buf ( g4307 , n4308  );
buf ( g4308 , n4309  );
buf ( g4309 , n4310  );
buf ( g4310 , n4311  );
buf ( g4311 , n4312  );
buf ( g4312 , n4313  );
buf ( g4313 , n4314  );
buf ( g4314 , n4315  );
buf ( g4315 , n4316  );
buf ( g4316 , n4317  );
buf ( g4317 , n4318  );
buf ( g4318 , n4319  );
buf ( g4319 , n4320  );
buf ( g4320 , n4321  );
buf ( g4321 , n4322  );
buf ( g4322 , n4323  );
buf ( g4323 , n4324  );
buf ( g4324 , n4325  );
buf ( g4325 , n4326  );
buf ( g4326 , n4327  );
buf ( g4327 , n4328  );
buf ( g4328 , n4329  );
buf ( g4329 , n4330  );
buf ( g4330 , n4331  );
buf ( g4331 , n4332  );
buf ( g4332 , n4333  );
buf ( g4333 , n4334  );
buf ( g4334 , n4335  );
buf ( g4335 , n4336  );
buf ( g4336 , n4337  );
buf ( g4337 , n4338  );
buf ( g4338 , n4339  );
buf ( g4339 , n4340  );
buf ( g4340 , n4341  );
buf ( g4341 , n4342  );
buf ( g4342 , n4343  );
buf ( g4343 , n4344  );
buf ( g4344 , n4345  );
buf ( g4345 , n4346  );
buf ( g4346 , n4347  );
buf ( g4347 , n4348  );
buf ( g4348 , n4349  );
buf ( g4349 , n4350  );
buf ( g4350 , n4351  );
buf ( g4351 , n4352  );
buf ( g4352 , n4353  );
buf ( g4353 , n4354  );
buf ( g4354 , n4355  );
buf ( g4355 , n4356  );
buf ( g4356 , n4357  );
buf ( g4357 , n4358  );
buf ( g4358 , n4359  );
buf ( g4359 , n4360  );
buf ( g4360 , n4361  );
buf ( g4361 , n4362  );
buf ( g4362 , n4363  );
buf ( g4363 , n4364  );
buf ( g4364 , n4365  );
buf ( g4365 , n4366  );
buf ( g4366 , n4367  );
buf ( g4367 , n4368  );
buf ( g4368 , n4369  );
buf ( g4369 , n4370  );
buf ( g4370 , n4371  );
buf ( g4371 , n4372  );
buf ( g4372 , n4373  );
buf ( g4373 , n4374  );
buf ( g4374 , n4375  );
buf ( g4375 , n4376  );
buf ( g4376 , n4377  );
buf ( g4377 , n4378  );
buf ( g4378 , n4379  );
buf ( g4379 , n4380  );
buf ( g4380 , n4381  );
buf ( g4381 , n4382  );
buf ( g4382 , n4383  );
buf ( g4383 , n4384  );
buf ( g4384 , n4385  );
buf ( g4385 , n4386  );
buf ( g4386 , n4387  );
buf ( g4387 , n4388  );
buf ( g4388 , n4389  );
buf ( g4389 , n4390  );
buf ( g4390 , n4391  );
buf ( g4391 , n4392  );
buf ( g4392 , n4393  );
buf ( g4393 , n4394  );
buf ( g4394 , n4395  );
buf ( g4395 , n4396  );
buf ( g4396 , n4397  );
buf ( g4397 , n4398  );
buf ( g4398 , n4399  );
buf ( g4399 , n4400  );
buf ( g4400 , n4401  );
buf ( g4401 , n4402  );
buf ( g4402 , n4403  );
buf ( g4403 , n4404  );
buf ( g4404 , n4405  );
buf ( g4405 , n4406  );
buf ( g4406 , n4407  );
buf ( g4407 , n4408  );
buf ( g4408 , n4409  );
buf ( g4409 , n4410  );
buf ( g4410 , n4411  );
buf ( g4411 , n4412  );
buf ( g4412 , n4413  );
buf ( g4413 , n4414  );
buf ( g4414 , n4415  );
buf ( g4415 , n4416  );
buf ( g4416 , n4417  );
buf ( g4417 , n4418  );
buf ( g4418 , n4419  );
buf ( g4419 , n4420  );
buf ( g4420 , n4421  );
buf ( g4421 , n4422  );
buf ( g4422 , n4423  );
buf ( g4423 , n4424  );
buf ( g4424 , n4425  );
buf ( g4425 , n4426  );
buf ( g4426 , n4427  );
buf ( g4427 , n4428  );
buf ( g4428 , n4429  );
buf ( g4429 , n4430  );
buf ( g4430 , n4431  );
buf ( g4431 , n4432  );
buf ( g4432 , n4433  );
buf ( g4433 , n4434  );
buf ( g4434 , n4435  );
buf ( g4435 , n4436  );
buf ( g4436 , n4437  );
buf ( g4437 , n4438  );
buf ( g4438 , n4439  );
buf ( g4439 , n4440  );
buf ( g4440 , n4441  );
buf ( g4441 , n4442  );
buf ( g4442 , n4443  );
buf ( g4443 , n4444  );
buf ( g4444 , n4445  );
buf ( g4445 , n4446  );
buf ( g4446 , n4447  );
buf ( g4447 , n4448  );
buf ( g4448 , n4449  );
buf ( g4449 , n4450  );
buf ( g4450 , n4451  );
buf ( g4451 , n4452  );
buf ( g4452 , n4453  );
buf ( g4453 , n4454  );
buf ( g4454 , n4455  );
buf ( g4455 , n4456  );
buf ( g4456 , n4457  );
buf ( g4457 , n4458  );
buf ( g4458 , n4459  );
buf ( g4459 , n4460  );
buf ( g4460 , n4461  );
buf ( g4461 , n4462  );
buf ( g4462 , n4463  );
buf ( g4463 , n4464  );
buf ( g4464 , n4465  );
buf ( g4465 , n4466  );
buf ( g4466 , n4467  );
buf ( g4467 , n4468  );
buf ( g4468 , n4469  );
buf ( g4469 , n4470  );
buf ( g4470 , n4471  );
buf ( g4471 , n4472  );
buf ( g4472 , n4473  );
buf ( g4473 , n4474  );
buf ( g4474 , n4475  );
buf ( g4475 , n4476  );
buf ( g4476 , n4477  );
buf ( g4477 , n4478  );
buf ( g4478 , n4479  );
buf ( g4479 , n4480  );
buf ( g4480 , n4481  );
buf ( g4481 , n4482  );
buf ( g4482 , n4483  );
buf ( g4483 , n4484  );
buf ( g4484 , n4485  );
buf ( g4485 , n4486  );
buf ( g4486 , n4487  );
buf ( g4487 , n4488  );
buf ( g4488 , n4489  );
buf ( g4489 , n4490  );
buf ( g4490 , n4491  );
buf ( g4491 , n4492  );
buf ( g4492 , n4493  );
buf ( g4493 , n4494  );
buf ( g4494 , n4495  );
buf ( g4495 , n4496  );
buf ( g4496 , n4497  );
buf ( g4497 , n4498  );
buf ( g4498 , n4499  );
buf ( g4499 , n4500  );
buf ( g4500 , n4501  );
buf ( g4501 , n4502  );
buf ( g4502 , n4503  );
buf ( g4503 , n4504  );
buf ( g4504 , n4505  );
buf ( g4505 , n4506  );
buf ( g4506 , n4507  );
buf ( g4507 , n4508  );
buf ( g4508 , n4509  );
buf ( g4509 , n4510  );
buf ( g4510 , n4511  );
buf ( g4511 , n4512  );
buf ( g4512 , n4513  );
buf ( g4513 , n4514  );
buf ( g4514 , n4515  );
buf ( g4515 , n4516  );
buf ( g4516 , n4517  );
buf ( g4517 , n4518  );
buf ( g4518 , n4519  );
buf ( g4519 , n4520  );
buf ( g4520 , n4521  );
buf ( g4521 , n4522  );
buf ( g4522 , n4523  );
buf ( g4523 , n4524  );
buf ( g4524 , n4525  );
buf ( g4525 , n4526  );
buf ( g4526 , n4527  );
buf ( g4527 , n4528  );
buf ( g4528 , n4529  );
buf ( g4529 , n4530  );
buf ( g4530 , n4531  );
buf ( g4531 , n4532  );
buf ( g4532 , n4533  );
buf ( g4533 , n4534  );
buf ( g4534 , n4535  );
buf ( g4535 , n4536  );
buf ( g4536 , n4537  );
buf ( g4537 , n4538  );
buf ( g4538 , n4539  );
buf ( g4539 , n4540  );
buf ( g4540 , n4541  );
buf ( g4541 , n4542  );
buf ( g4542 , n4543  );
buf ( g4543 , n4544  );
buf ( g4544 , n4545  );
buf ( g4545 , n4546  );
buf ( g4546 , n4547  );
buf ( g4547 , n4548  );
buf ( g4548 , n4549  );
buf ( g4549 , n4550  );
buf ( g4550 , n4551  );
buf ( g4551 , n4552  );
buf ( g4552 , n4553  );
buf ( g4553 , n4554  );
buf ( g4554 , n4555  );
buf ( g4555 , n4556  );
buf ( g4556 , n4557  );
buf ( g4557 , n4558  );
buf ( g4558 , n4559  );
buf ( g4559 , n4560  );
buf ( g4560 , n4561  );
buf ( g4561 , n4562  );
buf ( g4562 , n4563  );
buf ( g4563 , n4564  );
buf ( g4564 , n4565  );
buf ( g4565 , n4566  );
buf ( g4566 , n4567  );
buf ( g4567 , n4568  );
buf ( g4568 , n4569  );
buf ( g4569 , n4570  );
buf ( g4570 , n4571  );
buf ( g4571 , n4572  );
buf ( g4572 , n4573  );
buf ( g4573 , n4574  );
buf ( g4574 , n4575  );
buf ( g4575 , n4576  );
buf ( g4576 , n4577  );
buf ( g4577 , n4578  );
buf ( g4578 , n4579  );
buf ( g4579 , n4580  );
buf ( g4580 , n4581  );
buf ( g4581 , n4582  );
buf ( g4582 , n4583  );
buf ( g4583 , n4584  );
buf ( g4584 , n4585  );
buf ( g4585 , n4586  );
buf ( g4586 , n4587  );
buf ( g4587 , n4588  );
buf ( g4588 , n4589  );
buf ( g4589 , n4590  );
buf ( g4590 , n4591  );
buf ( g4591 , n4592  );
buf ( g4592 , n4593  );
buf ( g4593 , n4594  );
buf ( g4594 , n4595  );
buf ( g4595 , n4596  );
buf ( g4596 , n4597  );
buf ( g4597 , n4598  );
buf ( g4598 , n4599  );
buf ( g4599 , n4600  );
buf ( g4600 , n4601  );
buf ( g4601 , n4602  );
buf ( g4602 , n4603  );
buf ( g4603 , n4604  );
buf ( g4604 , n4605  );
buf ( g4605 , n4606  );
buf ( g4606 , n4607  );
buf ( g4607 , n4608  );
buf ( g4608 , n4609  );
buf ( g4609 , n4610  );
buf ( g4610 , n4611  );
buf ( g4611 , n4612  );
buf ( g4612 , n4613  );
buf ( g4613 , n4614  );
buf ( g4614 , n4615  );
buf ( g4615 , n4616  );
buf ( g4616 , n4617  );
buf ( g4617 , n4618  );
buf ( g4618 , n4619  );
buf ( g4619 , n4620  );
buf ( g4620 , n4621  );
buf ( g4621 , n4622  );
buf ( g4622 , n4623  );
buf ( g4623 , n4624  );
buf ( g4624 , n4625  );
buf ( g4625 , n4626  );
buf ( g4626 , n4627  );
buf ( g4627 , n4628  );
buf ( g4628 , n4629  );
buf ( g4629 , n4630  );
buf ( g4630 , n4631  );
buf ( g4631 , n4632  );
buf ( g4632 , n4633  );
buf ( g4633 , n4634  );
buf ( g4634 , n4635  );
buf ( g4635 , n4636  );
buf ( g4636 , n4637  );
buf ( g4637 , n4638  );
buf ( g4638 , n4639  );
buf ( g4639 , n4640  );
buf ( g4640 , n4641  );
buf ( g4641 , n4642  );
buf ( g4642 , n4643  );
buf ( g4643 , n4644  );
buf ( g4644 , n4645  );
buf ( g4645 , n4646  );
buf ( g4646 , n4647  );
buf ( g4647 , n4648  );
buf ( g4648 , n4649  );
buf ( g4649 , n4650  );
buf ( g4650 , n4651  );
buf ( g4651 , n4652  );
buf ( g4652 , n4653  );
buf ( g4653 , n4654  );
buf ( g4654 , n4655  );
buf ( g4655 , n4656  );
buf ( g4656 , n4657  );
buf ( g4657 , n4658  );
buf ( g4658 , n4659  );
buf ( g4659 , n4660  );
buf ( g4660 , n4661  );
buf ( g4661 , n4662  );
buf ( g4662 , n4663  );
buf ( g4663 , n4664  );
buf ( g4664 , n4665  );
buf ( g4665 , n4666  );
buf ( g4666 , n4667  );
buf ( g4667 , n4668  );
buf ( g4668 , n4669  );
buf ( g4669 , n4670  );
buf ( g4670 , n4671  );
buf ( g4671 , n4672  );
buf ( g4672 , n4673  );
buf ( g4673 , n4674  );
buf ( g4674 , n4675  );
buf ( g4675 , n4676  );
buf ( g4676 , n4677  );
buf ( g4677 , n4678  );
buf ( g4678 , n4679  );
buf ( g4679 , n4680  );
buf ( g4680 , n4681  );
buf ( g4681 , n4682  );
buf ( g4682 , n4683  );
buf ( g4683 , n4684  );
buf ( g4684 , n4685  );
buf ( g4685 , n4686  );
buf ( g4686 , n4687  );
buf ( g4687 , n4688  );
buf ( g4688 , n4689  );
buf ( g4689 , n4690  );
buf ( g4690 , n4691  );
buf ( g4691 , n4692  );
buf ( g4692 , n4693  );
buf ( g4693 , n4694  );
buf ( g4694 , n4695  );
buf ( g4695 , n4696  );
buf ( g4696 , n4697  );
buf ( g4697 , n4698  );
buf ( g4698 , n4699  );
buf ( g4699 , n4700  );
buf ( g4700 , n4701  );
buf ( g4701 , n4702  );
buf ( g4702 , n4703  );
buf ( g4703 , n4704  );
buf ( g4704 , n4705  );
buf ( g4705 , n4706  );
buf ( g4706 , n4707  );
buf ( g4707 , n4708  );
buf ( g4708 , n4709  );
buf ( g4709 , n4710  );
buf ( g4710 , n4711  );
buf ( g4711 , n4712  );
buf ( g4712 , n4713  );
buf ( g4713 , n4714  );
buf ( g4714 , n4715  );
buf ( g4715 , n4716  );
buf ( g4716 , n4717  );
buf ( g4717 , n4718  );
buf ( g4718 , n4719  );
buf ( g4719 , n4720  );
buf ( g4720 , n4721  );
buf ( g4721 , n4722  );
buf ( g4722 , n4723  );
buf ( g4723 , n4724  );
buf ( g4724 , n4725  );
buf ( g4725 , n4726  );
buf ( g4726 , n4727  );
buf ( g4727 , n4728  );
buf ( g4728 , n4729  );
buf ( g4729 , n4730  );
buf ( g4730 , n4731  );
buf ( g4731 , n4732  );
buf ( g4732 , n4733  );
buf ( g4733 , n4734  );
buf ( g4734 , n4735  );
buf ( g4735 , n4736  );
buf ( g4736 , n4737  );
buf ( g4737 , n4738  );
buf ( g4738 , n4739  );
buf ( g4739 , n4740  );
buf ( g4740 , n4741  );
buf ( g4741 , n4742  );
buf ( g4742 , n4743  );
buf ( g4743 , n4744  );
buf ( g4744 , n4745  );
buf ( g4745 , n4746  );
buf ( g4746 , n4747  );
buf ( g4747 , n4748  );
buf ( g4748 , n4749  );
buf ( g4749 , n4750  );
buf ( g4750 , n4751  );
buf ( g4751 , n4752  );
buf ( g4752 , n4753  );
buf ( g4753 , n4754  );
buf ( g4754 , n4755  );
buf ( g4755 , n4756  );
buf ( g4756 , n4757  );
buf ( g4757 , n4758  );
buf ( g4758 , n4759  );
buf ( g4759 , n4760  );
buf ( g4760 , n4761  );
buf ( g4761 , n4762  );
buf ( g4762 , n4763  );
buf ( g4763 , n4764  );
buf ( g4764 , n4765  );
buf ( g4765 , n4766  );
buf ( g4766 , n4767  );
buf ( g4767 , n4768  );
buf ( g4768 , n4769  );
buf ( g4769 , n4770  );
buf ( g4770 , n4771  );
buf ( g4771 , n4772  );
buf ( g4772 , n4773  );
buf ( g4773 , n4774  );
buf ( g4774 , n4775  );
buf ( g4775 , n4776  );
buf ( g4776 , n4777  );
buf ( g4777 , n4778  );
buf ( g4778 , n4779  );
buf ( g4779 , n4780  );
buf ( g4780 , n4781  );
buf ( g4781 , n4782  );
buf ( g4782 , n4783  );
buf ( g4783 , n4784  );
buf ( g4784 , n4785  );
buf ( g4785 , n4786  );
buf ( g4786 , n4787  );
buf ( g4787 , n4788  );
buf ( g4788 , n4789  );
buf ( g4789 , n4790  );
buf ( g4790 , n4791  );
buf ( g4791 , n4792  );
buf ( g4792 , n4793  );
buf ( g4793 , n4794  );
buf ( g4794 , n4795  );
buf ( g4795 , n4796  );
buf ( g4796 , n4797  );
buf ( g4797 , n4798  );
buf ( g4798 , n4799  );
buf ( g4799 , n4800  );
buf ( g4800 , n4801  );
buf ( g4801 , n4802  );
buf ( g4802 , n4803  );
buf ( g4803 , n4804  );
buf ( g4804 , n4805  );
buf ( g4805 , n4806  );
buf ( g4806 , n4807  );
buf ( g4807 , n4808  );
buf ( g4808 , n4809  );
buf ( g4809 , n4810  );
buf ( g4810 , n4811  );
buf ( g4811 , n4812  );
buf ( g4812 , n4813  );
buf ( g4813 , n4814  );
buf ( g4814 , n4815  );
buf ( g4815 , n4816  );
buf ( g4816 , n4817  );
buf ( g4817 , n4818  );
buf ( g4818 , n4819  );
buf ( g4819 , n4820  );
buf ( g4820 , n4821  );
buf ( g4821 , n4822  );
buf ( g4822 , n4823  );
buf ( g4823 , n4824  );
buf ( g4824 , n4825  );
buf ( g4825 , n4826  );
buf ( g4826 , n4827  );
buf ( g4827 , n4828  );
buf ( g4828 , n4829  );
buf ( g4829 , n4830  );
buf ( g4830 , n4831  );
buf ( g4831 , n4832  );
buf ( g4832 , n4833  );
buf ( g4833 , n4834  );
buf ( g4834 , n4835  );
buf ( g4835 , n4836  );
buf ( g4836 , n4837  );
buf ( g4837 , n4838  );
buf ( g4838 , n4839  );
buf ( g4839 , n4840  );
buf ( g4840 , n4841  );
buf ( g4841 , n4842  );
buf ( g4842 , n4843  );
buf ( g4843 , n4844  );
buf ( g4844 , n4845  );
buf ( g4845 , n4846  );
buf ( g4846 , n4847  );
buf ( g4847 , n4848  );
buf ( g4848 , n4849  );
buf ( g4849 , n4850  );
buf ( g4850 , n4851  );
buf ( g4851 , n4852  );
buf ( g4852 , n4853  );
buf ( g4853 , n4854  );
buf ( g4854 , n4855  );
buf ( g4855 , n4856  );
buf ( g4856 , n4857  );
buf ( g4857 , n4858  );
buf ( g4858 , n4859  );
buf ( g4859 , n4860  );
buf ( g4860 , n4861  );
buf ( g4861 , n4862  );
buf ( g4862 , n4863  );
buf ( g4863 , n4864  );
buf ( g4864 , n4865  );
buf ( g4865 , n4866  );
buf ( g4866 , n4867  );
buf ( g4867 , n4868  );
buf ( g4868 , n4869  );
buf ( g4869 , n4870  );
buf ( g4870 , n4871  );
buf ( g4871 , n4872  );
buf ( g4872 , n4873  );
buf ( g4873 , n4874  );
buf ( g4874 , n4875  );
buf ( g4875 , n4876  );
buf ( g4876 , n4877  );
buf ( g4877 , n4878  );
buf ( g4878 , n4879  );
buf ( g4879 , n4880  );
buf ( g4880 , n4881  );
buf ( g4881 , n4882  );
buf ( g4882 , n4883  );
buf ( g4883 , n4884  );
buf ( g4884 , n4885  );
buf ( g4885 , n4886  );
buf ( g4886 , n4887  );
buf ( g4887 , n4888  );
buf ( g4888 , n4889  );
buf ( g4889 , n4890  );
buf ( g4890 , n4891  );
buf ( g4891 , n4892  );
buf ( g4892 , n4893  );
buf ( g4893 , n4894  );
buf ( g4894 , n4895  );
buf ( g4895 , n4896  );
buf ( g4896 , n4897  );
buf ( g4897 , n4898  );
buf ( g4898 , n4899  );
buf ( g4899 , n4900  );
buf ( g4900 , n4901  );
buf ( g4901 , n4902  );
buf ( g4902 , n4903  );
buf ( g4903 , n4904  );
buf ( g4904 , n4905  );
buf ( g4905 , n4906  );
buf ( g4906 , n4907  );
buf ( g4907 , n4908  );
buf ( g4908 , n4909  );
buf ( g4909 , n4910  );
buf ( g4910 , n4911  );
buf ( g4911 , n4912  );
buf ( g4912 , n4913  );
buf ( g4913 , n4914  );
buf ( g4914 , n4915  );
buf ( g4915 , n4916  );
buf ( g4916 , n4917  );
buf ( g4917 , n4918  );
buf ( g4918 , n4919  );
buf ( g4919 , n4920  );
buf ( g4920 , n4921  );
buf ( g4921 , n4922  );
buf ( g4922 , n4923  );
buf ( g4923 , n4924  );
buf ( g4924 , n4925  );
buf ( g4925 , n4926  );
buf ( g4926 , n4927  );
buf ( g4927 , n4928  );
buf ( g4928 , n4929  );
buf ( g4929 , n4930  );
buf ( g4930 , n4931  );
buf ( g4931 , n4932  );
buf ( g4932 , n4933  );
buf ( g4933 , n4934  );
buf ( g4934 , n4935  );
buf ( g4935 , n4936  );
buf ( g4936 , n4937  );
buf ( g4937 , n4938  );
buf ( g4938 , n4939  );
buf ( g4939 , n4940  );
buf ( g4940 , n4941  );
buf ( g4941 , n4942  );
buf ( g4942 , n4943  );
buf ( g4943 , n4944  );
buf ( g4944 , n4945  );
buf ( g4945 , n4946  );
buf ( g4946 , n4947  );
buf ( g4947 , n4948  );
buf ( g4948 , n4949  );
buf ( g4949 , n4950  );
buf ( g4950 , n4951  );
buf ( g4951 , n4952  );
buf ( g4952 , n4953  );
buf ( g4953 , n4954  );
buf ( g4954 , n4955  );
buf ( g4955 , n4956  );
buf ( g4956 , n4957  );
buf ( g4957 , n4958  );
buf ( g4958 , n4959  );
buf ( g4959 , n4960  );
buf ( g4960 , n4961  );
buf ( g4961 , n4962  );
buf ( g4962 , n4963  );
buf ( g4963 , n4964  );
buf ( g4964 , n4965  );
buf ( g4965 , n4966  );
buf ( g4966 , n4967  );
buf ( g4967 , n4968  );
buf ( g4968 , n4969  );
buf ( g4969 , n4970  );
buf ( g4970 , n4971  );
buf ( g4971 , n4972  );
buf ( g4972 , n4973  );
buf ( g4973 , n4974  );
buf ( g4974 , n4975  );
buf ( g4975 , n4976  );
buf ( g4976 , n4977  );
buf ( g4977 , n4978  );
buf ( g4978 , n4979  );
buf ( g4979 , n4980  );
buf ( g4980 , n4981  );
buf ( g4981 , n4982  );
buf ( g4982 , n4983  );
buf ( g4983 , n4984  );
buf ( g4984 , n4985  );
buf ( g4985 , n4986  );
buf ( g4986 , n4987  );
buf ( g4987 , n4988  );
buf ( g4988 , n4989  );
buf ( g4989 , n4990  );
buf ( g4990 , n4991  );
buf ( g4991 , n4992  );
buf ( g4992 , n4993  );
buf ( g4993 , n4994  );
buf ( g4994 , n4995  );
buf ( g4995 , n4996  );
buf ( g4996 , n4997  );
buf ( g4997 , n4998  );
buf ( g4998 , n4999  );
buf ( g4999 , n5000  );
buf ( g5000 , n5001  );
buf ( g5001 , n5002  );
buf ( g5002 , n5003  );
buf ( g5003 , n5004  );
buf ( g5004 , n5005  );
buf ( g5005 , n5006  );
buf ( g5006 , n5007  );
buf ( g5007 , n5008  );
buf ( g5008 , n5009  );
buf ( g5009 , n5010  );
buf ( g5010 , n5011  );
buf ( g5011 , n5012  );
buf ( g5012 , n5013  );
buf ( g5013 , n5014  );
buf ( g5014 , n5015  );
buf ( g5015 , n5016  );
buf ( g5016 , n5017  );
buf ( g5017 , n5018  );
buf ( g5018 , n5019  );
buf ( g5019 , n5020  );
buf ( g5020 , n5021  );
buf ( g5021 , n5022  );
buf ( g5022 , n5023  );
buf ( g5023 , n5024  );
buf ( g5024 , n5025  );
buf ( g5025 , n5026  );
buf ( g5026 , n5027  );
buf ( g5027 , n5028  );
buf ( g5028 , n5029  );
buf ( g5029 , n5030  );
buf ( g5030 , n5031  );
buf ( g5031 , n5032  );
buf ( g5032 , n5033  );
buf ( g5033 , n5034  );
buf ( g5034 , n5035  );
buf ( g5035 , n5036  );
buf ( g5036 , n5037  );
buf ( g5037 , n5038  );
buf ( g5038 , n5039  );
buf ( g5039 , n5040  );
buf ( g5040 , n5041  );
buf ( g5041 , n5042  );
buf ( g5042 , n5043  );
buf ( g5043 , n5044  );
buf ( g5044 , n5045  );
buf ( g5045 , n5046  );
buf ( g5046 , n5047  );
buf ( g5047 , n5048  );
buf ( g5048 , n5049  );
buf ( g5049 , n5050  );
buf ( g5050 , n5051  );
buf ( g5051 , n5052  );
buf ( g5052 , n5053  );
buf ( g5053 , n5054  );
buf ( g5054 , n5055  );
buf ( g5055 , n5056  );
buf ( g5056 , n5057  );
buf ( g5057 , n5058  );
buf ( g5058 , n5059  );
buf ( g5059 , n5060  );
buf ( g5060 , n5061  );
buf ( g5061 , n5062  );
buf ( g5062 , n5063  );
buf ( g5063 , n5064  );
buf ( g5064 , n5065  );
buf ( g5065 , n5066  );
buf ( g5066 , n5067  );
buf ( g5067 , n5068  );
buf ( g5068 , n5069  );
buf ( g5069 , n5070  );
buf ( g5070 , n5071  );
buf ( g5071 , n5072  );
buf ( g5072 , n5073  );
buf ( g5073 , n5074  );
buf ( g5074 , n5075  );
buf ( g5075 , n5076  );
buf ( g5076 , n5077  );
buf ( g5077 , n5078  );
buf ( g5078 , n5079  );
buf ( g5079 , n5080  );
buf ( g5080 , n5081  );
buf ( g5081 , n5082  );
buf ( g5082 , n5083  );
buf ( g5083 , n5084  );
buf ( g5084 , n5085  );
buf ( g5085 , n5086  );
buf ( g5086 , n5087  );
buf ( g5087 , n5088  );
buf ( g5088 , n5089  );
buf ( g5089 , n5090  );
buf ( g5090 , n5091  );
buf ( g5091 , n5092  );
buf ( g5092 , n5093  );
buf ( g5093 , n5094  );
buf ( g5094 , n5095  );
buf ( g5095 , n5096  );
buf ( g5096 , n5097  );
buf ( g5097 , n5098  );
buf ( g5098 , n5099  );
buf ( g5099 , n5100  );
buf ( g5100 , n5101  );
buf ( g5101 , n5102  );
buf ( g5102 , n5103  );
buf ( g5103 , n5104  );
buf ( g5104 , n5105  );
buf ( g5105 , n5106  );
buf ( g5106 , n5107  );
buf ( g5107 , n5108  );
buf ( g5108 , n5109  );
buf ( g5109 , n5110  );
buf ( g5110 , n5111  );
buf ( g5111 , n5112  );
buf ( g5112 , n5113  );
buf ( g5113 , n5114  );
buf ( g5114 , n5115  );
buf ( g5115 , n5116  );
buf ( g5116 , n5117  );
buf ( g5117 , n5118  );
buf ( g5118 , n5119  );
buf ( g5119 , n5120  );
buf ( g5120 , n5121  );
buf ( g5121 , n5122  );
buf ( g5122 , n5123  );
buf ( g5123 , n5124  );
buf ( g5124 , n5125  );
buf ( g5125 , n5126  );
buf ( g5126 , n5127  );
buf ( g5127 , n5128  );
buf ( g5128 , n5129  );
buf ( g5129 , n5130  );
buf ( g5130 , n5131  );
buf ( g5131 , n5132  );
buf ( g5132 , n5133  );
buf ( g5133 , n5134  );
buf ( g5134 , n5135  );
buf ( g5135 , n5136  );
buf ( g5136 , n5137  );
buf ( g5137 , n5138  );
buf ( g5138 , n5139  );
buf ( g5139 , n5140  );
buf ( g5140 , n5141  );
buf ( g5141 , n5142  );
buf ( g5142 , n5143  );
buf ( g5143 , n5144  );
buf ( g5144 , n5145  );
buf ( g5145 , n5146  );
buf ( g5146 , n5147  );
buf ( g5147 , n5148  );
buf ( g5148 , n5149  );
buf ( g5149 , n5150  );
buf ( g5150 , n5151  );
buf ( g5151 , n5152  );
buf ( g5152 , n5153  );
buf ( g5153 , n5154  );
buf ( g5154 , n5155  );
buf ( g5155 , n5156  );
buf ( g5156 , n5157  );
buf ( g5157 , n5158  );
buf ( g5158 , n5159  );
buf ( g5159 , n5160  );
buf ( g5160 , n5161  );
buf ( g5161 , n5162  );
buf ( g5162 , n5163  );
buf ( g5163 , n5164  );
buf ( g5164 , n5165  );
buf ( g5165 , n5166  );
buf ( g5166 , n5167  );
buf ( g5167 , n5168  );
buf ( g5168 , n5169  );
buf ( g5169 , n5170  );
buf ( g5170 , n5171  );
buf ( g5171 , n5172  );
buf ( g5172 , n5173  );
buf ( g5173 , n5174  );
buf ( g5174 , n5175  );
buf ( g5175 , n5176  );
buf ( g5176 , n5177  );
buf ( g5177 , n5178  );
buf ( g5178 , n5179  );
buf ( g5179 , n5180  );
buf ( g5180 , n5181  );
buf ( g5181 , n5182  );
buf ( g5182 , n5183  );
buf ( g5183 , n5184  );
buf ( g5184 , n5185  );
buf ( g5185 , n5186  );
buf ( g5186 , n5187  );
buf ( g5187 , n5188  );
buf ( g5188 , n5189  );
buf ( g5189 , n5190  );
buf ( g5190 , n5191  );
buf ( g5191 , n5192  );
buf ( g5192 , n5193  );
buf ( g5193 , n5194  );
buf ( g5194 , n5195  );
buf ( g5195 , n5196  );
buf ( g5196 , n5197  );
buf ( g5197 , n5198  );
buf ( g5198 , n5199  );
buf ( g5199 , n5200  );
buf ( g5200 , n5201  );
buf ( g5201 , n5202  );
buf ( g5202 , n5203  );
buf ( g5203 , n5204  );
buf ( g5204 , n5205  );
buf ( g5205 , n5206  );
buf ( g5206 , n5207  );
buf ( g5207 , n5208  );
buf ( g5208 , n5209  );
buf ( g5209 , n5210  );
buf ( g5210 , n5211  );
buf ( g5211 , n5212  );
buf ( g5212 , n5213  );
buf ( g5213 , n5214  );
buf ( g5214 , n5215  );
buf ( g5215 , n5216  );
buf ( g5216 , n5217  );
buf ( g5217 , n5218  );
buf ( g5218 , n5219  );
buf ( g5219 , n5220  );
buf ( g5220 , n5221  );
buf ( g5221 , n5222  );
buf ( g5222 , n5223  );
buf ( g5223 , n5224  );
buf ( g5224 , n5225  );
buf ( g5225 , n5226  );
buf ( g5226 , n5227  );
buf ( g5227 , n5228  );
buf ( g5228 , n5229  );
buf ( g5229 , n5230  );
buf ( g5230 , n5231  );
buf ( g5231 , n5232  );
buf ( g5232 , n5233  );
buf ( g5233 , n5234  );
buf ( g5234 , n5235  );
buf ( g5235 , n5236  );
buf ( g5236 , n5237  );
buf ( g5237 , n5238  );
buf ( g5238 , n5239  );
buf ( g5239 , n5240  );
buf ( g5240 , n5241  );
buf ( g5241 , n5242  );
buf ( g5242 , n5243  );
buf ( g5243 , n5244  );
buf ( g5244 , n5245  );
buf ( g5245 , n5246  );
buf ( g5246 , n5247  );
buf ( g5247 , n5248  );
buf ( g5248 , n5249  );
buf ( g5249 , n5250  );
buf ( g5250 , n5251  );
buf ( g5251 , n5252  );
buf ( g5252 , n5253  );
buf ( g5253 , n5254  );
buf ( g5254 , n5255  );
buf ( g5255 , n5256  );
buf ( g5256 , n5257  );
buf ( g5257 , n5258  );
buf ( g5258 , n5259  );
buf ( g5259 , n5260  );
buf ( g5260 , n5261  );
buf ( g5261 , n5262  );
buf ( g5262 , n5263  );
buf ( g5263 , n5264  );
buf ( g5264 , n5265  );
buf ( g5265 , n5266  );
buf ( g5266 , n5267  );
buf ( g5267 , n5268  );
buf ( g5268 , n5269  );
buf ( g5269 , n5270  );
buf ( g5270 , n5271  );
buf ( g5271 , n5272  );
buf ( g5272 , n5273  );
buf ( g5273 , n5274  );
buf ( g5274 , n5275  );
buf ( g5275 , n5276  );
buf ( g5276 , n5277  );
buf ( g5277 , n5278  );
buf ( g5278 , n5279  );
buf ( g5279 , n5280  );
buf ( g5280 , n5281  );
buf ( g5281 , n5282  );
buf ( g5282 , n5283  );
buf ( g5283 , n5284  );
buf ( g5284 , n5285  );
buf ( g5285 , n5286  );
buf ( g5286 , n5287  );
buf ( g5287 , n5288  );
buf ( g5288 , n5289  );
buf ( g5289 , n5290  );
buf ( g5290 , n5291  );
buf ( g5291 , n5292  );
buf ( g5292 , n5293  );
buf ( g5293 , n5294  );
buf ( g5294 , n5295  );
buf ( g5295 , n5296  );
buf ( g5296 , n5297  );
buf ( g5297 , n5298  );
buf ( g5298 , n5299  );
buf ( g5299 , n5300  );
buf ( g5300 , n5301  );
buf ( g5301 , n5302  );
buf ( g5302 , n5303  );
buf ( g5303 , n5304  );
buf ( g5304 , n5305  );
buf ( g5305 , n5306  );
buf ( g5306 , n5307  );
buf ( g5307 , n5308  );
buf ( g5308 , n5309  );
buf ( g5309 , n5310  );
buf ( g5310 , n5311  );
buf ( g5311 , n5312  );
buf ( g5312 , n5313  );
buf ( g5313 , n5314  );
buf ( g5314 , n5315  );
buf ( g5315 , n5316  );
buf ( g5316 , n5317  );
buf ( g5317 , n5318  );
buf ( g5318 , n5319  );
buf ( g5319 , n5320  );
buf ( g5320 , n5321  );
buf ( g5321 , n5322  );
buf ( g5322 , n5323  );
buf ( g5323 , n5324  );
buf ( g5324 , n5325  );
buf ( g5325 , n5326  );
buf ( g5326 , n5327  );
buf ( g5327 , n5328  );
buf ( g5328 , n5329  );
buf ( g5329 , n5330  );
buf ( g5330 , n5331  );
buf ( g5331 , n5332  );
buf ( g5332 , n5333  );
buf ( g5333 , n5334  );
buf ( g5334 , n5335  );
buf ( g5335 , n5336  );
buf ( g5336 , n5337  );
buf ( g5337 , n5338  );
buf ( g5338 , n5339  );
buf ( g5339 , n5340  );
buf ( g5340 , n5341  );
buf ( g5341 , n5342  );
buf ( g5342 , n5343  );
buf ( g5343 , n5344  );
buf ( g5344 , n5345  );
buf ( g5345 , n5346  );
buf ( g5346 , n5347  );
buf ( g5347 , n5348  );
buf ( g5348 , n5349  );
buf ( g5349 , n5350  );
buf ( g5350 , n5351  );
buf ( g5351 , n5352  );
buf ( g5352 , n5353  );
buf ( g5353 , n5354  );
buf ( g5354 , n5355  );
buf ( g5355 , n5356  );
buf ( g5356 , n5357  );
buf ( g5357 , n5358  );
buf ( g5358 , n5359  );
buf ( g5359 , n5360  );
buf ( g5360 , n5361  );
buf ( g5361 , n5362  );
buf ( g5362 , n5363  );
buf ( g5363 , n5364  );
buf ( g5364 , n5365  );
buf ( g5365 , n5366  );
buf ( g5366 , n5367  );
buf ( g5367 , n5368  );
buf ( g5368 , n5369  );
buf ( g5369 , n5370  );
buf ( g5370 , n5371  );
buf ( g5371 , n5372  );
buf ( g5372 , n5373  );
buf ( g5373 , n5374  );
buf ( g5374 , n5375  );
buf ( g5375 , n5376  );
buf ( g5376 , n5377  );
buf ( g5377 , n5378  );
buf ( g5378 , n5379  );
buf ( g5379 , n5380  );
buf ( g5380 , n5381  );
buf ( g5381 , n5382  );
buf ( g5382 , n5383  );
buf ( g5383 , n5384  );
buf ( g5384 , n5385  );
buf ( g5385 , n5386  );
buf ( g5386 , n5387  );
buf ( g5387 , n5388  );
buf ( g5388 , n5389  );
buf ( g5389 , n5390  );
buf ( g5390 , n5391  );
buf ( g5391 , n5392  );
buf ( g5392 , n5393  );
buf ( g5393 , n5394  );
buf ( g5394 , n5395  );
buf ( g5395 , n5396  );
buf ( g5396 , n5397  );
buf ( g5397 , n5398  );
buf ( g5398 , n5399  );
buf ( g5399 , n5400  );
buf ( g5400 , n5401  );
buf ( g5401 , n5402  );
buf ( g5402 , n5403  );
buf ( g5403 , n5404  );
buf ( g5404 , n5405  );
buf ( g5405 , n5406  );
buf ( g5406 , n5407  );
buf ( g5407 , n5408  );
buf ( g5408 , n5409  );
buf ( g5409 , n5410  );
buf ( g5410 , n5411  );
buf ( g5411 , n5412  );
buf ( g5412 , n5413  );
buf ( g5413 , n5414  );
buf ( g5414 , n5415  );
buf ( g5415 , n5416  );
buf ( g5416 , n5417  );
buf ( g5417 , n5418  );
buf ( g5418 , n5419  );
buf ( g5419 , n5420  );
buf ( g5420 , n5421  );
buf ( g5421 , n5422  );
buf ( g5422 , n5423  );
buf ( g5423 , n5424  );
buf ( g5424 , n5425  );
buf ( g5425 , n5426  );
buf ( g5426 , n5427  );
buf ( g5427 , n5428  );
buf ( g5428 , n5429  );
buf ( g5429 , n5430  );
buf ( g5430 , n5431  );
buf ( g5431 , n5432  );
buf ( g5432 , n5433  );
buf ( g5433 , n5434  );
buf ( g5434 , n5435  );
buf ( g5435 , n5436  );
buf ( g5436 , n5437  );
buf ( g5437 , n5438  );
buf ( g5438 , n5439  );
buf ( g5439 , n5440  );
buf ( g5440 , n5441  );
buf ( g5441 , n5442  );
buf ( g5442 , n5443  );
buf ( g5443 , n5444  );
buf ( g5444 , n5445  );
buf ( g5445 , n5446  );
buf ( g5446 , n5447  );
buf ( g5447 , n5448  );
buf ( g5448 , n5449  );
buf ( g5449 , n5450  );
buf ( g5450 , n5451  );
buf ( g5451 , n5452  );
buf ( g5452 , n5453  );
buf ( g5453 , n5454  );
buf ( g5454 , n5455  );
buf ( g5455 , n5456  );
buf ( g5456 , n5457  );
buf ( g5457 , n5458  );
buf ( g5458 , n5459  );
buf ( g5459 , n5460  );
buf ( g5460 , n5461  );
buf ( g5461 , n5462  );
buf ( g5462 , n5463  );
buf ( g5463 , n5464  );
buf ( g5464 , n5465  );
buf ( g5465 , n5466  );
buf ( g5466 , n5467  );
buf ( g5467 , n5468  );
buf ( g5468 , n5469  );
buf ( g5469 , n5470  );
buf ( g5470 , n5471  );
buf ( g5471 , n5472  );
buf ( g5472 , n5473  );
buf ( g5473 , n5474  );
buf ( g5474 , n5475  );
buf ( g5475 , n5476  );
buf ( g5476 , n5477  );
buf ( g5477 , n5478  );
buf ( g5478 , n5479  );
buf ( g5479 , n5480  );
buf ( g5480 , n5481  );
buf ( g5481 , n5482  );
buf ( g5482 , n5483  );
buf ( g5483 , n5484  );
buf ( g5484 , n5485  );
buf ( g5485 , n5486  );
buf ( g5486 , n5487  );
buf ( g5487 , n5488  );
buf ( g5488 , n5489  );
buf ( g5489 , n5490  );
buf ( g5490 , n5491  );
buf ( g5491 , n5492  );
buf ( g5492 , n5493  );
buf ( g5493 , n5494  );
buf ( g5494 , n5495  );
buf ( g5495 , n5496  );
buf ( g5496 , n5497  );
buf ( g5497 , n5498  );
buf ( g5498 , n5499  );
buf ( g5499 , n5500  );
buf ( g5500 , n5501  );
buf ( g5501 , n5502  );
buf ( g5502 , n5503  );
buf ( g5503 , n5504  );
buf ( g5504 , n5505  );
buf ( g5505 , n5506  );
buf ( g5506 , n5507  );
buf ( g5507 , n5508  );
buf ( g5508 , n5509  );
buf ( g5509 , n5510  );
buf ( g5510 , n5511  );
buf ( g5511 , n5512  );
buf ( g5512 , n5513  );
buf ( g5513 , n5514  );
buf ( g5514 , n5515  );
buf ( g5515 , n5516  );
buf ( g5516 , n5517  );
buf ( g5517 , n5518  );
buf ( g5518 , n5519  );
buf ( g5519 , n5520  );
buf ( g5520 , n5521  );
buf ( g5521 , n5522  );
buf ( g5522 , n5523  );
buf ( g5523 , n5524  );
buf ( g5524 , n5525  );
buf ( g5525 , n5526  );
buf ( g5526 , n5527  );
buf ( g5527 , n5528  );
buf ( g5528 , n5529  );
buf ( g5529 , n5530  );
buf ( g5530 , n5531  );
buf ( g5531 , n5532  );
buf ( g5532 , n5533  );
buf ( g5533 , n5534  );
buf ( g5534 , n5535  );
buf ( g5535 , n5536  );
buf ( g5536 , n5537  );
buf ( g5537 , n5538  );
buf ( g5538 , n5539  );
buf ( g5539 , n5540  );
buf ( g5540 , n5541  );
buf ( g5541 , n5542  );
buf ( g5542 , n5543  );
buf ( g5543 , n5544  );
buf ( g5544 , n5545  );
buf ( g5545 , n5546  );
buf ( g5546 , n5547  );
buf ( g5547 , n5548  );
buf ( g5548 , n5549  );
buf ( g5549 , n5550  );
buf ( g5550 , n5551  );
buf ( g5551 , n5552  );
buf ( g5552 , n5553  );
buf ( g5553 , n5554  );
buf ( g5554 , n5555  );
buf ( g5555 , n5556  );
buf ( g5556 , n5557  );
buf ( g5557 , n5558  );
buf ( g5558 , n5559  );
buf ( g5559 , n5560  );
buf ( g5560 , n5561  );
buf ( g5561 , n5562  );
buf ( g5562 , n5563  );
buf ( g5563 , n5564  );
buf ( g5564 , n5565  );
buf ( g5565 , n5566  );
buf ( g5566 , n5567  );
buf ( g5567 , n5568  );
buf ( g5568 , n5569  );
buf ( g5569 , n5570  );
buf ( g5570 , n5571  );
buf ( g5571 , n5572  );
buf ( g5572 , n5573  );
buf ( g5573 , n5574  );
buf ( g5574 , n5575  );
buf ( g5575 , n5576  );
buf ( g5576 , n5577  );
buf ( g5577 , n5578  );
buf ( g5578 , n5579  );
buf ( g5579 , n5580  );
buf ( g5580 , n5581  );
buf ( g5581 , n5582  );
buf ( g5582 , n5583  );
buf ( g5583 , n5584  );
buf ( g5584 , n5585  );
buf ( g5585 , n5586  );
buf ( g5586 , n5587  );
buf ( g5587 , n5588  );
buf ( g5588 , n5589  );
buf ( g5589 , n5590  );
buf ( g5590 , n5591  );
buf ( g5591 , n5592  );
buf ( g5592 , n5593  );
buf ( g5593 , n5594  );
buf ( g5594 , n5595  );
buf ( g5595 , n5596  );
buf ( g5596 , n5597  );
buf ( g5597 , n5598  );
buf ( g5598 , n5599  );
buf ( g5599 , n5600  );
buf ( g5600 , n5601  );
buf ( g5601 , n5602  );
buf ( g5602 , n5603  );
buf ( g5603 , n5604  );
buf ( g5604 , n5605  );
buf ( g5605 , n5606  );
buf ( g5606 , n5607  );
buf ( g5607 , n5608  );
buf ( g5608 , n5609  );
buf ( g5609 , n5610  );
buf ( g5610 , n5611  );
buf ( g5611 , n5612  );
buf ( g5612 , n5613  );
buf ( g5613 , n5614  );
buf ( g5614 , n5615  );
buf ( g5615 , n5616  );
buf ( g5616 , n5617  );
buf ( g5617 , n5618  );
buf ( g5618 , n5619  );
buf ( g5619 , n5620  );
buf ( g5620 , n5621  );
buf ( g5621 , n5622  );
buf ( g5622 , n5623  );
buf ( g5623 , n5624  );
buf ( g5624 , n5625  );
buf ( g5625 , n5626  );
buf ( g5626 , n5627  );
buf ( g5627 , n5628  );
buf ( g5628 , n5629  );
buf ( g5629 , n5630  );
buf ( g5630 , n5631  );
buf ( g5631 , n5632  );
buf ( g5632 , n5633  );
buf ( g5633 , n5634  );
buf ( g5634 , n5635  );
buf ( g5635 , n5636  );
buf ( g5636 , n5637  );
buf ( g5637 , n5638  );
buf ( g5638 , n5639  );
buf ( g5639 , n5640  );
buf ( g5640 , n5641  );
buf ( g5641 , n5642  );
buf ( g5642 , n5643  );
buf ( g5643 , n5644  );
buf ( g5644 , n5645  );
buf ( g5645 , n5646  );
buf ( g5646 , n5647  );
buf ( g5647 , n5648  );
buf ( g5648 , n5649  );
buf ( g5649 , n5650  );
buf ( g5650 , n5651  );
buf ( g5651 , n5652  );
buf ( g5652 , n5653  );
buf ( g5653 , n5654  );
buf ( g5654 , n5655  );
buf ( g5655 , n5656  );
buf ( g5656 , n5657  );
buf ( g5657 , n5658  );
buf ( g5658 , n5659  );
buf ( g5659 , n5660  );
buf ( g5660 , n5661  );
buf ( g5661 , n5662  );
buf ( g5662 , n5663  );
buf ( g5663 , n5664  );
buf ( g5664 , n5665  );
buf ( g5665 , n5666  );
buf ( g5666 , n5667  );
buf ( g5667 , n5668  );
buf ( g5668 , n5669  );
buf ( g5669 , n5670  );
buf ( g5670 , n5671  );
buf ( g5671 , n5672  );
buf ( g5672 , n5673  );
buf ( g5673 , n5674  );
buf ( g5674 , n5675  );
buf ( g5675 , n5676  );
buf ( g5676 , n5677  );
buf ( g5677 , n5678  );
buf ( g5678 , n5679  );
buf ( g5679 , n5680  );
buf ( g5680 , n5681  );
buf ( g5681 , n5682  );
buf ( g5682 , n5683  );
buf ( g5683 , n5684  );
buf ( g5684 , n5685  );
buf ( g5685 , n5686  );
buf ( g5686 , n5687  );
buf ( g5687 , n5688  );
buf ( g5688 , n5689  );
buf ( g5689 , n5690  );
buf ( g5690 , n5691  );
buf ( g5691 , n5692  );
buf ( g5692 , n5693  );
buf ( g5693 , n5694  );
buf ( g5694 , n5695  );
buf ( g5695 , n5696  );
buf ( g5696 , n5697  );
buf ( g5697 , n5698  );
buf ( g5698 , n5699  );
buf ( g5699 , n5700  );
buf ( g5700 , n5701  );
buf ( g5701 , n5702  );
buf ( g5702 , n5703  );
buf ( g5703 , n5704  );
buf ( g5704 , n5705  );
buf ( g5705 , n5706  );
buf ( g5706 , n5707  );
buf ( g5707 , n5708  );
buf ( g5708 , n5709  );
buf ( g5709 , n5710  );
buf ( g5710 , n5711  );
buf ( g5711 , n5712  );
buf ( g5712 , n5713  );
buf ( g5713 , n5714  );
buf ( g5714 , n5715  );
buf ( g5715 , n5716  );
buf ( g5716 , n5717  );
buf ( g5717 , n5718  );
buf ( g5718 , n5719  );
buf ( g5719 , n5720  );
buf ( g5720 , n5721  );
buf ( g5721 , n5722  );
buf ( g5722 , n5723  );
buf ( g5723 , n5724  );
buf ( g5724 , n5725  );
buf ( g5725 , n5726  );
buf ( g5726 , n5727  );
buf ( g5727 , n5728  );
buf ( g5728 , n5729  );
buf ( g5729 , n5730  );
buf ( g5730 , n5731  );
buf ( g5731 , n5732  );
buf ( g5732 , n5733  );
buf ( g5733 , n5734  );
buf ( g5734 , n5735  );
buf ( g5735 , n5736  );
buf ( g5736 , n5737  );
buf ( g5737 , n5738  );
buf ( g5738 , n5739  );
buf ( g5739 , n5740  );
buf ( g5740 , n5741  );
buf ( g5741 , n5742  );
buf ( g5742 , n5743  );
buf ( g5743 , n5744  );
buf ( g5744 , n5745  );
buf ( g5745 , n5746  );
buf ( g5746 , n5747  );
buf ( g5747 , n5748  );
buf ( g5748 , n5749  );
buf ( g5749 , n5750  );
buf ( g5750 , n5751  );
buf ( g5751 , n5752  );
buf ( g5752 , n5753  );
buf ( g5753 , n5754  );
buf ( g5754 , n5755  );
buf ( g5755 , n5756  );
buf ( g5756 , n5757  );
buf ( g5757 , n5758  );
buf ( g5758 , n5759  );
buf ( g5759 , n5760  );
buf ( g5760 , n5761  );
buf ( g5761 , n5762  );
buf ( g5762 , n5763  );
buf ( g5763 , n5764  );
buf ( g5764 , n5765  );
buf ( g5765 , n5766  );
buf ( g5766 , n5767  );
buf ( g5767 , n5768  );
buf ( g5768 , n5769  );
buf ( g5769 , n5770  );
buf ( g5770 , n5771  );
buf ( g5771 , n5772  );
buf ( g5772 , n5773  );
buf ( g5773 , n5774  );
buf ( g5774 , n5775  );
buf ( g5775 , n5776  );
buf ( g5776 , n5777  );
buf ( g5777 , n5778  );
buf ( g5778 , n5779  );
buf ( g5779 , n5780  );
buf ( g5780 , n5781  );
buf ( g5781 , n5782  );
buf ( g5782 , n5783  );
buf ( g5783 , n5784  );
buf ( g5784 , n5785  );
buf ( g5785 , n5786  );
buf ( g5786 , n5787  );
buf ( g5787 , n5788  );
buf ( g5788 , n5789  );
buf ( g5789 , n5790  );
buf ( g5790 , n5791  );
buf ( g5791 , n5792  );
buf ( g5792 , n5793  );
buf ( g5793 , n5794  );
buf ( g5794 , n5795  );
buf ( g5795 , n5796  );
buf ( g5796 , n5797  );
buf ( g5797 , n5798  );
buf ( g5798 , n5799  );
buf ( g5799 , n5800  );
buf ( g5800 , n5801  );
buf ( g5801 , n5802  );
buf ( g5802 , n5803  );
buf ( g5803 , n5804  );
buf ( g5804 , n5805  );
buf ( g5805 , n5806  );
buf ( g5806 , n5807  );
buf ( g5807 , n5808  );
buf ( g5808 , n5809  );
buf ( g5809 , n5810  );
buf ( g5810 , n5811  );
buf ( g5811 , n5812  );
buf ( g5812 , n5813  );
buf ( g5813 , n5814  );
buf ( g5814 , n5815  );
buf ( g5815 , n5816  );
buf ( g5816 , n5817  );
buf ( g5817 , n5818  );
buf ( g5818 , n5819  );
buf ( g5819 , n5820  );
buf ( g5820 , n5821  );
buf ( g5821 , n5822  );
buf ( g5822 , n5823  );
buf ( g5823 , n5824  );
buf ( g5824 , n5825  );
buf ( g5825 , n5826  );
buf ( g5826 , n5827  );
buf ( g5827 , n5828  );
buf ( g5828 , n5829  );
buf ( g5829 , n5830  );
buf ( g5830 , n5831  );
buf ( g5831 , n5832  );
buf ( g5832 , n5833  );
buf ( g5833 , n5834  );
buf ( g5834 , n5835  );
buf ( g5835 , n5836  );
buf ( g5836 , n5837  );
buf ( g5837 , n5838  );
buf ( g5838 , n5839  );
buf ( g5839 , n5840  );
buf ( g5840 , n5841  );
buf ( g5841 , n5842  );
buf ( g5842 , n5843  );
buf ( g5843 , n5844  );
buf ( g5844 , n5845  );
buf ( g5845 , n5846  );
buf ( g5846 , n5847  );
buf ( g5847 , n5848  );
buf ( g5848 , n5849  );
buf ( g5849 , n5850  );
buf ( g5850 , n5851  );
buf ( g5851 , n5852  );
buf ( g5852 , n5853  );
buf ( g5853 , n5854  );
buf ( g5854 , n5855  );
buf ( g5855 , n5856  );
buf ( g5856 , n5857  );
buf ( g5857 , n5858  );
buf ( g5858 , n5859  );
buf ( g5859 , n5860  );
buf ( g5860 , n5861  );
buf ( g5861 , n5862  );
buf ( g5862 , n5863  );
buf ( g5863 , n5864  );
buf ( g5864 , n5865  );
buf ( g5865 , n5866  );
buf ( g5866 , n5867  );
buf ( g5867 , n5868  );
buf ( g5868 , n5869  );
buf ( g5869 , n5870  );
buf ( g5870 , n5871  );
buf ( g5871 , n5872  );
buf ( g5872 , n5873  );
buf ( g5873 , n5874  );
buf ( g5874 , n5875  );
buf ( g5875 , n5876  );
buf ( g5876 , n5877  );
buf ( g5877 , n5878  );
buf ( g5878 , n5879  );
buf ( g5879 , n5880  );
buf ( g5880 , n5881  );
buf ( g5881 , n5882  );
buf ( g5882 , n5883  );
buf ( g5883 , n5884  );
buf ( g5884 , n5885  );
buf ( g5885 , n5886  );
buf ( g5886 , n5887  );
buf ( g5887 , n5888  );
buf ( g5888 , n5889  );
buf ( g5889 , n5890  );
buf ( g5890 , n5891  );
buf ( g5891 , n5892  );
buf ( g5892 , n5893  );
buf ( g5893 , n5894  );
buf ( g5894 , n5895  );
buf ( g5895 , n5896  );
buf ( g5896 , n5897  );
buf ( g5897 , n5898  );
buf ( g5898 , n5899  );
buf ( g5899 , n5900  );
buf ( g5900 , n5901  );
buf ( g5901 , n5902  );
buf ( g5902 , n5903  );
buf ( g5903 , n5904  );
buf ( g5904 , n5905  );
buf ( g5905 , n5906  );
buf ( g5906 , n5907  );
buf ( g5907 , n5908  );
buf ( g5908 , n5909  );
buf ( g5909 , n5910  );
buf ( g5910 , n5911  );
buf ( g5911 , n5912  );
buf ( g5912 , n5913  );
buf ( g5913 , n5914  );
buf ( g5914 , n5915  );
buf ( g5915 , n5916  );
buf ( g5916 , n5917  );
buf ( g5917 , n5918  );
buf ( g5918 , n5919  );
buf ( g5919 , n5920  );
buf ( g5920 , n5921  );
buf ( g5921 , n5922  );
buf ( g5922 , n5923  );
buf ( g5923 , n5924  );
buf ( g5924 , n5925  );
buf ( g5925 , n5926  );
buf ( g5926 , n5927  );
buf ( g5927 , n5928  );
buf ( g5928 , n5929  );
buf ( g5929 , n5930  );
buf ( g5930 , n5931  );
buf ( g5931 , n5932  );
buf ( g5932 , n5933  );
buf ( g5933 , n5934  );
buf ( g5934 , n5935  );
buf ( g5935 , n5936  );
buf ( g5936 , n5937  );
buf ( g5937 , n5938  );
buf ( g5938 , n5939  );
buf ( g5939 , n5940  );
buf ( g5940 , n5941  );
buf ( g5941 , n5942  );
buf ( g5942 , n5943  );
buf ( g5943 , n5944  );
buf ( g5944 , n5945  );
buf ( g5945 , n5946  );
buf ( g5946 , n5947  );
buf ( g5947 , n5948  );
buf ( g5948 , n5949  );
buf ( g5949 , n5950  );
buf ( g5950 , n5951  );
buf ( g5951 , n5952  );
buf ( g5952 , n5953  );
buf ( g5953 , n5954  );
buf ( g5954 , n5955  );
buf ( g5955 , n5956  );
buf ( g5956 , n5957  );
buf ( g5957 , n5958  );
buf ( g5958 , n5959  );
buf ( g5959 , n5960  );
buf ( g5960 , n5961  );
buf ( g5961 , n5962  );
buf ( g5962 , n5963  );
buf ( g5963 , n5964  );
buf ( g5964 , n5965  );
buf ( g5965 , n5966  );
buf ( g5966 , n5967  );
buf ( g5967 , n5968  );
buf ( g5968 , n5969  );
buf ( g5969 , n5970  );
buf ( g5970 , n5971  );
buf ( g5971 , n5972  );
buf ( g5972 , n5973  );
buf ( g5973 , n5974  );
buf ( g5974 , n5975  );
buf ( g5975 , n5976  );
buf ( g5976 , n5977  );
buf ( g5977 , n5978  );
buf ( g5978 , n5979  );
buf ( g5979 , n5980  );
buf ( g5980 , n5981  );
buf ( g5981 , n5982  );
buf ( g5982 , n5983  );
buf ( g5983 , n5984  );
buf ( g5984 , n5985  );
buf ( g5985 , n5986  );
buf ( g5986 , n5987  );
buf ( g5987 , n5988  );
buf ( g5988 , n5989  );
buf ( g5989 , n5990  );
buf ( g5990 , n5991  );
buf ( g5991 , n5992  );
buf ( g5992 , n5993  );
buf ( g5993 , n5994  );
buf ( g5994 , n5995  );
buf ( g5995 , n5996  );
buf ( g5996 , n5997  );
buf ( g5997 , n5998  );
buf ( g5998 , n5999  );
buf ( g5999 , n6000  );
buf ( g6000 , n6001  );
buf ( g6001 , n6002  );
buf ( g6002 , n6003  );
buf ( g6003 , n6004  );
buf ( g6004 , n6005  );
buf ( g6005 , n6006  );
buf ( g6006 , n6007  );
buf ( g6007 , n6008  );
buf ( g6008 , n6009  );
buf ( g6009 , n6010  );
buf ( g6010 , n6011  );
buf ( g6011 , n6012  );
buf ( g6012 , n6013  );
buf ( g6013 , n6014  );
buf ( g6014 , n6015  );
buf ( g6015 , n6016  );
buf ( g6016 , n6017  );
buf ( g6017 , n6018  );
buf ( g6018 , n6019  );
buf ( g6019 , n6020  );
buf ( g6020 , n6021  );
buf ( g6021 , n6022  );
buf ( g6022 , n6023  );
buf ( g6023 , n6024  );
buf ( g6024 , n6025  );
buf ( g6025 , n6026  );
buf ( g6026 , n6027  );
buf ( g6027 , n6028  );
buf ( g6028 , n6029  );
buf ( g6029 , n6030  );
buf ( g6030 , n6031  );
buf ( g6031 , n6032  );
buf ( g6032 , n6033  );
buf ( g6033 , n6034  );
buf ( g6034 , n6035  );
buf ( g6035 , n6036  );
buf ( g6036 , n6037  );
buf ( g6037 , n6038  );
buf ( g6038 , n6039  );
buf ( g6039 , n6040  );
buf ( g6040 , n6041  );
buf ( g6041 , n6042  );
buf ( g6042 , n6043  );
buf ( g6043 , n6044  );
buf ( g6044 , n6045  );
buf ( g6045 , n6046  );
buf ( g6046 , n6047  );
buf ( g6047 , n6048  );
buf ( g6048 , n6049  );
buf ( g6049 , n6050  );
buf ( g6050 , n6051  );
buf ( g6051 , n6052  );
buf ( g6052 , n6053  );
buf ( g6053 , n6054  );
buf ( g6054 , n6055  );
buf ( g6055 , n6056  );
buf ( g6056 , n6057  );
buf ( g6057 , n6058  );
buf ( g6058 , n6059  );
buf ( g6059 , n6060  );
buf ( g6060 , n6061  );
buf ( g6061 , n6062  );
buf ( g6062 , n6063  );
buf ( g6063 , n6064  );
buf ( g6064 , n6065  );
buf ( g6065 , n6066  );
buf ( g6066 , n6067  );
buf ( g6067 , n6068  );
buf ( g6068 , n6069  );
buf ( g6069 , n6070  );
buf ( g6070 , n6071  );
buf ( g6071 , n6072  );
buf ( g6072 , n6073  );
buf ( g6073 , n6074  );
buf ( g6074 , n6075  );
buf ( g6075 , n6076  );
buf ( g6076 , n6077  );
buf ( g6077 , n6078  );
buf ( g6078 , n6079  );
buf ( g6079 , n6080  );
buf ( g6080 , n6081  );
buf ( g6081 , n6082  );
buf ( g6082 , n6083  );
buf ( g6083 , n6084  );
buf ( g6084 , n6085  );
buf ( g6085 , n6086  );
buf ( g6086 , n6087  );
buf ( g6087 , n6088  );
buf ( g6088 , n6089  );
buf ( g6089 , n6090  );
buf ( g6090 , n6091  );
buf ( g6091 , n6092  );
buf ( g6092 , n6093  );
buf ( g6093 , n6094  );
buf ( g6094 , n6095  );
buf ( g6095 , n6096  );
buf ( g6096 , n6097  );
buf ( g6097 , n6098  );
buf ( g6098 , n6099  );
buf ( g6099 , n6100  );
buf ( g6100 , n6101  );
buf ( g6101 , n6102  );
buf ( g6102 , n6103  );
buf ( g6103 , n6104  );
buf ( g6104 , n6105  );
buf ( g6105 , n6106  );
buf ( g6106 , n6107  );
buf ( g6107 , n6108  );
buf ( g6108 , n6109  );
buf ( g6109 , n6110  );
buf ( g6110 , n6111  );
buf ( g6111 , n6112  );
buf ( g6112 , n6113  );
buf ( g6113 , n6114  );
buf ( g6114 , n6115  );
buf ( g6115 , n6116  );
buf ( g6116 , n6117  );
buf ( g6117 , n6118  );
buf ( g6118 , n6119  );
buf ( g6119 , n6120  );
buf ( g6120 , n6121  );
buf ( g6121 , n6122  );
buf ( g6122 , n6123  );
buf ( g6123 , n6124  );
buf ( g6124 , n6125  );
buf ( g6125 , n6126  );
buf ( g6126 , n6127  );
buf ( g6127 , n6128  );
buf ( g6128 , n6129  );
buf ( g6129 , n6130  );
buf ( g6130 , n6131  );
buf ( g6131 , n6132  );
buf ( g6132 , n6133  );
buf ( g6133 , n6134  );
buf ( g6134 , n6135  );
buf ( g6135 , n6136  );
buf ( g6136 , n6137  );
buf ( g6137 , n6138  );
buf ( g6138 , n6139  );
buf ( g6139 , n6140  );
buf ( g6140 , n6141  );
buf ( g6141 , n6142  );
buf ( g6142 , n6143  );
buf ( g6143 , n6144  );
buf ( g6144 , n6145  );
buf ( g6145 , n6146  );
buf ( g6146 , n6147  );
buf ( g6147 , n6148  );
buf ( g6148 , n6149  );
buf ( g6149 , n6150  );
buf ( g6150 , n6151  );
buf ( g6151 , n6152  );
buf ( g6152 , n6153  );
buf ( g6153 , n6154  );
buf ( g6154 , n6155  );
buf ( g6155 , n6156  );
buf ( g6156 , n6157  );
buf ( g6157 , n6158  );
buf ( g6158 , n6159  );
buf ( g6159 , n6160  );
buf ( g6160 , n6161  );
buf ( g6161 , n6162  );
buf ( g6162 , n6163  );
buf ( g6163 , n6164  );
buf ( g6164 , n6165  );
buf ( g6165 , n6166  );
buf ( g6166 , n6167  );
buf ( g6167 , n6168  );
buf ( g6168 , n6169  );
buf ( g6169 , n6170  );
buf ( g6170 , n6171  );
buf ( g6171 , n6172  );
buf ( g6172 , n6173  );
buf ( g6173 , n6174  );
buf ( g6174 , n6175  );
buf ( g6175 , n6176  );
buf ( g6176 , n6177  );
buf ( g6177 , n6178  );
buf ( g6178 , n6179  );
buf ( g6179 , n6180  );
buf ( g6180 , n6181  );
buf ( g6181 , n6182  );
buf ( g6182 , n6183  );
buf ( g6183 , n6184  );
buf ( g6184 , n6185  );
buf ( g6185 , n6186  );
buf ( g6186 , n6187  );
buf ( g6187 , n6188  );
buf ( g6188 , n6189  );
buf ( g6189 , n6190  );
buf ( g6190 , n6191  );
buf ( g6191 , n6192  );
buf ( g6192 , n6193  );
buf ( g6193 , n6194  );
buf ( g6194 , n6195  );
buf ( g6195 , n6196  );
buf ( g6196 , n6197  );
buf ( g6197 , n6198  );
buf ( g6198 , n6199  );
buf ( g6199 , n6200  );
buf ( g6200 , n6201  );
buf ( g6201 , n6202  );
buf ( g6202 , n6203  );
buf ( g6203 , n6204  );
buf ( g6204 , n6205  );
buf ( g6205 , n6206  );
buf ( g6206 , n6207  );
buf ( g6207 , n6208  );
buf ( g6208 , n6209  );
buf ( g6209 , n6210  );
buf ( g6210 , n6211  );
buf ( g6211 , n6212  );
buf ( g6212 , n6213  );
buf ( g6213 , n6214  );
buf ( g6214 , n6215  );
buf ( g6215 , n6216  );
buf ( g6216 , n6217  );
buf ( g6217 , n6218  );
buf ( g6218 , n6219  );
buf ( g6219 , n6220  );
buf ( g6220 , n6221  );
buf ( g6221 , n6222  );
buf ( g6222 , n6223  );
buf ( g6223 , n6224  );
buf ( g6224 , n6225  );
buf ( g6225 , n6226  );
buf ( g6226 , n6227  );
buf ( g6227 , n6228  );
buf ( g6228 , n6229  );
buf ( g6229 , n6230  );
buf ( g6230 , n6231  );
buf ( g6231 , n6232  );
buf ( g6232 , n6233  );
buf ( g6233 , n6234  );
buf ( g6234 , n6235  );
buf ( g6235 , n6236  );
buf ( g6236 , n6237  );
buf ( g6237 , n6238  );
buf ( g6238 , n6239  );
buf ( g6239 , n6240  );
buf ( g6240 , n6241  );
buf ( g6241 , n6242  );
buf ( g6242 , n6243  );
buf ( g6243 , n6244  );
buf ( g6244 , n6245  );
buf ( g6245 , n6246  );
buf ( g6246 , n6247  );
buf ( g6247 , n6248  );
buf ( g6248 , n6249  );
buf ( g6249 , n6250  );
buf ( g6250 , n6251  );
buf ( g6251 , n6252  );
buf ( g6252 , n6253  );
buf ( g6253 , n6254  );
buf ( g6254 , n6255  );
buf ( g6255 , n6256  );
buf ( g6256 , n6257  );
buf ( g6257 , n6258  );
buf ( g6258 , n6259  );
buf ( g6259 , n6260  );
buf ( g6260 , n6261  );
buf ( g6261 , n6262  );
buf ( g6262 , n6263  );
buf ( g6263 , n6264  );
buf ( g6264 , n6265  );
buf ( g6265 , n6266  );
buf ( g6266 , n6267  );
buf ( g6267 , n6268  );
buf ( g6268 , n6269  );
buf ( g6269 , n6270  );
buf ( g6270 , n6271  );
buf ( g6271 , n6272  );
buf ( g6272 , n6273  );
buf ( g6273 , n6274  );
buf ( g6274 , n6275  );
buf ( g6275 , n6276  );
buf ( g6276 , n6277  );
buf ( g6277 , n6278  );
buf ( g6278 , n6279  );
buf ( g6279 , n6280  );
buf ( g6280 , n6281  );
buf ( g6281 , n6282  );
buf ( g6282 , n6283  );
buf ( g6283 , n6284  );
buf ( g6284 , n6285  );
buf ( g6285 , n6286  );
buf ( g6286 , n6287  );
buf ( g6287 , n6288  );
buf ( g6288 , n6289  );
buf ( g6289 , n6290  );
buf ( g6290 , n6291  );
buf ( g6291 , n6292  );
buf ( g6292 , n6293  );
buf ( g6293 , n6294  );
buf ( g6294 , n6295  );
buf ( g6295 , n6296  );
buf ( g6296 , n6297  );
buf ( g6297 , n6298  );
buf ( g6298 , n6299  );
buf ( g6299 , n6300  );
buf ( g6300 , n6301  );
buf ( g6301 , n6302  );
buf ( g6302 , n6303  );
buf ( g6303 , n6304  );
buf ( g6304 , n6305  );
buf ( g6305 , n6306  );
buf ( g6306 , n6307  );
buf ( g6307 , n6308  );
buf ( g6308 , n6309  );
buf ( g6309 , n6310  );
buf ( g6310 , n6311  );
buf ( g6311 , n6312  );
buf ( g6312 , n6313  );
buf ( g6313 , n6314  );
buf ( g6314 , n6315  );
buf ( g6315 , n6316  );
buf ( g6316 , n6317  );
buf ( g6317 , n6318  );
buf ( g6318 , n6319  );
buf ( g6319 , n6320  );
buf ( g6320 , n6321  );
buf ( g6321 , n6322  );
buf ( g6322 , n6323  );
buf ( g6323 , n6324  );
buf ( g6324 , n6325  );
buf ( g6325 , n6326  );
buf ( g6326 , n6327  );
buf ( g6327 , n6328  );
buf ( g6328 , n6329  );
buf ( g6329 , n6330  );
buf ( g6330 , n6331  );
buf ( g6331 , n6332  );
buf ( g6332 , n6333  );
buf ( g6333 , n6334  );
buf ( g6334 , n6335  );
buf ( g6335 , n6336  );
buf ( g6336 , n6337  );
buf ( g6337 , n6338  );
buf ( g6338 , n6339  );
buf ( g6339 , n6340  );
buf ( g6340 , n6341  );
buf ( g6341 , n6342  );
buf ( g6342 , n6343  );
buf ( g6343 , n6344  );
buf ( g6344 , n6345  );
buf ( g6345 , n6346  );
buf ( g6346 , n6347  );
buf ( g6347 , n6348  );
buf ( g6348 , n6349  );
buf ( g6349 , n6350  );
buf ( g6350 , n6351  );
buf ( g6351 , n6352  );
buf ( g6352 , n6353  );
buf ( g6353 , n6354  );
buf ( g6354 , n6355  );
buf ( g6355 , n6356  );
buf ( g6356 , n6357  );
buf ( g6357 , n6358  );
buf ( g6358 , n6359  );
buf ( g6359 , n6360  );
buf ( g6360 , n6361  );
buf ( g6361 , n6362  );
buf ( g6362 , n6363  );
buf ( g6363 , n6364  );
buf ( g6364 , n6365  );
buf ( g6365 , n6366  );
buf ( g6366 , n6367  );
buf ( g6367 , n6368  );
buf ( g6368 , n6369  );
buf ( g6369 , n6370  );
buf ( g6370 , n6371  );
buf ( g6371 , n6372  );
buf ( g6372 , n6373  );
buf ( g6373 , n6374  );
buf ( g6374 , n6375  );
buf ( g6375 , n6376  );
buf ( g6376 , n6377  );
buf ( g6377 , n6378  );
buf ( g6378 , n6379  );
buf ( g6379 , n6380  );
buf ( g6380 , n6381  );
buf ( g6381 , n6382  );
buf ( g6382 , n6383  );
buf ( g6383 , n6384  );
buf ( g6384 , n6385  );
buf ( g6385 , n6386  );
buf ( g6386 , n6387  );
buf ( g6387 , n6388  );
buf ( g6388 , n6389  );
buf ( g6389 , n6390  );
buf ( g6390 , n6391  );
buf ( g6391 , n6392  );
buf ( g6392 , n6393  );
buf ( g6393 , n6394  );
buf ( g6394 , n6395  );
buf ( g6395 , n6396  );
buf ( g6396 , n6397  );
buf ( g6397 , n6398  );
buf ( g6398 , n6399  );
buf ( g6399 , n6400  );
buf ( g6400 , n6401  );
buf ( g6401 , n6402  );
buf ( g6402 , n6403  );
buf ( g6403 , n6404  );
buf ( g6404 , n6405  );
buf ( g6405 , n6406  );
buf ( g6406 , n6407  );
buf ( g6407 , n6408  );
buf ( g6408 , n6409  );
buf ( g6409 , n6410  );
buf ( g6410 , n6411  );
buf ( g6411 , n6412  );
buf ( g6412 , n6413  );
buf ( g6413 , n6414  );
buf ( g6414 , n6415  );
buf ( g6415 , n6416  );
buf ( g6416 , n6417  );
buf ( g6417 , n6418  );
buf ( g6418 , n6419  );
buf ( g6419 , n6420  );
buf ( g6420 , n6421  );
buf ( g6421 , n6422  );
buf ( g6422 , n6423  );
buf ( g6423 , n6424  );
buf ( g6424 , n6425  );
buf ( g6425 , n6426  );
buf ( g6426 , n6427  );
buf ( g6427 , n6428  );
buf ( g6428 , n6429  );
buf ( g6429 , n6430  );
buf ( g6430 , n6431  );
buf ( g6431 , n6432  );
buf ( g6432 , n6433  );
buf ( g6433 , n6434  );
buf ( g6434 , n6435  );
buf ( g6435 , n6436  );
buf ( g6436 , n6437  );
buf ( g6437 , n6438  );
buf ( g6438 , n6439  );
buf ( g6439 , n6440  );
buf ( g6440 , n6441  );
buf ( g6441 , n6442  );
buf ( g6442 , n6443  );
buf ( g6443 , n6444  );
buf ( g6444 , n6445  );
buf ( g6445 , n6446  );
buf ( g6446 , n6447  );
buf ( g6447 , n6448  );
buf ( g6448 , n6449  );
buf ( g6449 , n6450  );
buf ( g6450 , n6451  );
buf ( g6451 , n6452  );
buf ( g6452 , n6453  );
buf ( g6453 , n6454  );
buf ( g6454 , n6455  );
buf ( g6455 , n6456  );
buf ( g6456 , n6457  );
buf ( g6457 , n6458  );
buf ( g6458 , n6459  );
buf ( g6459 , n6460  );
buf ( g6460 , n6461  );
buf ( g6461 , n6462  );
buf ( g6462 , n6463  );
buf ( g6463 , n6464  );
buf ( g6464 , n6465  );
buf ( g6465 , n6466  );
buf ( g6466 , n6467  );
buf ( g6467 , n6468  );
buf ( g6468 , n6469  );
buf ( g6469 , n6470  );
buf ( g6470 , n6471  );
buf ( g6471 , n6472  );
buf ( g6472 , n6473  );
buf ( g6473 , n6474  );
buf ( g6474 , n6475  );
buf ( g6475 , n6476  );
buf ( g6476 , n6477  );
buf ( g6477 , n6478  );
buf ( g6478 , n6479  );
buf ( g6479 , n6480  );
buf ( g6480 , n6481  );
buf ( g6481 , n6482  );
buf ( g6482 , n6483  );
buf ( g6483 , n6484  );
buf ( g6484 , n6485  );
buf ( g6485 , n6486  );
buf ( g6486 , n6487  );
buf ( g6487 , n6488  );
buf ( g6488 , n6489  );
buf ( g6489 , n6490  );
buf ( g6490 , n6491  );
buf ( g6491 , n6492  );
buf ( g6492 , n6493  );
buf ( g6493 , n6494  );
buf ( g6494 , n6495  );
buf ( g6495 , n6496  );
buf ( g6496 , n6497  );
buf ( g6497 , n6498  );
buf ( g6498 , n6499  );
buf ( g6499 , n6500  );
buf ( g6500 , n6501  );
buf ( g6501 , n6502  );
buf ( g6502 , n6503  );
buf ( g6503 , n6504  );
buf ( g6504 , n6505  );
buf ( g6505 , n6506  );
buf ( g6506 , n6507  );
buf ( g6507 , n6508  );
buf ( g6508 , n6509  );
buf ( g6509 , n6510  );
buf ( g6510 , n6511  );
buf ( g6511 , n6512  );
buf ( g6512 , n6513  );
buf ( g6513 , n6514  );
buf ( g6514 , n6515  );
buf ( g6515 , n6516  );
buf ( g6516 , n6517  );
buf ( g6517 , n6518  );
buf ( g6518 , n6519  );
buf ( g6519 , n6520  );
buf ( g6520 , n6521  );
buf ( g6521 , n6522  );
buf ( g6522 , n6523  );
buf ( g6523 , n6524  );
buf ( g6524 , n6525  );
buf ( g6525 , n6526  );
buf ( g6526 , n6527  );
buf ( g6527 , n6528  );
buf ( g6528 , n6529  );
buf ( g6529 , n6530  );
buf ( g6530 , n6531  );
buf ( g6531 , n6532  );
buf ( g6532 , n6533  );
buf ( g6533 , n6534  );
buf ( g6534 , n6535  );
buf ( g6535 , n6536  );
buf ( g6536 , n6537  );
buf ( g6537 , n6538  );
buf ( g6538 , n6539  );
buf ( g6539 , n6540  );
buf ( g6540 , n6541  );
buf ( g6541 , n6542  );
buf ( g6542 , n6543  );
buf ( g6543 , n6544  );
buf ( g6544 , n6545  );
buf ( g6545 , n6546  );
buf ( g6546 , n6547  );
buf ( g6547 , n6548  );
buf ( g6548 , n6549  );
buf ( g6549 , n6550  );
buf ( g6550 , n6551  );
buf ( g6551 , n6552  );
buf ( g6552 , n6553  );
buf ( g6553 , n6554  );
buf ( g6554 , n6555  );
buf ( g6555 , n6556  );
buf ( g6556 , n6557  );
buf ( g6557 , n6558  );
buf ( g6558 , n6559  );
buf ( g6559 , n6560  );
buf ( g6560 , n6561  );
buf ( g6561 , n6562  );
buf ( g6562 , n6563  );
buf ( g6563 , n6564  );
buf ( g6564 , n6565  );
buf ( g6565 , n6566  );
buf ( g6566 , n6567  );
buf ( g6567 , n6568  );
buf ( g6568 , n6569  );
buf ( g6569 , n6570  );
buf ( g6570 , n6571  );
buf ( g6571 , n6572  );
buf ( g6572 , n6573  );
buf ( g6573 , n6574  );
buf ( g6574 , n6575  );
buf ( g6575 , n6576  );
buf ( g6576 , n6577  );
buf ( g6577 , n6578  );
buf ( g6578 , n6579  );
buf ( g6579 , n6580  );
buf ( g6580 , n6581  );
buf ( g6581 , n6582  );
buf ( g6582 , n6583  );
buf ( g6583 , n6584  );
buf ( g6584 , n6585  );
buf ( g6585 , n6586  );
buf ( g6586 , n6587  );
buf ( g6587 , n6588  );
buf ( g6588 , n6589  );
buf ( g6589 , n6590  );
buf ( g6590 , n6591  );
buf ( g6591 , n6592  );
buf ( g6592 , n6593  );
buf ( g6593 , n6594  );
buf ( g6594 , n6595  );
buf ( g6595 , n6596  );
buf ( g6596 , n6597  );
buf ( g6597 , n6598  );
buf ( g6598 , n6599  );
buf ( g6599 , n6600  );
buf ( g6600 , n6601  );
buf ( g6601 , n6602  );
buf ( g6602 , n6603  );
buf ( g6603 , n6604  );
buf ( g6604 , n6605  );
buf ( g6605 , n6606  );
buf ( g6606 , n6607  );
buf ( g6607 , n6608  );
buf ( g6608 , n6609  );
buf ( g6609 , n6610  );
buf ( g6610 , n6611  );
buf ( g6611 , n6612  );
buf ( g6612 , n6613  );
buf ( g6613 , n6614  );
buf ( g6614 , n6615  );
buf ( g6615 , n6616  );
buf ( g6616 , n6617  );
buf ( g6617 , n6618  );
buf ( g6618 , n6619  );
buf ( g6619 , n6620  );
buf ( g6620 , n6621  );
buf ( g6621 , n6622  );
buf ( g6622 , n6623  );
buf ( g6623 , n6624  );
buf ( g6624 , n6625  );
buf ( g6625 , n6626  );
buf ( g6626 , n6627  );
buf ( g6627 , n6628  );
buf ( g6628 , n6629  );
buf ( g6629 , n6630  );
buf ( g6630 , n6631  );
buf ( g6631 , n6632  );
buf ( g6632 , n6633  );
buf ( g6633 , n6634  );
buf ( g6634 , n6635  );
buf ( g6635 , n6636  );
buf ( g6636 , n6637  );
buf ( g6637 , n6638  );
buf ( g6638 , n6639  );
buf ( g6639 , n6640  );
buf ( g6640 , n6641  );
buf ( g6641 , n6642  );
buf ( g6642 , n6643  );
buf ( g6643 , n6644  );
buf ( g6644 , n6645  );
buf ( g6645 , n6646  );
buf ( g6646 , n6647  );
buf ( g6647 , n6648  );
buf ( g6648 , n6649  );
buf ( g6649 , n6650  );
buf ( g6650 , n6651  );
buf ( g6651 , n6652  );
buf ( g6652 , n6653  );
buf ( g6653 , n6654  );
buf ( g6654 , n6655  );
buf ( g6655 , n6656  );
buf ( g6656 , n6657  );
buf ( g6657 , n6658  );
buf ( g6658 , n6659  );
buf ( g6659 , n6660  );
buf ( g6660 , n6661  );
buf ( g6661 , n6662  );
buf ( g6662 , n6663  );
buf ( g6663 , n6664  );
buf ( g6664 , n6665  );
buf ( g6665 , n6666  );
buf ( g6666 , n6667  );
buf ( g6667 , n6668  );
buf ( g6668 , n6669  );
buf ( g6669 , n6670  );
buf ( g6670 , n6671  );
buf ( g6671 , n6672  );
buf ( g6672 , n6673  );
buf ( g6673 , n6674  );
buf ( g6674 , n6675  );
buf ( g6675 , n6676  );
buf ( g6676 , n6677  );
buf ( g6677 , n6678  );
buf ( g6678 , n6679  );
buf ( g6679 , n6680  );
buf ( g6680 , n6681  );
buf ( g6681 , n6682  );
buf ( g6682 , n6683  );
buf ( g6683 , n6684  );
buf ( g6684 , n6685  );
buf ( g6685 , n6686  );
buf ( g6686 , n6687  );
buf ( g6687 , n6688  );
buf ( g6688 , n6689  );
buf ( g6689 , n6690  );
buf ( g6690 , n6691  );
buf ( g6691 , n6692  );
buf ( g6692 , n6693  );
buf ( g6693 , n6694  );
buf ( g6694 , n6695  );
buf ( g6695 , n6696  );
buf ( g6696 , n6697  );
buf ( g6697 , n6698  );
buf ( g6698 , n6699  );
buf ( g6699 , n6700  );
buf ( g6700 , n6701  );
buf ( g6701 , n6702  );
buf ( g6702 , n6703  );
buf ( g6703 , n6704  );
buf ( g6704 , n6705  );
buf ( g6705 , n6706  );
buf ( g6706 , n6707  );
buf ( g6707 , n6708  );
buf ( g6708 , n6709  );
buf ( g6709 , n6710  );
buf ( g6710 , n6711  );
buf ( g6711 , n6712  );
buf ( g6712 , n6713  );
buf ( g6713 , n6714  );
buf ( g6714 , n6715  );
buf ( g6715 , n6716  );
buf ( g6716 , n6717  );
buf ( g6717 , n6718  );
buf ( g6718 , n6719  );
buf ( g6719 , n6720  );
buf ( g6720 , n6721  );
buf ( g6721 , n6722  );
buf ( g6722 , n6723  );
buf ( g6723 , n6724  );
buf ( g6724 , n6725  );
buf ( g6725 , n6726  );
buf ( g6726 , n6727  );
buf ( g6727 , n6728  );
buf ( g6728 , n6729  );
buf ( g6729 , n6730  );
buf ( g6730 , n6731  );
buf ( g6731 , n6732  );
buf ( g6732 , n6733  );
buf ( g6733 , n6734  );
buf ( g6734 , n6735  );
buf ( g6735 , n6736  );
buf ( g6736 , n6737  );
buf ( g6737 , n6738  );
buf ( g6738 , n6739  );
buf ( g6739 , n6740  );
buf ( g6740 , n6741  );
buf ( g6741 , n6742  );
buf ( g6742 , n6743  );
buf ( g6743 , n6744  );
buf ( g6744 , n6745  );
buf ( g6745 , n6746  );
buf ( g6746 , n6747  );
buf ( g6747 , n6748  );
buf ( g6748 , n6749  );
buf ( g6749 , n6750  );
buf ( g6750 , n6751  );
buf ( g6751 , n6752  );
buf ( g6752 , n6753  );
buf ( g6753 , n6754  );
buf ( g6754 , n6755  );
buf ( g6755 , n6756  );
buf ( g6756 , n6757  );
buf ( g6757 , n6758  );
buf ( g6758 , n6759  );
buf ( g6759 , n6760  );
buf ( g6760 , n6761  );
buf ( g6761 , n6762  );
buf ( g6762 , n6763  );
buf ( g6763 , n6764  );
buf ( g6764 , n6765  );
buf ( g6765 , n6766  );
buf ( g6766 , n6767  );
buf ( g6767 , n6768  );
buf ( g6768 , n6769  );
buf ( g6769 , n6770  );
buf ( g6770 , n6771  );
buf ( g6771 , n6772  );
buf ( g6772 , n6773  );
buf ( g6773 , n6774  );
buf ( g6774 , n6775  );
buf ( g6775 , n6776  );
buf ( g6776 , n6777  );
buf ( g6777 , n6778  );
buf ( g6778 , n6779  );
buf ( g6779 , n6780  );
buf ( g6780 , n6781  );
buf ( g6781 , n6782  );
buf ( g6782 , n6783  );
buf ( g6783 , n6784  );
buf ( g6784 , n6785  );
buf ( g6785 , n6786  );
buf ( g6786 , n6787  );
buf ( g6787 , n6788  );
buf ( g6788 , n6789  );
buf ( g6789 , n6790  );
buf ( g6790 , n6791  );
buf ( g6791 , n6792  );
buf ( g6792 , n6793  );
buf ( g6793 , n6794  );
buf ( g6794 , n6795  );
buf ( g6795 , n6796  );
buf ( g6796 , n6797  );
buf ( g6797 , n6798  );
buf ( g6798 , n6799  );
buf ( g6799 , n6800  );
buf ( g6800 , n6801  );
buf ( g6801 , n6802  );
buf ( g6802 , n6803  );
buf ( g6803 , n6804  );
buf ( g6804 , n6805  );
buf ( g6805 , n6806  );
buf ( g6806 , n6807  );
buf ( g6807 , n6808  );
buf ( g6808 , n6809  );
buf ( g6809 , n6810  );
buf ( g6810 , n6811  );
buf ( g6811 , n6812  );
buf ( g6812 , n6813  );
buf ( g6813 , n6814  );
buf ( g6814 , n6815  );
buf ( g6815 , n6816  );
buf ( g6816 , n6817  );
buf ( g6817 , n6818  );
buf ( g6818 , n6819  );
buf ( g6819 , n6820  );
buf ( g6820 , n6821  );
buf ( g6821 , n6822  );
buf ( g6822 , n6823  );
buf ( g6823 , n6824  );
buf ( g6824 , n6825  );
buf ( g6825 , n6826  );
buf ( g6826 , n6827  );
buf ( g6827 , n6828  );
buf ( g6828 , n6829  );
buf ( g6829 , n6830  );
buf ( g6830 , n6831  );
buf ( g6831 , n6832  );
buf ( g6832 , n6833  );
buf ( g6833 , n6834  );
buf ( g6834 , n6835  );
buf ( g6835 , n6836  );
buf ( g6836 , n6837  );
buf ( g6837 , n6838  );
buf ( g6838 , n6839  );
buf ( g6839 , n6840  );
buf ( g6840 , n6841  );
buf ( g6841 , n6842  );
buf ( g6842 , n6843  );
buf ( g6843 , n6844  );
buf ( g6844 , n6845  );
buf ( g6845 , n6846  );
buf ( g6846 , n6847  );
buf ( g6847 , n6848  );
buf ( g6848 , n6849  );
buf ( g6849 , n6850  );
buf ( g6850 , n6851  );
buf ( g6851 , n6852  );
buf ( g6852 , n6853  );
buf ( g6853 , n6854  );
buf ( g6854 , n6855  );
buf ( g6855 , n6856  );
buf ( g6856 , n6857  );
buf ( g6857 , n6858  );
buf ( g6858 , n6859  );
buf ( g6859 , n6860  );
buf ( g6860 , n6861  );
buf ( g6861 , n6862  );
buf ( g6862 , n6863  );
buf ( g6863 , n6864  );
buf ( g6864 , n6865  );
buf ( g6865 , n6866  );
buf ( g6866 , n6867  );
buf ( g6867 , n6868  );
buf ( g6868 , n6869  );
buf ( g6869 , n6870  );
buf ( g6870 , n6871  );
buf ( g6871 , n6872  );
buf ( g6872 , n6873  );
buf ( g6873 , n6874  );
buf ( g6874 , n6875  );
buf ( g6875 , n6876  );
buf ( g6876 , n6877  );
buf ( g6877 , n6878  );
buf ( g6878 , n6879  );
buf ( g6879 , n6880  );
buf ( g6880 , n6881  );
buf ( g6881 , n6882  );
buf ( g6882 , n6883  );
buf ( g6883 , n6884  );
buf ( g6884 , n6885  );
buf ( g6885 , n6886  );
buf ( g6886 , n6887  );
buf ( g6887 , n6888  );
buf ( g6888 , n6889  );
buf ( g6889 , n6890  );
buf ( g6890 , n6891  );
buf ( g6891 , n6892  );
buf ( g6892 , n6893  );
buf ( g6893 , n6894  );
buf ( g6894 , n6895  );
buf ( g6895 , n6896  );
buf ( g6896 , n6897  );
buf ( g6897 , n6898  );
buf ( g6898 , n6899  );
buf ( g6899 , n6900  );
buf ( g6900 , n6901  );
buf ( g6901 , n6902  );
buf ( g6902 , n6903  );
buf ( g6903 , n6904  );
buf ( g6904 , n6905  );
buf ( g6905 , n6906  );
buf ( g6906 , n6907  );
buf ( g6907 , n6908  );
buf ( g6908 , n6909  );
buf ( g6909 , n6910  );
buf ( g6910 , n6911  );
buf ( g6911 , n6912  );
buf ( g6912 , n6913  );
buf ( g6913 , n6914  );
buf ( g6914 , n6915  );
buf ( g6915 , n6916  );
buf ( g6916 , n6917  );
buf ( g6917 , n6918  );
buf ( g6918 , n6919  );
buf ( g6919 , n6920  );
buf ( g6920 , n6921  );
buf ( g6921 , n6922  );
buf ( g6922 , n6923  );
buf ( g6923 , n6924  );
buf ( g6924 , n6925  );
buf ( g6925 , n6926  );
buf ( g6926 , n6927  );
buf ( g6927 , n6928  );
buf ( g6928 , n6929  );
buf ( g6929 , n6930  );
buf ( g6930 , n6931  );
buf ( g6931 , n6932  );
buf ( g6932 , n6933  );
buf ( g6933 , n6934  );
buf ( g6934 , n6935  );
buf ( g6935 , n6936  );
buf ( g6936 , n6937  );
buf ( g6937 , n6938  );
buf ( g6938 , n6939  );
buf ( g6939 , n6940  );
buf ( g6940 , n6941  );
buf ( g6941 , n6942  );
buf ( g6942 , n6943  );
buf ( g6943 , n6944  );
buf ( g6944 , n6945  );
buf ( g6945 , n6946  );
buf ( g6946 , n6947  );
buf ( g6947 , n6948  );
buf ( g6948 , n6949  );
buf ( g6949 , n6950  );
buf ( g6950 , n6951  );
buf ( g6951 , n6952  );
buf ( g6952 , n6953  );
buf ( g6953 , n6954  );
buf ( g6954 , n6955  );
buf ( g6955 , n6956  );
buf ( g6956 , n6957  );
buf ( g6957 , n6958  );
buf ( g6958 , n6959  );
buf ( g6959 , n6960  );
buf ( g6960 , n6961  );
buf ( g6961 , n6962  );
buf ( g6962 , n6963  );
buf ( g6963 , n6964  );
buf ( g6964 , n6965  );
buf ( g6965 , n6966  );
buf ( g6966 , n6967  );
buf ( g6967 , n6968  );
buf ( g6968 , n6969  );
buf ( g6969 , n6970  );
buf ( g6970 , n6971  );
buf ( g6971 , n6972  );
buf ( g6972 , n6973  );
buf ( g6973 , n6974  );
buf ( g6974 , n6975  );
buf ( g6975 , n6976  );
buf ( g6976 , n6977  );
buf ( g6977 , n6978  );
buf ( g6978 , n6979  );
buf ( g6979 , n6980  );
buf ( g6980 , n6981  );
buf ( g6981 , n6982  );
buf ( g6982 , n6983  );
buf ( g6983 , n6984  );
buf ( g6984 , n6985  );
buf ( g6985 , n6986  );
buf ( g6986 , n6987  );
buf ( g6987 , n6988  );
buf ( g6988 , n6989  );
buf ( g6989 , n6990  );
buf ( g6990 , n6991  );
buf ( g6991 , n6992  );
buf ( g6992 , n6993  );
buf ( g6993 , n6994  );
buf ( g6994 , n6995  );
buf ( g6995 , n6996  );
buf ( g6996 , n6997  );
buf ( g6997 , n6998  );
buf ( g6998 , n6999  );
buf ( g6999 , n7000  );
buf ( g7000 , n7001  );
buf ( g7001 , n7002  );
buf ( g7002 , n7003  );
buf ( g7003 , n7004  );
buf ( g7004 , n7005  );
buf ( g7005 , n7006  );
buf ( g7006 , n7007  );
buf ( g7007 , n7008  );
buf ( g7008 , n7009  );
buf ( g7009 , n7010  );
buf ( g7010 , n7011  );
buf ( g7011 , n7012  );
buf ( g7012 , n7013  );
buf ( g7013 , n7014  );
buf ( g7014 , n7015  );
buf ( g7015 , n7016  );
buf ( g7016 , n7017  );
buf ( g7017 , n7018  );
buf ( g7018 , n7019  );
buf ( g7019 , n7020  );
buf ( g7020 , n7021  );
buf ( g7021 , n7022  );
buf ( g7022 , n7023  );
buf ( g7023 , n7024  );
buf ( g7024 , n7025  );
buf ( g7025 , n7026  );
buf ( g7026 , n7027  );
buf ( g7027 , n7028  );
buf ( g7028 , n7029  );
buf ( g7029 , n7030  );
buf ( g7030 , n7031  );
buf ( g7031 , n7032  );
buf ( g7032 , n7033  );
buf ( g7033 , n7034  );
buf ( g7034 , n7035  );
buf ( g7035 , n7036  );
buf ( g7036 , n7037  );
buf ( g7037 , n7038  );
buf ( g7038 , n7039  );
buf ( g7039 , n7040  );
buf ( g7040 , n7041  );
buf ( g7041 , n7042  );
buf ( g7042 , n7043  );
buf ( g7043 , n7044  );
buf ( g7044 , n7045  );
buf ( g7045 , n7046  );
buf ( g7046 , n7047  );
buf ( g7047 , n7048  );
buf ( g7048 , n7049  );
buf ( g7049 , n7050  );
buf ( g7050 , n7051  );
buf ( g7051 , n7052  );
buf ( g7052 , n7053  );
buf ( g7053 , n7054  );
buf ( g7054 , n7055  );
buf ( g7055 , n7056  );
buf ( g7056 , n7057  );
buf ( g7057 , n7058  );
buf ( g7058 , n7059  );
buf ( g7059 , n7060  );
buf ( g7060 , n7061  );
buf ( g7061 , n7062  );
buf ( g7062 , n7063  );
buf ( g7063 , n7064  );
buf ( g7064 , n7065  );
buf ( g7065 , n7066  );
buf ( g7066 , n7067  );
buf ( g7067 , n7068  );
buf ( g7068 , n7069  );
buf ( g7069 , n7070  );
buf ( g7070 , n7071  );
buf ( g7071 , n7072  );
buf ( g7072 , n7073  );
buf ( g7073 , n7074  );
buf ( g7074 , n7075  );
buf ( g7075 , n7076  );
buf ( g7076 , n7077  );
buf ( g7077 , n7078  );
buf ( g7078 , n7079  );
buf ( g7079 , n7080  );
buf ( g7080 , n7081  );
buf ( g7081 , n7082  );
buf ( g7082 , n7083  );
buf ( g7083 , n7084  );
buf ( g7084 , n7085  );
buf ( g7085 , n7086  );
buf ( g7086 , n7087  );
buf ( g7087 , n7088  );
buf ( g7088 , n7089  );
buf ( g7089 , n7090  );
buf ( g7090 , n7091  );
buf ( g7091 , n7092  );
buf ( g7092 , n7093  );
buf ( g7093 , n7094  );
buf ( g7094 , n7095  );
buf ( g7095 , n7096  );
buf ( g7096 , n7097  );
buf ( g7097 , n7098  );
buf ( g7098 , n7099  );
buf ( g7099 , n7100  );
buf ( g7100 , n7101  );
buf ( g7101 , n7102  );
buf ( g7102 , n7103  );
buf ( g7103 , n7104  );
buf ( g7104 , n7105  );
buf ( g7105 , n7106  );
buf ( g7106 , n7107  );
buf ( g7107 , n7108  );
buf ( g7108 , n7109  );
buf ( g7109 , n7110  );
buf ( g7110 , n7111  );
buf ( g7111 , n7112  );
buf ( g7112 , n7113  );
buf ( g7113 , n7114  );
buf ( g7114 , n7115  );
buf ( g7115 , n7116  );
buf ( g7116 , n7117  );
buf ( g7117 , n7118  );
buf ( g7118 , n7119  );
buf ( g7119 , n7120  );
buf ( g7120 , n7121  );
buf ( g7121 , n7122  );
buf ( g7122 , n7123  );
buf ( g7123 , n7124  );
buf ( g7124 , n7125  );
buf ( g7125 , n7126  );
buf ( g7126 , n7127  );
buf ( g7127 , n7128  );
buf ( g7128 , n7129  );
buf ( g7129 , n7130  );
buf ( g7130 , n7131  );
buf ( g7131 , n7132  );
buf ( g7132 , n7133  );
buf ( g7133 , n7134  );
buf ( g7134 , n7135  );
buf ( g7135 , n7136  );
buf ( g7136 , n7137  );
buf ( g7137 , n7138  );
buf ( g7138 , n7139  );
buf ( g7139 , n7140  );
buf ( g7140 , n7141  );
buf ( g7141 , n7142  );
buf ( g7142 , n7143  );
buf ( g7143 , n7144  );
buf ( g7144 , n7145  );
buf ( g7145 , n7146  );
buf ( g7146 , n7147  );
buf ( g7147 , n7148  );
buf ( g7148 , n7149  );
buf ( g7149 , n7150  );
buf ( g7150 , n7151  );
buf ( g7151 , n7152  );
buf ( g7152 , n7153  );
buf ( g7153 , n7154  );
buf ( g7154 , n7155  );
buf ( g7155 , n7156  );
buf ( g7156 , n7157  );
buf ( g7157 , n7158  );
buf ( g7158 , n7159  );
buf ( g7159 , n7160  );
buf ( g7160 , n7161  );
buf ( g7161 , n7162  );
buf ( g7162 , n7163  );
buf ( g7163 , n7164  );
buf ( g7164 , n7165  );
buf ( g7165 , n7166  );
buf ( g7166 , n7167  );
buf ( g7167 , n7168  );
buf ( g7168 , n7169  );
buf ( g7169 , n7170  );
buf ( g7170 , n7171  );
buf ( g7171 , n7172  );
buf ( g7172 , n7173  );
buf ( g7173 , n7174  );
buf ( g7174 , n7175  );
buf ( g7175 , n7176  );
buf ( g7176 , n7177  );
buf ( g7177 , n7178  );
buf ( g7178 , n7179  );
buf ( g7179 , n7180  );
buf ( g7180 , n7181  );
buf ( g7181 , n7182  );
buf ( g7182 , n7183  );
buf ( g7183 , n7184  );
buf ( g7184 , n7185  );
buf ( g7185 , n7186  );
buf ( g7186 , n7187  );
buf ( g7187 , n7188  );
buf ( g7188 , n7189  );
buf ( g7189 , n7190  );
buf ( g7190 , n7191  );
buf ( g7191 , n7192  );
buf ( g7192 , n7193  );
buf ( g7193 , n7194  );
buf ( g7194 , n7195  );
buf ( g7195 , n7196  );
buf ( g7196 , n7197  );
buf ( g7197 , n7198  );
buf ( g7198 , n7199  );
buf ( g7199 , n7200  );
buf ( g7200 , n7201  );
buf ( g7201 , n7202  );
buf ( g7202 , n7203  );
buf ( g7203 , n7204  );
buf ( g7204 , n7205  );
buf ( g7205 , n7206  );
buf ( g7206 , n7207  );
buf ( g7207 , n7208  );
buf ( g7208 , n7209  );
buf ( g7209 , n7210  );
buf ( g7210 , n7211  );
buf ( g7211 , n7212  );
buf ( g7212 , n7213  );
buf ( g7213 , n7214  );
buf ( g7214 , n7215  );
buf ( g7215 , n7216  );
buf ( g7216 , n7217  );
buf ( g7217 , n7218  );
buf ( g7218 , n7219  );
buf ( g7219 , n7220  );
buf ( g7220 , n7221  );
buf ( g7221 , n7222  );
buf ( g7222 , n7223  );
buf ( g7223 , n7224  );
buf ( g7224 , n7225  );
buf ( g7225 , n7226  );
buf ( g7226 , n7227  );
buf ( g7227 , n7228  );
buf ( g7228 , n7229  );
buf ( g7229 , n7230  );
buf ( g7230 , n7231  );
buf ( g7231 , n7232  );
buf ( g7232 , n7233  );
buf ( g7233 , n7234  );
buf ( g7234 , n7235  );
buf ( g7235 , n7236  );
buf ( g7236 , n7237  );
buf ( g7237 , n7238  );
buf ( g7238 , n7239  );
buf ( g7239 , n7240  );
buf ( g7240 , n7241  );
buf ( g7241 , n7242  );
buf ( g7242 , n7243  );
buf ( g7243 , n7244  );
buf ( g7244 , n7245  );
buf ( g7245 , n7246  );
buf ( g7246 , n7247  );
buf ( g7247 , n7248  );
buf ( g7248 , n7249  );
buf ( g7249 , n7250  );
buf ( g7250 , n7251  );
buf ( g7251 , n7252  );
buf ( g7252 , n7253  );
buf ( g7253 , n7254  );
buf ( g7254 , n7255  );
buf ( g7255 , n7256  );
buf ( g7256 , n7257  );
buf ( g7257 , n7258  );
buf ( g7258 , n7259  );
buf ( g7259 , n7260  );
buf ( g7260 , n7261  );
buf ( g7261 , n7262  );
buf ( g7262 , n7263  );
buf ( g7263 , n7264  );
buf ( g7264 , n7265  );
buf ( g7265 , n7266  );
buf ( g7266 , n7267  );
buf ( g7267 , n7268  );
buf ( g7268 , n7269  );
buf ( g7269 , n7270  );
buf ( g7270 , n7271  );
buf ( g7271 , n7272  );
buf ( g7272 , n7273  );
buf ( g7273 , n7274  );
buf ( g7274 , n7275  );
buf ( g7275 , n7276  );
buf ( g7276 , n7277  );
buf ( g7277 , n7278  );
buf ( g7278 , n7279  );
buf ( g7279 , n7280  );
buf ( g7280 , n7281  );
buf ( g7281 , n7282  );
buf ( g7282 , n7283  );
buf ( g7283 , n7284  );
buf ( g7284 , n7285  );
buf ( g7285 , n7286  );
buf ( g7286 , n7287  );
buf ( g7287 , n7288  );
buf ( g7288 , n7289  );
buf ( g7289 , n7290  );
buf ( g7290 , n7291  );
buf ( g7291 , n7292  );
buf ( g7292 , n7293  );
buf ( g7293 , n7294  );
buf ( g7294 , n7295  );
buf ( g7295 , n7296  );
buf ( g7296 , n7297  );
buf ( g7297 , n7298  );
buf ( g7298 , n7299  );
buf ( g7299 , n7300  );
buf ( g7300 , n7301  );
buf ( g7301 , n7302  );
buf ( g7302 , n7303  );
buf ( g7303 , n7304  );
buf ( g7304 , n7305  );
buf ( g7305 , n7306  );
buf ( g7306 , n7307  );
buf ( g7307 , n7308  );
buf ( g7308 , n7309  );
buf ( g7309 , n7310  );
buf ( g7310 , n7311  );
buf ( g7311 , n7312  );
buf ( g7312 , n7313  );
buf ( g7313 , n7314  );
buf ( g7314 , n7315  );
buf ( g7315 , n7316  );
buf ( g7316 , n7317  );
buf ( g7317 , n7318  );
buf ( g7318 , n7319  );
buf ( g7319 , n7320  );
buf ( g7320 , n7321  );
buf ( g7321 , n7322  );
buf ( g7322 , n7323  );
buf ( g7323 , n7324  );
buf ( g7324 , n7325  );
buf ( g7325 , n7326  );
buf ( g7326 , n7327  );
buf ( g7327 , n7328  );
buf ( g7328 , n7329  );
buf ( g7329 , n7330  );
buf ( g7330 , n7331  );
buf ( g7331 , n7332  );
buf ( g7332 , n7333  );
buf ( g7333 , n7334  );
buf ( g7334 , n7335  );
buf ( g7335 , n7336  );
buf ( g7336 , n7337  );
buf ( g7337 , n7338  );
buf ( g7338 , n7339  );
buf ( g7339 , n7340  );
buf ( g7340 , n7341  );
buf ( g7341 , n7342  );
buf ( g7342 , n7343  );
buf ( g7343 , n7344  );
buf ( g7344 , n7345  );
buf ( g7345 , n7346  );
buf ( g7346 , n7347  );
buf ( g7347 , n7348  );
buf ( g7348 , n7349  );
buf ( g7349 , n7350  );
buf ( g7350 , n7351  );
buf ( g7351 , n7352  );
buf ( g7352 , n7353  );
buf ( g7353 , n7354  );
buf ( g7354 , n7355  );
buf ( g7355 , n7356  );
buf ( g7356 , n7357  );
buf ( g7357 , n7358  );
buf ( g7358 , n7359  );
buf ( g7359 , n7360  );
buf ( g7360 , n7361  );
buf ( g7361 , n7362  );
buf ( g7362 , n7363  );
buf ( g7363 , n7364  );
buf ( g7364 , n7365  );
buf ( g7365 , n7366  );
buf ( g7366 , n7367  );
buf ( g7367 , n7368  );
buf ( g7368 , n7369  );
buf ( g7369 , n7370  );
buf ( g7370 , n7371  );
buf ( g7371 , n7372  );
buf ( g7372 , n7373  );
buf ( g7373 , n7374  );
buf ( g7374 , n7375  );
buf ( g7375 , n7376  );
buf ( g7376 , n7377  );
buf ( g7377 , n7378  );
buf ( g7378 , n7379  );
buf ( g7379 , n7380  );
buf ( g7380 , n7381  );
buf ( g7381 , n7382  );
buf ( g7382 , n7383  );
buf ( g7383 , n7384  );
buf ( g7384 , n7385  );
buf ( g7385 , n7386  );
buf ( g7386 , n7387  );
buf ( g7387 , n7388  );
buf ( g7388 , n7389  );
buf ( g7389 , n7390  );
buf ( g7390 , n7391  );
buf ( g7391 , n7392  );
buf ( g7392 , n7393  );
buf ( g7393 , n7394  );
buf ( g7394 , n7395  );
buf ( g7395 , n7396  );
buf ( g7396 , n7397  );
buf ( g7397 , n7398  );
buf ( g7398 , n7399  );
buf ( g7399 , n7400  );
buf ( g7400 , n7401  );
buf ( g7401 , n7402  );
buf ( g7402 , n7403  );
buf ( g7403 , n7404  );
buf ( g7404 , n7405  );
buf ( g7405 , n7406  );
buf ( g7406 , n7407  );
buf ( g7407 , n7408  );
buf ( g7408 , n7409  );
buf ( g7409 , n7410  );
buf ( g7410 , n7411  );
buf ( g7411 , n7412  );
buf ( g7412 , n7413  );
buf ( g7413 , n7414  );
buf ( g7414 , n7415  );
buf ( g7415 , n7416  );
buf ( g7416 , n7417  );
buf ( g7417 , n7418  );
buf ( g7418 , n7419  );
buf ( g7419 , n7420  );
buf ( g7420 , n7421  );
buf ( g7421 , n7422  );
buf ( g7422 , n7423  );
buf ( g7423 , n7424  );
buf ( g7424 , n7425  );
buf ( g7425 , n7426  );
buf ( g7426 , n7427  );
buf ( g7427 , n7428  );
buf ( g7428 , n7429  );
buf ( g7429 , n7430  );
buf ( g7430 , n7431  );
buf ( g7431 , n7432  );
buf ( g7432 , n7433  );
buf ( g7433 , n7434  );
buf ( g7434 , n7435  );
buf ( g7435 , n7436  );
buf ( g7436 , n7437  );
buf ( g7437 , n7438  );
buf ( g7438 , n7439  );
buf ( g7439 , n7440  );
buf ( g7440 , n7441  );
buf ( g7441 , n7442  );
buf ( g7442 , n7443  );
buf ( g7443 , n7444  );
buf ( g7444 , n7445  );
buf ( g7445 , n7446  );
buf ( g7446 , n7447  );
buf ( g7447 , n7448  );
buf ( g7448 , n7449  );
buf ( g7449 , n7450  );
buf ( g7450 , n7451  );
buf ( g7451 , n7452  );
buf ( g7452 , n7453  );
buf ( g7453 , n7454  );
buf ( g7454 , n7455  );
buf ( g7455 , n7456  );
buf ( g7456 , n7457  );
buf ( g7457 , n7458  );
buf ( g7458 , n7459  );
buf ( g7459 , n7460  );
buf ( g7460 , n7461  );
buf ( g7461 , n7462  );
buf ( g7462 , n7463  );
buf ( g7463 , n7464  );
buf ( g7464 , n7465  );
buf ( g7465 , n7466  );
buf ( g7466 , n7467  );
buf ( g7467 , n7468  );
buf ( g7468 , n7469  );
buf ( g7469 , n7470  );
buf ( g7470 , n7471  );
buf ( g7471 , n7472  );
buf ( g7472 , n7473  );
buf ( g7473 , n7474  );
buf ( g7474 , n7475  );
buf ( g7475 , n7476  );
buf ( g7476 , n7477  );
buf ( g7477 , n7478  );
buf ( g7478 , n7479  );
buf ( g7479 , n7480  );
buf ( g7480 , n7481  );
buf ( g7481 , n7482  );
buf ( g7482 , n7483  );
buf ( g7483 , n7484  );
buf ( g7484 , n7485  );
buf ( g7485 , n7486  );
buf ( g7486 , n7487  );
buf ( g7487 , n7488  );
buf ( g7488 , n7489  );
buf ( g7489 , n7490  );
buf ( g7490 , n7491  );
buf ( g7491 , n7492  );
buf ( g7492 , n7493  );
buf ( g7493 , n7494  );
buf ( g7494 , n7495  );
buf ( g7495 , n7496  );
buf ( g7496 , n7497  );
buf ( g7497 , n7498  );
buf ( g7498 , n7499  );
buf ( g7499 , n7500  );
buf ( g7500 , n7501  );
buf ( g7501 , n7502  );
buf ( g7502 , n7503  );
buf ( g7503 , n7504  );
buf ( g7504 , n7505  );
buf ( g7505 , n7506  );
buf ( g7506 , n7507  );
buf ( g7507 , n7508  );
buf ( g7508 , n7509  );
buf ( g7509 , n7510  );
buf ( g7510 , n7511  );
buf ( g7511 , n7512  );
buf ( g7512 , n7513  );
buf ( g7513 , n7514  );
buf ( g7514 , n7515  );
buf ( g7515 , n7516  );
buf ( g7516 , n7517  );
buf ( g7517 , n7518  );
buf ( g7518 , n7519  );
buf ( g7519 , n7520  );
buf ( g7520 , n7521  );
buf ( g7521 , n7522  );
buf ( g7522 , n7523  );
buf ( g7523 , n7524  );
buf ( g7524 , n7525  );
buf ( g7525 , n7526  );
buf ( g7526 , n7527  );
buf ( g7527 , n7528  );
buf ( g7528 , n7529  );
buf ( g7529 , n7530  );
buf ( g7530 , n7531  );
buf ( g7531 , n7532  );
buf ( g7532 , n7533  );
buf ( g7533 , n7534  );
buf ( g7534 , n7535  );
buf ( g7535 , n7536  );
buf ( g7536 , n7537  );
buf ( g7537 , n7538  );
buf ( g7538 , n7539  );
buf ( g7539 , n7540  );
buf ( g7540 , n7541  );
buf ( g7541 , n7542  );
buf ( g7542 , n7543  );
buf ( g7543 , n7544  );
buf ( g7544 , n7545  );
buf ( g7545 , n7546  );
buf ( g7546 , n7547  );
buf ( g7547 , n7548  );
buf ( g7548 , n7549  );
buf ( g7549 , n7550  );
buf ( g7550 , n7551  );
buf ( g7551 , n7552  );
buf ( g7552 , n7553  );
buf ( g7553 , n7554  );
buf ( g7554 , n7555  );
buf ( g7555 , n7556  );
buf ( g7556 , n7557  );
buf ( g7557 , n7558  );
buf ( g7558 , n7559  );
buf ( g7559 , n7560  );
buf ( g7560 , n7561  );
buf ( g7561 , n7562  );
buf ( g7562 , n7563  );
buf ( g7563 , n7564  );
buf ( g7564 , n7565  );
buf ( g7565 , n7566  );
buf ( g7566 , n7567  );
buf ( g7567 , n7568  );
buf ( g7568 , n7569  );
buf ( g7569 , n7570  );
buf ( g7570 , n7571  );
buf ( g7571 , n7572  );
buf ( g7572 , n7573  );
buf ( g7573 , n7574  );
buf ( g7574 , n7575  );
buf ( g7575 , n7576  );
buf ( g7576 , n7577  );
buf ( g7577 , n7578  );
buf ( g7578 , n7579  );
buf ( g7579 , n7580  );
buf ( g7580 , n7581  );
buf ( g7581 , n7582  );
buf ( g7582 , n7583  );
buf ( g7583 , n7584  );
buf ( g7584 , n7585  );
buf ( g7585 , n7586  );
buf ( g7586 , n7587  );
buf ( g7587 , n7588  );
buf ( g7588 , n7589  );
buf ( g7589 , n7590  );
buf ( g7590 , n7591  );
buf ( g7591 , n7592  );
buf ( g7592 , n7593  );
buf ( g7593 , n7594  );
buf ( g7594 , n7595  );
buf ( g7595 , n7596  );
buf ( g7596 , n7597  );
buf ( g7597 , n7598  );
buf ( g7598 , n7599  );
buf ( g7599 , n7600  );
buf ( g7600 , n7601  );
buf ( g7601 , n7602  );
buf ( g7602 , n7603  );
buf ( g7603 , n7604  );
buf ( g7604 , n7605  );
buf ( g7605 , n7606  );
buf ( g7606 , n7607  );
buf ( g7607 , n7608  );
buf ( g7608 , n7609  );
buf ( g7609 , n7610  );
buf ( g7610 , n7611  );
buf ( g7611 , n7612  );
buf ( g7612 , n7613  );
buf ( g7613 , n7614  );
buf ( g7614 , n7615  );
buf ( g7615 , n7616  );
buf ( g7616 , n7617  );
buf ( g7617 , n7618  );
buf ( g7618 , n7619  );
buf ( g7619 , n7620  );
buf ( g7620 , n7621  );
buf ( g7621 , n7622  );
buf ( g7622 , n7623  );
buf ( g7623 , n7624  );
buf ( g7624 , n7625  );
buf ( g7625 , n7626  );
buf ( g7626 , n7627  );
buf ( g7627 , n7628  );
buf ( g7628 , n7629  );
buf ( g7629 , n7630  );
buf ( g7630 , n7631  );
buf ( g7631 , n7632  );
buf ( g7632 , n7633  );
buf ( g7633 , n7634  );
buf ( g7634 , n7635  );
buf ( g7635 , n7636  );
buf ( g7636 , n7637  );
buf ( g7637 , n7638  );
buf ( g7638 , n7639  );
buf ( g7639 , n7640  );
buf ( g7640 , n7641  );
buf ( g7641 , n7642  );
buf ( g7642 , n7643  );
buf ( g7643 , n7644  );
buf ( g7644 , n7645  );
buf ( g7645 , n7646  );
buf ( g7646 , n7647  );
buf ( g7647 , n7648  );
buf ( g7648 , n7649  );
buf ( g7649 , n7650  );
buf ( g7650 , n7651  );
buf ( g7651 , n7652  );
buf ( g7652 , n7653  );
buf ( g7653 , n7654  );
buf ( g7654 , n7655  );
buf ( g7655 , n7656  );
buf ( g7656 , n7657  );
buf ( g7657 , n7658  );
buf ( g7658 , n7659  );
buf ( g7659 , n7660  );
buf ( g7660 , n7661  );
buf ( g7661 , n7662  );
buf ( g7662 , n7663  );
buf ( g7663 , n7664  );
buf ( g7664 , n7665  );
buf ( g7665 , n7666  );
buf ( g7666 , n7667  );
buf ( g7667 , n7668  );
buf ( g7668 , n7669  );
buf ( g7669 , n7670  );
buf ( g7670 , n7671  );
buf ( g7671 , n7672  );
buf ( g7672 , n7673  );
buf ( g7673 , n7674  );
buf ( g7674 , n7675  );
buf ( g7675 , n7676  );
buf ( g7676 , n7677  );
buf ( g7677 , n7678  );
buf ( g7678 , n7679  );
buf ( g7679 , n7680  );
buf ( g7680 , n7681  );
buf ( g7681 , n7682  );
buf ( g7682 , n7683  );
buf ( g7683 , n7684  );
buf ( g7684 , n7685  );
buf ( g7685 , n7686  );
buf ( g7686 , n7687  );
buf ( g7687 , n7688  );
buf ( g7688 , n7689  );
buf ( g7689 , n7690  );
buf ( g7690 , n7691  );
buf ( g7691 , n7692  );
buf ( g7692 , n7693  );
buf ( g7693 , n7694  );
buf ( g7694 , n7695  );
buf ( g7695 , n7696  );
buf ( g7696 , n7697  );
buf ( g7697 , n7698  );
buf ( g7698 , n7699  );
buf ( g7699 , n7700  );
buf ( g7700 , n7701  );
buf ( g7701 , n7702  );
buf ( g7702 , n7703  );
buf ( g7703 , n7704  );
buf ( g7704 , n7705  );
buf ( g7705 , n7706  );
buf ( g7706 , n7707  );
buf ( g7707 , n7708  );
buf ( g7708 , n7709  );
buf ( g7709 , n7710  );
buf ( g7710 , n7711  );
buf ( g7711 , n7712  );
buf ( g7712 , n7713  );
buf ( g7713 , n7714  );
buf ( g7714 , n7715  );
buf ( g7715 , n7716  );
buf ( g7716 , n7717  );
buf ( g7717 , n7718  );
buf ( g7718 , n7719  );
buf ( g7719 , n7720  );
buf ( g7720 , n7721  );
buf ( g7721 , n7722  );
buf ( g7722 , n7723  );
buf ( g7723 , n7724  );
buf ( g7724 , n7725  );
buf ( g7725 , n7726  );
buf ( g7726 , n7727  );
buf ( g7727 , n7728  );
buf ( g7728 , n7729  );
buf ( g7729 , n7730  );
buf ( g7730 , n7731  );
buf ( g7731 , n7732  );
buf ( g7732 , n7733  );
buf ( g7733 , n7734  );
buf ( g7734 , n7735  );
buf ( g7735 , n7736  );
buf ( g7736 , n7737  );
buf ( g7737 , n7738  );
buf ( g7738 , n7739  );
buf ( g7739 , n7740  );
buf ( g7740 , n7741  );
buf ( g7741 , n7742  );
buf ( g7742 , n7743  );
buf ( g7743 , n7744  );
buf ( g7744 , n7745  );
buf ( g7745 , n7746  );
buf ( g7746 , n7747  );
buf ( g7747 , n7748  );
buf ( g7748 , n7749  );
buf ( g7749 , n7750  );
buf ( g7750 , n7751  );
buf ( g7751 , n7752  );
buf ( g7752 , n7753  );
buf ( g7753 , n7754  );
buf ( g7754 , n7755  );
buf ( g7755 , n7756  );
buf ( g7756 , n7757  );
buf ( g7757 , n7758  );
buf ( g7758 , n7759  );
buf ( g7759 , n7760  );
buf ( g7760 , n7761  );
buf ( g7761 , n7762  );
buf ( g7762 , n7763  );
buf ( g7763 , n7764  );
buf ( g7764 , n7765  );
buf ( g7765 , n7766  );
buf ( g7766 , n7767  );
buf ( g7767 , n7768  );
buf ( g7768 , n7769  );
buf ( g7769 , n7770  );
buf ( g7770 , n7771  );
buf ( g7771 , n7772  );
buf ( g7772 , n7773  );
buf ( g7773 , n7774  );
buf ( g7774 , n7775  );
buf ( g7775 , n7776  );
buf ( g7776 , n7777  );
buf ( g7777 , n7778  );
buf ( g7778 , n7779  );
buf ( g7779 , n7780  );
buf ( g7780 , n7781  );
buf ( g7781 , n7782  );
buf ( g7782 , n7783  );
buf ( g7783 , n7784  );
buf ( g7784 , n7785  );
buf ( g7785 , n7786  );
buf ( g7786 , n7787  );
buf ( g7787 , n7788  );
buf ( g7788 , n7789  );
buf ( g7789 , n7790  );
buf ( g7790 , n7791  );
buf ( g7791 , n7792  );
buf ( g7792 , n7793  );
buf ( g7793 , n7794  );
buf ( g7794 , n7795  );
buf ( g7795 , n7796  );
buf ( g7796 , n7797  );
buf ( g7797 , n7798  );
buf ( g7798 , n7799  );
buf ( g7799 , n7800  );
buf ( g7800 , n7801  );
buf ( g7801 , n7802  );
buf ( g7802 , n7803  );
buf ( g7803 , n7804  );
buf ( g7804 , n7805  );
buf ( g7805 , n7806  );
buf ( g7806 , n7807  );
buf ( g7807 , n7808  );
buf ( g7808 , n7809  );
buf ( g7809 , n7810  );
buf ( g7810 , n7811  );
buf ( g7811 , n7812  );
buf ( g7812 , n7813  );
buf ( g7813 , n7814  );
buf ( g7814 , n7815  );
buf ( g7815 , n7816  );
buf ( g7816 , n7817  );
buf ( g7817 , n7818  );
buf ( g7818 , n7819  );
buf ( g7819 , n7820  );
buf ( g7820 , n7821  );
buf ( g7821 , n7822  );
buf ( g7822 , n7823  );
buf ( g7823 , n7824  );
buf ( g7824 , n7825  );
buf ( g7825 , n7826  );
buf ( g7826 , n7827  );
buf ( g7827 , n7828  );
buf ( g7828 , n7829  );
buf ( g7829 , n7830  );
buf ( g7830 , n7831  );
buf ( g7831 , n7832  );
buf ( g7832 , n7833  );
buf ( g7833 , n7834  );
buf ( g7834 , n7835  );
buf ( g7835 , n7836  );
buf ( g7836 , n7837  );
buf ( g7837 , n7838  );
buf ( g7838 , n7839  );
buf ( g7839 , n7840  );
buf ( g7840 , n7841  );
buf ( g7841 , n7842  );
buf ( g7842 , n7843  );
buf ( g7843 , n7844  );
buf ( g7844 , n7845  );
buf ( g7845 , n7846  );
buf ( g7846 , n7847  );
buf ( g7847 , n7848  );
buf ( g7848 , n7849  );
buf ( g7849 , n7850  );
buf ( g7850 , n7851  );
buf ( g7851 , n7852  );
buf ( g7852 , n7853  );
buf ( g7853 , n7854  );
buf ( g7854 , n7855  );
buf ( g7855 , n7856  );
buf ( g7856 , n7857  );
buf ( g7857 , n7858  );
buf ( g7858 , n7859  );
buf ( g7859 , n7860  );
buf ( g7860 , n7861  );
buf ( g7861 , n7862  );
buf ( g7862 , n7863  );
buf ( g7863 , n7864  );
buf ( g7864 , n7865  );
buf ( g7865 , n7866  );
buf ( g7866 , n7867  );
buf ( g7867 , n7868  );
buf ( g7868 , n7869  );
buf ( g7869 , n7870  );
buf ( g7870 , n7871  );
buf ( g7871 , n7872  );
buf ( g7872 , n7873  );
buf ( g7873 , n7874  );
buf ( g7874 , n7875  );
buf ( g7875 , n7876  );
buf ( g7876 , n7877  );
buf ( g7877 , n7878  );
buf ( g7878 , n7879  );
buf ( g7879 , n7880  );
buf ( g7880 , n7881  );
buf ( g7881 , n7882  );
buf ( g7882 , n7883  );
buf ( g7883 , n7884  );
buf ( g7884 , n7885  );
buf ( g7885 , n7886  );
buf ( g7886 , n7887  );
buf ( g7887 , n7888  );
buf ( g7888 , n7889  );
buf ( g7889 , n7890  );
buf ( g7890 , n7891  );
buf ( g7891 , n7892  );
buf ( g7892 , n7893  );
buf ( g7893 , n7894  );
buf ( g7894 , n7895  );
buf ( g7895 , n7896  );
buf ( g7896 , n7897  );
buf ( g7897 , n7898  );
buf ( g7898 , n7899  );
buf ( g7899 , n7900  );
buf ( g7900 , n7901  );
buf ( g7901 , n7902  );
buf ( g7902 , n7903  );
buf ( g7903 , n7904  );
buf ( g7904 , n7905  );
buf ( g7905 , n7906  );
buf ( g7906 , n7907  );
buf ( g7907 , n7908  );
buf ( g7908 , n7909  );
buf ( g7909 , n7910  );
buf ( g7910 , n7911  );
buf ( g7911 , n7912  );
buf ( g7912 , n7913  );
buf ( g7913 , n7914  );
buf ( g7914 , n7915  );
buf ( g7915 , n7916  );
buf ( g7916 , n7917  );
buf ( g7917 , n7918  );
buf ( g7918 , n7919  );
buf ( g7919 , n7920  );
buf ( g7920 , n7921  );
buf ( g7921 , n7922  );
buf ( g7922 , n7923  );
buf ( g7923 , n7924  );
buf ( g7924 , n7925  );
buf ( g7925 , n7926  );
buf ( g7926 , n7927  );
buf ( g7927 , n7928  );
buf ( g7928 , n7929  );
buf ( g7929 , n7930  );
buf ( g7930 , n7931  );
buf ( g7931 , n7932  );
buf ( g7932 , n7933  );
buf ( g7933 , n7934  );
buf ( g7934 , n7935  );
buf ( g7935 , n7936  );
buf ( g7936 , n7937  );
buf ( g7937 , n7938  );
buf ( g7938 , n7939  );
buf ( g7939 , n7940  );
buf ( g7940 , n7941  );
buf ( g7941 , n7942  );
buf ( g7942 , n7943  );
buf ( g7943 , n7944  );
buf ( g7944 , n7945  );
buf ( g7945 , n7946  );
buf ( g7946 , n7947  );
buf ( g7947 , n7948  );
buf ( g7948 , n7949  );
buf ( g7949 , n7950  );
buf ( g7950 , n7951  );
buf ( g7951 , n7952  );
buf ( g7952 , n7953  );
buf ( g7953 , n7954  );
buf ( g7954 , n7955  );
buf ( g7955 , n7956  );
buf ( g7956 , n7957  );
buf ( g7957 , n7958  );
buf ( g7958 , n7959  );
buf ( g7959 , n7960  );
buf ( g7960 , n7961  );
buf ( g7961 , n7962  );
buf ( g7962 , n7963  );
buf ( g7963 , n7964  );
buf ( g7964 , n7965  );
buf ( g7965 , n7966  );
buf ( g7966 , n7967  );
buf ( g7967 , n7968  );
buf ( g7968 , n7969  );
buf ( g7969 , n7970  );
buf ( g7970 , n7971  );
buf ( g7971 , n7972  );
buf ( g7972 , n7973  );
buf ( g7973 , n7974  );
buf ( g7974 , n7975  );
buf ( g7975 , n7976  );
buf ( g7976 , n7977  );
buf ( g7977 , n7978  );
buf ( g7978 , n7979  );
buf ( g7979 , n7980  );
buf ( g7980 , n7981  );
buf ( g7981 , n7982  );
buf ( g7982 , n7983  );
buf ( g7983 , n7984  );
buf ( g7984 , n7985  );
buf ( g7985 , n7986  );
buf ( g7986 , n7987  );
buf ( g7987 , n7988  );
buf ( g7988 , n7989  );
buf ( g7989 , n7990  );
buf ( g7990 , n7991  );
buf ( g7991 , n7992  );
buf ( g7992 , n7993  );
buf ( g7993 , n7994  );
buf ( g7994 , n7995  );
buf ( g7995 , n7996  );
buf ( g7996 , n7997  );
buf ( g7997 , n7998  );
buf ( g7998 , n7999  );
buf ( g7999 , n8000  );
buf ( g8000 , n8001  );
buf ( g8001 , n8002  );
buf ( g8002 , n8003  );
buf ( g8003 , n8004  );
buf ( g8004 , n8005  );
buf ( g8005 , n8006  );
buf ( g8006 , n8007  );
buf ( g8007 , n8008  );
buf ( g8008 , n8009  );
buf ( g8009 , n8010  );
buf ( g8010 , n8011  );
buf ( g8011 , n8012  );
buf ( g8012 , n8013  );
buf ( g8013 , n8014  );
buf ( g8014 , n8015  );
buf ( g8015 , n8016  );
buf ( g8016 , n8017  );
buf ( g8017 , n8018  );
buf ( g8018 , n8019  );
buf ( g8019 , n8020  );
buf ( g8020 , n8021  );
buf ( g8021 , n8022  );
buf ( g8022 , n8023  );
buf ( g8023 , n8024  );
buf ( g8024 , n8025  );
buf ( g8025 , n8026  );
buf ( g8026 , n8027  );
buf ( g8027 , n8028  );
buf ( g8028 , n8029  );
buf ( g8029 , n8030  );
buf ( g8030 , n8031  );
buf ( g8031 , n8032  );
buf ( g8032 , n8033  );
buf ( g8033 , n8034  );
buf ( g8034 , n8035  );
buf ( g8035 , n8036  );
buf ( g8036 , n8037  );
buf ( g8037 , n8038  );
buf ( g8038 , n8039  );
buf ( g8039 , n8040  );
buf ( g8040 , n8041  );
buf ( g8041 , n8042  );
buf ( g8042 , n8043  );
buf ( g8043 , n8044  );
buf ( g8044 , n8045  );
buf ( g8045 , n8046  );
buf ( g8046 , n8047  );
buf ( g8047 , n8048  );
buf ( g8048 , n8049  );
buf ( g8049 , n8050  );
buf ( g8050 , n8051  );
buf ( g8051 , n8052  );
buf ( g8052 , n8053  );
buf ( g8053 , n8054  );
buf ( g8054 , n8055  );
buf ( g8055 , n8056  );
buf ( g8056 , n8057  );
buf ( g8057 , n8058  );
buf ( g8058 , n8059  );
buf ( g8059 , n8060  );
buf ( g8060 , n8061  );
buf ( g8061 , n8062  );
buf ( g8062 , n8063  );
buf ( g8063 , n8064  );
buf ( g8064 , n8065  );
buf ( g8065 , n8066  );
buf ( g8066 , n8067  );
buf ( g8067 , n8068  );
buf ( g8068 , n8069  );
buf ( g8069 , n8070  );
buf ( g8070 , n8071  );
buf ( g8071 , n8072  );
buf ( g8072 , n8073  );
buf ( g8073 , n8074  );
buf ( g8074 , n8075  );
buf ( g8075 , n8076  );
buf ( g8076 , n8077  );
buf ( g8077 , n8078  );
buf ( g8078 , n8079  );
buf ( g8079 , n8080  );
buf ( g8080 , n8081  );
buf ( g8081 , n8082  );
buf ( g8082 , n8083  );
buf ( g8083 , n8084  );
buf ( g8084 , n8085  );
buf ( g8085 , n8086  );
buf ( g8086 , n8087  );
buf ( g8087 , n8088  );
buf ( g8088 , n8089  );
buf ( g8089 , n8090  );
buf ( g8090 , n8091  );
buf ( g8091 , n8092  );
buf ( g8092 , n8093  );
buf ( g8093 , n8094  );
buf ( g8094 , n8095  );
buf ( g8095 , n8096  );
buf ( g8096 , n8097  );
buf ( g8097 , n8098  );
buf ( g8098 , n8099  );
buf ( g8099 , n8100  );
buf ( g8100 , n8101  );
buf ( g8101 , n8102  );
buf ( g8102 , n8103  );
buf ( g8103 , n8104  );
buf ( g8104 , n8105  );
buf ( g8105 , n8106  );
buf ( g8106 , n8107  );
buf ( g8107 , n8108  );
buf ( g8108 , n8109  );
buf ( g8109 , n8110  );
buf ( g8110 , n8111  );
buf ( g8111 , n8112  );
buf ( g8112 , n8113  );
buf ( g8113 , n8114  );
buf ( g8114 , n8115  );
buf ( g8115 , n8116  );
buf ( g8116 , n8117  );
buf ( g8117 , n8118  );
buf ( g8118 , n8119  );
buf ( g8119 , n8120  );
buf ( g8120 , n8121  );
buf ( g8121 , n8122  );
buf ( g8122 , n8123  );
buf ( g8123 , n8124  );
buf ( g8124 , n8125  );
buf ( g8125 , n8126  );
buf ( g8126 , n8127  );
buf ( g8127 , n8128  );
buf ( g8128 , n8129  );
buf ( g8129 , n8130  );
buf ( g8130 , n8131  );
buf ( g8131 , n8132  );
buf ( g8132 , n8133  );
buf ( g8133 , n8134  );
buf ( g8134 , n8135  );
buf ( g8135 , n8136  );
buf ( g8136 , n8137  );
buf ( g8137 , n8138  );
buf ( g8138 , n8139  );
buf ( g8139 , n8140  );
buf ( g8140 , n8141  );
buf ( g8141 , n8142  );
buf ( g8142 , n8143  );
buf ( g8143 , n8144  );
buf ( g8144 , n8145  );
buf ( g8145 , n8146  );
buf ( g8146 , n8147  );
buf ( g8147 , n8148  );
buf ( g8148 , n8149  );
buf ( g8149 , n8150  );
buf ( g8150 , n8151  );
buf ( g8151 , n8152  );
buf ( g8152 , n8153  );
buf ( g8153 , n8154  );
buf ( g8154 , n8155  );
buf ( g8155 , n8156  );
buf ( g8156 , n8157  );
buf ( g8157 , n8158  );
buf ( g8158 , n8159  );
buf ( g8159 , n8160  );
buf ( g8160 , n8161  );
buf ( g8161 , n8162  );
buf ( g8162 , n8163  );
buf ( g8163 , n8164  );
buf ( g8164 , n8165  );
buf ( g8165 , n8166  );
buf ( g8166 , n8167  );
buf ( g8167 , n8168  );
buf ( g8168 , n8169  );
buf ( g8169 , n8170  );
buf ( g8170 , n8171  );
buf ( g8171 , n8172  );
buf ( g8172 , n8173  );
buf ( g8173 , n8174  );
buf ( g8174 , n8175  );
buf ( g8175 , n8176  );
buf ( g8176 , n8177  );
buf ( g8177 , n8178  );
buf ( g8178 , n8179  );
buf ( g8179 , n8180  );
buf ( g8180 , n8181  );
buf ( g8181 , n8182  );
buf ( g8182 , n8183  );
buf ( g8183 , n8184  );
buf ( g8184 , n8185  );
buf ( g8185 , n8186  );
buf ( g8186 , n8187  );
buf ( g8187 , n8188  );
buf ( g8188 , n8189  );
buf ( g8189 , n8190  );
buf ( g8190 , n8191  );
buf ( g8191 , n8192  );
buf ( g8192 , n8193  );
buf ( g8193 , n8194  );
buf ( g8194 , n8195  );
buf ( g8195 , n8196  );
buf ( g8196 , n8197  );
buf ( g8197 , n8198  );
buf ( g8198 , n8199  );
buf ( g8199 , n8200  );
buf ( g8200 , n8201  );
buf ( g8201 , n8202  );
buf ( g8202 , n8203  );
buf ( g8203 , n8204  );
buf ( g8204 , n8205  );
buf ( g8205 , n8206  );
buf ( g8206 , n8207  );
buf ( g8207 , n8208  );
buf ( g8208 , n8209  );
buf ( g8209 , n8210  );
buf ( g8210 , n8211  );
buf ( g8211 , n8212  );
buf ( g8212 , n8213  );
buf ( g8213 , n8214  );
buf ( g8214 , n8215  );
buf ( g8215 , n8216  );
buf ( g8216 , n8217  );
buf ( g8217 , n8218  );
buf ( g8218 , n8219  );
buf ( g8219 , n8220  );
buf ( g8220 , n8221  );
buf ( g8221 , n8222  );
buf ( g8222 , n8223  );
buf ( g8223 , n8224  );
buf ( g8224 , n8225  );
buf ( g8225 , n8226  );
buf ( g8226 , n8227  );
buf ( g8227 , n8228  );
buf ( g8228 , n8229  );
buf ( g8229 , n8230  );
buf ( g8230 , n8231  );
buf ( g8231 , n8232  );
buf ( g8232 , n8233  );
buf ( g8233 , n8234  );
buf ( g8234 , n8235  );
buf ( g8235 , n8236  );
buf ( g8236 , n8237  );
buf ( g8237 , n8238  );
buf ( g8238 , n8239  );
buf ( g8239 , n8240  );
buf ( g8240 , n8241  );
buf ( g8241 , n8242  );
buf ( g8242 , n8243  );
buf ( g8243 , n8244  );
buf ( g8244 , n8245  );
buf ( g8245 , n8246  );
buf ( g8246 , n8247  );
buf ( g8247 , n8248  );
buf ( g8248 , n8249  );
buf ( g8249 , n8250  );
buf ( g8250 , n8251  );
buf ( g8251 , n8252  );
buf ( g8252 , n8253  );
buf ( g8253 , n8254  );
buf ( g8254 , n8255  );
buf ( g8255 , n8256  );
buf ( g8256 , n8257  );
buf ( g8257 , n8258  );
buf ( g8258 , n8259  );
buf ( g8259 , n8260  );
buf ( g8260 , n8261  );
buf ( g8261 , n8262  );
buf ( g8262 , n8263  );
buf ( g8263 , n8264  );
buf ( g8264 , n8265  );
buf ( g8265 , n8266  );
buf ( g8266 , n8267  );
buf ( g8267 , n8268  );
buf ( g8268 , n8269  );
buf ( g8269 , n8270  );
buf ( g8270 , n8271  );
buf ( g8271 , n8272  );
buf ( g8272 , n8273  );
buf ( g8273 , n8274  );
buf ( g8274 , n8275  );
buf ( g8275 , n8276  );
buf ( g8276 , n8277  );
buf ( g8277 , n8278  );
buf ( g8278 , n8279  );
buf ( g8279 , n8280  );
buf ( g8280 , n8281  );
buf ( g8281 , n8282  );
buf ( g8282 , n8283  );
buf ( g8283 , n8284  );
buf ( g8284 , n8285  );
buf ( g8285 , n8286  );
buf ( g8286 , n8287  );
buf ( g8287 , n8288  );
buf ( g8288 , n8289  );
buf ( g8289 , n8290  );
buf ( g8290 , n8291  );
buf ( g8291 , n8292  );
buf ( g8292 , n8293  );
buf ( g8293 , n8294  );
buf ( g8294 , n8295  );
buf ( g8295 , n8296  );
buf ( g8296 , n8297  );
buf ( g8297 , n8298  );
buf ( g8298 , n8299  );
buf ( g8299 , n8300  );
buf ( g8300 , n8301  );
buf ( g8301 , n8302  );
buf ( g8302 , n8303  );
buf ( g8303 , n8304  );
buf ( g8304 , n8305  );
buf ( g8305 , n8306  );
buf ( g8306 , n8307  );
buf ( g8307 , n8308  );
buf ( g8308 , n8309  );
buf ( g8309 , n8310  );
buf ( g8310 , n8311  );
buf ( g8311 , n8312  );
buf ( g8312 , n8313  );
buf ( g8313 , n8314  );
buf ( g8314 , n8315  );
buf ( g8315 , n8316  );
buf ( g8316 , n8317  );
buf ( g8317 , n8318  );
buf ( g8318 , n8319  );
buf ( g8319 , n8320  );
buf ( g8320 , n8321  );
buf ( g8321 , n8322  );
buf ( g8322 , n8323  );
buf ( g8323 , n8324  );
buf ( g8324 , n8325  );
buf ( g8325 , n8326  );
buf ( g8326 , n8327  );
buf ( g8327 , n8328  );
buf ( g8328 , n8329  );
buf ( g8329 , n8330  );
buf ( g8330 , n8331  );
buf ( g8331 , n8332  );
buf ( g8332 , n8333  );
buf ( g8333 , n8334  );
buf ( g8334 , n8335  );
buf ( g8335 , n8336  );
buf ( g8336 , n8337  );
buf ( g8337 , n8338  );
buf ( g8338 , n8339  );
buf ( g8339 , n8340  );
buf ( g8340 , n8341  );
buf ( g8341 , n8342  );
buf ( g8342 , n8343  );
buf ( g8343 , n8344  );
buf ( g8344 , n8345  );
buf ( g8345 , n8346  );
buf ( g8346 , n8347  );
buf ( g8347 , n8348  );
buf ( g8348 , n8349  );
buf ( g8349 , n8350  );
buf ( g8350 , n8351  );
buf ( g8351 , n8352  );
buf ( g8352 , n8353  );
buf ( g8353 , n8354  );
buf ( g8354 , n8355  );
buf ( g8355 , n8356  );
buf ( g8356 , n8357  );
buf ( g8357 , n8358  );
buf ( g8358 , n8359  );
buf ( g8359 , n8360  );
buf ( g8360 , n8361  );
buf ( g8361 , n8362  );
buf ( g8362 , n8363  );
buf ( g8363 , n8364  );
buf ( g8364 , n8365  );
buf ( g8365 , n8366  );
buf ( g8366 , n8367  );
buf ( g8367 , n8368  );
buf ( g8368 , n8369  );
buf ( g8369 , n8370  );
buf ( g8370 , n8371  );
buf ( g8371 , n8372  );
buf ( g8372 , n8373  );
buf ( g8373 , n8374  );
buf ( g8374 , n8375  );
buf ( g8375 , n8376  );
buf ( g8376 , n8377  );
buf ( g8377 , n8378  );
buf ( g8378 , n8379  );
buf ( g8379 , n8380  );
buf ( g8380 , n8381  );
buf ( g8381 , n8382  );
buf ( g8382 , n8383  );
buf ( g8383 , n8384  );
buf ( g8384 , n8385  );
buf ( g8385 , n8386  );
buf ( g8386 , n8387  );
buf ( g8387 , n8388  );
buf ( g8388 , n8389  );
buf ( g8389 , n8390  );
buf ( g8390 , n8391  );
buf ( g8391 , n8392  );
buf ( g8392 , n8393  );
buf ( g8393 , n8394  );
buf ( g8394 , n8395  );
buf ( g8395 , n8396  );
buf ( g8396 , n8397  );
buf ( g8397 , n8398  );
buf ( g8398 , n8399  );
buf ( g8399 , n8400  );
buf ( g8400 , n8401  );
buf ( g8401 , n8402  );
buf ( g8402 , n8403  );
buf ( g8403 , n8404  );
buf ( g8404 , n8405  );
buf ( g8405 , n8406  );
buf ( g8406 , n8407  );
buf ( g8407 , n8408  );
buf ( g8408 , n8409  );
buf ( g8409 , n8410  );
buf ( g8410 , n8411  );
buf ( g8411 , n8412  );
buf ( g8412 , n8413  );
buf ( g8413 , n8414  );
buf ( g8414 , n8415  );
buf ( g8415 , n8416  );
buf ( g8416 , n8417  );
buf ( g8417 , n8418  );
buf ( g8418 , n8419  );
buf ( g8419 , n8420  );
buf ( g8420 , n8421  );
buf ( g8421 , n8422  );
buf ( g8422 , n8423  );
buf ( g8423 , n8424  );
buf ( g8424 , n8425  );
buf ( g8425 , n8426  );
buf ( g8426 , n8427  );
buf ( g8427 , n8428  );
buf ( g8428 , n8429  );
buf ( g8429 , n8430  );
buf ( g8430 , n8431  );
buf ( g8431 , n8432  );
buf ( g8432 , n8433  );
buf ( g8433 , n8434  );
buf ( g8434 , n8435  );
buf ( g8435 , n8436  );
buf ( g8436 , n8437  );
buf ( g8437 , n8438  );
buf ( g8438 , n8439  );
buf ( g8439 , n8440  );
buf ( g8440 , n8441  );
buf ( g8441 , n8442  );
buf ( g8442 , n8443  );
buf ( g8443 , n8444  );
buf ( g8444 , n8445  );
buf ( g8445 , n8446  );
buf ( g8446 , n8447  );
buf ( g8447 , n8448  );
buf ( g8448 , n8449  );
buf ( g8449 , n8450  );
buf ( g8450 , n8451  );
buf ( g8451 , n8452  );
buf ( g8452 , n8453  );
buf ( g8453 , n8454  );
buf ( g8454 , n8455  );
buf ( g8455 , n8456  );
buf ( g8456 , n8457  );
buf ( g8457 , n8458  );
buf ( g8458 , n8459  );
buf ( g8459 , n8460  );
buf ( g8460 , n8461  );
buf ( g8461 , n8462  );
buf ( g8462 , n8463  );
buf ( g8463 , n8464  );
buf ( g8464 , n8465  );
buf ( g8465 , n8466  );
buf ( g8466 , n8467  );
buf ( g8467 , n8468  );
buf ( g8468 , n8469  );
buf ( g8469 , n8470  );
buf ( g8470 , n8471  );
buf ( g8471 , n8472  );
buf ( g8472 , n8473  );
buf ( g8473 , n8474  );
buf ( g8474 , n8475  );
buf ( g8475 , n8476  );
buf ( g8476 , n8477  );
buf ( g8477 , n8478  );
buf ( g8478 , n8479  );
buf ( g8479 , n8480  );
buf ( g8480 , n8481  );
buf ( g8481 , n8482  );
buf ( g8482 , n8483  );
buf ( g8483 , n8484  );
buf ( g8484 , n8485  );
buf ( g8485 , n8486  );
buf ( g8486 , n8487  );
buf ( g8487 , n8488  );
buf ( g8488 , n8489  );
buf ( g8489 , n8490  );
buf ( g8490 , n8491  );
buf ( g8491 , n8492  );
buf ( g8492 , n8493  );
buf ( g8493 , n8494  );
buf ( g8494 , n8495  );
buf ( g8495 , n8496  );
buf ( g8496 , n8497  );
buf ( g8497 , n8498  );
buf ( g8498 , n8499  );
buf ( g8499 , n8500  );
buf ( g8500 , n8501  );
buf ( g8501 , n8502  );
buf ( g8502 , n8503  );
buf ( g8503 , n8504  );
buf ( g8504 , n8505  );
buf ( g8505 , n8506  );
buf ( g8506 , n8507  );
buf ( g8507 , n8508  );
buf ( g8508 , n8509  );
buf ( g8509 , n8510  );
buf ( g8510 , n8511  );
buf ( g8511 , n8512  );
buf ( g8512 , n8513  );
buf ( g8513 , n8514  );
buf ( g8514 , n8515  );
buf ( g8515 , n8516  );
buf ( g8516 , n8517  );
buf ( g8517 , n8518  );
buf ( g8518 , n8519  );
buf ( g8519 , n8520  );
buf ( g8520 , n8521  );
buf ( g8521 , n8522  );
buf ( g8522 , n8523  );
buf ( g8523 , n8524  );
buf ( g8524 , n8525  );
buf ( g8525 , n8526  );
buf ( g8526 , n8527  );
buf ( g8527 , n8528  );
buf ( g8528 , n8529  );
buf ( g8529 , n8530  );
buf ( g8530 , n8531  );
buf ( g8531 , n8532  );
buf ( g8532 , n8533  );
buf ( g8533 , n8534  );
buf ( g8534 , n8535  );
buf ( g8535 , n8536  );
buf ( g8536 , n8537  );
buf ( g8537 , n8538  );
buf ( g8538 , n8539  );
buf ( g8539 , n8540  );
buf ( g8540 , n8541  );
buf ( g8541 , n8542  );
buf ( g8542 , n8543  );
buf ( g8543 , n8544  );
buf ( g8544 , n8545  );
buf ( g8545 , n8546  );
buf ( g8546 , n8547  );
buf ( g8547 , n8548  );
buf ( g8548 , n8549  );
buf ( g8549 , n8550  );
buf ( g8550 , n8551  );
buf ( g8551 , n8552  );
buf ( g8552 , n8553  );
buf ( g8553 , n8554  );
buf ( g8554 , n8555  );
buf ( g8555 , n8556  );
buf ( g8556 , n8557  );
buf ( g8557 , n8558  );
buf ( g8558 , n8559  );
buf ( g8559 , n8560  );
buf ( g8560 , n8561  );
buf ( g8561 , n8562  );
buf ( g8562 , n8563  );
buf ( g8563 , n8564  );
buf ( g8564 , n8565  );
buf ( g8565 , n8566  );
buf ( g8566 , n8567  );
buf ( g8567 , n8568  );
buf ( g8568 , n8569  );
buf ( g8569 , n8570  );
buf ( g8570 , n8571  );
buf ( g8571 , n8572  );
buf ( g8572 , n8573  );
buf ( g8573 , n8574  );
buf ( g8574 , n8575  );
buf ( g8575 , n8576  );
buf ( g8576 , n8577  );
buf ( g8577 , n8578  );
buf ( g8578 , n8579  );
buf ( g8579 , n8580  );
buf ( g8580 , n8581  );
buf ( g8581 , n8582  );
buf ( g8582 , n8583  );
buf ( g8583 , n8584  );
buf ( g8584 , n8585  );
buf ( g8585 , n8586  );
buf ( g8586 , n8587  );
buf ( g8587 , n8588  );
buf ( g8588 , n8589  );
buf ( g8589 , n8590  );
buf ( g8590 , n8591  );
buf ( g8591 , n8592  );
buf ( g8592 , n8593  );
buf ( g8593 , n8594  );
buf ( g8594 , n8595  );
buf ( g8595 , n8596  );
buf ( g8596 , n8597  );
buf ( g8597 , n8598  );
buf ( g8598 , n8599  );
buf ( g8599 , n8600  );
buf ( g8600 , n8601  );
buf ( g8601 , n8602  );
buf ( g8602 , n8603  );
buf ( g8603 , n8604  );
buf ( g8604 , n8605  );
buf ( g8605 , n8606  );
buf ( g8606 , n8607  );
buf ( g8607 , n8608  );
buf ( g8608 , n8609  );
buf ( g8609 , n8610  );
buf ( g8610 , n8611  );
buf ( g8611 , n8612  );
buf ( g8612 , n8613  );
buf ( g8613 , n8614  );
buf ( g8614 , n8615  );
buf ( g8615 , n8616  );
buf ( g8616 , n8617  );
buf ( g8617 , n8618  );
buf ( g8618 , n8619  );
buf ( g8619 , n8620  );
buf ( g8620 , n8621  );
buf ( g8621 , n8622  );
buf ( g8622 , n8623  );
buf ( g8623 , n8624  );
buf ( g8624 , n8625  );
buf ( g8625 , n8626  );
buf ( g8626 , n8627  );
buf ( g8627 , n8628  );
buf ( g8628 , n8629  );
buf ( g8629 , n8630  );
buf ( g8630 , n8631  );
buf ( g8631 , n8632  );
buf ( g8632 , n8633  );
buf ( g8633 , n8634  );
buf ( g8634 , n8635  );
buf ( g8635 , n8636  );
buf ( g8636 , n8637  );
buf ( g8637 , n8638  );
buf ( g8638 , n8639  );
buf ( g8639 , n8640  );
buf ( g8640 , n8641  );
buf ( g8641 , n8642  );
buf ( g8642 , n8643  );
buf ( g8643 , n8644  );
buf ( g8644 , n8645  );
buf ( g8645 , n8646  );
buf ( g8646 , n8647  );
buf ( g8647 , n8648  );
buf ( g8648 , n8649  );
buf ( g8649 , n8650  );
buf ( g8650 , n8651  );
buf ( g8651 , n8652  );
buf ( g8652 , n8653  );
buf ( g8653 , n8654  );
buf ( g8654 , n8655  );
buf ( g8655 , n8656  );
buf ( g8656 , n8657  );
buf ( g8657 , n8658  );
buf ( g8658 , n8659  );
buf ( g8659 , n8660  );
buf ( g8660 , n8661  );
buf ( g8661 , n8662  );
buf ( g8662 , n8663  );
buf ( g8663 , n8664  );
buf ( g8664 , n8665  );
buf ( g8665 , n8666  );
buf ( g8666 , n8667  );
buf ( g8667 , n8668  );
buf ( g8668 , n8669  );
buf ( g8669 , n8670  );
buf ( g8670 , n8671  );
buf ( g8671 , n8672  );
buf ( g8672 , n8673  );
buf ( g8673 , n8674  );
buf ( g8674 , n8675  );
buf ( g8675 , n8676  );
buf ( g8676 , n8677  );
buf ( g8677 , n8678  );
buf ( g8678 , n8679  );
buf ( g8679 , n8680  );
buf ( g8680 , n8681  );
buf ( g8681 , n8682  );
buf ( g8682 , n8683  );
buf ( g8683 , n8684  );
buf ( g8684 , n8685  );
buf ( g8685 , n8686  );
buf ( g8686 , n8687  );
buf ( g8687 , n8688  );
buf ( g8688 , n8689  );
buf ( g8689 , n8690  );
buf ( g8690 , n8691  );
buf ( g8691 , n8692  );
buf ( g8692 , n8693  );
buf ( g8693 , n8694  );
buf ( g8694 , n8695  );
buf ( g8695 , n8696  );
buf ( g8696 , n8697  );
buf ( g8697 , n8698  );
buf ( g8698 , n8699  );
buf ( g8699 , n8700  );
buf ( g8700 , n8701  );
buf ( g8701 , n8702  );
buf ( g8702 , n8703  );
buf ( g8703 , n8704  );
buf ( g8704 , n8705  );
buf ( g8705 , n8706  );
buf ( g8706 , n8707  );
buf ( g8707 , n8708  );
buf ( g8708 , n8709  );
buf ( g8709 , n8710  );
buf ( g8710 , n8711  );
buf ( g8711 , n8712  );
buf ( g8712 , n8713  );
buf ( g8713 , n8714  );
buf ( g8714 , n8715  );
buf ( g8715 , n8716  );
buf ( g8716 , n8717  );
buf ( g8717 , n8718  );
buf ( g8718 , n8719  );
buf ( g8719 , n8720  );
buf ( g8720 , n8721  );
buf ( g8721 , n8722  );
buf ( g8722 , n8723  );
buf ( g8723 , n8724  );
buf ( g8724 , n8725  );
buf ( g8725 , n8726  );
buf ( g8726 , n8727  );
buf ( g8727 , n8728  );
buf ( g8728 , n8729  );
buf ( g8729 , n8730  );
buf ( g8730 , n8731  );
buf ( g8731 , n8732  );
buf ( g8732 , n8733  );
buf ( g8733 , n8734  );
buf ( g8734 , n8735  );
buf ( g8735 , n8736  );
buf ( g8736 , n8737  );
buf ( g8737 , n8738  );
buf ( g8738 , n8739  );
buf ( g8739 , n8740  );
buf ( g8740 , n8741  );
buf ( g8741 , n8742  );
buf ( g8742 , n8743  );
buf ( g8743 , n8744  );
buf ( g8744 , n8745  );
buf ( g8745 , n8746  );
buf ( g8746 , n8747  );
buf ( g8747 , n8748  );
buf ( g8748 , n8749  );
buf ( g8749 , n8750  );
buf ( g8750 , n8751  );
buf ( g8751 , n8752  );
buf ( g8752 , n8753  );
buf ( g8753 , n8754  );
buf ( g8754 , n8755  );
buf ( g8755 , n8756  );
buf ( g8756 , n8757  );
buf ( g8757 , n8758  );
buf ( g8758 , n8759  );
buf ( g8759 , n8760  );
buf ( g8760 , n8761  );
buf ( g8761 , n8762  );
buf ( g8762 , n8763  );
buf ( g8763 , n8764  );
buf ( g8764 , n8765  );
buf ( g8765 , n8766  );
buf ( g8766 , n8767  );
buf ( g8767 , n8768  );
buf ( g8768 , n8769  );
buf ( g8769 , n8770  );
buf ( g8770 , n8771  );
buf ( g8771 , n8772  );
buf ( g8772 , n8773  );
buf ( g8773 , n8774  );
buf ( g8774 , n8775  );
buf ( g8775 , n8776  );
buf ( g8776 , n8777  );
buf ( g8777 , n8778  );
buf ( g8778 , n8779  );
buf ( g8779 , n8780  );
buf ( g8780 , n8781  );
buf ( g8781 , n8782  );
buf ( g8782 , n8783  );
buf ( g8783 , n8784  );
buf ( g8784 , n8785  );
buf ( g8785 , n8786  );
buf ( g8786 , n8787  );
buf ( g8787 , n8788  );
buf ( g8788 , n8789  );
buf ( g8789 , n8790  );
buf ( g8790 , n8791  );
buf ( g8791 , n8792  );
buf ( g8792 , n8793  );
buf ( g8793 , n8794  );
buf ( g8794 , n8795  );
buf ( g8795 , n8796  );
buf ( g8796 , n8797  );
buf ( g8797 , n8798  );
buf ( g8798 , n8799  );
buf ( g8799 , n8800  );
buf ( g8800 , n8801  );
buf ( g8801 , n8802  );
buf ( g8802 , n8803  );
buf ( g8803 , n8804  );
buf ( g8804 , n8805  );
buf ( g8805 , n8806  );
buf ( g8806 , n8807  );
buf ( g8807 , n8808  );
buf ( g8808 , n8809  );
buf ( g8809 , n8810  );
buf ( g8810 , n8811  );
buf ( g8811 , n8812  );
buf ( g8812 , n8813  );
buf ( g8813 , n8814  );
buf ( g8814 , n8815  );
buf ( g8815 , n8816  );
buf ( g8816 , n8817  );
buf ( g8817 , n8818  );
buf ( g8818 , n8819  );
buf ( g8819 , n8820  );
buf ( g8820 , n8821  );
buf ( g8821 , n8822  );
buf ( g8822 , n8823  );
buf ( g8823 , n8824  );
buf ( g8824 , n8825  );
buf ( g8825 , n8826  );
buf ( g8826 , n8827  );
buf ( g8827 , n8828  );
buf ( g8828 , n8829  );
buf ( g8829 , n8830  );
buf ( g8830 , n8831  );
buf ( g8831 , n8832  );
buf ( g8832 , n8833  );
buf ( g8833 , n8834  );
buf ( g8834 , n8835  );
buf ( g8835 , n8836  );
buf ( g8836 , n8837  );
buf ( g8837 , n8838  );
buf ( g8838 , n8839  );
buf ( g8839 , n8840  );
buf ( g8840 , n8841  );
buf ( g8841 , n8842  );
buf ( g8842 , n8843  );
buf ( g8843 , n8844  );
buf ( g8844 , n8845  );
buf ( g8845 , n8846  );
buf ( g8846 , n8847  );
buf ( g8847 , n8848  );
buf ( g8848 , n8849  );
buf ( g8849 , n8850  );
buf ( g8850 , n8851  );
buf ( g8851 , n8852  );
buf ( g8852 , n8853  );
buf ( g8853 , n8854  );
buf ( g8854 , n8855  );
buf ( g8855 , n8856  );
buf ( g8856 , n8857  );
buf ( g8857 , n8858  );
buf ( g8858 , n8859  );
buf ( g8859 , n8860  );
buf ( g8860 , n8861  );
buf ( g8861 , n8862  );
buf ( g8862 , n8863  );
buf ( g8863 , n8864  );
buf ( g8864 , n8865  );
buf ( g8865 , n8866  );
buf ( g8866 , n8867  );
buf ( g8867 , n8868  );
buf ( g8868 , n8869  );
buf ( g8869 , n8870  );
buf ( g8870 , n8871  );
buf ( g8871 , n8872  );
buf ( g8872 , n8873  );
buf ( g8873 , n8874  );
buf ( g8874 , n8875  );
buf ( g8875 , n8876  );
buf ( g8876 , n8877  );
buf ( g8877 , n8878  );
buf ( g8878 , n8879  );
buf ( g8879 , n8880  );
buf ( g8880 , n8881  );
buf ( g8881 , n8882  );
buf ( g8882 , n8883  );
buf ( g8883 , n8884  );
buf ( g8884 , n8885  );
buf ( g8885 , n8886  );
buf ( g8886 , n8887  );
buf ( g8887 , n8888  );
buf ( g8888 , n8889  );
buf ( g8889 , n8890  );
buf ( g8890 , n8891  );
buf ( g8891 , n8892  );
buf ( g8892 , n8893  );
buf ( g8893 , n8894  );
buf ( g8894 , n8895  );
buf ( g8895 , n8896  );
buf ( g8896 , n8897  );
buf ( g8897 , n8898  );
buf ( g8898 , n8899  );
buf ( g8899 , n8900  );
buf ( g8900 , n8901  );
buf ( g8901 , n8902  );
buf ( g8902 , n8903  );
buf ( g8903 , n8904  );
buf ( g8904 , n8905  );
buf ( g8905 , n8906  );
buf ( g8906 , n8907  );
buf ( g8907 , n8908  );
buf ( g8908 , n8909  );
buf ( g8909 , n8910  );
buf ( g8910 , n8911  );
buf ( g8911 , n8912  );
buf ( g8912 , n8913  );
buf ( g8913 , n8914  );
buf ( g8914 , n8915  );
buf ( g8915 , n8916  );
buf ( g8916 , n8917  );
buf ( g8917 , n8918  );
buf ( g8918 , n8919  );
buf ( g8919 , n8920  );
buf ( g8920 , n8921  );
buf ( g8921 , n8922  );
buf ( g8922 , n8923  );
buf ( g8923 , n8924  );
buf ( g8924 , n8925  );
buf ( g8925 , n8926  );
buf ( g8926 , n8927  );
buf ( g8927 , n8928  );
buf ( g8928 , n8929  );
buf ( g8929 , n8930  );
buf ( g8930 , n8931  );
buf ( g8931 , n8932  );
buf ( g8932 , n8933  );
buf ( g8933 , n8934  );
buf ( g8934 , n8935  );
buf ( g8935 , n8936  );
buf ( g8936 , n8937  );
buf ( g8937 , n8938  );
buf ( g8938 , n8939  );
buf ( g8939 , n8940  );
buf ( g8940 , n8941  );
buf ( g8941 , n8942  );
buf ( g8942 , n8943  );
buf ( g8943 , n8944  );
buf ( g8944 , n8945  );
buf ( g8945 , n8946  );
buf ( g8946 , n8947  );
buf ( g8947 , n8948  );
buf ( g8948 , n8949  );
buf ( g8949 , n8950  );
buf ( g8950 , n8951  );
buf ( g8951 , n8952  );
buf ( g8952 , n8953  );
buf ( g8953 , n8954  );
buf ( g8954 , n8955  );
buf ( g8955 , n8956  );
buf ( g8956 , n8957  );
buf ( g8957 , n8958  );
buf ( g8958 , n8959  );
buf ( g8959 , n8960  );
buf ( g8960 , n8961  );
buf ( g8961 , n8962  );
buf ( g8962 , n8963  );
buf ( g8963 , n8964  );
buf ( g8964 , n8965  );
buf ( g8965 , n8966  );
buf ( g8966 , n8967  );
buf ( g8967 , n8968  );
buf ( g8968 , n8969  );
buf ( g8969 , n8970  );
buf ( g8970 , n8971  );
buf ( g8971 , n8972  );
buf ( g8972 , n8973  );
buf ( g8973 , n8974  );
buf ( g8974 , n8975  );
buf ( g8975 , n8976  );
buf ( g8976 , n8977  );
buf ( g8977 , n8978  );
buf ( g8978 , n8979  );
buf ( n1875 , n1081 );
buf ( n1876 , n1080 );
buf ( n1877 , n1085 );
buf ( n1878 , n1036 );
buf ( n1879 , n1084 );
buf ( n1880 , n1017 );
buf ( n1881 , n1011 );
buf ( n1882 , n1035 );
buf ( n1883 , n898 );
buf ( n1884 , n910 );
buf ( n1885 , n1037 );
buf ( n1886 , n1038 );
buf ( n1887 , n1039 );
buf ( n1888 , n1042 );
buf ( n1889 , n1043 );
buf ( n1890 , n1034 );
buf ( n1891 , n1118 );
buf ( n1892 , n1355 );
buf ( n1893 , n1117 );
buf ( n1894 , n1093 );
buf ( n1895 , n1090 );
buf ( n1896 , n1101 );
buf ( n1897 , n1091 );
buf ( n1898 , n913 );
buf ( n1899 , n911 );
buf ( n1900 , n1040 );
buf ( n1901 , n1041 );
buf ( n1902 , n1031 );
buf ( n1903 , n772 );
buf ( n1904 , n795 );
buf ( n1905 , n690 );
buf ( n1906 , n790 );
buf ( n1907 , n385 );
buf ( n1908 , n1149 );
buf ( n1909 , n1144 );
buf ( n1910 , 1'b0 );
buf ( n1911 , 1'b0 );
buf ( n1912 , 1'b0 );
buf ( n1913 , 1'b0 );
buf ( n1914 , 1'b0 );
buf ( n1915 , 1'b0 );
buf ( n1916 , 1'b0 );
buf ( n1917 , 1'b0 );
buf ( n1918 , 1'b0 );
buf ( n1919 , 1'b0 );
buf ( n1920 , 1'b0 );
buf ( n1921 , 1'b0 );
buf ( n1922 , n216 );
buf ( n1923 , n213 );
buf ( n1924 , n201 );
buf ( n1925 , n214 );
buf ( n1926 , n1830 );
buf ( n1927 , n2 );
buf ( n1928 , n130 );
buf ( n1929 , n132 );
buf ( n1930 , n155 );
buf ( n1931 , n146 );
buf ( n1932 , n129 );
buf ( n1933 , n131 );
buf ( n1934 , n149 );
buf ( n1935 , n150 );
buf ( n1936 , n176 );
buf ( n1937 , n1104 );
buf ( n1938 , n1029 );
buf ( n1939 , n30025 );
buf ( n1940 , n1105 );
buf ( n1941 , n1114 );
buf ( n1942 , n1836 );
buf ( n1943 , n1835 );
buf ( n1944 , n1839 );
buf ( n1945 , n1844 );
buf ( n1946 , n1837 );
buf ( n1947 , n16040 );
buf ( n1948 , n15908 );
buf ( n1949 , n15913 );
buf ( n1950 , n15917 );
buf ( n1951 , n15922 );
buf ( n1952 , n15926 );
buf ( n1953 , n15930 );
buf ( n1954 , n15934 );
buf ( n1955 , n15938 );
buf ( n1956 , n15942 );
buf ( n1957 , n15946 );
buf ( n1958 , n15950 );
buf ( n1959 , n15956 );
buf ( n1960 , n15960 );
buf ( n1961 , n15964 );
buf ( n1962 , n15968 );
buf ( n1963 , n15972 );
buf ( n1964 , n15976 );
buf ( n1965 , n16068 );
buf ( n1966 , n15980 );
buf ( n1967 , n15984 );
buf ( n1968 , n15988 );
buf ( n1969 , n15992 );
buf ( n1970 , n15996 );
buf ( n1971 , n16000 );
buf ( n1972 , n16004 );
buf ( n1973 , n16008 );
buf ( n1974 , n16012 );
buf ( n1975 , n16016 );
buf ( n1976 , n16020 );
buf ( n1977 , n16024 );
buf ( n1978 , n16028 );
buf ( n1979 , n16032 );
buf ( n1980 , n16036 );
buf ( n1981 , n16084 );
buf ( n1982 , n16044 );
buf ( n1983 , n16048 );
buf ( n1984 , n16052 );
buf ( n1985 , n16056 );
buf ( n1986 , n16060 );
buf ( n1987 , n15904 );
buf ( n1988 , n16064 );
buf ( n1989 , n16088 );
buf ( n1990 , n16072 );
buf ( n1991 , n16076 );
buf ( n1992 , n16080 );
buf ( n1993 , n16092 );
buf ( n1994 , 1'b1 );
buf ( n1995 , n15287 );
buf ( n1996 , 1'b0 );
buf ( n1997 , 1'b0 );
buf ( n1998 , n30355 );
buf ( n1999 , n14878 );
buf ( n2000 , 1'b0 );
buf ( n2001 , 1'b0 );
buf ( n2002 , n30357 );
buf ( n2003 , n16112 );
buf ( n2004 , 1'b0 );
buf ( n2005 , 1'b0 );
buf ( n2006 , n30375 );
buf ( n2007 , n14900 );
buf ( n2008 , 1'b0 );
buf ( n2009 , 1'b0 );
buf ( n2010 , n30340 );
buf ( n2011 , n14919 );
buf ( n2012 , 1'b0 );
buf ( n2013 , 1'b0 );
buf ( n2014 , n30348 );
buf ( n2015 , n20612 );
buf ( n2016 , 1'b0 );
buf ( n2017 , 1'b0 );
buf ( n2018 , n30374 );
buf ( n2019 , n26524 );
buf ( n2020 , 1'b0 );
buf ( n2021 , 1'b0 );
buf ( n2022 , n30355 );
buf ( n2023 , n20620 );
buf ( n2024 , 1'b0 );
buf ( n2025 , 1'b0 );
buf ( n2026 , n30372 );
buf ( n2027 , n12824 );
buf ( n2028 , 1'b0 );
buf ( n2029 , 1'b0 );
buf ( n2030 , n30358 );
buf ( n2031 , n21784 );
buf ( n2032 , 1'b0 );
buf ( n2033 , 1'b0 );
buf ( n2034 , n30358 );
buf ( n2035 , n13201 );
buf ( n2036 , 1'b0 );
buf ( n2037 , 1'b0 );
buf ( n2038 , n30355 );
buf ( n2039 , n13851 );
buf ( n2040 , 1'b0 );
buf ( n2041 , 1'b0 );
buf ( n2042 , n30345 );
buf ( n2043 , n12729 );
buf ( n2044 , 1'b0 );
buf ( n2045 , 1'b0 );
buf ( n2046 , n30347 );
buf ( n2047 , n28007 );
buf ( n2048 , 1'b0 );
buf ( n2049 , 1'b0 );
buf ( n2050 , n30347 );
buf ( n2051 , n13515 );
buf ( n2052 , 1'b0 );
buf ( n2053 , 1'b0 );
buf ( n2054 , n30375 );
buf ( n2055 , n13460 );
buf ( n2056 , 1'b0 );
buf ( n2057 , 1'b0 );
buf ( n2058 , n30378 );
buf ( n2059 , n12764 );
buf ( n2060 , 1'b0 );
buf ( n2061 , 1'b0 );
buf ( n2062 , n30375 );
buf ( n2063 , n13922 );
buf ( n2064 , 1'b0 );
buf ( n2065 , 1'b0 );
buf ( n2066 , n30347 );
buf ( n2067 , n16483 );
buf ( n2068 , 1'b0 );
buf ( n2069 , 1'b0 );
buf ( n2070 , n30378 );
buf ( n2071 , n13443 );
buf ( n2072 , 1'b0 );
buf ( n2073 , 1'b0 );
buf ( n2074 , n30374 );
buf ( n2075 , n13936 );
buf ( n2076 , 1'b0 );
buf ( n2077 , 1'b0 );
buf ( n2078 , n30376 );
buf ( n2079 , n14823 );
buf ( n2080 , 1'b0 );
buf ( n2081 , 1'b0 );
buf ( n2082 , n30345 );
buf ( n2083 , n15304 );
buf ( n2084 , 1'b0 );
buf ( n2085 , 1'b0 );
buf ( n2086 , n30375 );
buf ( n2087 , n13978 );
buf ( n2088 , 1'b0 );
buf ( n2089 , 1'b0 );
buf ( n2090 , n30358 );
buf ( n2091 , n14394 );
buf ( n2092 , 1'b0 );
buf ( n2093 , 1'b0 );
buf ( n2094 , n30372 );
buf ( n2095 , n18866 );
buf ( n2096 , 1'b0 );
buf ( n2097 , 1'b0 );
buf ( n2098 , n30358 );
buf ( n2099 , n13993 );
buf ( n2100 , 1'b0 );
buf ( n2101 , 1'b0 );
buf ( n2102 , n30347 );
buf ( n2103 , n16497 );
buf ( n2104 , 1'b0 );
buf ( n2105 , 1'b0 );
buf ( n2106 , n30374 );
buf ( n2107 , n14003 );
buf ( n2108 , 1'b0 );
buf ( n2109 , 1'b0 );
buf ( n2110 , n30345 );
buf ( n2111 , n14626 );
buf ( n2112 , 1'b0 );
buf ( n2113 , 1'b0 );
buf ( n2114 , n30345 );
buf ( n2115 , n29066 );
buf ( n2116 , 1'b0 );
buf ( n2117 , 1'b0 );
buf ( n2118 , n30347 );
buf ( n2119 , n14405 );
buf ( n2120 , 1'b0 );
buf ( n2121 , 1'b0 );
buf ( n2122 , n30345 );
buf ( n2123 , n14633 );
buf ( n2124 , 1'b0 );
buf ( n2125 , 1'b0 );
buf ( n2126 , n30345 );
buf ( n2127 , n14639 );
buf ( n2128 , 1'b0 );
buf ( n2129 , 1'b0 );
buf ( n2130 , n30376 );
buf ( n2131 , n14645 );
buf ( n2132 , 1'b0 );
buf ( n2133 , 1'b0 );
buf ( n2134 , n30345 );
buf ( n2135 , n14408 );
buf ( n2136 , 1'b0 );
buf ( n2137 , 1'b0 );
buf ( n2138 , n30345 );
buf ( n2139 , n14650 );
buf ( n2140 , 1'b0 );
buf ( n2141 , 1'b0 );
buf ( n2142 , n30347 );
buf ( n2143 , n14654 );
buf ( n2144 , 1'b0 );
buf ( n2145 , 1'b0 );
buf ( n2146 , n30358 );
buf ( n2147 , n14658 );
buf ( n2148 , 1'b0 );
buf ( n2149 , 1'b0 );
buf ( n2150 , n30376 );
buf ( n2151 , n14662 );
buf ( n2152 , 1'b0 );
buf ( n2153 , 1'b0 );
buf ( n2154 , n30372 );
buf ( n2155 , n14418 );
buf ( n2156 , 1'b0 );
buf ( n2157 , 1'b0 );
buf ( n2158 , n30358 );
buf ( n2159 , n14411 );
buf ( n2160 , 1'b0 );
buf ( n2161 , 1'b0 );
buf ( n2162 , n30376 );
buf ( n2163 , n14414 );
buf ( n2164 , 1'b0 );
buf ( n2165 , 1'b0 );
buf ( n2166 , n30375 );
buf ( n2167 , n14668 );
buf ( n2168 , 1'b0 );
buf ( n2169 , 1'b0 );
buf ( n2170 , n30355 );
buf ( n2171 , n14672 );
buf ( n2172 , 1'b0 );
buf ( n2173 , 1'b0 );
buf ( n2174 , n30358 );
buf ( n2175 , n14384 );
buf ( n2176 , 1'b0 );
buf ( n2177 , 1'b0 );
buf ( n2178 , n30375 );
buf ( n2179 , n14676 );
buf ( n2180 , 1'b0 );
buf ( n2181 , 1'b0 );
buf ( n2182 , n30347 );
buf ( n2183 , n14932 );
buf ( n2184 , 1'b0 );
buf ( n2185 , 1'b0 );
buf ( n2186 , n30376 );
buf ( n2187 , n26537 );
buf ( n2188 , 1'b0 );
buf ( n2189 , 1'b0 );
buf ( n2190 , n30358 );
buf ( n2191 , n14150 );
buf ( n2192 , 1'b0 );
buf ( n2193 , 1'b0 );
buf ( n2194 , n30347 );
buf ( n2195 , n16518 );
buf ( n2196 , 1'b0 );
buf ( n2197 , 1'b0 );
buf ( n2198 , n30352 );
buf ( n2199 , n14427 );
buf ( n2200 , 1'b0 );
buf ( n2201 , 1'b0 );
buf ( n2202 , n30358 );
buf ( n2203 , n14837 );
buf ( n2204 , 1'b0 );
buf ( n2205 , 1'b0 );
buf ( n2206 , n30374 );
buf ( n2207 , n14687 );
buf ( n2208 , 1'b0 );
buf ( n2209 , 1'b0 );
buf ( n2210 , n30347 );
buf ( n2211 , n14444 );
buf ( n2212 , 1'b0 );
buf ( n2213 , 1'b0 );
buf ( n2214 , n30347 );
buf ( n2215 , n14853 );
buf ( n2216 , 1'b0 );
buf ( n2217 , 1'b0 );
buf ( n2218 , n30355 );
buf ( n2219 , n28701 );
buf ( n2220 , 1'b0 );
buf ( n2221 , 1'b0 );
buf ( n2222 , n30355 );
buf ( n2223 , n17255 );
buf ( n2224 , 1'b0 );
buf ( n2225 , 1'b0 );
buf ( n2226 , n30352 );
buf ( n2227 , n18014 );
buf ( n2228 , 1'b0 );
buf ( n2229 , 1'b0 );
buf ( n2230 , n30345 );
buf ( n2231 , n191 );
buf ( n2232 , 1'b0 );
buf ( n2233 , 1'b0 );
buf ( n2234 , n30351 );
buf ( n2235 , n27723 );
buf ( n2236 , 1'b0 );
buf ( n2237 , 1'b0 );
buf ( n2238 , n30352 );
buf ( n2239 , n14704 );
buf ( n2240 , 1'b0 );
buf ( n2241 , 1'b0 );
buf ( n2242 , n30358 );
buf ( n2243 , n28907 );
buf ( n2244 , 1'b0 );
buf ( n2245 , 1'b0 );
buf ( n2246 , n30345 );
buf ( n2247 , n27989 );
buf ( n2248 , 1'b0 );
buf ( n2249 , 1'b0 );
buf ( n2250 , n30352 );
buf ( n2251 , n30336 );
buf ( n2252 , 1'b0 );
buf ( n2253 , 1'b0 );
buf ( n2254 , n30358 );
buf ( n2255 , n21793 );
buf ( n2256 , 1'b0 );
buf ( n2257 , 1'b0 );
buf ( n2258 , n30353 );
buf ( n2259 , n29688 );
buf ( n2260 , 1'b0 );
buf ( n2261 , 1'b0 );
buf ( n2262 , n30352 );
buf ( n2263 , n28012 );
buf ( n2264 , 1'b0 );
buf ( n2265 , 1'b0 );
buf ( n2266 , n30355 );
buf ( n2267 , n15562 );
buf ( n2268 , 1'b0 );
buf ( n2269 , 1'b0 );
buf ( n2270 , n30347 );
buf ( n2271 , n29886 );
buf ( n2272 , 1'b0 );
buf ( n2273 , 1'b0 );
buf ( n2274 , n30345 );
buf ( n2275 , n14016 );
buf ( n2276 , 1'b0 );
buf ( n2277 , 1'b0 );
buf ( n2278 , n30376 );
buf ( n2279 , n14168 );
buf ( n2280 , 1'b0 );
buf ( n2281 , 1'b0 );
buf ( n2282 , n30345 );
buf ( n2283 , n14029 );
buf ( n2284 , 1'b0 );
buf ( n2285 , 1'b0 );
buf ( n2286 , n1 );
buf ( n2287 , n28696 );
buf ( n2288 , 1'b0 );
buf ( n2289 , 1'b0 );
buf ( n2290 , n30355 );
buf ( n2291 , n13834 );
buf ( n2292 , 1'b0 );
buf ( n2293 , 1'b0 );
buf ( n2294 , n30376 );
buf ( n2295 , n14044 );
buf ( n2296 , 1'b0 );
buf ( n2297 , 1'b0 );
buf ( n2298 , n30358 );
buf ( n2299 , n14058 );
buf ( n2300 , 1'b0 );
buf ( n2301 , 1'b0 );
buf ( n2302 , n30355 );
buf ( n2303 , n13860 );
buf ( n2304 , 1'b0 );
buf ( n2305 , 1'b0 );
buf ( n2306 , n30372 );
buf ( n2307 , n14140 );
buf ( n2308 , 1'b0 );
buf ( n2309 , 1'b0 );
buf ( n2310 , n30358 );
buf ( n2311 , n14072 );
buf ( n2312 , 1'b0 );
buf ( n2313 , 1'b0 );
buf ( n2314 , n30376 );
buf ( n2315 , n14087 );
buf ( n2316 , 1'b0 );
buf ( n2317 , 1'b0 );
buf ( n2318 , n30353 );
buf ( n2319 , n13878 );
buf ( n2320 , 1'b0 );
buf ( n2321 , 1'b0 );
buf ( n2322 , n30356 );
buf ( n2323 , n13910 );
buf ( n2324 , 1'b0 );
buf ( n2325 , 1'b0 );
buf ( n2326 , n30347 );
buf ( n2327 , n13964 );
buf ( n2328 , 1'b0 );
buf ( n2329 , 1'b0 );
buf ( n2330 , n30355 );
buf ( n2331 , n13705 );
buf ( n2332 , 1'b0 );
buf ( n2333 , 1'b0 );
buf ( n2334 , n1 );
buf ( n2335 , n28685 );
buf ( n2336 , 1'b0 );
buf ( n2337 , 1'b0 );
buf ( n2338 , n1 );
buf ( n2339 , n28674 );
buf ( n2340 , 1'b0 );
buf ( n2341 , 1'b0 );
buf ( n2342 , n30378 );
buf ( n2343 , n14534 );
buf ( n2344 , 1'b0 );
buf ( n2345 , 1'b0 );
buf ( n2346 , n1 );
buf ( n2347 , n28663 );
buf ( n2348 , 1'b0 );
buf ( n2349 , 1'b0 );
buf ( n2350 , n30351 );
buf ( n2351 , n16531 );
buf ( n2352 , 1'b0 );
buf ( n2353 , 1'b0 );
buf ( n2354 , n30376 );
buf ( n2355 , n16547 );
buf ( n2356 , 1'b0 );
buf ( n2357 , 1'b0 );
buf ( n2358 , n30355 );
buf ( n2359 , n13745 );
buf ( n2360 , 1'b0 );
buf ( n2361 , 1'b0 );
buf ( n2362 , n30353 );
buf ( n2363 , n13410 );
buf ( n2364 , 1'b0 );
buf ( n2365 , 1'b0 );
buf ( n2366 , n30376 );
buf ( n2367 , n16125 );
buf ( n2368 , 1'b0 );
buf ( n2369 , 1'b0 );
buf ( n2370 , n30351 );
buf ( n2371 , n19406 );
buf ( n2372 , 1'b0 );
buf ( n2373 , 1'b0 );
buf ( n2374 , n30374 );
buf ( n2375 , n20340 );
buf ( n2376 , 1'b0 );
buf ( n2377 , 1'b0 );
buf ( n2378 , n30345 );
buf ( n2379 , n16563 );
buf ( n2380 , 1'b0 );
buf ( n2381 , 1'b0 );
buf ( n2382 , n30351 );
buf ( n2383 , n20340 );
buf ( n2384 , 1'b0 );
buf ( n2385 , 1'b0 );
buf ( n2386 , n30378 );
buf ( n2387 , n20130 );
buf ( n2388 , 1'b0 );
buf ( n2389 , 1'b0 );
buf ( n2390 , n30345 );
buf ( n2391 , n14104 );
buf ( n2392 , 1'b0 );
buf ( n2393 , 1'b0 );
buf ( n2394 , n30378 );
buf ( n2395 , n14109 );
buf ( n2396 , 1'b0 );
buf ( n2397 , 1'b0 );
buf ( n2398 , n30374 );
buf ( n2399 , n14092 );
buf ( n2400 , 1'b0 );
buf ( n2401 , 1'b0 );
buf ( n2402 , n30345 );
buf ( n2403 , n13943 );
buf ( n2404 , 1'b0 );
buf ( n2405 , 1'b0 );
buf ( n2406 , n30355 );
buf ( n2407 , n14099 );
buf ( n2408 , 1'b0 );
buf ( n2409 , 1'b0 );
buf ( n2410 , n30353 );
buf ( n2411 , n13767 );
buf ( n2412 , 1'b0 );
buf ( n2413 , 1'b0 );
buf ( n2414 , n30355 );
buf ( n2415 , n13778 );
buf ( n2416 , 1'b0 );
buf ( n2417 , 1'b0 );
buf ( n2418 , n30352 );
buf ( n2419 , n13892 );
buf ( n2420 , 1'b0 );
buf ( n2421 , 1'b0 );
buf ( n2422 , n30355 );
buf ( n2423 , n13793 );
buf ( n2424 , 1'b0 );
buf ( n2425 , 1'b0 );
buf ( n2426 , n30374 );
buf ( n2427 , n13803 );
buf ( n2428 , 1'b0 );
buf ( n2429 , 1'b0 );
buf ( n2430 , n30345 );
buf ( n2431 , n16469 );
buf ( n2432 , 1'b0 );
buf ( n2433 , 1'b0 );
buf ( n2434 , n30372 );
buf ( n2435 , n16600 );
buf ( n2436 , 1'b0 );
buf ( n2437 , 1'b0 );
buf ( n2438 , n30376 );
buf ( n2439 , n16581 );
buf ( n2440 , 1'b0 );
buf ( n2441 , 1'b0 );
buf ( n2442 , n30378 );
buf ( n2443 , n16588 );
buf ( n2444 , 1'b0 );
buf ( n2445 , 1'b0 );
buf ( n2446 , n30345 );
buf ( n2447 , n16593 );
buf ( n2448 , 1'b0 );
buf ( n2449 , 1'b0 );
buf ( n2450 , n30374 );
buf ( n2451 , n14784 );
buf ( n2452 , 1'b0 );
buf ( n2453 , 1'b0 );
buf ( n2454 , n30372 );
buf ( n2455 , n29993 );
buf ( n2456 , 1'b0 );
buf ( n2457 , 1'b0 );
buf ( n2458 , n30345 );
buf ( n2459 , n29903 );
buf ( n2460 , 1'b0 );
buf ( n2461 , 1'b0 );
buf ( n2462 , n30374 );
buf ( n2463 , n29990 );
buf ( n2464 , 1'b0 );
buf ( n2465 , 1'b0 );
buf ( n2466 , n30356 );
buf ( n2467 , n13813 );
buf ( n2468 , 1'b0 );
buf ( n2469 , 1'b0 );
buf ( n2470 , n30378 );
buf ( n2471 , n29981 );
buf ( n2472 , 1'b0 );
buf ( n2473 , 1'b0 );
buf ( n2474 , n30345 );
buf ( n2475 , n13825 );
buf ( n2476 , 1'b0 );
buf ( n2477 , 1'b0 );
buf ( n2478 , n30353 );
buf ( n2479 , n14175 );
buf ( n2480 , 1'b0 );
buf ( n2481 , 1'b0 );
buf ( n2482 , n30355 );
buf ( n2483 , n13578 );
buf ( n2484 , 1'b0 );
buf ( n2485 , 1'b0 );
buf ( n2486 , n30343 );
buf ( n2487 , n14126 );
buf ( n2488 , 1'b0 );
buf ( n2489 , 1'b0 );
buf ( n2490 , n30376 );
buf ( n2491 , n14535 );
buf ( n2492 , 1'b0 );
buf ( n2493 , 1'b0 );
buf ( n2494 , n30345 );
buf ( n2495 , n30168 );
buf ( n2496 , 1'b0 );
buf ( n2497 , 1'b0 );
buf ( n2498 , n30374 );
buf ( n2499 , n20631 );
buf ( n2500 , 1'b0 );
buf ( n2501 , 1'b0 );
buf ( n2502 , n30378 );
buf ( n2503 , n14536 );
buf ( n2504 , 1'b0 );
buf ( n2505 , 1'b0 );
buf ( n2506 , n30376 );
buf ( n2507 , n14537 );
buf ( n2508 , 1'b0 );
buf ( n2509 , 1'b0 );
buf ( n2510 , n30355 );
buf ( n2511 , n29976 );
buf ( n2512 , 1'b0 );
buf ( n2513 , 1'b0 );
buf ( n2514 , n30356 );
buf ( n2515 , n29967 );
buf ( n2516 , 1'b0 );
buf ( n2517 , 1'b0 );
buf ( n2518 , n30355 );
buf ( n2519 , n29970 );
buf ( n2520 , 1'b0 );
buf ( n2521 , 1'b0 );
buf ( n2522 , n30376 );
buf ( n2523 , n29973 );
buf ( n2524 , 1'b0 );
buf ( n2525 , 1'b0 );
buf ( n2526 , n30378 );
buf ( n2527 , n13898 );
buf ( n2528 , 1'b0 );
buf ( n2529 , 1'b0 );
buf ( n2530 , n30353 );
buf ( n2531 , n13867 );
buf ( n2532 , 1'b0 );
buf ( n2533 , 1'b0 );
buf ( n2534 , n30376 );
buf ( n2535 , n13950 );
buf ( n2536 , 1'b0 );
buf ( n2537 , 1'b0 );
buf ( n2538 , n30374 );
buf ( n2539 , n13703 );
buf ( n2540 , 1'b0 );
buf ( n2541 , 1'b0 );
buf ( n2542 , n1 );
buf ( n2543 , n29907 );
buf ( n2544 , 1'b0 );
buf ( n2545 , 1'b0 );
buf ( n2546 , n1 );
buf ( n2547 , n19480 );
buf ( n2548 , 1'b0 );
buf ( n2549 , 1'b0 );
buf ( n2550 , n30353 );
buf ( n2551 , n15570 );
buf ( n2552 , 1'b0 );
buf ( n2553 , 1'b0 );
buf ( n2554 , n30356 );
buf ( n2555 , n14940 );
buf ( n2556 , 1'b0 );
buf ( n2557 , 1'b0 );
buf ( n2558 , n30355 );
buf ( n2559 , n15576 );
buf ( n2560 , 1'b0 );
buf ( n2561 , 1'b0 );
buf ( n2562 , n30345 );
buf ( n2563 , n30329 );
buf ( n2564 , 1'b0 );
buf ( n2565 , 1'b0 );
buf ( n2566 , n1 );
buf ( n2567 , n19553 );
buf ( n2568 , 1'b0 );
buf ( n2569 , 1'b0 );
buf ( n2570 , n1 );
buf ( n2571 , n19625 );
buf ( n2572 , 1'b0 );
buf ( n2573 , 1'b0 );
buf ( n2574 , n30371 );
buf ( n2575 , n30323 );
buf ( n2576 , 1'b0 );
buf ( n2577 , 1'b0 );
buf ( n2578 , n30355 );
buf ( n2579 , n30216 );
buf ( n2580 , 1'b0 );
buf ( n2581 , 1'b0 );
buf ( n2582 , n30356 );
buf ( n2583 , n30073 );
buf ( n2584 , 1'b0 );
buf ( n2585 , 1'b0 );
buf ( n2586 , n30374 );
buf ( n2587 , n30220 );
buf ( n2588 , 1'b0 );
buf ( n2589 , 1'b0 );
buf ( n2590 , n30355 );
buf ( n2591 , n13773 );
buf ( n2592 , 1'b0 );
buf ( n2593 , 1'b0 );
buf ( n2594 , n30356 );
buf ( n2595 , n13788 );
buf ( n2596 , 1'b0 );
buf ( n2597 , 1'b0 );
buf ( n2598 , n30374 );
buf ( n2599 , n14615 );
buf ( n2600 , 1'b0 );
buf ( n2601 , 1'b0 );
buf ( n2602 , n30353 );
buf ( n2603 , n13799 );
buf ( n2604 , 1'b0 );
buf ( n2605 , 1'b0 );
buf ( n2606 , n30374 );
buf ( n2607 , n27383 );
buf ( n2608 , 1'b0 );
buf ( n2609 , 1'b0 );
buf ( n2610 , n30353 );
buf ( n2611 , n29422 );
buf ( n2612 , 1'b0 );
buf ( n2613 , 1'b0 );
buf ( n2614 , n30374 );
buf ( n2615 , n30224 );
buf ( n2616 , 1'b0 );
buf ( n2617 , 1'b0 );
buf ( n2618 , n30352 );
buf ( n2619 , n30160 );
buf ( n2620 , 1'b0 );
buf ( n2621 , 1'b0 );
buf ( n2622 , n30343 );
buf ( n2623 , n30228 );
buf ( n2624 , 1'b0 );
buf ( n2625 , 1'b0 );
buf ( n2626 , n30374 );
buf ( n2627 , n30232 );
buf ( n2628 , 1'b0 );
buf ( n2629 , 1'b0 );
buf ( n2630 , n30371 );
buf ( n2631 , n30248 );
buf ( n2632 , 1'b0 );
buf ( n2633 , 1'b0 );
buf ( n2634 , n30353 );
buf ( n2635 , n30176 );
buf ( n2636 , 1'b0 );
buf ( n2637 , 1'b0 );
buf ( n2638 , n30374 );
buf ( n2639 , n30319 );
buf ( n2640 , 1'b0 );
buf ( n2641 , 1'b0 );
buf ( n2642 , n30343 );
buf ( n2643 , n30236 );
buf ( n2644 , 1'b0 );
buf ( n2645 , 1'b0 );
buf ( n2646 , n30374 );
buf ( n2647 , n30315 );
buf ( n2648 , 1'b0 );
buf ( n2649 , 1'b0 );
buf ( n2650 , n30355 );
buf ( n2651 , n30045 );
buf ( n2652 , 1'b0 );
buf ( n2653 , 1'b0 );
buf ( n2654 , n30343 );
buf ( n2655 , n30180 );
buf ( n2656 , 1'b0 );
buf ( n2657 , 1'b0 );
buf ( n2658 , n30351 );
buf ( n2659 , n30164 );
buf ( n2660 , 1'b0 );
buf ( n2661 , 1'b0 );
buf ( n2662 , n30345 );
buf ( n2663 , n30311 );
buf ( n2664 , 1'b0 );
buf ( n2665 , 1'b0 );
buf ( n2666 , n30352 );
buf ( n2667 , n30152 );
buf ( n2668 , 1'b0 );
buf ( n2669 , 1'b0 );
buf ( n2670 , n30371 );
buf ( n2671 , n30140 );
buf ( n2672 , 1'b0 );
buf ( n2673 , 1'b0 );
buf ( n2674 , n30355 );
buf ( n2675 , n30061 );
buf ( n2676 , 1'b0 );
buf ( n2677 , 1'b0 );
buf ( n2678 , n30374 );
buf ( n2679 , n30307 );
buf ( n2680 , 1'b0 );
buf ( n2681 , 1'b0 );
buf ( n2682 , n30376 );
buf ( n2683 , n30128 );
buf ( n2684 , 1'b0 );
buf ( n2685 , 1'b0 );
buf ( n2686 , n30358 );
buf ( n2687 , n30298 );
buf ( n2688 , 1'b0 );
buf ( n2689 , 1'b0 );
buf ( n2690 , n30356 );
buf ( n2691 , n30290 );
buf ( n2692 , 1'b0 );
buf ( n2693 , 1'b0 );
buf ( n2694 , n30358 );
buf ( n2695 , n30294 );
buf ( n2696 , 1'b0 );
buf ( n2697 , 1'b0 );
buf ( n2698 , n30343 );
buf ( n2699 , n30120 );
buf ( n2700 , 1'b0 );
buf ( n2701 , 1'b0 );
buf ( n2702 , n30355 );
buf ( n2703 , n30204 );
buf ( n2704 , 1'b0 );
buf ( n2705 , 1'b0 );
buf ( n2706 , n30355 );
buf ( n2707 , n30132 );
buf ( n2708 , 1'b0 );
buf ( n2709 , 1'b0 );
buf ( n2710 , n30356 );
buf ( n2711 , n30057 );
buf ( n2712 , 1'b0 );
buf ( n2713 , 1'b0 );
buf ( n2714 , n30358 );
buf ( n2715 , n30270 );
buf ( n2716 , 1'b0 );
buf ( n2717 , 1'b0 );
buf ( n2718 , n30355 );
buf ( n2719 , n30274 );
buf ( n2720 , 1'b0 );
buf ( n2721 , 1'b0 );
buf ( n2722 , n30371 );
buf ( n2723 , n30112 );
buf ( n2724 , 1'b0 );
buf ( n2725 , 1'b0 );
buf ( n2726 , n30355 );
buf ( n2727 , n30282 );
buf ( n2728 , 1'b0 );
buf ( n2729 , 1'b0 );
buf ( n2730 , n30374 );
buf ( n2731 , n16613 );
buf ( n2732 , 1'b0 );
buf ( n2733 , 1'b0 );
buf ( n2734 , n1 );
buf ( n2735 , n19699 );
buf ( n2736 , 1'b0 );
buf ( n2737 , 1'b0 );
buf ( n2738 , n30343 );
buf ( n2739 , n28724 );
buf ( n2740 , 1'b0 );
buf ( n2741 , 1'b0 );
buf ( n2742 , n30371 );
buf ( n2743 , n29863 );
buf ( n2744 , 1'b0 );
buf ( n2745 , 1'b0 );
buf ( n2746 , n30356 );
buf ( n2747 , n13762 );
buf ( n2748 , 1'b0 );
buf ( n2749 , 1'b0 );
buf ( n2750 , n30356 );
buf ( n2751 , n13808 );
buf ( n2752 , 1'b0 );
buf ( n2753 , 1'b0 );
buf ( n2754 , n30371 );
buf ( n2755 , n13819 );
buf ( n2756 , 1'b0 );
buf ( n2757 , 1'b0 );
buf ( n2758 , n30356 );
buf ( n2759 , n14744 );
buf ( n2760 , 1'b0 );
buf ( n2761 , 1'b0 );
buf ( n2762 , n30356 );
buf ( n2763 , n14743 );
buf ( n2764 , 1'b0 );
buf ( n2765 , 1'b0 );
buf ( n2766 , n30371 );
buf ( n2767 , n14745 );
buf ( n2768 , 1'b0 );
buf ( n2769 , 1'b0 );
buf ( n2770 , n30374 );
buf ( n2771 , n26542 );
buf ( n2772 , 1'b0 );
buf ( n2773 , 1'b0 );
buf ( n2774 , n30343 );
buf ( n2775 , n30368 );
buf ( n2776 , 1'b0 );
buf ( n2777 , 1'b0 );
buf ( n2778 , n30343 );
buf ( n2779 , n28921 );
buf ( n2780 , 1'b0 );
buf ( n2781 , 1'b0 );
buf ( n2782 , n30371 );
buf ( n2783 , n30262 );
buf ( n2784 , 1'b0 );
buf ( n2785 , 1'b0 );
buf ( n2786 , n30358 );
buf ( n2787 , n28030 );
buf ( n2788 , 1'b0 );
buf ( n2789 , 1'b0 );
buf ( n2790 , n30374 );
buf ( n2791 , n27734 );
buf ( n2792 , 1'b0 );
buf ( n2793 , 1'b0 );
buf ( n2794 , n30371 );
buf ( n2795 , n27740 );
buf ( n2796 , 1'b0 );
buf ( n2797 , 1'b0 );
buf ( n2798 , n30343 );
buf ( n2799 , n14765 );
buf ( n2800 , 1'b0 );
buf ( n2801 , 1'b0 );
buf ( n2802 , n30342 );
buf ( n2803 , n28045 );
buf ( n2804 , 1'b0 );
buf ( n2805 , 1'b0 );
buf ( n2806 , n30356 );
buf ( n2807 , n28059 );
buf ( n2808 , 1'b0 );
buf ( n2809 , 1'b0 );
buf ( n2810 , n30371 );
buf ( n2811 , n28072 );
buf ( n2812 , 1'b0 );
buf ( n2813 , 1'b0 );
buf ( n2814 , n30371 );
buf ( n2815 , n28085 );
buf ( n2816 , 1'b0 );
buf ( n2817 , 1'b0 );
buf ( n2818 , n30353 );
buf ( n2819 , n28098 );
buf ( n2820 , 1'b0 );
buf ( n2821 , 1'b0 );
buf ( n2822 , n30351 );
buf ( n2823 , n28115 );
buf ( n2824 , 1'b0 );
buf ( n2825 , 1'b0 );
buf ( n2826 , n30353 );
buf ( n2827 , n28129 );
buf ( n2828 , 1'b0 );
buf ( n2829 , 1'b0 );
buf ( n2830 , n30343 );
buf ( n2831 , n28501 );
buf ( n2832 , 1'b0 );
buf ( n2833 , 1'b0 );
buf ( n2834 , n30356 );
buf ( n2835 , n28467 );
buf ( n2836 , 1'b0 );
buf ( n2837 , 1'b0 );
buf ( n2838 , n30358 );
buf ( n2839 , n28479 );
buf ( n2840 , 1'b0 );
buf ( n2841 , 1'b0 );
buf ( n2842 , n30342 );
buf ( n2843 , n28455 );
buf ( n2844 , 1'b0 );
buf ( n2845 , 1'b0 );
buf ( n2846 , n30343 );
buf ( n2847 , n28443 );
buf ( n2848 , 1'b0 );
buf ( n2849 , 1'b0 );
buf ( n2850 , n30356 );
buf ( n2851 , n28431 );
buf ( n2852 , 1'b0 );
buf ( n2853 , 1'b0 );
buf ( n2854 , n30342 );
buf ( n2855 , n28419 );
buf ( n2856 , 1'b0 );
buf ( n2857 , 1'b0 );
buf ( n2858 , n30358 );
buf ( n2859 , n16767 );
buf ( n2860 , 1'b0 );
buf ( n2861 , 1'b0 );
buf ( n2862 , n30342 );
buf ( n2863 , n16620 );
buf ( n2864 , 1'b0 );
buf ( n2865 , 1'b0 );
buf ( n2866 , n30343 );
buf ( n2867 , n28404 );
buf ( n2868 , 1'b0 );
buf ( n2869 , 1'b0 );
buf ( n2870 , n30346 );
buf ( n2871 , n14742 );
buf ( n2872 , 1'b0 );
buf ( n2873 , 1'b0 );
buf ( n2874 , n30356 );
buf ( n2875 , n28143 );
buf ( n2876 , 1'b0 );
buf ( n2877 , 1'b0 );
buf ( n2878 , n30371 );
buf ( n2879 , n28156 );
buf ( n2880 , 1'b0 );
buf ( n2881 , 1'b0 );
buf ( n2882 , n30351 );
buf ( n2883 , n28166 );
buf ( n2884 , 1'b0 );
buf ( n2885 , 1'b0 );
buf ( n2886 , n1 );
buf ( n2887 , n396 );
buf ( n2888 , 1'b0 );
buf ( n2889 , 1'b0 );
buf ( n2890 , n30353 );
buf ( n2891 , n30015 );
buf ( n2892 , 1'b0 );
buf ( n2893 , 1'b0 );
buf ( n2894 , n30342 );
buf ( n2895 , n25287 );
buf ( n2896 , 1'b0 );
buf ( n2897 , 1'b0 );
buf ( n2898 , n30371 );
buf ( n2899 , n28179 );
buf ( n2900 , 1'b0 );
buf ( n2901 , 1'b0 );
buf ( n2902 , n30353 );
buf ( n2903 , n28192 );
buf ( n2904 , 1'b0 );
buf ( n2905 , 1'b0 );
buf ( n2906 , n30375 );
buf ( n2907 , n28205 );
buf ( n2908 , 1'b0 );
buf ( n2909 , 1'b0 );
buf ( n2910 , n30352 );
buf ( n2911 , n28218 );
buf ( n2912 , 1'b0 );
buf ( n2913 , 1'b0 );
buf ( n2914 , n30353 );
buf ( n2915 , n28738 );
buf ( n2916 , 1'b0 );
buf ( n2917 , 1'b0 );
buf ( n2918 , n30353 );
buf ( n2919 , n28751 );
buf ( n2920 , 1'b0 );
buf ( n2921 , 1'b0 );
buf ( n2922 , n30356 );
buf ( n2923 , n28764 );
buf ( n2924 , 1'b0 );
buf ( n2925 , 1'b0 );
buf ( n2926 , n30353 );
buf ( n2927 , n28777 );
buf ( n2928 , 1'b0 );
buf ( n2929 , 1'b0 );
buf ( n2930 , n30351 );
buf ( n2931 , n28843 );
buf ( n2932 , 1'b0 );
buf ( n2933 , 1'b0 );
buf ( n2934 , n30375 );
buf ( n2935 , n28790 );
buf ( n2936 , 1'b0 );
buf ( n2937 , 1'b0 );
buf ( n2938 , n30376 );
buf ( n2939 , n28803 );
buf ( n2940 , 1'b0 );
buf ( n2941 , 1'b0 );
buf ( n2942 , n30352 );
buf ( n2943 , n20653 );
buf ( n2944 , 1'b0 );
buf ( n2945 , 1'b0 );
buf ( n2946 , n30375 );
buf ( n2947 , n29173 );
buf ( n2948 , 1'b0 );
buf ( n2949 , 1'b0 );
buf ( n2950 , n30346 );
buf ( n2951 , n29078 );
buf ( n2952 , 1'b0 );
buf ( n2953 , 1'b0 );
buf ( n2954 , n30376 );
buf ( n2955 , n28522 );
buf ( n2956 , 1'b0 );
buf ( n2957 , 1'b0 );
buf ( n2958 , n30371 );
buf ( n2959 , n28389 );
buf ( n2960 , 1'b0 );
buf ( n2961 , 1'b0 );
buf ( n2962 , n30351 );
buf ( n2963 , n27389 );
buf ( n2964 , 1'b0 );
buf ( n2965 , 1'b0 );
buf ( n2966 , n30351 );
buf ( n2967 , n26552 );
buf ( n2968 , 1'b0 );
buf ( n2969 , 1'b0 );
buf ( n2970 , n30353 );
buf ( n2971 , n27400 );
buf ( n2972 , 1'b0 );
buf ( n2973 , 1'b0 );
buf ( n2974 , n30375 );
buf ( n2975 , n14614 );
buf ( n2976 , 1'b0 );
buf ( n2977 , 1'b0 );
buf ( n2978 , n30346 );
buf ( n2979 , n14947 );
buf ( n2980 , 1'b0 );
buf ( n2981 , 1'b0 );
buf ( n2982 , n30375 );
buf ( n2983 , n28231 );
buf ( n2984 , 1'b0 );
buf ( n2985 , 1'b0 );
buf ( n2986 , n30371 );
buf ( n2987 , n28816 );
buf ( n2988 , 1'b0 );
buf ( n2989 , 1'b0 );
buf ( n2990 , n30356 );
buf ( n2991 , n28244 );
buf ( n2992 , 1'b0 );
buf ( n2993 , 1'b0 );
buf ( n2994 , n30378 );
buf ( n2995 , n25348 );
buf ( n2996 , 1'b0 );
buf ( n2997 , 1'b0 );
buf ( n2998 , n30343 );
buf ( n2999 , n29789 );
buf ( n3000 , 1'b0 );
buf ( n3001 , 1'b0 );
buf ( n3002 , n30378 );
buf ( n3003 , n29784 );
buf ( n3004 , 1'b0 );
buf ( n3005 , 1'b0 );
buf ( n3006 , n30375 );
buf ( n3007 , n29736 );
buf ( n3008 , 1'b0 );
buf ( n3009 , 1'b0 );
buf ( n3010 , n30352 );
buf ( n3011 , n29779 );
buf ( n3012 , 1'b0 );
buf ( n3013 , 1'b0 );
buf ( n3014 , n30352 );
buf ( n3015 , n30020 );
buf ( n3016 , 1'b0 );
buf ( n3017 , 1'b0 );
buf ( n3018 , n30375 );
buf ( n3019 , n29741 );
buf ( n3020 , 1'b0 );
buf ( n3021 , 1'b0 );
buf ( n3022 , n1 );
buf ( n3023 , n30103 );
buf ( n3024 , 1'b0 );
buf ( n3025 , 1'b0 );
buf ( n3026 , n30375 );
buf ( n3027 , n29340 );
buf ( n3028 , 1'b0 );
buf ( n3029 , 1'b0 );
buf ( n3030 , n30356 );
buf ( n3031 , n28251 );
buf ( n3032 , 1'b0 );
buf ( n3033 , 1'b0 );
buf ( n3034 , n30346 );
buf ( n3035 , n27403 );
buf ( n3036 , 1'b0 );
buf ( n3037 , 1'b0 );
buf ( n3038 , n30375 );
buf ( n3039 , n20153 );
buf ( n3040 , 1'b0 );
buf ( n3041 , 1'b0 );
buf ( n3042 , n30342 );
buf ( n3043 , n29335 );
buf ( n3044 , 1'b0 );
buf ( n3045 , 1'b0 );
buf ( n3046 , n30346 );
buf ( n3047 , n15695 );
buf ( n3048 , 1'b0 );
buf ( n3049 , 1'b0 );
buf ( n3050 , n30351 );
buf ( n3051 , n29774 );
buf ( n3052 , 1'b0 );
buf ( n3053 , 1'b0 );
buf ( n3054 , n30345 );
buf ( n3055 , n25409 );
buf ( n3056 , 1'b0 );
buf ( n3057 , 1'b0 );
buf ( n3058 , n30372 );
buf ( n3059 , n25470 );
buf ( n3060 , 1'b0 );
buf ( n3061 , 1'b0 );
buf ( n3062 , n30353 );
buf ( n3063 , n25528 );
buf ( n3064 , 1'b0 );
buf ( n3065 , 1'b0 );
buf ( n3066 , n30375 );
buf ( n3067 , n16624 );
buf ( n3068 , 1'b0 );
buf ( n3069 , 1'b0 );
buf ( n3070 , n30371 );
buf ( n3071 , n29743 );
buf ( n3072 , 1'b0 );
buf ( n3073 , 1'b0 );
buf ( n3074 , n30353 );
buf ( n3075 , n29769 );
buf ( n3076 , 1'b0 );
buf ( n3077 , 1'b0 );
buf ( n3078 , n30371 );
buf ( n3079 , n29748 );
buf ( n3080 , 1'b0 );
buf ( n3081 , 1'b0 );
buf ( n3082 , n30352 );
buf ( n3083 , n29759 );
buf ( n3084 , 1'b0 );
buf ( n3085 , 1'b0 );
buf ( n3086 , n30352 );
buf ( n3087 , n29764 );
buf ( n3088 , 1'b0 );
buf ( n3089 , 1'b0 );
buf ( n3090 , n30356 );
buf ( n3091 , n29754 );
buf ( n3092 , 1'b0 );
buf ( n3093 , 1'b0 );
buf ( n3094 , n30345 );
buf ( n3095 , n29424 );
buf ( n3096 , 1'b0 );
buf ( n3097 , 1'b0 );
buf ( n3098 , n30346 );
buf ( n3099 , n29168 );
buf ( n3100 , 1'b0 );
buf ( n3101 , 1'b0 );
buf ( n3102 , n30356 );
buf ( n3103 , n16141 );
buf ( n3104 , 1'b0 );
buf ( n3105 , 1'b0 );
buf ( n3106 , n30371 );
buf ( n3107 , n16456 );
buf ( n3108 , 1'b0 );
buf ( n3109 , 1'b0 );
buf ( n3110 , n30371 );
buf ( n3111 , n16456 );
buf ( n3112 , 1'b0 );
buf ( n3113 , 1'b0 );
buf ( n3114 , n30358 );
buf ( n3115 , n16130 );
buf ( n3116 , 1'b0 );
buf ( n3117 , 1'b0 );
buf ( n3118 , n30371 );
buf ( n3119 , n15702 );
buf ( n3120 , 1'b0 );
buf ( n3121 , 1'b0 );
buf ( n3122 , n30353 );
buf ( n3123 , n14972 );
buf ( n3124 , 1'b0 );
buf ( n3125 , 1'b0 );
buf ( n3126 , n30371 );
buf ( n3127 , n18033 );
buf ( n3128 , 1'b0 );
buf ( n3129 , 1'b0 );
buf ( n3130 , n30342 );
buf ( n3131 , n16155 );
buf ( n3132 , 1'b0 );
buf ( n3133 , 1'b0 );
buf ( n3134 , n30352 );
buf ( n3135 , n16630 );
buf ( n3136 , 1'b0 );
buf ( n3137 , 1'b0 );
buf ( n3138 , n30371 );
buf ( n3139 , n28825 );
buf ( n3140 , 1'b0 );
buf ( n3141 , 1'b0 );
buf ( n3142 , n30346 );
buf ( n3143 , n30124 );
buf ( n3144 , 1'b0 );
buf ( n3145 , 1'b0 );
buf ( n3146 , n30346 );
buf ( n3147 , n16160 );
buf ( n3148 , 1'b0 );
buf ( n3149 , 1'b0 );
buf ( n3150 , n30353 );
buf ( n3151 , n16164 );
buf ( n3152 , 1'b0 );
buf ( n3153 , 1'b0 );
buf ( n3154 , n30346 );
buf ( n3155 , n16169 );
buf ( n3156 , 1'b0 );
buf ( n3157 , 1'b0 );
buf ( n3158 , n30371 );
buf ( n3159 , n16174 );
buf ( n3160 , 1'b0 );
buf ( n3161 , 1'b0 );
buf ( n3162 , n30353 );
buf ( n3163 , n16179 );
buf ( n3164 , 1'b0 );
buf ( n3165 , 1'b0 );
buf ( n3166 , n30346 );
buf ( n3167 , n16186 );
buf ( n3168 , 1'b0 );
buf ( n3169 , 1'b0 );
buf ( n3170 , n30342 );
buf ( n3171 , n16192 );
buf ( n3172 , 1'b0 );
buf ( n3173 , 1'b0 );
buf ( n3174 , n30342 );
buf ( n3175 , n16193 );
buf ( n3176 , 1'b0 );
buf ( n3177 , 1'b0 );
buf ( n3178 , n30346 );
buf ( n3179 , n16200 );
buf ( n3180 , 1'b0 );
buf ( n3181 , 1'b0 );
buf ( n3182 , n30378 );
buf ( n3183 , n16210 );
buf ( n3184 , 1'b0 );
buf ( n3185 , 1'b0 );
buf ( n3186 , n30345 );
buf ( n3187 , n16218 );
buf ( n3188 , 1'b0 );
buf ( n3189 , 1'b0 );
buf ( n3190 , n30346 );
buf ( n3191 , n16226 );
buf ( n3192 , 1'b0 );
buf ( n3193 , 1'b0 );
buf ( n3194 , n30346 );
buf ( n3195 , n30010 );
buf ( n3196 , 1'b0 );
buf ( n3197 , 1'b0 );
buf ( n3198 , n30342 );
buf ( n3199 , n16635 );
buf ( n3200 , 1'b0 );
buf ( n3201 , 1'b0 );
buf ( n3202 , n30371 );
buf ( n3203 , n16608 );
buf ( n3204 , 1'b0 );
buf ( n3205 , 1'b0 );
buf ( n3206 , n30342 );
buf ( n3207 , n16640 );
buf ( n3208 , 1'b0 );
buf ( n3209 , 1'b0 );
buf ( n3210 , n30343 );
buf ( n3211 , n16652 );
buf ( n3212 , 1'b0 );
buf ( n3213 , 1'b0 );
buf ( n3214 , n30343 );
buf ( n3215 , n16577 );
buf ( n3216 , 1'b0 );
buf ( n3217 , 1'b0 );
buf ( n3218 , n30343 );
buf ( n3219 , n16712 );
buf ( n3220 , 1'b0 );
buf ( n3221 , 1'b0 );
buf ( n3222 , n30351 );
buf ( n3223 , n16646 );
buf ( n3224 , 1'b0 );
buf ( n3225 , 1'b0 );
buf ( n3226 , n30342 );
buf ( n3227 , n16232 );
buf ( n3228 , 1'b0 );
buf ( n3229 , 1'b0 );
buf ( n3230 , n30358 );
buf ( n3231 , n16240 );
buf ( n3232 , 1'b0 );
buf ( n3233 , 1'b0 );
buf ( n3234 , n30351 );
buf ( n3235 , n20206 );
buf ( n3236 , 1'b0 );
buf ( n3237 , 1'b0 );
buf ( n3238 , n30343 );
buf ( n3239 , n30286 );
buf ( n3240 , 1'b0 );
buf ( n3241 , 1'b0 );
buf ( n3242 , n30342 );
buf ( n3243 , n21832 );
buf ( n3244 , 1'b0 );
buf ( n3245 , 1'b0 );
buf ( n3246 , n30346 );
buf ( n3247 , n21846 );
buf ( n3248 , 1'b0 );
buf ( n3249 , 1'b0 );
buf ( n3250 , n30358 );
buf ( n3251 , n21857 );
buf ( n3252 , 1'b0 );
buf ( n3253 , 1'b0 );
buf ( n3254 , n30342 );
buf ( n3255 , n21872 );
buf ( n3256 , 1'b0 );
buf ( n3257 , 1'b0 );
buf ( n3258 , n30351 );
buf ( n3259 , n21884 );
buf ( n3260 , 1'b0 );
buf ( n3261 , 1'b0 );
buf ( n3262 , n30352 );
buf ( n3263 , n21897 );
buf ( n3264 , 1'b0 );
buf ( n3265 , 1'b0 );
buf ( n3266 , n30351 );
buf ( n3267 , n21906 );
buf ( n3268 , 1'b0 );
buf ( n3269 , 1'b0 );
buf ( n3270 , n30352 );
buf ( n3271 , n25535 );
buf ( n3272 , 1'b0 );
buf ( n3273 , 1'b0 );
buf ( n3274 , n30346 );
buf ( n3275 , n21915 );
buf ( n3276 , 1'b0 );
buf ( n3277 , 1'b0 );
buf ( n3278 , n30351 );
buf ( n3279 , n21927 );
buf ( n3280 , 1'b0 );
buf ( n3281 , 1'b0 );
buf ( n3282 , n30342 );
buf ( n3283 , n21937 );
buf ( n3284 , 1'b0 );
buf ( n3285 , 1'b0 );
buf ( n3286 , n30346 );
buf ( n3287 , n25541 );
buf ( n3288 , 1'b0 );
buf ( n3289 , 1'b0 );
buf ( n3290 , n30342 );
buf ( n3291 , n25548 );
buf ( n3292 , 1'b0 );
buf ( n3293 , 1'b0 );
buf ( n3294 , n30351 );
buf ( n3295 , n21947 );
buf ( n3296 , 1'b0 );
buf ( n3297 , 1'b0 );
buf ( n3298 , n30346 );
buf ( n3299 , n25554 );
buf ( n3300 , 1'b0 );
buf ( n3301 , 1'b0 );
buf ( n3302 , n30342 );
buf ( n3303 , n23614 );
buf ( n3304 , 1'b0 );
buf ( n3305 , 1'b0 );
buf ( n3306 , n30343 );
buf ( n3307 , n23622 );
buf ( n3308 , 1'b0 );
buf ( n3309 , 1'b0 );
buf ( n3310 , n30342 );
buf ( n3311 , n23629 );
buf ( n3312 , 1'b0 );
buf ( n3313 , 1'b0 );
buf ( n3314 , n30342 );
buf ( n3315 , n25560 );
buf ( n3316 , 1'b0 );
buf ( n3317 , 1'b0 );
buf ( n3318 , n30346 );
buf ( n3319 , n23634 );
buf ( n3320 , 1'b0 );
buf ( n3321 , 1'b0 );
buf ( n3322 , n30346 );
buf ( n3323 , n29749 );
buf ( n3324 , 1'b0 );
buf ( n3325 , 1'b0 );
buf ( n3326 , n30342 );
buf ( n3327 , n30003 );
buf ( n3328 , 1'b0 );
buf ( n3329 , 1'b0 );
buf ( n3330 , n30346 );
buf ( n3331 , n17262 );
buf ( n3332 , 1'b0 );
buf ( n3333 , 1'b0 );
buf ( n3334 , n30346 );
buf ( n3335 , n23640 );
buf ( n3336 , 1'b0 );
buf ( n3337 , 1'b0 );
buf ( n3338 , n30352 );
buf ( n3339 , n25565 );
buf ( n3340 , 1'b0 );
buf ( n3341 , 1'b0 );
buf ( n3342 , n30378 );
buf ( n3343 , n23652 );
buf ( n3344 , 1'b0 );
buf ( n3345 , 1'b0 );
buf ( n3346 , n30346 );
buf ( n3347 , n21958 );
buf ( n3348 , 1'b0 );
buf ( n3349 , 1'b0 );
buf ( n3350 , n30343 );
buf ( n3351 , n21967 );
buf ( n3352 , 1'b0 );
buf ( n3353 , 1'b0 );
buf ( n3354 , n30378 );
buf ( n3355 , n21975 );
buf ( n3356 , 1'b0 );
buf ( n3357 , 1'b0 );
buf ( n3358 , n30378 );
buf ( n3359 , n21985 );
buf ( n3360 , 1'b0 );
buf ( n3361 , 1'b0 );
buf ( n3362 , n30346 );
buf ( n3363 , n21994 );
buf ( n3364 , 1'b0 );
buf ( n3365 , 1'b0 );
buf ( n3366 , n30343 );
buf ( n3367 , n22003 );
buf ( n3368 , 1'b0 );
buf ( n3369 , 1'b0 );
buf ( n3370 , n30352 );
buf ( n3371 , n22012 );
buf ( n3372 , 1'b0 );
buf ( n3373 , 1'b0 );
buf ( n3374 , n30351 );
buf ( n3375 , n22022 );
buf ( n3376 , 1'b0 );
buf ( n3377 , 1'b0 );
buf ( n3378 , n30346 );
buf ( n3379 , n23659 );
buf ( n3380 , 1'b0 );
buf ( n3381 , 1'b0 );
buf ( n3382 , n30352 );
buf ( n3383 , n22031 );
buf ( n3384 , 1'b0 );
buf ( n3385 , 1'b0 );
buf ( n3386 , n30352 );
buf ( n3387 , n22040 );
buf ( n3388 , 1'b0 );
buf ( n3389 , 1'b0 );
buf ( n3390 , n30352 );
buf ( n3391 , n22049 );
buf ( n3392 , 1'b0 );
buf ( n3393 , 1'b0 );
buf ( n3394 , n30343 );
buf ( n3395 , n22058 );
buf ( n3396 , 1'b0 );
buf ( n3397 , 1'b0 );
buf ( n3398 , n30378 );
buf ( n3399 , n22073 );
buf ( n3400 , 1'b0 );
buf ( n3401 , 1'b0 );
buf ( n3402 , n30378 );
buf ( n3403 , n22082 );
buf ( n3404 , 1'b0 );
buf ( n3405 , 1'b0 );
buf ( n3406 , n30346 );
buf ( n3407 , n15567 );
buf ( n3408 , 1'b0 );
buf ( n3409 , 1'b0 );
buf ( n3410 , n30342 );
buf ( n3411 , n16248 );
buf ( n3412 , 1'b0 );
buf ( n3413 , 1'b0 );
buf ( n3414 , n1 );
buf ( n3415 , n563 );
buf ( n3416 , 1'b0 );
buf ( n3417 , 1'b0 );
buf ( n3418 , n30346 );
buf ( n3419 , n16256 );
buf ( n3420 , 1'b0 );
buf ( n3421 , 1'b0 );
buf ( n3422 , n30342 );
buf ( n3423 , n22091 );
buf ( n3424 , 1'b0 );
buf ( n3425 , 1'b0 );
buf ( n3426 , n30342 );
buf ( n3427 , n23666 );
buf ( n3428 , 1'b0 );
buf ( n3429 , 1'b0 );
buf ( n3430 , n30346 );
buf ( n3431 , n15202 );
buf ( n3432 , 1'b0 );
buf ( n3433 , 1'b0 );
buf ( n3434 , n30342 );
buf ( n3435 , n16370 );
buf ( n3436 , 1'b0 );
buf ( n3437 , 1'b0 );
buf ( n3438 , n30346 );
buf ( n3439 , n23671 );
buf ( n3440 , 1'b0 );
buf ( n3441 , 1'b0 );
buf ( n3442 , n30352 );
buf ( n3443 , n22098 );
buf ( n3444 , 1'b0 );
buf ( n3445 , 1'b0 );
buf ( n3446 , n30351 );
buf ( n3447 , n22107 );
buf ( n3448 , 1'b0 );
buf ( n3449 , 1'b0 );
buf ( n3450 , n30351 );
buf ( n3451 , n22115 );
buf ( n3452 , 1'b0 );
buf ( n3453 , 1'b0 );
buf ( n3454 , n30342 );
buf ( n3455 , n22124 );
buf ( n3456 , 1'b0 );
buf ( n3457 , 1'b0 );
buf ( n3458 , n30342 );
buf ( n3459 , n22132 );
buf ( n3460 , 1'b0 );
buf ( n3461 , 1'b0 );
buf ( n3462 , n30343 );
buf ( n3463 , n23677 );
buf ( n3464 , 1'b0 );
buf ( n3465 , 1'b0 );
buf ( n3466 , n30358 );
buf ( n3467 , n22141 );
buf ( n3468 , 1'b0 );
buf ( n3469 , 1'b0 );
buf ( n3470 , n30342 );
buf ( n3471 , n22149 );
buf ( n3472 , 1'b0 );
buf ( n3473 , 1'b0 );
buf ( n3474 , n30342 );
buf ( n3475 , n23683 );
buf ( n3476 , 1'b0 );
buf ( n3477 , 1'b0 );
buf ( n3478 , n30371 );
buf ( n3479 , n22170 );
buf ( n3480 , 1'b0 );
buf ( n3481 , 1'b0 );
buf ( n3482 , n30346 );
buf ( n3483 , n22178 );
buf ( n3484 , 1'b0 );
buf ( n3485 , 1'b0 );
buf ( n3486 , n30346 );
buf ( n3487 , n22187 );
buf ( n3488 , 1'b0 );
buf ( n3489 , 1'b0 );
buf ( n3490 , n30346 );
buf ( n3491 , n22194 );
buf ( n3492 , 1'b0 );
buf ( n3493 , 1'b0 );
buf ( n3494 , n30342 );
buf ( n3495 , n23689 );
buf ( n3496 , 1'b0 );
buf ( n3497 , 1'b0 );
buf ( n3498 , n30346 );
buf ( n3499 , n22201 );
buf ( n3500 , 1'b0 );
buf ( n3501 , 1'b0 );
buf ( n3502 , n30353 );
buf ( n3503 , n23695 );
buf ( n3504 , 1'b0 );
buf ( n3505 , 1'b0 );
buf ( n3506 , n30346 );
buf ( n3507 , n23701 );
buf ( n3508 , 1'b0 );
buf ( n3509 , 1'b0 );
buf ( n3510 , n30346 );
buf ( n3511 , n23706 );
buf ( n3512 , 1'b0 );
buf ( n3513 , 1'b0 );
buf ( n3514 , n30352 );
buf ( n3515 , n15088 );
buf ( n3516 , 1'b0 );
buf ( n3517 , 1'b0 );
buf ( n3518 , n30342 );
buf ( n3519 , n16411 );
buf ( n3520 , 1'b0 );
buf ( n3521 , 1'b0 );
buf ( n3522 , n30371 );
buf ( n3523 , n15900 );
buf ( n3524 , 1'b0 );
buf ( n3525 , 1'b0 );
buf ( n3526 , n30358 );
buf ( n3527 , n17161 );
buf ( n3528 , 1'b0 );
buf ( n3529 , 1'b0 );
buf ( n3530 , n30371 );
buf ( n3531 , n17343 );
buf ( n3532 , 1'b0 );
buf ( n3533 , 1'b0 );
buf ( n3534 , n30356 );
buf ( n3535 , n18070 );
buf ( n3536 , 1'b0 );
buf ( n3537 , 1'b0 );
buf ( n3538 , n30371 );
buf ( n3539 , n20663 );
buf ( n3540 , 1'b0 );
buf ( n3541 , 1'b0 );
buf ( n3542 , n30375 );
buf ( n3543 , n18086 );
buf ( n3544 , 1'b0 );
buf ( n3545 , 1'b0 );
buf ( n3546 , n30372 );
buf ( n3547 , n18508 );
buf ( n3548 , 1'b0 );
buf ( n3549 , 1'b0 );
buf ( n3550 , n30345 );
buf ( n3551 , n18528 );
buf ( n3552 , 1'b0 );
buf ( n3553 , 1'b0 );
buf ( n3554 , n30342 );
buf ( n3555 , n23712 );
buf ( n3556 , 1'b0 );
buf ( n3557 , 1'b0 );
buf ( n3558 , n30375 );
buf ( n3559 , n25571 );
buf ( n3560 , 1'b0 );
buf ( n3561 , 1'b0 );
buf ( n3562 , n30356 );
buf ( n3563 , n23718 );
buf ( n3564 , 1'b0 );
buf ( n3565 , 1'b0 );
buf ( n3566 , n30375 );
buf ( n3567 , n23723 );
buf ( n3568 , 1'b0 );
buf ( n3569 , 1'b0 );
buf ( n3570 , n30375 );
buf ( n3571 , n25577 );
buf ( n3572 , 1'b0 );
buf ( n3573 , 1'b0 );
buf ( n3574 , n30378 );
buf ( n3575 , n23728 );
buf ( n3576 , 1'b0 );
buf ( n3577 , 1'b0 );
buf ( n3578 , n30378 );
buf ( n3579 , n25583 );
buf ( n3580 , 1'b0 );
buf ( n3581 , 1'b0 );
buf ( n3582 , n30356 );
buf ( n3583 , n23733 );
buf ( n3584 , 1'b0 );
buf ( n3585 , 1'b0 );
buf ( n3586 , n30346 );
buf ( n3587 , n23738 );
buf ( n3588 , 1'b0 );
buf ( n3589 , 1'b0 );
buf ( n3590 , n30375 );
buf ( n3591 , n23744 );
buf ( n3592 , 1'b0 );
buf ( n3593 , 1'b0 );
buf ( n3594 , n30351 );
buf ( n3595 , n23749 );
buf ( n3596 , 1'b0 );
buf ( n3597 , 1'b0 );
buf ( n3598 , n30351 );
buf ( n3599 , n23755 );
buf ( n3600 , 1'b0 );
buf ( n3601 , 1'b0 );
buf ( n3602 , n30352 );
buf ( n3603 , n23760 );
buf ( n3604 , 1'b0 );
buf ( n3605 , 1'b0 );
buf ( n3606 , n30376 );
buf ( n3607 , n23765 );
buf ( n3608 , 1'b0 );
buf ( n3609 , 1'b0 );
buf ( n3610 , n30351 );
buf ( n3611 , n23770 );
buf ( n3612 , 1'b0 );
buf ( n3613 , 1'b0 );
buf ( n3614 , n30353 );
buf ( n3615 , n23780 );
buf ( n3616 , 1'b0 );
buf ( n3617 , 1'b0 );
buf ( n3618 , n30353 );
buf ( n3619 , n23775 );
buf ( n3620 , 1'b0 );
buf ( n3621 , 1'b0 );
buf ( n3622 , n30352 );
buf ( n3623 , n22207 );
buf ( n3624 , 1'b0 );
buf ( n3625 , 1'b0 );
buf ( n3626 , n30353 );
buf ( n3627 , n23786 );
buf ( n3628 , 1'b0 );
buf ( n3629 , 1'b0 );
buf ( n3630 , n30371 );
buf ( n3631 , n27757 );
buf ( n3632 , 1'b0 );
buf ( n3633 , 1'b0 );
buf ( n3634 , n30371 );
buf ( n3635 , n23797 );
buf ( n3636 , 1'b0 );
buf ( n3637 , 1'b0 );
buf ( n3638 , n30356 );
buf ( n3639 , n27749 );
buf ( n3640 , 1'b0 );
buf ( n3641 , 1'b0 );
buf ( n3642 , n30343 );
buf ( n3643 , n27768 );
buf ( n3644 , 1'b0 );
buf ( n3645 , 1'b0 );
buf ( n3646 , n30342 );
buf ( n3647 , n25597 );
buf ( n3648 , 1'b0 );
buf ( n3649 , 1'b0 );
buf ( n3650 , n30356 );
buf ( n3651 , n22223 );
buf ( n3652 , 1'b0 );
buf ( n3653 , 1'b0 );
buf ( n3654 , n30343 );
buf ( n3655 , n22233 );
buf ( n3656 , 1'b0 );
buf ( n3657 , 1'b0 );
buf ( n3658 , n30358 );
buf ( n3659 , n22243 );
buf ( n3660 , 1'b0 );
buf ( n3661 , 1'b0 );
buf ( n3662 , n30356 );
buf ( n3663 , n22251 );
buf ( n3664 , 1'b0 );
buf ( n3665 , 1'b0 );
buf ( n3666 , n30371 );
buf ( n3667 , n23805 );
buf ( n3668 , 1'b0 );
buf ( n3669 , 1'b0 );
buf ( n3670 , n30356 );
buf ( n3671 , n22259 );
buf ( n3672 , 1'b0 );
buf ( n3673 , 1'b0 );
buf ( n3674 , n30343 );
buf ( n3675 , n22267 );
buf ( n3676 , 1'b0 );
buf ( n3677 , 1'b0 );
buf ( n3678 , n30371 );
buf ( n3679 , n22276 );
buf ( n3680 , 1'b0 );
buf ( n3681 , 1'b0 );
buf ( n3682 , n30371 );
buf ( n3683 , n22284 );
buf ( n3684 , 1'b0 );
buf ( n3685 , 1'b0 );
buf ( n3686 , n30343 );
buf ( n3687 , n22293 );
buf ( n3688 , 1'b0 );
buf ( n3689 , 1'b0 );
buf ( n3690 , n30374 );
buf ( n3691 , n23812 );
buf ( n3692 , 1'b0 );
buf ( n3693 , 1'b0 );
buf ( n3694 , n30371 );
buf ( n3695 , n22302 );
buf ( n3696 , 1'b0 );
buf ( n3697 , 1'b0 );
buf ( n3698 , n30356 );
buf ( n3699 , n22311 );
buf ( n3700 , 1'b0 );
buf ( n3701 , 1'b0 );
buf ( n3702 , n30356 );
buf ( n3703 , n23820 );
buf ( n3704 , 1'b0 );
buf ( n3705 , 1'b0 );
buf ( n3706 , n30343 );
buf ( n3707 , n22323 );
buf ( n3708 , 1'b0 );
buf ( n3709 , 1'b0 );
buf ( n3710 , n30374 );
buf ( n3711 , n22335 );
buf ( n3712 , 1'b0 );
buf ( n3713 , 1'b0 );
buf ( n3714 , n30355 );
buf ( n3715 , n17844 );
buf ( n3716 , 1'b0 );
buf ( n3717 , 1'b0 );
buf ( n3718 , n30358 );
buf ( n3719 , n23825 );
buf ( n3720 , 1'b0 );
buf ( n3721 , 1'b0 );
buf ( n3722 , n30355 );
buf ( n3723 , n16774 );
buf ( n3724 , 1'b0 );
buf ( n3725 , 1'b0 );
buf ( n3726 , n30355 );
buf ( n3727 , n23838 );
buf ( n3728 , 1'b0 );
buf ( n3729 , 1'b0 );
buf ( n3730 , n30376 );
buf ( n3731 , n28914 );
buf ( n3732 , 1'b0 );
buf ( n3733 , 1'b0 );
buf ( n3734 , n1 );
buf ( n3735 , n759 );
buf ( n3736 , 1'b0 );
buf ( n3737 , 1'b0 );
buf ( n3738 , n30374 );
buf ( n3739 , n22353 );
buf ( n3740 , 1'b0 );
buf ( n3741 , 1'b0 );
buf ( n3742 , n30371 );
buf ( n3743 , n22362 );
buf ( n3744 , 1'b0 );
buf ( n3745 , 1'b0 );
buf ( n3746 , n30352 );
buf ( n3747 , n23846 );
buf ( n3748 , 1'b0 );
buf ( n3749 , 1'b0 );
buf ( n3750 , n30343 );
buf ( n3751 , n22371 );
buf ( n3752 , 1'b0 );
buf ( n3753 , 1'b0 );
buf ( n3754 , n30355 );
buf ( n3755 , n22380 );
buf ( n3756 , 1'b0 );
buf ( n3757 , 1'b0 );
buf ( n3758 , n30343 );
buf ( n3759 , n22387 );
buf ( n3760 , 1'b0 );
buf ( n3761 , 1'b0 );
buf ( n3762 , n30374 );
buf ( n3763 , n17889 );
buf ( n3764 , 1'b0 );
buf ( n3765 , 1'b0 );
buf ( n3766 , n30343 );
buf ( n3767 , n20224 );
buf ( n3768 , 1'b0 );
buf ( n3769 , 1'b0 );
buf ( n3770 , n30352 );
buf ( n3771 , n23852 );
buf ( n3772 , 1'b0 );
buf ( n3773 , 1'b0 );
buf ( n3774 , n30353 );
buf ( n3775 , n21600 );
buf ( n3776 , 1'b0 );
buf ( n3777 , 1'b0 );
buf ( n3778 , n30374 );
buf ( n3779 , n22401 );
buf ( n3780 , 1'b0 );
buf ( n3781 , 1'b0 );
buf ( n3782 , n30356 );
buf ( n3783 , n22406 );
buf ( n3784 , 1'b0 );
buf ( n3785 , 1'b0 );
buf ( n3786 , n30355 );
buf ( n3787 , n22418 );
buf ( n3788 , 1'b0 );
buf ( n3789 , 1'b0 );
buf ( n3790 , n30356 );
buf ( n3791 , n27773 );
buf ( n3792 , 1'b0 );
buf ( n3793 , 1'b0 );
buf ( n3794 , n30355 );
buf ( n3795 , n22430 );
buf ( n3796 , 1'b0 );
buf ( n3797 , 1'b0 );
buf ( n3798 , n30376 );
buf ( n3799 , n22439 );
buf ( n3800 , 1'b0 );
buf ( n3801 , 1'b0 );
buf ( n3802 , n30353 );
buf ( n3803 , n22448 );
buf ( n3804 , 1'b0 );
buf ( n3805 , 1'b0 );
buf ( n3806 , n30376 );
buf ( n3807 , n22456 );
buf ( n3808 , 1'b0 );
buf ( n3809 , 1'b0 );
buf ( n3810 , n30355 );
buf ( n3811 , n22464 );
buf ( n3812 , 1'b0 );
buf ( n3813 , 1'b0 );
buf ( n3814 , n30376 );
buf ( n3815 , n23867 );
buf ( n3816 , 1'b0 );
buf ( n3817 , 1'b0 );
buf ( n3818 , n30378 );
buf ( n3819 , n23875 );
buf ( n3820 , 1'b0 );
buf ( n3821 , 1'b0 );
buf ( n3822 , n30345 );
buf ( n3823 , n23881 );
buf ( n3824 , 1'b0 );
buf ( n3825 , 1'b0 );
buf ( n3826 , n30376 );
buf ( n3827 , n23890 );
buf ( n3828 , 1'b0 );
buf ( n3829 , 1'b0 );
buf ( n3830 , n30345 );
buf ( n3831 , n22476 );
buf ( n3832 , 1'b0 );
buf ( n3833 , 1'b0 );
buf ( n3834 , n30378 );
buf ( n3835 , n23898 );
buf ( n3836 , 1'b0 );
buf ( n3837 , 1'b0 );
buf ( n3838 , n30374 );
buf ( n3839 , n23904 );
buf ( n3840 , 1'b0 );
buf ( n3841 , 1'b0 );
buf ( n3842 , n30345 );
buf ( n3843 , n23911 );
buf ( n3844 , 1'b0 );
buf ( n3845 , 1'b0 );
buf ( n3846 , n30345 );
buf ( n3847 , n23917 );
buf ( n3848 , 1'b0 );
buf ( n3849 , 1'b0 );
buf ( n3850 , n30378 );
buf ( n3851 , n23924 );
buf ( n3852 , 1'b0 );
buf ( n3853 , 1'b0 );
buf ( n3854 , n30372 );
buf ( n3855 , n23931 );
buf ( n3856 , 1'b0 );
buf ( n3857 , 1'b0 );
buf ( n3858 , n30345 );
buf ( n3859 , n20241 );
buf ( n3860 , 1'b0 );
buf ( n3861 , 1'b0 );
buf ( n3862 , n30353 );
buf ( n3863 , n16706 );
buf ( n3864 , 1'b0 );
buf ( n3865 , 1'b0 );
buf ( n3866 , n30355 );
buf ( n3867 , n25604 );
buf ( n3868 , 1'b0 );
buf ( n3869 , 1'b0 );
buf ( n3870 , n30374 );
buf ( n3871 , n15807 );
buf ( n3872 , 1'b0 );
buf ( n3873 , 1'b0 );
buf ( n3874 , n30378 );
buf ( n3875 , n29678 );
buf ( n3876 , 1'b0 );
buf ( n3877 , 1'b0 );
buf ( n3878 , n30351 );
buf ( n3879 , n17458 );
buf ( n3880 , 1'b0 );
buf ( n3881 , 1'b0 );
buf ( n3882 , n30345 );
buf ( n3883 , n17424 );
buf ( n3884 , 1'b0 );
buf ( n3885 , 1'b0 );
buf ( n3886 , n30351 );
buf ( n3887 , n18123 );
buf ( n3888 , 1'b0 );
buf ( n3889 , 1'b0 );
buf ( n3890 , n30376 );
buf ( n3891 , n22488 );
buf ( n3892 , 1'b0 );
buf ( n3893 , 1'b0 );
buf ( n3894 , n30351 );
buf ( n3895 , n29367 );
buf ( n3896 , 1'b0 );
buf ( n3897 , 1'b0 );
buf ( n3898 , n30378 );
buf ( n3899 , n28830 );
buf ( n3900 , 1'b0 );
buf ( n3901 , 1'b0 );
buf ( n3902 , n30347 );
buf ( n3903 , n28256 );
buf ( n3904 , 1'b0 );
buf ( n3905 , 1'b0 );
buf ( n3906 , n30356 );
buf ( n3907 , n27778 );
buf ( n3908 , 1'b0 );
buf ( n3909 , 1'b0 );
buf ( n3910 , n30358 );
buf ( n3911 , n22505 );
buf ( n3912 , 1'b0 );
buf ( n3913 , 1'b0 );
buf ( n3914 , n30372 );
buf ( n3915 , n25611 );
buf ( n3916 , 1'b0 );
buf ( n3917 , 1'b0 );
buf ( n3918 , n30358 );
buf ( n3919 , n18548 );
buf ( n3920 , 1'b0 );
buf ( n3921 , 1'b0 );
buf ( n3922 , n30376 );
buf ( n3923 , n18154 );
buf ( n3924 , 1'b0 );
buf ( n3925 , 1'b0 );
buf ( n3926 , n30355 );
buf ( n3927 , n20677 );
buf ( n3928 , 1'b0 );
buf ( n3929 , 1'b0 );
buf ( n3930 , n30352 );
buf ( n3931 , n18170 );
buf ( n3932 , 1'b0 );
buf ( n3933 , 1'b0 );
buf ( n3934 , n30358 );
buf ( n3935 , n18888 );
buf ( n3936 , 1'b0 );
buf ( n3937 , 1'b0 );
buf ( n3938 , n30352 );
buf ( n3939 , n19716 );
buf ( n3940 , 1'b0 );
buf ( n3941 , 1'b0 );
buf ( n3942 , n30352 );
buf ( n3943 , n18568 );
buf ( n3944 , 1'b0 );
buf ( n3945 , 1'b0 );
buf ( n3946 , n30351 );
buf ( n3947 , n22512 );
buf ( n3948 , 1'b0 );
buf ( n3949 , 1'b0 );
buf ( n3950 , n30352 );
buf ( n3951 , n23937 );
buf ( n3952 , 1'b0 );
buf ( n3953 , 1'b0 );
buf ( n3954 , n30355 );
buf ( n3955 , n22517 );
buf ( n3956 , 1'b0 );
buf ( n3957 , 1'b0 );
buf ( n3958 , n30374 );
buf ( n3959 , n22523 );
buf ( n3960 , 1'b0 );
buf ( n3961 , 1'b0 );
buf ( n3962 , n30358 );
buf ( n3963 , n22528 );
buf ( n3964 , 1'b0 );
buf ( n3965 , 1'b0 );
buf ( n3966 , n30347 );
buf ( n3967 , n22535 );
buf ( n3968 , 1'b0 );
buf ( n3969 , 1'b0 );
buf ( n3970 , n30358 );
buf ( n3971 , n22542 );
buf ( n3972 , 1'b0 );
buf ( n3973 , 1'b0 );
buf ( n3974 , n30375 );
buf ( n3975 , n23943 );
buf ( n3976 , 1'b0 );
buf ( n3977 , 1'b0 );
buf ( n3978 , n30358 );
buf ( n3979 , n23949 );
buf ( n3980 , 1'b0 );
buf ( n3981 , 1'b0 );
buf ( n3982 , n30375 );
buf ( n3983 , n22548 );
buf ( n3984 , 1'b0 );
buf ( n3985 , 1'b0 );
buf ( n3986 , n30376 );
buf ( n3987 , n22563 );
buf ( n3988 , 1'b0 );
buf ( n3989 , 1'b0 );
buf ( n3990 , n30347 );
buf ( n3991 , n22568 );
buf ( n3992 , 1'b0 );
buf ( n3993 , 1'b0 );
buf ( n3994 , n30345 );
buf ( n3995 , n23955 );
buf ( n3996 , 1'b0 );
buf ( n3997 , 1'b0 );
buf ( n3998 , n30376 );
buf ( n3999 , n22573 );
buf ( n4000 , 1'b0 );
buf ( n4001 , 1'b0 );
buf ( n4002 , n30345 );
buf ( n4003 , n23961 );
buf ( n4004 , 1'b0 );
buf ( n4005 , 1'b0 );
buf ( n4006 , n30345 );
buf ( n4007 , n23967 );
buf ( n4008 , 1'b0 );
buf ( n4009 , 1'b0 );
buf ( n4010 , n30345 );
buf ( n4011 , n22578 );
buf ( n4012 , 1'b0 );
buf ( n4013 , 1'b0 );
buf ( n4014 , n30347 );
buf ( n4015 , n23973 );
buf ( n4016 , 1'b0 );
buf ( n4017 , 1'b0 );
buf ( n4018 , n30358 );
buf ( n4019 , n23978 );
buf ( n4020 , 1'b0 );
buf ( n4021 , 1'b0 );
buf ( n4022 , n30345 );
buf ( n4023 , n28264 );
buf ( n4024 , 1'b0 );
buf ( n4025 , 1'b0 );
buf ( n4026 , n30376 );
buf ( n4027 , n27417 );
buf ( n4028 , 1'b0 );
buf ( n4029 , 1'b0 );
buf ( n4030 , n30378 );
buf ( n4031 , n22593 );
buf ( n4032 , 1'b0 );
buf ( n4033 , 1'b0 );
buf ( n4034 , n30347 );
buf ( n4035 , n20692 );
buf ( n4036 , 1'b0 );
buf ( n4037 , 1'b0 );
buf ( n4038 , n30375 );
buf ( n4039 , n20259 );
buf ( n4040 , 1'b0 );
buf ( n4041 , 1'b0 );
buf ( n4042 , n30347 );
buf ( n4043 , n28272 );
buf ( n4044 , 1'b0 );
buf ( n4045 , 1'b0 );
buf ( n4046 , n30345 );
buf ( n4047 , n27789 );
buf ( n4048 , 1'b0 );
buf ( n4049 , 1'b0 );
buf ( n4050 , n30355 );
buf ( n4051 , n25624 );
buf ( n4052 , 1'b0 );
buf ( n4053 , 1'b0 );
buf ( n4054 , n30376 );
buf ( n4055 , n22608 );
buf ( n4056 , 1'b0 );
buf ( n4057 , 1'b0 );
buf ( n4058 , n30372 );
buf ( n4059 , n22629 );
buf ( n4060 , 1'b0 );
buf ( n4061 , 1'b0 );
buf ( n4062 , n30340 );
buf ( n4063 , n23989 );
buf ( n4064 , 1'b0 );
buf ( n4065 , 1'b0 );
buf ( n4066 , n30356 );
buf ( n4067 , n23997 );
buf ( n4068 , 1'b0 );
buf ( n4069 , 1'b0 );
buf ( n4070 , n30376 );
buf ( n4071 , n22638 );
buf ( n4072 , 1'b0 );
buf ( n4073 , 1'b0 );
buf ( n4074 , n30372 );
buf ( n4075 , n24013 );
buf ( n4076 , 1'b0 );
buf ( n4077 , 1'b0 );
buf ( n4078 , n30375 );
buf ( n4079 , n24006 );
buf ( n4080 , 1'b0 );
buf ( n4081 , 1'b0 );
buf ( n4082 , n30352 );
buf ( n4083 , n22650 );
buf ( n4084 , 1'b0 );
buf ( n4085 , 1'b0 );
buf ( n4086 , n30343 );
buf ( n4087 , n22658 );
buf ( n4088 , 1'b0 );
buf ( n4089 , 1'b0 );
buf ( n4090 , n30348 );
buf ( n4091 , n22667 );
buf ( n4092 , 1'b0 );
buf ( n4093 , 1'b0 );
buf ( n4094 , n30372 );
buf ( n4095 , n22675 );
buf ( n4096 , 1'b0 );
buf ( n4097 , 1'b0 );
buf ( n4098 , n30340 );
buf ( n4099 , n22684 );
buf ( n4100 , 1'b0 );
buf ( n4101 , 1'b0 );
buf ( n4102 , n30357 );
buf ( n4103 , n22695 );
buf ( n4104 , 1'b0 );
buf ( n4105 , 1'b0 );
buf ( n4106 , n30340 );
buf ( n4107 , n22703 );
buf ( n4108 , 1'b0 );
buf ( n4109 , 1'b0 );
buf ( n4110 , n30340 );
buf ( n4111 , n22713 );
buf ( n4112 , 1'b0 );
buf ( n4113 , 1'b0 );
buf ( n4114 , n30357 );
buf ( n4115 , n24021 );
buf ( n4116 , 1'b0 );
buf ( n4117 , 1'b0 );
buf ( n4118 , n30348 );
buf ( n4119 , n22721 );
buf ( n4120 , 1'b0 );
buf ( n4121 , 1'b0 );
buf ( n4122 , n30354 );
buf ( n4123 , n24029 );
buf ( n4124 , 1'b0 );
buf ( n4125 , 1'b0 );
buf ( n4126 , n30340 );
buf ( n4127 , n24034 );
buf ( n4128 , 1'b0 );
buf ( n4129 , 1'b0 );
buf ( n4130 , n30375 );
buf ( n4131 , n17244 );
buf ( n4132 , 1'b0 );
buf ( n4133 , 1'b0 );
buf ( n4134 , n30357 );
buf ( n4135 , n22729 );
buf ( n4136 , 1'b0 );
buf ( n4137 , 1'b0 );
buf ( n4138 , n30357 );
buf ( n4139 , n27438 );
buf ( n4140 , 1'b0 );
buf ( n4141 , 1'b0 );
buf ( n4142 , n30347 );
buf ( n4143 , n22737 );
buf ( n4144 , 1'b0 );
buf ( n4145 , 1'b0 );
buf ( n4146 , n30357 );
buf ( n4147 , n24040 );
buf ( n4148 , 1'b0 );
buf ( n4149 , 1'b0 );
buf ( n4150 , n30357 );
buf ( n4151 , n24046 );
buf ( n4152 , 1'b0 );
buf ( n4153 , 1'b0 );
buf ( n4154 , n30354 );
buf ( n4155 , n24051 );
buf ( n4156 , 1'b0 );
buf ( n4157 , 1'b0 );
buf ( n4158 , n30357 );
buf ( n4159 , n24057 );
buf ( n4160 , 1'b0 );
buf ( n4161 , 1'b0 );
buf ( n4162 , n30340 );
buf ( n4163 , n20277 );
buf ( n4164 , 1'b0 );
buf ( n4165 , 1'b0 );
buf ( n4166 , n30340 );
buf ( n4167 , n22750 );
buf ( n4168 , 1'b0 );
buf ( n4169 , 1'b0 );
buf ( n4170 , n30375 );
buf ( n4171 , n24063 );
buf ( n4172 , 1'b0 );
buf ( n4173 , 1'b0 );
buf ( n4174 , n30347 );
buf ( n4175 , n22761 );
buf ( n4176 , 1'b0 );
buf ( n4177 , 1'b0 );
buf ( n4178 , n30348 );
buf ( n4179 , n18894 );
buf ( n4180 , 1'b0 );
buf ( n4181 , 1'b0 );
buf ( n4182 , n30357 );
buf ( n4183 , n24073 );
buf ( n4184 , 1'b0 );
buf ( n4185 , 1'b0 );
buf ( n4186 , n30357 );
buf ( n4187 , n22789 );
buf ( n4188 , 1'b0 );
buf ( n4189 , 1'b0 );
buf ( n4190 , n30357 );
buf ( n4191 , n22769 );
buf ( n4192 , 1'b0 );
buf ( n4193 , 1'b0 );
buf ( n4194 , n30373 );
buf ( n4195 , n18584 );
buf ( n4196 , 1'b0 );
buf ( n4197 , 1'b0 );
buf ( n4198 , n30348 );
buf ( n4199 , n22780 );
buf ( n4200 , 1'b0 );
buf ( n4201 , 1'b0 );
buf ( n4202 , n30375 );
buf ( n4203 , n22797 );
buf ( n4204 , 1'b0 );
buf ( n4205 , 1'b0 );
buf ( n4206 , n30340 );
buf ( n4207 , n18207 );
buf ( n4208 , 1'b0 );
buf ( n4209 , 1'b0 );
buf ( n4210 , n30373 );
buf ( n4211 , n22808 );
buf ( n4212 , 1'b0 );
buf ( n4213 , 1'b0 );
buf ( n4214 , n30357 );
buf ( n4215 , n22819 );
buf ( n4216 , 1'b0 );
buf ( n4217 , 1'b0 );
buf ( n4218 , n30357 );
buf ( n4219 , n22828 );
buf ( n4220 , 1'b0 );
buf ( n4221 , 1'b0 );
buf ( n4222 , n30347 );
buf ( n4223 , n22837 );
buf ( n4224 , 1'b0 );
buf ( n4225 , 1'b0 );
buf ( n4226 , n30347 );
buf ( n4227 , n22846 );
buf ( n4228 , 1'b0 );
buf ( n4229 , 1'b0 );
buf ( n4230 , n30348 );
buf ( n4231 , n22856 );
buf ( n4232 , 1'b0 );
buf ( n4233 , 1'b0 );
buf ( n4234 , n30375 );
buf ( n4235 , n22864 );
buf ( n4236 , 1'b0 );
buf ( n4237 , 1'b0 );
buf ( n4238 , n30348 );
buf ( n4239 , n17936 );
buf ( n4240 , 1'b0 );
buf ( n4241 , 1'b0 );
buf ( n4242 , n1 );
buf ( n4243 , n30208 );
buf ( n4244 , 1'b0 );
buf ( n4245 , 1'b0 );
buf ( n4246 , n30348 );
buf ( n4247 , n17211 );
buf ( n4248 , 1'b0 );
buf ( n4249 , 1'b0 );
buf ( n4250 , n30357 );
buf ( n4251 , n17688 );
buf ( n4252 , 1'b0 );
buf ( n4253 , 1'b0 );
buf ( n4254 , n30354 );
buf ( n4255 , n18238 );
buf ( n4256 , 1'b0 );
buf ( n4257 , 1'b0 );
buf ( n4258 , n30348 );
buf ( n4259 , n20715 );
buf ( n4260 , 1'b0 );
buf ( n4261 , 1'b0 );
buf ( n4262 , n30347 );
buf ( n4263 , n18253 );
buf ( n4264 , 1'b0 );
buf ( n4265 , 1'b0 );
buf ( n4266 , n30347 );
buf ( n4267 , n20296 );
buf ( n4268 , 1'b0 );
buf ( n4269 , 1'b0 );
buf ( n4270 , n30377 );
buf ( n4271 , n18604 );
buf ( n4272 , 1'b0 );
buf ( n4273 , 1'b0 );
buf ( n4274 , n30348 );
buf ( n4275 , n18618 );
buf ( n4276 , 1'b0 );
buf ( n4277 , 1'b0 );
buf ( n4278 , n30347 );
buf ( n4279 , n24079 );
buf ( n4280 , 1'b0 );
buf ( n4281 , 1'b0 );
buf ( n4282 , n30357 );
buf ( n4283 , n24085 );
buf ( n4284 , 1'b0 );
buf ( n4285 , 1'b0 );
buf ( n4286 , n30348 );
buf ( n4287 , n24091 );
buf ( n4288 , 1'b0 );
buf ( n4289 , 1'b0 );
buf ( n4290 , n30349 );
buf ( n4291 , n24096 );
buf ( n4292 , 1'b0 );
buf ( n4293 , 1'b0 );
buf ( n4294 , n30348 );
buf ( n4295 , n24103 );
buf ( n4296 , 1'b0 );
buf ( n4297 , 1'b0 );
buf ( n4298 , n30373 );
buf ( n4299 , n24108 );
buf ( n4300 , 1'b0 );
buf ( n4301 , 1'b0 );
buf ( n4302 , n30354 );
buf ( n4303 , n24113 );
buf ( n4304 , 1'b0 );
buf ( n4305 , 1'b0 );
buf ( n4306 , n30348 );
buf ( n4307 , n24119 );
buf ( n4308 , 1'b0 );
buf ( n4309 , 1'b0 );
buf ( n4310 , n30377 );
buf ( n4311 , n24124 );
buf ( n4312 , 1'b0 );
buf ( n4313 , 1'b0 );
buf ( n4314 , n30347 );
buf ( n4315 , n24129 );
buf ( n4316 , 1'b0 );
buf ( n4317 , 1'b0 );
buf ( n4318 , n30354 );
buf ( n4319 , n24134 );
buf ( n4320 , 1'b0 );
buf ( n4321 , 1'b0 );
buf ( n4322 , n30348 );
buf ( n4323 , n24140 );
buf ( n4324 , 1'b0 );
buf ( n4325 , 1'b0 );
buf ( n4326 , n30349 );
buf ( n4327 , n24145 );
buf ( n4328 , 1'b0 );
buf ( n4329 , 1'b0 );
buf ( n4330 , n30377 );
buf ( n4331 , n24150 );
buf ( n4332 , 1'b0 );
buf ( n4333 , 1'b0 );
buf ( n4334 , n30354 );
buf ( n4335 , n24156 );
buf ( n4336 , 1'b0 );
buf ( n4337 , 1'b0 );
buf ( n4338 , n30373 );
buf ( n4339 , n24161 );
buf ( n4340 , 1'b0 );
buf ( n4341 , 1'b0 );
buf ( n4342 , n30354 );
buf ( n4343 , n28280 );
buf ( n4344 , 1'b0 );
buf ( n4345 , 1'b0 );
buf ( n4346 , n30375 );
buf ( n4347 , n25650 );
buf ( n4348 , 1'b0 );
buf ( n4349 , 1'b0 );
buf ( n4350 , n30377 );
buf ( n4351 , n20313 );
buf ( n4352 , 1'b0 );
buf ( n4353 , 1'b0 );
buf ( n4354 , n30354 );
buf ( n4355 , n27713 );
buf ( n4356 , 1'b0 );
buf ( n4357 , 1'b0 );
buf ( n4358 , n30373 );
buf ( n4359 , n25663 );
buf ( n4360 , 1'b0 );
buf ( n4361 , 1'b0 );
buf ( n4362 , n30340 );
buf ( n4363 , n22879 );
buf ( n4364 , 1'b0 );
buf ( n4365 , 1'b0 );
buf ( n4366 , n30348 );
buf ( n4367 , n27420 );
buf ( n4368 , 1'b0 );
buf ( n4369 , 1'b0 );
buf ( n4370 , n30349 );
buf ( n4371 , n22887 );
buf ( n4372 , 1'b0 );
buf ( n4373 , 1'b0 );
buf ( n4374 , n30377 );
buf ( n4375 , n27998 );
buf ( n4376 , 1'b0 );
buf ( n4377 , 1'b0 );
buf ( n4378 , n30373 );
buf ( n4379 , n22895 );
buf ( n4380 , 1'b0 );
buf ( n4381 , 1'b0 );
buf ( n4382 , n30377 );
buf ( n4383 , n22907 );
buf ( n4384 , 1'b0 );
buf ( n4385 , 1'b0 );
buf ( n4386 , n30377 );
buf ( n4387 , n22915 );
buf ( n4388 , 1'b0 );
buf ( n4389 , 1'b0 );
buf ( n4390 , n30354 );
buf ( n4391 , n22924 );
buf ( n4392 , 1'b0 );
buf ( n4393 , 1'b0 );
buf ( n4394 , n30373 );
buf ( n4395 , n24169 );
buf ( n4396 , 1'b0 );
buf ( n4397 , 1'b0 );
buf ( n4398 , n30348 );
buf ( n4399 , n22932 );
buf ( n4400 , 1'b0 );
buf ( n4401 , 1'b0 );
buf ( n4402 , n30354 );
buf ( n4403 , n22943 );
buf ( n4404 , 1'b0 );
buf ( n4405 , 1'b0 );
buf ( n4406 , n30373 );
buf ( n4407 , n22951 );
buf ( n4408 , 1'b0 );
buf ( n4409 , 1'b0 );
buf ( n4410 , n30373 );
buf ( n4411 , n22959 );
buf ( n4412 , 1'b0 );
buf ( n4413 , 1'b0 );
buf ( n4414 , n30354 );
buf ( n4415 , n22968 );
buf ( n4416 , 1'b0 );
buf ( n4417 , 1'b0 );
buf ( n4418 , n30357 );
buf ( n4419 , n22985 );
buf ( n4420 , 1'b0 );
buf ( n4421 , 1'b0 );
buf ( n4422 , n30377 );
buf ( n4423 , n24176 );
buf ( n4424 , 1'b0 );
buf ( n4425 , 1'b0 );
buf ( n4426 , n30373 );
buf ( n4427 , n24184 );
buf ( n4428 , 1'b0 );
buf ( n4429 , 1'b0 );
buf ( n4430 , n30349 );
buf ( n4431 , n22993 );
buf ( n4432 , 1'b0 );
buf ( n4433 , 1'b0 );
buf ( n4434 , n30377 );
buf ( n4435 , n24197 );
buf ( n4436 , 1'b0 );
buf ( n4437 , 1'b0 );
buf ( n4438 , n30357 );
buf ( n4439 , n23001 );
buf ( n4440 , 1'b0 );
buf ( n4441 , 1'b0 );
buf ( n4442 , n30357 );
buf ( n4443 , n24205 );
buf ( n4444 , 1'b0 );
buf ( n4445 , 1'b0 );
buf ( n4446 , n30354 );
buf ( n4447 , n24213 );
buf ( n4448 , 1'b0 );
buf ( n4449 , 1'b0 );
buf ( n4450 , n30373 );
buf ( n4451 , n23009 );
buf ( n4452 , 1'b0 );
buf ( n4453 , 1'b0 );
buf ( n4454 , n30349 );
buf ( n4455 , n23017 );
buf ( n4456 , 1'b0 );
buf ( n4457 , 1'b0 );
buf ( n4458 , n30349 );
buf ( n4459 , n27337 );
buf ( n4460 , 1'b0 );
buf ( n4461 , 1'b0 );
buf ( n4462 , n30373 );
buf ( n4463 , n23025 );
buf ( n4464 , 1'b0 );
buf ( n4465 , 1'b0 );
buf ( n4466 , n30357 );
buf ( n4467 , n27340 );
buf ( n4468 , 1'b0 );
buf ( n4469 , 1'b0 );
buf ( n4470 , n30377 );
buf ( n4471 , n26583 );
buf ( n4472 , 1'b0 );
buf ( n4473 , 1'b0 );
buf ( n4474 , n30357 );
buf ( n4475 , n26588 );
buf ( n4476 , 1'b0 );
buf ( n4477 , 1'b0 );
buf ( n4478 , n30354 );
buf ( n4479 , n17895 );
buf ( n4480 , 1'b0 );
buf ( n4481 , 1'b0 );
buf ( n4482 , n30349 );
buf ( n4483 , n15853 );
buf ( n4484 , 1'b0 );
buf ( n4485 , 1'b0 );
buf ( n4486 , n30349 );
buf ( n4487 , n20730 );
buf ( n4488 , 1'b0 );
buf ( n4489 , 1'b0 );
buf ( n4490 , n30348 );
buf ( n4491 , n16825 );
buf ( n4492 , 1'b0 );
buf ( n4493 , 1'b0 );
buf ( n4494 , n30349 );
buf ( n4495 , n25677 );
buf ( n4496 , 1'b0 );
buf ( n4497 , 1'b0 );
buf ( n4498 , n30373 );
buf ( n4499 , n28644 );
buf ( n4500 , 1'b0 );
buf ( n4501 , 1'b0 );
buf ( n4502 , n30348 );
buf ( n4503 , n24226 );
buf ( n4504 , 1'b0 );
buf ( n4505 , 1'b0 );
buf ( n4506 , n30373 );
buf ( n4507 , n20331 );
buf ( n4508 , 1'b0 );
buf ( n4509 , 1'b0 );
buf ( n4510 , n30357 );
buf ( n4511 , n25687 );
buf ( n4512 , 1'b0 );
buf ( n4513 , 1'b0 );
buf ( n4514 , n30349 );
buf ( n4515 , n24236 );
buf ( n4516 , 1'b0 );
buf ( n4517 , 1'b0 );
buf ( n4518 , n1 );
buf ( n4519 , n19721 );
buf ( n4520 , 1'b0 );
buf ( n4521 , 1'b0 );
buf ( n4522 , n30348 );
buf ( n4523 , n20744 );
buf ( n4524 , 1'b0 );
buf ( n4525 , 1'b0 );
buf ( n4526 , n30372 );
buf ( n4527 , n23476 );
buf ( n4528 , 1'b0 );
buf ( n4529 , 1'b0 );
buf ( n4530 , n30354 );
buf ( n4531 , n25693 );
buf ( n4532 , 1'b0 );
buf ( n4533 , 1'b0 );
buf ( n4534 , n30349 );
buf ( n4535 , n20336 );
buf ( n4536 , 1'b0 );
buf ( n4537 , 1'b0 );
buf ( n4538 , n30354 );
buf ( n4539 , n25698 );
buf ( n4540 , 1'b0 );
buf ( n4541 , 1'b0 );
buf ( n4542 , n30348 );
buf ( n4543 , n25707 );
buf ( n4544 , 1'b0 );
buf ( n4545 , 1'b0 );
buf ( n4546 , n30373 );
buf ( n4547 , n25714 );
buf ( n4548 , 1'b0 );
buf ( n4549 , 1'b0 );
buf ( n4550 , n30373 );
buf ( n4551 , n25721 );
buf ( n4552 , 1'b0 );
buf ( n4553 , 1'b0 );
buf ( n4554 , n30354 );
buf ( n4555 , n25729 );
buf ( n4556 , 1'b0 );
buf ( n4557 , 1'b0 );
buf ( n4558 , n30348 );
buf ( n4559 , n23033 );
buf ( n4560 , 1'b0 );
buf ( n4561 , 1'b0 );
buf ( n4562 , n30349 );
buf ( n4563 , n25735 );
buf ( n4564 , 1'b0 );
buf ( n4565 , 1'b0 );
buf ( n4566 , n30354 );
buf ( n4567 , n17791 );
buf ( n4568 , 1'b0 );
buf ( n4569 , 1'b0 );
buf ( n4570 , n1 );
buf ( n4571 , n30069 );
buf ( n4572 , 1'b0 );
buf ( n4573 , 1'b0 );
buf ( n4574 , n1 );
buf ( n4575 , n29923 );
buf ( n4576 , 1'b0 );
buf ( n4577 , 1'b0 );
buf ( n4578 , n30349 );
buf ( n4579 , n17493 );
buf ( n4580 , 1'b0 );
buf ( n4581 , 1'b0 );
buf ( n4582 , n30354 );
buf ( n4583 , n18619 );
buf ( n4584 , 1'b0 );
buf ( n4585 , 1'b0 );
buf ( n4586 , n30373 );
buf ( n4587 , n17750 );
buf ( n4588 , 1'b0 );
buf ( n4589 , 1'b0 );
buf ( n4590 , n30348 );
buf ( n4591 , n18635 );
buf ( n4592 , 1'b0 );
buf ( n4593 , 1'b0 );
buf ( n4594 , n30372 );
buf ( n4595 , n18284 );
buf ( n4596 , 1'b0 );
buf ( n4597 , 1'b0 );
buf ( n4598 , n30373 );
buf ( n4599 , n19739 );
buf ( n4600 , 1'b0 );
buf ( n4601 , 1'b0 );
buf ( n4602 , n30373 );
buf ( n4603 , n25742 );
buf ( n4604 , 1'b0 );
buf ( n4605 , 1'b0 );
buf ( n4606 , n30349 );
buf ( n4607 , n25748 );
buf ( n4608 , 1'b0 );
buf ( n4609 , 1'b0 );
buf ( n4610 , n30348 );
buf ( n4611 , n25273 );
buf ( n4612 , 1'b0 );
buf ( n4613 , 1'b0 );
buf ( n4614 , n30340 );
buf ( n4615 , n20775 );
buf ( n4616 , 1'b0 );
buf ( n4617 , 1'b0 );
buf ( n4618 , n30354 );
buf ( n4619 , n20147 );
buf ( n4620 , 1'b0 );
buf ( n4621 , 1'b0 );
buf ( n4622 , n30354 );
buf ( n4623 , n23041 );
buf ( n4624 , 1'b0 );
buf ( n4625 , 1'b0 );
buf ( n4626 , n30377 );
buf ( n4627 , n23049 );
buf ( n4628 , 1'b0 );
buf ( n4629 , 1'b0 );
buf ( n4630 , n30354 );
buf ( n4631 , n23057 );
buf ( n4632 , 1'b0 );
buf ( n4633 , 1'b0 );
buf ( n4634 , n30357 );
buf ( n4635 , n23065 );
buf ( n4636 , 1'b0 );
buf ( n4637 , 1'b0 );
buf ( n4638 , n30349 );
buf ( n4639 , n24247 );
buf ( n4640 , 1'b0 );
buf ( n4641 , 1'b0 );
buf ( n4642 , n1 );
buf ( n4643 , n30085 );
buf ( n4644 , 1'b0 );
buf ( n4645 , 1'b0 );
buf ( n4646 , n30372 );
buf ( n4647 , n27435 );
buf ( n4648 , 1'b0 );
buf ( n4649 , 1'b0 );
buf ( n4650 , n30349 );
buf ( n4651 , n18320 );
buf ( n4652 , 1'b0 );
buf ( n4653 , 1'b0 );
buf ( n4654 , n30372 );
buf ( n4655 , n17527 );
buf ( n4656 , 1'b0 );
buf ( n4657 , 1'b0 );
buf ( n4658 , n30354 );
buf ( n4659 , n16453 );
buf ( n4660 , 1'b0 );
buf ( n4661 , 1'b0 );
buf ( n4662 , n1 );
buf ( n4663 , n30097 );
buf ( n4664 , 1'b0 );
buf ( n4665 , 1'b0 );
buf ( n4666 , n30354 );
buf ( n4667 , n25755 );
buf ( n4668 , 1'b0 );
buf ( n4669 , 1'b0 );
buf ( n4670 , n30377 );
buf ( n4671 , n25761 );
buf ( n4672 , 1'b0 );
buf ( n4673 , 1'b0 );
buf ( n4674 , n30349 );
buf ( n4675 , n23080 );
buf ( n4676 , 1'b0 );
buf ( n4677 , 1'b0 );
buf ( n4678 , n30377 );
buf ( n4679 , n25767 );
buf ( n4680 , 1'b0 );
buf ( n4681 , 1'b0 );
buf ( n4682 , n30377 );
buf ( n4683 , n25773 );
buf ( n4684 , 1'b0 );
buf ( n4685 , 1'b0 );
buf ( n4686 , n30349 );
buf ( n4687 , n20840 );
buf ( n4688 , 1'b0 );
buf ( n4689 , 1'b0 );
buf ( n4690 , n30377 );
buf ( n4691 , n20129 );
buf ( n4692 , 1'b0 );
buf ( n4693 , 1'b0 );
buf ( n4694 , n30373 );
buf ( n4695 , n17605 );
buf ( n4696 , 1'b0 );
buf ( n4697 , 1'b0 );
buf ( n4698 , n30354 );
buf ( n4699 , n18335 );
buf ( n4700 , 1'b0 );
buf ( n4701 , 1'b0 );
buf ( n4702 , n1 );
buf ( n4703 , n19814 );
buf ( n4704 , 1'b0 );
buf ( n4705 , 1'b0 );
buf ( n4706 , n30357 );
buf ( n4707 , n18904 );
buf ( n4708 , 1'b0 );
buf ( n4709 , 1'b0 );
buf ( n4710 , n30377 );
buf ( n4711 , n18917 );
buf ( n4712 , 1'b0 );
buf ( n4713 , 1'b0 );
buf ( n4714 , n30372 );
buf ( n4715 , n18655 );
buf ( n4716 , 1'b0 );
buf ( n4717 , 1'b0 );
buf ( n4718 , n30377 );
buf ( n4719 , n25779 );
buf ( n4720 , 1'b0 );
buf ( n4721 , 1'b0 );
buf ( n4722 , n30373 );
buf ( n4723 , n25784 );
buf ( n4724 , 1'b0 );
buf ( n4725 , 1'b0 );
buf ( n4726 , n30349 );
buf ( n4727 , n25790 );
buf ( n4728 , 1'b0 );
buf ( n4729 , 1'b0 );
buf ( n4730 , n30377 );
buf ( n4731 , n25796 );
buf ( n4732 , 1'b0 );
buf ( n4733 , 1'b0 );
buf ( n4734 , n30377 );
buf ( n4735 , n25802 );
buf ( n4736 , 1'b0 );
buf ( n4737 , 1'b0 );
buf ( n4738 , n30372 );
buf ( n4739 , n25808 );
buf ( n4740 , 1'b0 );
buf ( n4741 , 1'b0 );
buf ( n4742 , n30377 );
buf ( n4743 , n25819 );
buf ( n4744 , 1'b0 );
buf ( n4745 , 1'b0 );
buf ( n4746 , n30373 );
buf ( n4747 , n25909 );
buf ( n4748 , 1'b0 );
buf ( n4749 , 1'b0 );
buf ( n4750 , n30372 );
buf ( n4751 , n25915 );
buf ( n4752 , 1'b0 );
buf ( n4753 , 1'b0 );
buf ( n4754 , n30377 );
buf ( n4755 , n25920 );
buf ( n4756 , 1'b0 );
buf ( n4757 , 1'b0 );
buf ( n4758 , n30349 );
buf ( n4759 , n25926 );
buf ( n4760 , 1'b0 );
buf ( n4761 , 1'b0 );
buf ( n4762 , n30372 );
buf ( n4763 , n25932 );
buf ( n4764 , 1'b0 );
buf ( n4765 , 1'b0 );
buf ( n4766 , n30372 );
buf ( n4767 , n25999 );
buf ( n4768 , 1'b0 );
buf ( n4769 , 1'b0 );
buf ( n4770 , n30349 );
buf ( n4771 , n26004 );
buf ( n4772 , 1'b0 );
buf ( n4773 , 1'b0 );
buf ( n4774 , n30372 );
buf ( n4775 , n26009 );
buf ( n4776 , 1'b0 );
buf ( n4777 , 1'b0 );
buf ( n4778 , n30373 );
buf ( n4779 , n18934 );
buf ( n4780 , 1'b0 );
buf ( n4781 , 1'b0 );
buf ( n4782 , n30373 );
buf ( n4783 , n18678 );
buf ( n4784 , 1'b0 );
buf ( n4785 , 1'b0 );
buf ( n4786 , n30349 );
buf ( n4787 , n26700 );
buf ( n4788 , 1'b0 );
buf ( n4789 , 1'b0 );
buf ( n4790 , n30372 );
buf ( n4791 , n26711 );
buf ( n4792 , 1'b0 );
buf ( n4793 , 1'b0 );
buf ( n4794 , n30349 );
buf ( n4795 , n26023 );
buf ( n4796 , 1'b0 );
buf ( n4797 , 1'b0 );
buf ( n4798 , n30377 );
buf ( n4799 , n27301 );
buf ( n4800 , 1'b0 );
buf ( n4801 , 1'b0 );
buf ( n4802 , n30377 );
buf ( n4803 , n30384 );
buf ( n4804 , 1'b0 );
buf ( n4805 , 1'b0 );
buf ( n4806 , n30372 );
buf ( n4807 , n19822 );
buf ( n4808 , 1'b0 );
buf ( n4809 , 1'b0 );
buf ( n4810 , n30377 );
buf ( n4811 , n26029 );
buf ( n4812 , 1'b0 );
buf ( n4813 , 1'b0 );
buf ( n4814 , n30349 );
buf ( n4815 , n26035 );
buf ( n4816 , 1'b0 );
buf ( n4817 , 1'b0 );
buf ( n4818 , n30377 );
buf ( n4819 , n17842 );
buf ( n4820 , 1'b0 );
buf ( n4821 , 1'b0 );
buf ( n4822 , n30357 );
buf ( n4823 , n17842 );
buf ( n4824 , 1'b0 );
buf ( n4825 , 1'b0 );
buf ( n4826 , n30373 );
buf ( n4827 , n20122 );
buf ( n4828 , 1'b0 );
buf ( n4829 , 1'b0 );
buf ( n4830 , n30377 );
buf ( n4831 , n20857 );
buf ( n4832 , 1'b0 );
buf ( n4833 , 1'b0 );
buf ( n4834 , n30377 );
buf ( n4835 , n17733 );
buf ( n4836 , 1'b0 );
buf ( n4837 , 1'b0 );
buf ( n4838 , n30349 );
buf ( n4839 , n20104 );
buf ( n4840 , 1'b0 );
buf ( n4841 , 1'b0 );
buf ( n4842 , n1 );
buf ( n4843 , n19896 );
buf ( n4844 , 1'b0 );
buf ( n4845 , 1'b0 );
buf ( n4846 , n30354 );
buf ( n4847 , n16761 );
buf ( n4848 , 1'b0 );
buf ( n4849 , 1'b0 );
buf ( n4850 , n1 );
buf ( n4851 , n19024 );
buf ( n4852 , 1'b0 );
buf ( n4853 , 1'b0 );
buf ( n4854 , n30354 );
buf ( n4855 , n18948 );
buf ( n4856 , 1'b0 );
buf ( n4857 , 1'b0 );
buf ( n4858 , n30377 );
buf ( n4859 , n18366 );
buf ( n4860 , 1'b0 );
buf ( n4861 , 1'b0 );
buf ( n4862 , n30354 );
buf ( n4863 , n18691 );
buf ( n4864 , 1'b0 );
buf ( n4865 , 1'b0 );
buf ( n4866 , n30340 );
buf ( n4867 , n19914 );
buf ( n4868 , 1'b0 );
buf ( n4869 , 1'b0 );
buf ( n4870 , n30348 );
buf ( n4871 , n26725 );
buf ( n4872 , 1'b0 );
buf ( n4873 , 1'b0 );
buf ( n4874 , n30373 );
buf ( n4875 , n26051 );
buf ( n4876 , 1'b0 );
buf ( n4877 , 1'b0 );
buf ( n4878 , n30372 );
buf ( n4879 , n20871 );
buf ( n4880 , 1'b0 );
buf ( n4881 , 1'b0 );
buf ( n4882 , n1 );
buf ( n4883 , n19106 );
buf ( n4884 , 1'b0 );
buf ( n4885 , 1'b0 );
buf ( n4886 , n30373 );
buf ( n4887 , n18413 );
buf ( n4888 , 1'b0 );
buf ( n4889 , 1'b0 );
buf ( n4890 , n30354 );
buf ( n4891 , n19112 );
buf ( n4892 , 1'b0 );
buf ( n4893 , 1'b0 );
buf ( n4894 , n30348 );
buf ( n4895 , n19925 );
buf ( n4896 , 1'b0 );
buf ( n4897 , 1'b0 );
buf ( n4898 , n30354 );
buf ( n4899 , n30380 );
buf ( n4900 , 1'b0 );
buf ( n4901 , 1'b0 );
buf ( n4902 , n30373 );
buf ( n4903 , n23468 );
buf ( n4904 , 1'b0 );
buf ( n4905 , 1'b0 );
buf ( n4906 , n30348 );
buf ( n4907 , n18450 );
buf ( n4908 , 1'b0 );
buf ( n4909 , 1'b0 );
buf ( n4910 , n1 );
buf ( n4911 , n29943 );
buf ( n4912 , 1'b0 );
buf ( n4913 , 1'b0 );
buf ( n4914 , n30354 );
buf ( n4915 , n18470 );
buf ( n4916 , 1'b0 );
buf ( n4917 , 1'b0 );
buf ( n4918 , n30372 );
buf ( n4919 , n19118 );
buf ( n4920 , 1'b0 );
buf ( n4921 , 1'b0 );
buf ( n4922 , n30349 );
buf ( n4923 , n19124 );
buf ( n4924 , 1'b0 );
buf ( n4925 , 1'b0 );
buf ( n4926 , n30357 );
buf ( n4927 , n19130 );
buf ( n4928 , 1'b0 );
buf ( n4929 , 1'b0 );
buf ( n4930 , n30348 );
buf ( n4931 , n18480 );
buf ( n4932 , 1'b0 );
buf ( n4933 , 1'b0 );
buf ( n4934 , n30349 );
buf ( n4935 , n19134 );
buf ( n4936 , 1'b0 );
buf ( n4937 , 1'b0 );
buf ( n4938 , n30354 );
buf ( n4939 , n18490 );
buf ( n4940 , 1'b0 );
buf ( n4941 , 1'b0 );
buf ( n4942 , n30357 );
buf ( n4943 , n18027 );
buf ( n4944 , 1'b0 );
buf ( n4945 , 1'b0 );
buf ( n4946 , n30373 );
buf ( n4947 , n17997 );
buf ( n4948 , 1'b0 );
buf ( n4949 , 1'b0 );
buf ( n4950 , n30349 );
buf ( n4951 , n17974 );
buf ( n4952 , 1'b0 );
buf ( n4953 , 1'b0 );
buf ( n4954 , n30373 );
buf ( n4955 , n1141 );
buf ( n4956 , 1'b0 );
buf ( n4957 , 1'b0 );
buf ( n4958 , n30354 );
buf ( n4959 , n1130 );
buf ( n4960 , 1'b0 );
buf ( n4961 , 1'b0 );
buf ( n4962 , n30349 );
buf ( n4963 , n1134 );
buf ( n4964 , 1'b0 );
buf ( n4965 , 1'b0 );
buf ( n4966 , n30373 );
buf ( n4967 , n1135 );
buf ( n4968 , 1'b0 );
buf ( n4969 , 1'b0 );
buf ( n4970 , n30357 );
buf ( n4971 , n19997 );
buf ( n4972 , 1'b0 );
buf ( n4973 , 1'b0 );
buf ( n4974 , n30354 );
buf ( n4975 , n19140 );
buf ( n4976 , 1'b0 );
buf ( n4977 , 1'b0 );
buf ( n4978 , n30354 );
buf ( n4979 , n17961 );
buf ( n4980 , 1'b0 );
buf ( n4981 , 1'b0 );
buf ( n4982 , n30348 );
buf ( n4983 , n18870 );
buf ( n4984 , 1'b0 );
buf ( n4985 , 1'b0 );
buf ( n4986 , n30354 );
buf ( n4987 , n20889 );
buf ( n4988 , 1'b0 );
buf ( n4989 , 1'b0 );
buf ( n4990 , n30377 );
buf ( n4991 , n20900 );
buf ( n4992 , 1'b0 );
buf ( n4993 , 1'b0 );
buf ( n4994 , n30340 );
buf ( n4995 , n20882 );
buf ( n4996 , 1'b0 );
buf ( n4997 , 1'b0 );
buf ( n4998 , n30373 );
buf ( n4999 , n20909 );
buf ( n5000 , 1'b0 );
buf ( n5001 , 1'b0 );
buf ( n5002 , n30377 );
buf ( n5003 , n20920 );
buf ( n5004 , 1'b0 );
buf ( n5005 , 1'b0 );
buf ( n5006 , n30375 );
buf ( n5007 , n20934 );
buf ( n5008 , 1'b0 );
buf ( n5009 , 1'b0 );
buf ( n5010 , n1 );
buf ( n5011 , n26773 );
buf ( n5012 , 1'b0 );
buf ( n5013 , 1'b0 );
buf ( n5014 , n30354 );
buf ( n5015 , n20437 );
buf ( n5016 , 1'b0 );
buf ( n5017 , 1'b0 );
buf ( n5018 , n30377 );
buf ( n5019 , n20943 );
buf ( n5020 , 1'b0 );
buf ( n5021 , 1'b0 );
buf ( n5022 , n30348 );
buf ( n5023 , n20951 );
buf ( n5024 , 1'b0 );
buf ( n5025 , 1'b0 );
buf ( n5026 , n30354 );
buf ( n5027 , n20760 );
buf ( n5028 , 1'b0 );
buf ( n5029 , 1'b0 );
buf ( n5030 , n30354 );
buf ( n5031 , n20701 );
buf ( n5032 , 1'b0 );
buf ( n5033 , 1'b0 );
buf ( n5034 , n30373 );
buf ( n5035 , n20959 );
buf ( n5036 , 1'b0 );
buf ( n5037 , 1'b0 );
buf ( n5038 , n30349 );
buf ( n5039 , n24270 );
buf ( n5040 , 1'b0 );
buf ( n5041 , 1'b0 );
buf ( n5042 , n30348 );
buf ( n5043 , n20001 );
buf ( n5044 , 1'b0 );
buf ( n5045 , 1'b0 );
buf ( n5046 , n30348 );
buf ( n5047 , n20968 );
buf ( n5048 , 1'b0 );
buf ( n5049 , 1'b0 );
buf ( n5050 , n30377 );
buf ( n5051 , n20010 );
buf ( n5052 , 1'b0 );
buf ( n5053 , 1'b0 );
buf ( n5054 , n30347 );
buf ( n5055 , n20014 );
buf ( n5056 , 1'b0 );
buf ( n5057 , 1'b0 );
buf ( n5058 , n30348 );
buf ( n5059 , n20018 );
buf ( n5060 , 1'b0 );
buf ( n5061 , 1'b0 );
buf ( n5062 , n30375 );
buf ( n5063 , n20022 );
buf ( n5064 , 1'b0 );
buf ( n5065 , 1'b0 );
buf ( n5066 , n30348 );
buf ( n5067 , n20976 );
buf ( n5068 , 1'b0 );
buf ( n5069 , 1'b0 );
buf ( n5070 , n30347 );
buf ( n5071 , n22496 );
buf ( n5072 , 1'b0 );
buf ( n5073 , 1'b0 );
buf ( n5074 , n1 );
buf ( n5075 , n30244 );
buf ( n5076 , 1'b0 );
buf ( n5077 , 1'b0 );
buf ( n5078 , n30357 );
buf ( n5079 , n22976 );
buf ( n5080 , 1'b0 );
buf ( n5081 , 1'b0 );
buf ( n5082 , n30340 );
buf ( n5083 , n22558 );
buf ( n5084 , 1'b0 );
buf ( n5085 , 1'b0 );
buf ( n5086 , n30375 );
buf ( n5087 , n20453 );
buf ( n5088 , 1'b0 );
buf ( n5089 , 1'b0 );
buf ( n5090 , n30373 );
buf ( n5091 , n24285 );
buf ( n5092 , 1'b0 );
buf ( n5093 , 1'b0 );
buf ( n5094 , n30357 );
buf ( n5095 , n1129 );
buf ( n5096 , 1'b0 );
buf ( n5097 , 1'b0 );
buf ( n5098 , n30347 );
buf ( n5099 , n1133 );
buf ( n5100 , 1'b0 );
buf ( n5101 , 1'b0 );
buf ( n5102 , n30375 );
buf ( n5103 , n24348 );
buf ( n5104 , 1'b0 );
buf ( n5105 , 1'b0 );
buf ( n5106 , n30340 );
buf ( n5107 , n20982 );
buf ( n5108 , 1'b0 );
buf ( n5109 , 1'b0 );
buf ( n5110 , n30357 );
buf ( n5111 , n20988 );
buf ( n5112 , 1'b0 );
buf ( n5113 , 1'b0 );
buf ( n5114 , n30357 );
buf ( n5115 , n20994 );
buf ( n5116 , 1'b0 );
buf ( n5117 , 1'b0 );
buf ( n5118 , n30347 );
buf ( n5119 , n21002 );
buf ( n5120 , 1'b0 );
buf ( n5121 , 1'b0 );
buf ( n5122 , n1 );
buf ( n5123 , n30192 );
buf ( n5124 , 1'b0 );
buf ( n5125 , 1'b0 );
buf ( n5126 , n1 );
buf ( n5127 , n30093 );
buf ( n5128 , 1'b0 );
buf ( n5129 , 1'b0 );
buf ( n5130 , n30357 );
buf ( n5131 , n19703 );
buf ( n5132 , 1'b0 );
buf ( n5133 , 1'b0 );
buf ( n5134 , n1 );
buf ( n5135 , n30136 );
buf ( n5136 , 1'b0 );
buf ( n5137 , 1'b0 );
buf ( n5138 , n30375 );
buf ( n5139 , n20460 );
buf ( n5140 , 1'b0 );
buf ( n5141 , 1'b0 );
buf ( n5142 , n1 );
buf ( n5143 , n29897 );
buf ( n5144 , 1'b0 );
buf ( n5145 , 1'b0 );
buf ( n5146 , n30372 );
buf ( n5147 , n19395 );
buf ( n5148 , 1'b0 );
buf ( n5149 , 1'b0 );
buf ( n5150 , n30348 );
buf ( n5151 , n20086 );
buf ( n5152 , 1'b0 );
buf ( n5153 , 1'b0 );
buf ( n5154 , n30352 );
buf ( n5155 , n18697 );
buf ( n5156 , 1'b0 );
buf ( n5157 , 1'b0 );
buf ( n5158 , n30375 );
buf ( n5159 , n20026 );
buf ( n5160 , 1'b0 );
buf ( n5161 , 1'b0 );
buf ( n5162 , n30356 );
buf ( n5163 , n20027 );
buf ( n5164 , 1'b0 );
buf ( n5165 , 1'b0 );
buf ( n5166 , n30340 );
buf ( n5167 , n20030 );
buf ( n5168 , 1'b0 );
buf ( n5169 , 1'b0 );
buf ( n5170 , n30376 );
buf ( n5171 , n20038 );
buf ( n5172 , 1'b0 );
buf ( n5173 , 1'b0 );
buf ( n5174 , n1 );
buf ( n5175 , n29889 );
buf ( n5176 , 1'b0 );
buf ( n5177 , 1'b0 );
buf ( n5178 , n30372 );
buf ( n5179 , n21023 );
buf ( n5180 , 1'b0 );
buf ( n5181 , 1'b0 );
buf ( n5182 , n30376 );
buf ( n5183 , n21011 );
buf ( n5184 , 1'b0 );
buf ( n5185 , 1'b0 );
buf ( n5186 , n30376 );
buf ( n5187 , n20471 );
buf ( n5188 , 1'b0 );
buf ( n5189 , 1'b0 );
buf ( n5190 , n30349 );
buf ( n5191 , n22395 );
buf ( n5192 , 1'b0 );
buf ( n5193 , 1'b0 );
buf ( n5194 , n30376 );
buf ( n5195 , n21492 );
buf ( n5196 , 1'b0 );
buf ( n5197 , 1'b0 );
buf ( n5198 , n30378 );
buf ( n5199 , n20480 );
buf ( n5200 , 1'b0 );
buf ( n5201 , 1'b0 );
buf ( n5202 , n30375 );
buf ( n5203 , n21728 );
buf ( n5204 , 1'b0 );
buf ( n5205 , 1'b0 );
buf ( n5206 , n30372 );
buf ( n5207 , n21736 );
buf ( n5208 , 1'b0 );
buf ( n5209 , 1'b0 );
buf ( n5210 , n30372 );
buf ( n5211 , n22343 );
buf ( n5212 , 1'b0 );
buf ( n5213 , 1'b0 );
buf ( n5214 , n30375 );
buf ( n5215 , n21776 );
buf ( n5216 , 1'b0 );
buf ( n5217 , 1'b0 );
buf ( n5218 , n30375 );
buf ( n5219 , n20491 );
buf ( n5220 , 1'b0 );
buf ( n5221 , 1'b0 );
buf ( n5222 , n30355 );
buf ( n5223 , n21031 );
buf ( n5224 , 1'b0 );
buf ( n5225 , 1'b0 );
buf ( n5226 , n30375 );
buf ( n5227 , n21039 );
buf ( n5228 , 1'b0 );
buf ( n5229 , 1'b0 );
buf ( n5230 , n30375 );
buf ( n5231 , n23501 );
buf ( n5232 , 1'b0 );
buf ( n5233 , 1'b0 );
buf ( n5234 , n30378 );
buf ( n5235 , n21047 );
buf ( n5236 , 1'b0 );
buf ( n5237 , 1'b0 );
buf ( n5238 , n30347 );
buf ( n5239 , n21056 );
buf ( n5240 , 1'b0 );
buf ( n5241 , 1'b0 );
buf ( n5242 , n30347 );
buf ( n5243 , n20504 );
buf ( n5244 , 1'b0 );
buf ( n5245 , 1'b0 );
buf ( n5246 , n30345 );
buf ( n5247 , n21066 );
buf ( n5248 , 1'b0 );
buf ( n5249 , 1'b0 );
buf ( n5250 , n30378 );
buf ( n5251 , n21556 );
buf ( n5252 , 1'b0 );
buf ( n5253 , 1'b0 );
buf ( n5254 , n30347 );
buf ( n5255 , n21074 );
buf ( n5256 , 1'b0 );
buf ( n5257 , 1'b0 );
buf ( n5258 , n30347 );
buf ( n5259 , n21082 );
buf ( n5260 , 1'b0 );
buf ( n5261 , 1'b0 );
buf ( n5262 , n30378 );
buf ( n5263 , n21091 );
buf ( n5264 , 1'b0 );
buf ( n5265 , 1'b0 );
buf ( n5266 , n30378 );
buf ( n5267 , n21100 );
buf ( n5268 , 1'b0 );
buf ( n5269 , 1'b0 );
buf ( n5270 , n30375 );
buf ( n5271 , n21108 );
buf ( n5272 , 1'b0 );
buf ( n5273 , 1'b0 );
buf ( n5274 , n30374 );
buf ( n5275 , n21117 );
buf ( n5276 , 1'b0 );
buf ( n5277 , 1'b0 );
buf ( n5278 , n30358 );
buf ( n5279 , n21126 );
buf ( n5280 , 1'b0 );
buf ( n5281 , 1'b0 );
buf ( n5282 , n30358 );
buf ( n5283 , n21564 );
buf ( n5284 , 1'b0 );
buf ( n5285 , 1'b0 );
buf ( n5286 , n30347 );
buf ( n5287 , n21135 );
buf ( n5288 , 1'b0 );
buf ( n5289 , 1'b0 );
buf ( n5290 , n30358 );
buf ( n5291 , n21143 );
buf ( n5292 , 1'b0 );
buf ( n5293 , 1'b0 );
buf ( n5294 , n30347 );
buf ( n5295 , n23509 );
buf ( n5296 , 1'b0 );
buf ( n5297 , 1'b0 );
buf ( n5298 , n30372 );
buf ( n5299 , n21151 );
buf ( n5300 , 1'b0 );
buf ( n5301 , 1'b0 );
buf ( n5302 , n30358 );
buf ( n5303 , n21159 );
buf ( n5304 , 1'b0 );
buf ( n5305 , 1'b0 );
buf ( n5306 , n30358 );
buf ( n5307 , n21168 );
buf ( n5308 , 1'b0 );
buf ( n5309 , 1'b0 );
buf ( n5310 , n30374 );
buf ( n5311 , n21178 );
buf ( n5312 , 1'b0 );
buf ( n5313 , 1'b0 );
buf ( n5314 , n30372 );
buf ( n5315 , n21548 );
buf ( n5316 , 1'b0 );
buf ( n5317 , 1'b0 );
buf ( n5318 , n30358 );
buf ( n5319 , n20513 );
buf ( n5320 , 1'b0 );
buf ( n5321 , 1'b0 );
buf ( n5322 , n30358 );
buf ( n5323 , n21187 );
buf ( n5324 , 1'b0 );
buf ( n5325 , 1'b0 );
buf ( n5326 , n30374 );
buf ( n5327 , n21196 );
buf ( n5328 , 1'b0 );
buf ( n5329 , 1'b0 );
buf ( n5330 , n30374 );
buf ( n5331 , n21516 );
buf ( n5332 , 1'b0 );
buf ( n5333 , 1'b0 );
buf ( n5334 , n30347 );
buf ( n5335 , n21204 );
buf ( n5336 , 1'b0 );
buf ( n5337 , 1'b0 );
buf ( n5338 , n30356 );
buf ( n5339 , n21212 );
buf ( n5340 , 1'b0 );
buf ( n5341 , 1'b0 );
buf ( n5342 , n30374 );
buf ( n5343 , n21221 );
buf ( n5344 , 1'b0 );
buf ( n5345 , 1'b0 );
buf ( n5346 , n30345 );
buf ( n5347 , n21508 );
buf ( n5348 , 1'b0 );
buf ( n5349 , 1'b0 );
buf ( n5350 , n30376 );
buf ( n5351 , n23457 );
buf ( n5352 , 1'b0 );
buf ( n5353 , 1'b0 );
buf ( n5354 , n30376 );
buf ( n5355 , n21720 );
buf ( n5356 , 1'b0 );
buf ( n5357 , 1'b0 );
buf ( n5358 , n30351 );
buf ( n5359 , n20523 );
buf ( n5360 , 1'b0 );
buf ( n5361 , 1'b0 );
buf ( n5362 , n30351 );
buf ( n5363 , n21229 );
buf ( n5364 , 1'b0 );
buf ( n5365 , 1'b0 );
buf ( n5366 , n30347 );
buf ( n5367 , n21712 );
buf ( n5368 , 1'b0 );
buf ( n5369 , 1'b0 );
buf ( n5370 , n30355 );
buf ( n5371 , n21237 );
buf ( n5372 , 1'b0 );
buf ( n5373 , 1'b0 );
buf ( n5374 , n30351 );
buf ( n5375 , n23484 );
buf ( n5376 , 1'b0 );
buf ( n5377 , 1'b0 );
buf ( n5378 , n30351 );
buf ( n5379 , n21245 );
buf ( n5380 , 1'b0 );
buf ( n5381 , 1'b0 );
buf ( n5382 , n30356 );
buf ( n5383 , n21253 );
buf ( n5384 , 1'b0 );
buf ( n5385 , 1'b0 );
buf ( n5386 , n30345 );
buf ( n5387 , n21277 );
buf ( n5388 , 1'b0 );
buf ( n5389 , 1'b0 );
buf ( n5390 , n30353 );
buf ( n5391 , n21261 );
buf ( n5392 , 1'b0 );
buf ( n5393 , 1'b0 );
buf ( n5394 , n30378 );
buf ( n5395 , n21269 );
buf ( n5396 , 1'b0 );
buf ( n5397 , 1'b0 );
buf ( n5398 , n30374 );
buf ( n5399 , n21285 );
buf ( n5400 , 1'b0 );
buf ( n5401 , 1'b0 );
buf ( n5402 , n30374 );
buf ( n5403 , n21704 );
buf ( n5404 , 1'b0 );
buf ( n5405 , 1'b0 );
buf ( n5406 , n30353 );
buf ( n5407 , n21500 );
buf ( n5408 , 1'b0 );
buf ( n5409 , 1'b0 );
buf ( n5410 , n30353 );
buf ( n5411 , n20534 );
buf ( n5412 , 1'b0 );
buf ( n5413 , 1'b0 );
buf ( n5414 , n30378 );
buf ( n5415 , n21293 );
buf ( n5416 , 1'b0 );
buf ( n5417 , 1'b0 );
buf ( n5418 , n30343 );
buf ( n5419 , n23449 );
buf ( n5420 , 1'b0 );
buf ( n5421 , 1'b0 );
buf ( n5422 , n30353 );
buf ( n5423 , n20603 );
buf ( n5424 , 1'b0 );
buf ( n5425 , 1'b0 );
buf ( n5426 , n30376 );
buf ( n5427 , n20542 );
buf ( n5428 , 1'b0 );
buf ( n5429 , 1'b0 );
buf ( n5430 , n30376 );
buf ( n5431 , n21340 );
buf ( n5432 , 1'b0 );
buf ( n5433 , 1'b0 );
buf ( n5434 , n30376 );
buf ( n5435 , n20550 );
buf ( n5436 , 1'b0 );
buf ( n5437 , 1'b0 );
buf ( n5438 , n30345 );
buf ( n5439 , n20558 );
buf ( n5440 , 1'b0 );
buf ( n5441 , 1'b0 );
buf ( n5442 , n30376 );
buf ( n5443 , n29591 );
buf ( n5444 , 1'b0 );
buf ( n5445 , 1'b0 );
buf ( n5446 , n30378 );
buf ( n5447 , n29431 );
buf ( n5448 , 1'b0 );
buf ( n5449 , 1'b0 );
buf ( n5450 , n30378 );
buf ( n5451 , n29470 );
buf ( n5452 , 1'b0 );
buf ( n5453 , 1'b0 );
buf ( n5454 , n30376 );
buf ( n5455 , n1142 );
buf ( n5456 , 1'b0 );
buf ( n5457 , 1'b0 );
buf ( n5458 , n30376 );
buf ( n5459 , n1131 );
buf ( n5460 , 1'b0 );
buf ( n5461 , 1'b0 );
buf ( n5462 , n30353 );
buf ( n5463 , n1132 );
buf ( n5464 , 1'b0 );
buf ( n5465 , 1'b0 );
buf ( n5466 , n30374 );
buf ( n5467 , n1137 );
buf ( n5468 , 1'b0 );
buf ( n5469 , 1'b0 );
buf ( n5470 , n30376 );
buf ( n5471 , n1138 );
buf ( n5472 , 1'b0 );
buf ( n5473 , 1'b0 );
buf ( n5474 , n30356 );
buf ( n5475 , n1139 );
buf ( n5476 , 1'b0 );
buf ( n5477 , 1'b0 );
buf ( n5478 , n30374 );
buf ( n5479 , n21696 );
buf ( n5480 , 1'b0 );
buf ( n5481 , 1'b0 );
buf ( n5482 , n30374 );
buf ( n5483 , n21301 );
buf ( n5484 , 1'b0 );
buf ( n5485 , 1'b0 );
buf ( n5486 , n30343 );
buf ( n5487 , n21309 );
buf ( n5488 , 1'b0 );
buf ( n5489 , 1'b0 );
buf ( n5490 , n30343 );
buf ( n5491 , n20567 );
buf ( n5492 , 1'b0 );
buf ( n5493 , 1'b0 );
buf ( n5494 , n30353 );
buf ( n5495 , n1103 );
buf ( n5496 , 1'b0 );
buf ( n5497 , 1'b0 );
buf ( n5498 , n30374 );
buf ( n5499 , n1140 );
buf ( n5500 , 1'b0 );
buf ( n5501 , 1'b0 );
buf ( n5502 , n30343 );
buf ( n5503 , n29382 );
buf ( n5504 , 1'b0 );
buf ( n5505 , 1'b0 );
buf ( n5506 , n30343 );
buf ( n5507 , n23088 );
buf ( n5508 , 1'b0 );
buf ( n5509 , 1'b0 );
buf ( n5510 , n30374 );
buf ( n5511 , n21315 );
buf ( n5512 , 1'b0 );
buf ( n5513 , 1'b0 );
buf ( n5514 , n30345 );
buf ( n5515 , n21323 );
buf ( n5516 , 1'b0 );
buf ( n5517 , 1'b0 );
buf ( n5518 , n30353 );
buf ( n5519 , n21331 );
buf ( n5520 , 1'b0 );
buf ( n5521 , 1'b0 );
buf ( n5522 , n30351 );
buf ( n5523 , n18794 );
buf ( n5524 , 1'b0 );
buf ( n5525 , 1'b0 );
buf ( n5526 , n1 );
buf ( n5527 , n30077 );
buf ( n5528 , 1'b0 );
buf ( n5529 , 1'b0 );
buf ( n5530 , n1 );
buf ( n5531 , n26691 );
buf ( n5532 , 1'b0 );
buf ( n5533 , 1'b0 );
buf ( n5534 , n30374 );
buf ( n5535 , n18789 );
buf ( n5536 , 1'b0 );
buf ( n5537 , 1'b0 );
buf ( n5538 , n1 );
buf ( n5539 , n26644 );
buf ( n5540 , 1'b0 );
buf ( n5541 , 1'b0 );
buf ( n5542 , n1 );
buf ( n5543 , n26821 );
buf ( n5544 , 1'b0 );
buf ( n5545 , 1'b0 );
buf ( n5546 , n30374 );
buf ( n5547 , n18701 );
buf ( n5548 , 1'b0 );
buf ( n5549 , 1'b0 );
buf ( n5550 , n1 );
buf ( n5551 , n30260 );
buf ( n5552 , 1'b0 );
buf ( n5553 , 1'b0 );
buf ( n5554 , n30351 );
buf ( n5555 , n18704 );
buf ( n5556 , 1'b0 );
buf ( n5557 , 1'b0 );
buf ( n5558 , n30376 );
buf ( n5559 , n18708 );
buf ( n5560 , 1'b0 );
buf ( n5561 , 1'b0 );
buf ( n5562 , n30358 );
buf ( n5563 , n24368 );
buf ( n5564 , 1'b0 );
buf ( n5565 , 1'b0 );
buf ( n5566 , n30358 );
buf ( n5567 , n24371 );
buf ( n5568 , 1'b0 );
buf ( n5569 , 1'b0 );
buf ( n5570 , n1 );
buf ( n5571 , n17841 );
buf ( n5572 , 1'b0 );
buf ( n5573 , 1'b0 );
buf ( n5574 , n30376 );
buf ( n5575 , n21688 );
buf ( n5576 , 1'b0 );
buf ( n5577 , 1'b0 );
buf ( n5578 , n30376 );
buf ( n5579 , n1126 );
buf ( n5580 , 1'b0 );
buf ( n5581 , 1'b0 );
buf ( n5582 , n30356 );
buf ( n5583 , n27476 );
buf ( n5584 , 1'b0 );
buf ( n5585 , 1'b0 );
buf ( n5586 , n30371 );
buf ( n5587 , n26190 );
buf ( n5588 , 1'b0 );
buf ( n5589 , 1'b0 );
buf ( n5590 , n30376 );
buf ( n5591 , n27513 );
buf ( n5592 , 1'b0 );
buf ( n5593 , 1'b0 );
buf ( n5594 , n30376 );
buf ( n5595 , n27378 );
buf ( n5596 , 1'b0 );
buf ( n5597 , 1'b0 );
buf ( n5598 , n30356 );
buf ( n5599 , n21665 );
buf ( n5600 , 1'b0 );
buf ( n5601 , 1'b0 );
buf ( n5602 , n1 );
buf ( n5603 , n29987 );
buf ( n5604 , 1'b0 );
buf ( n5605 , 1'b0 );
buf ( n5606 , n1 );
buf ( n5607 , n30053 );
buf ( n5608 , 1'b0 );
buf ( n5609 , 1'b0 );
buf ( n5610 , n30371 );
buf ( n5611 , n24374 );
buf ( n5612 , 1'b0 );
buf ( n5613 , 1'b0 );
buf ( n5614 , n30343 );
buf ( n5615 , n24377 );
buf ( n5616 , 1'b0 );
buf ( n5617 , 1'b0 );
buf ( n5618 , n1 );
buf ( n5619 , n30089 );
buf ( n5620 , 1'b0 );
buf ( n5621 , 1'b0 );
buf ( n5622 , n1 );
buf ( n5623 , n30196 );
buf ( n5624 , 1'b0 );
buf ( n5625 , 1'b0 );
buf ( n5626 , n1 );
buf ( n5627 , n30184 );
buf ( n5628 , 1'b0 );
buf ( n5629 , 1'b0 );
buf ( n5630 , n1 );
buf ( n5631 , n30302 );
buf ( n5632 , 1'b0 );
buf ( n5633 , 1'b0 );
buf ( n5634 , n1 );
buf ( n5635 , n30144 );
buf ( n5636 , 1'b0 );
buf ( n5637 , 1'b0 );
buf ( n5638 , n1 );
buf ( n5639 , n30148 );
buf ( n5640 , 1'b0 );
buf ( n5641 , 1'b0 );
buf ( n5642 , n1 );
buf ( n5643 , n30049 );
buf ( n5644 , 1'b0 );
buf ( n5645 , 1'b0 );
buf ( n5646 , n1 );
buf ( n5647 , n30107 );
buf ( n5648 , 1'b0 );
buf ( n5649 , 1'b0 );
buf ( n5650 , n1 );
buf ( n5651 , n30156 );
buf ( n5652 , 1'b0 );
buf ( n5653 , 1'b0 );
buf ( n5654 , n1 );
buf ( n5655 , n30256 );
buf ( n5656 , 1'b0 );
buf ( n5657 , 1'b0 );
buf ( n5658 , n1 );
buf ( n5659 , n29913 );
buf ( n5660 , 1'b0 );
buf ( n5661 , 1'b0 );
buf ( n5662 , n30352 );
buf ( n5663 , n21540 );
buf ( n5664 , 1'b0 );
buf ( n5665 , 1'b0 );
buf ( n5666 , n30351 );
buf ( n5667 , n18784 );
buf ( n5668 , 1'b0 );
buf ( n5669 , 1'b0 );
buf ( n5670 , n30351 );
buf ( n5671 , n18711 );
buf ( n5672 , 1'b0 );
buf ( n5673 , 1'b0 );
buf ( n5674 , n30352 );
buf ( n5675 , n20065 );
buf ( n5676 , 1'b0 );
buf ( n5677 , 1'b0 );
buf ( n5678 , n30352 );
buf ( n5679 , n18714 );
buf ( n5680 , 1'b0 );
buf ( n5681 , 1'b0 );
buf ( n5682 , n30371 );
buf ( n5683 , n20075 );
buf ( n5684 , 1'b0 );
buf ( n5685 , 1'b0 );
buf ( n5686 , n30343 );
buf ( n5687 , n18717 );
buf ( n5688 , 1'b0 );
buf ( n5689 , 1'b0 );
buf ( n5690 , n30346 );
buf ( n5691 , n18495 );
buf ( n5692 , 1'b0 );
buf ( n5693 , 1'b0 );
buf ( n5694 , n30375 );
buf ( n5695 , n18757 );
buf ( n5696 , 1'b0 );
buf ( n5697 , 1'b0 );
buf ( n5698 , n30342 );
buf ( n5699 , n18780 );
buf ( n5700 , 1'b0 );
buf ( n5701 , 1'b0 );
buf ( n5702 , n30342 );
buf ( n5703 , n18775 );
buf ( n5704 , 1'b0 );
buf ( n5705 , 1'b0 );
buf ( n5706 , n30342 );
buf ( n5707 , n18769 );
buf ( n5708 , 1'b0 );
buf ( n5709 , 1'b0 );
buf ( n5710 , n30375 );
buf ( n5711 , n18764 );
buf ( n5712 , 1'b0 );
buf ( n5713 , 1'b0 );
buf ( n5714 , n30352 );
buf ( n5715 , n19366 );
buf ( n5716 , 1'b0 );
buf ( n5717 , 1'b0 );
buf ( n5718 , n30352 );
buf ( n5719 , n19145 );
buf ( n5720 , 1'b0 );
buf ( n5721 , 1'b0 );
buf ( n5722 , n30342 );
buf ( n5723 , n19150 );
buf ( n5724 , 1'b0 );
buf ( n5725 , 1'b0 );
buf ( n5726 , n30342 );
buf ( n5727 , n19175 );
buf ( n5728 , 1'b0 );
buf ( n5729 , 1'b0 );
buf ( n5730 , n30346 );
buf ( n5731 , n19155 );
buf ( n5732 , 1'b0 );
buf ( n5733 , 1'b0 );
buf ( n5734 , n30346 );
buf ( n5735 , n19160 );
buf ( n5736 , 1'b0 );
buf ( n5737 , 1'b0 );
buf ( n5738 , n30351 );
buf ( n5739 , n19165 );
buf ( n5740 , 1'b0 );
buf ( n5741 , 1'b0 );
buf ( n5742 , n30351 );
buf ( n5743 , n19170 );
buf ( n5744 , 1'b0 );
buf ( n5745 , 1'b0 );
buf ( n5746 , n30353 );
buf ( n5747 , n26422 );
buf ( n5748 , 1'b0 );
buf ( n5749 , 1'b0 );
buf ( n5750 , n30371 );
buf ( n5751 , n29653 );
buf ( n5752 , 1'b0 );
buf ( n5753 , 1'b0 );
buf ( n5754 , n30352 );
buf ( n5755 , n29438 );
buf ( n5756 , 1'b0 );
buf ( n5757 , 1'b0 );
buf ( n5758 , n30356 );
buf ( n5759 , n1128 );
buf ( n5760 , 1'b0 );
buf ( n5761 , 1'b0 );
buf ( n5762 , n30342 );
buf ( n5763 , n29630 );
buf ( n5764 , 1'b0 );
buf ( n5765 , 1'b0 );
buf ( n5766 , n30342 );
buf ( n5767 , n29444 );
buf ( n5768 , 1'b0 );
buf ( n5769 , 1'b0 );
buf ( n5770 , n30378 );
buf ( n5771 , n19180 );
buf ( n5772 , 1'b0 );
buf ( n5773 , 1'b0 );
buf ( n5774 , n30356 );
buf ( n5775 , n19185 );
buf ( n5776 , 1'b0 );
buf ( n5777 , 1'b0 );
buf ( n5778 , n30375 );
buf ( n5779 , n1136 );
buf ( n5780 , 1'b0 );
buf ( n5781 , 1'b0 );
buf ( n5782 , n30375 );
buf ( n5783 , n1127 );
buf ( n5784 , 1'b0 );
buf ( n5785 , 1'b0 );
buf ( n5786 , n30351 );
buf ( n5787 , n16898 );
buf ( n5788 , 1'b0 );
buf ( n5789 , 1'b0 );
buf ( n5790 , n30351 );
buf ( n5791 , n16969 );
buf ( n5792 , 1'b0 );
buf ( n5793 , 1'b0 );
buf ( n5794 , n30352 );
buf ( n5795 , n17040 );
buf ( n5796 , 1'b0 );
buf ( n5797 , 1'b0 );
buf ( n5798 , n30342 );
buf ( n5799 , n17110 );
buf ( n5800 , 1'b0 );
buf ( n5801 , 1'b0 );
buf ( n5802 , n1 );
buf ( n5803 , n30278 );
buf ( n5804 , 1'b0 );
buf ( n5805 , 1'b0 );
buf ( n5806 , n1 );
buf ( n5807 , n30266 );
buf ( n5808 , 1'b0 );
buf ( n5809 , 1'b0 );
buf ( n5810 , n30351 );
buf ( n5811 , n30240 );
buf ( n5812 , 1'b0 );
buf ( n5813 , 1'b0 );
buf ( n5814 , n30352 );
buf ( n5815 , n21358 );
buf ( n5816 , 1'b0 );
buf ( n5817 , 1'b0 );
buf ( n5818 , n1 );
buf ( n5819 , n30172 );
buf ( n5820 , 1'b0 );
buf ( n5821 , 1'b0 );
buf ( n5822 , n1 );
buf ( n5823 , n30065 );
buf ( n5824 , 1'b0 );
buf ( n5825 , 1'b0 );
buf ( n5826 , n30353 );
buf ( n5827 , n20585 );
buf ( n5828 , 1'b0 );
buf ( n5829 , 1'b0 );
buf ( n5830 , n30353 );
buf ( n5831 , n20575 );
buf ( n5832 , 1'b0 );
buf ( n5833 , 1'b0 );
buf ( n5834 , n30346 );
buf ( n5835 , n20580 );
buf ( n5836 , 1'b0 );
buf ( n5837 , 1'b0 );
buf ( n5838 , n30346 );
buf ( n5839 , n21359 );
buf ( n5840 , 1'b0 );
buf ( n5841 , 1'b0 );
buf ( n5842 , n1 );
buf ( n5843 , n30101 );
buf ( n5844 , 1'b0 );
buf ( n5845 , 1'b0 );
buf ( n5846 , n1 );
buf ( n5847 , n30200 );
buf ( n5848 , 1'b0 );
buf ( n5849 , 1'b0 );
buf ( n5850 , n30352 );
buf ( n5851 , n20080 );
buf ( n5852 , 1'b0 );
buf ( n5853 , 1'b0 );
buf ( n5854 , n1 );
buf ( n5855 , n30212 );
buf ( n5856 , 1'b0 );
buf ( n5857 , 1'b0 );
buf ( n5858 , n30371 );
buf ( n5859 , n29916 );
buf ( n5860 , 1'b0 );
buf ( n5861 , 1'b0 );
buf ( n5862 , n30346 );
buf ( n5863 , n26205 );
buf ( n5864 , 1'b0 );
buf ( n5865 , 1'b0 );
buf ( n5866 , n30346 );
buf ( n5867 , n29417 );
buf ( n5868 , 1'b0 );
buf ( n5869 , 1'b0 );
buf ( n5870 , n30342 );
buf ( n5871 , n29411 );
buf ( n5872 , 1'b0 );
buf ( n5873 , 1'b0 );
buf ( n5874 , n30345 );
buf ( n5875 , n29450 );
buf ( n5876 , 1'b0 );
buf ( n5877 , 1'b0 );
buf ( n5878 , n30371 );
buf ( n5879 , n20590 );
buf ( n5880 , 1'b0 );
buf ( n5881 , 1'b0 );
buf ( n5882 , n30378 );
buf ( n5883 , n24397 );
buf ( n5884 , 1'b0 );
buf ( n5885 , 1'b0 );
buf ( n5886 , n1 );
buf ( n5887 , n30188 );
buf ( n5888 , 1'b0 );
buf ( n5889 , 1'b0 );
buf ( n5890 , n30342 );
buf ( n5891 , n29389 );
buf ( n5892 , 1'b0 );
buf ( n5893 , 1'b0 );
buf ( n5894 , n30342 );
buf ( n5895 , n20082 );
buf ( n5896 , 1'b0 );
buf ( n5897 , 1'b0 );
buf ( n5898 , n30378 );
buf ( n5899 , n26843 );
buf ( n5900 , 1'b0 );
buf ( n5901 , 1'b0 );
buf ( n5902 , n30342 );
buf ( n5903 , n27793 );
buf ( n5904 , 1'b0 );
buf ( n5905 , 1'b0 );
buf ( n5906 , n1 );
buf ( n5907 , n29953 );
buf ( n5908 , 1'b0 );
buf ( n5909 , 1'b0 );
buf ( n5910 , n30343 );
buf ( n5911 , n21621 );
buf ( n5912 , 1'b0 );
buf ( n5913 , 1'b0 );
buf ( n5914 , n30343 );
buf ( n5915 , n21378 );
buf ( n5916 , 1'b0 );
buf ( n5917 , 1'b0 );
buf ( n5918 , n30371 );
buf ( n5919 , n21397 );
buf ( n5920 , 1'b0 );
buf ( n5921 , 1'b0 );
buf ( n5922 , n30371 );
buf ( n5923 , n21417 );
buf ( n5924 , 1'b0 );
buf ( n5925 , 1'b0 );
buf ( n5926 , n30343 );
buf ( n5927 , n24428 );
buf ( n5928 , 1'b0 );
buf ( n5929 , 1'b0 );
buf ( n5930 , n30342 );
buf ( n5931 , n21457 );
buf ( n5932 , 1'b0 );
buf ( n5933 , 1'b0 );
buf ( n5934 , n30371 );
buf ( n5935 , n27971 );
buf ( n5936 , 1'b0 );
buf ( n5937 , 1'b0 );
buf ( n5938 , n30371 );
buf ( n5939 , n27526 );
buf ( n5940 , 1'b0 );
buf ( n5941 , 1'b0 );
buf ( n5942 , n1 );
buf ( n5943 , n29957 );
buf ( n5944 , 1'b0 );
buf ( n5945 , 1'b0 );
buf ( n5946 , n1 );
buf ( n5947 , n29961 );
buf ( n5948 , 1'b0 );
buf ( n5949 , 1'b0 );
buf ( n5950 , n1 );
buf ( n5951 , n30081 );
buf ( n5952 , 1'b0 );
buf ( n5953 , 1'b0 );
buf ( n5954 , n1 );
buf ( n5955 , n30333 );
buf ( n5956 , 1'b0 );
buf ( n5957 , 1'b0 );
buf ( n5958 , n30351 );
buf ( n5959 , n29964 );
buf ( n5960 , 1'b0 );
buf ( n5961 , 1'b0 );
buf ( n5962 , n30342 );
buf ( n5963 , n28286 );
buf ( n5964 , 1'b0 );
buf ( n5965 , 1'b0 );
buf ( n5966 , n30346 );
buf ( n5967 , n29647 );
buf ( n5968 , 1'b0 );
buf ( n5969 , 1'b0 );
buf ( n5970 , n30378 );
buf ( n5971 , n29457 );
buf ( n5972 , 1'b0 );
buf ( n5973 , 1'b0 );
buf ( n5974 , n30346 );
buf ( n5975 , n29641 );
buf ( n5976 , 1'b0 );
buf ( n5977 , 1'b0 );
buf ( n5978 , n30343 );
buf ( n5979 , n26848 );
buf ( n5980 , 1'b0 );
buf ( n5981 , 1'b0 );
buf ( n5982 , n30346 );
buf ( n5983 , n26849 );
buf ( n5984 , 1'b0 );
buf ( n5985 , 1'b0 );
buf ( n5986 , n30342 );
buf ( n5987 , n24440 );
buf ( n5988 , 1'b0 );
buf ( n5989 , 1'b0 );
buf ( n5990 , n30351 );
buf ( n5991 , n24445 );
buf ( n5992 , 1'b0 );
buf ( n5993 , 1'b0 );
buf ( n5994 , n30342 );
buf ( n5995 , n24450 );
buf ( n5996 , 1'b0 );
buf ( n5997 , 1'b0 );
buf ( n5998 , n30352 );
buf ( n5999 , n24455 );
buf ( n6000 , 1'b0 );
buf ( n6001 , 1'b0 );
buf ( n6002 , n30358 );
buf ( n6003 , n24460 );
buf ( n6004 , 1'b0 );
buf ( n6005 , 1'b0 );
buf ( n6006 , n30351 );
buf ( n6007 , n24465 );
buf ( n6008 , 1'b0 );
buf ( n6009 , 1'b0 );
buf ( n6010 , n30351 );
buf ( n6011 , n24471 );
buf ( n6012 , 1'b0 );
buf ( n6013 , 1'b0 );
buf ( n6014 , n30342 );
buf ( n6015 , n24476 );
buf ( n6016 , 1'b0 );
buf ( n6017 , 1'b0 );
buf ( n6018 , n30345 );
buf ( n6019 , n24481 );
buf ( n6020 , 1'b0 );
buf ( n6021 , 1'b0 );
buf ( n6022 , n30342 );
buf ( n6023 , n24486 );
buf ( n6024 , 1'b0 );
buf ( n6025 , 1'b0 );
buf ( n6026 , n30371 );
buf ( n6027 , n24491 );
buf ( n6028 , 1'b0 );
buf ( n6029 , 1'b0 );
buf ( n6030 , n30371 );
buf ( n6031 , n24496 );
buf ( n6032 , 1'b0 );
buf ( n6033 , 1'b0 );
buf ( n6034 , n30371 );
buf ( n6035 , n24501 );
buf ( n6036 , 1'b0 );
buf ( n6037 , 1'b0 );
buf ( n6038 , n30371 );
buf ( n6039 , n24512 );
buf ( n6040 , 1'b0 );
buf ( n6041 , 1'b0 );
buf ( n6042 , n30346 );
buf ( n6043 , n24517 );
buf ( n6044 , 1'b0 );
buf ( n6045 , 1'b0 );
buf ( n6046 , n30353 );
buf ( n6047 , n24522 );
buf ( n6048 , 1'b0 );
buf ( n6049 , 1'b0 );
buf ( n6050 , n30351 );
buf ( n6051 , n24527 );
buf ( n6052 , 1'b0 );
buf ( n6053 , 1'b0 );
buf ( n6054 , n30346 );
buf ( n6055 , n29464 );
buf ( n6056 , 1'b0 );
buf ( n6057 , 1'b0 );
buf ( n6058 , n1 );
buf ( n6059 , n29052 );
buf ( n6060 , 1'b0 );
buf ( n6061 , 1'b0 );
buf ( n6062 , n30375 );
buf ( n6063 , n26861 );
buf ( n6064 , 1'b0 );
buf ( n6065 , 1'b0 );
buf ( n6066 , n30343 );
buf ( n6067 , n24540 );
buf ( n6068 , 1'b0 );
buf ( n6069 , 1'b0 );
buf ( n6070 , n30371 );
buf ( n6071 , n27533 );
buf ( n6072 , 1'b0 );
buf ( n6073 , 1'b0 );
buf ( n6074 , n30353 );
buf ( n6075 , n26306 );
buf ( n6076 , 1'b0 );
buf ( n6077 , 1'b0 );
buf ( n6078 , n1 );
buf ( n6079 , n29035 );
buf ( n6080 , 1'b0 );
buf ( n6081 , 1'b0 );
buf ( n6082 , n30371 );
buf ( n6083 , n26870 );
buf ( n6084 , 1'b0 );
buf ( n6085 , 1'b0 );
buf ( n6086 , n30375 );
buf ( n6087 , n24546 );
buf ( n6088 , 1'b0 );
buf ( n6089 , 1'b0 );
buf ( n6090 , n30356 );
buf ( n6091 , n24551 );
buf ( n6092 , 1'b0 );
buf ( n6093 , 1'b0 );
buf ( n6094 , n30375 );
buf ( n6095 , n24557 );
buf ( n6096 , 1'b0 );
buf ( n6097 , 1'b0 );
buf ( n6098 , n30342 );
buf ( n6099 , n24562 );
buf ( n6100 , 1'b0 );
buf ( n6101 , 1'b0 );
buf ( n6102 , n30346 );
buf ( n6103 , n24354 );
buf ( n6104 , 1'b0 );
buf ( n6105 , 1'b0 );
buf ( n6106 , n30358 );
buf ( n6107 , n24567 );
buf ( n6108 , 1'b0 );
buf ( n6109 , 1'b0 );
buf ( n6110 , n30342 );
buf ( n6111 , n24572 );
buf ( n6112 , 1'b0 );
buf ( n6113 , 1'b0 );
buf ( n6114 , n30343 );
buf ( n6115 , n24577 );
buf ( n6116 , 1'b0 );
buf ( n6117 , 1'b0 );
buf ( n6118 , n30342 );
buf ( n6119 , n24364 );
buf ( n6120 , 1'b0 );
buf ( n6121 , 1'b0 );
buf ( n6122 , n30374 );
buf ( n6123 , n24582 );
buf ( n6124 , 1'b0 );
buf ( n6125 , 1'b0 );
buf ( n6126 , n30343 );
buf ( n6127 , n24588 );
buf ( n6128 , 1'b0 );
buf ( n6129 , 1'b0 );
buf ( n6130 , n30356 );
buf ( n6131 , n24593 );
buf ( n6132 , 1'b0 );
buf ( n6133 , 1'b0 );
buf ( n6134 , n30371 );
buf ( n6135 , n23588 );
buf ( n6136 , 1'b0 );
buf ( n6137 , 1'b0 );
buf ( n6138 , n30355 );
buf ( n6139 , n28289 );
buf ( n6140 , 1'b0 );
buf ( n6141 , 1'b0 );
buf ( n6142 , n30356 );
buf ( n6143 , n23090 );
buf ( n6144 , 1'b0 );
buf ( n6145 , 1'b0 );
buf ( n6146 , n30343 );
buf ( n6147 , n28283 );
buf ( n6148 , 1'b0 );
buf ( n6149 , 1'b0 );
buf ( n6150 , n30355 );
buf ( n6151 , n27808 );
buf ( n6152 , 1'b0 );
buf ( n6153 , 1'b0 );
buf ( n6154 , n30345 );
buf ( n6155 , n24598 );
buf ( n6156 , 1'b0 );
buf ( n6157 , 1'b0 );
buf ( n6158 , n30374 );
buf ( n6159 , n24603 );
buf ( n6160 , 1'b0 );
buf ( n6161 , 1'b0 );
buf ( n6162 , n30353 );
buf ( n6163 , n24608 );
buf ( n6164 , 1'b0 );
buf ( n6165 , 1'b0 );
buf ( n6166 , n30374 );
buf ( n6167 , n24613 );
buf ( n6168 , 1'b0 );
buf ( n6169 , 1'b0 );
buf ( n6170 , n30353 );
buf ( n6171 , n24618 );
buf ( n6172 , 1'b0 );
buf ( n6173 , 1'b0 );
buf ( n6174 , n30374 );
buf ( n6175 , n24623 );
buf ( n6176 , 1'b0 );
buf ( n6177 , 1'b0 );
buf ( n6178 , n30371 );
buf ( n6179 , n28294 );
buf ( n6180 , 1'b0 );
buf ( n6181 , 1'b0 );
buf ( n6182 , n30378 );
buf ( n6183 , n27541 );
buf ( n6184 , 1'b0 );
buf ( n6185 , 1'b0 );
buf ( n6186 , n30356 );
buf ( n6187 , n26871 );
buf ( n6188 , 1'b0 );
buf ( n6189 , 1'b0 );
buf ( n6190 , n30374 );
buf ( n6191 , n29919 );
buf ( n6192 , 1'b0 );
buf ( n6193 , 1'b0 );
buf ( n6194 , n30343 );
buf ( n6195 , n24628 );
buf ( n6196 , 1'b0 );
buf ( n6197 , 1'b0 );
buf ( n6198 , n30356 );
buf ( n6199 , n25227 );
buf ( n6200 , 1'b0 );
buf ( n6201 , 1'b0 );
buf ( n6202 , n30372 );
buf ( n6203 , n24633 );
buf ( n6204 , 1'b0 );
buf ( n6205 , 1'b0 );
buf ( n6206 , n30376 );
buf ( n6207 , n24639 );
buf ( n6208 , 1'b0 );
buf ( n6209 , 1'b0 );
buf ( n6210 , n30374 );
buf ( n6211 , n23578 );
buf ( n6212 , 1'b0 );
buf ( n6213 , 1'b0 );
buf ( n6214 , n30345 );
buf ( n6215 , n24644 );
buf ( n6216 , 1'b0 );
buf ( n6217 , 1'b0 );
buf ( n6218 , n30345 );
buf ( n6219 , n24646 );
buf ( n6220 , 1'b0 );
buf ( n6221 , 1'b0 );
buf ( n6222 , n30374 );
buf ( n6223 , n23092 );
buf ( n6224 , 1'b0 );
buf ( n6225 , 1'b0 );
buf ( n6226 , n30353 );
buf ( n6227 , n23094 );
buf ( n6228 , 1'b0 );
buf ( n6229 , 1'b0 );
buf ( n6230 , n30355 );
buf ( n6231 , n29018 );
buf ( n6232 , 1'b0 );
buf ( n6233 , 1'b0 );
buf ( n6234 , n1 );
buf ( n6235 , n26909 );
buf ( n6236 , 1'b0 );
buf ( n6237 , 1'b0 );
buf ( n6238 , n1 );
buf ( n6239 , n26941 );
buf ( n6240 , 1'b0 );
buf ( n6241 , 1'b0 );
buf ( n6242 , n1 );
buf ( n6243 , n26974 );
buf ( n6244 , 1'b0 );
buf ( n6245 , 1'b0 );
buf ( n6246 , n30353 );
buf ( n6247 , n24649 );
buf ( n6248 , 1'b0 );
buf ( n6249 , 1'b0 );
buf ( n6250 , n30355 );
buf ( n6251 , n24651 );
buf ( n6252 , 1'b0 );
buf ( n6253 , 1'b0 );
buf ( n6254 , n30355 );
buf ( n6255 , n24654 );
buf ( n6256 , 1'b0 );
buf ( n6257 , 1'b0 );
buf ( n6258 , n30353 );
buf ( n6259 , n24657 );
buf ( n6260 , 1'b0 );
buf ( n6261 , 1'b0 );
buf ( n6262 , n30345 );
buf ( n6263 , n23096 );
buf ( n6264 , 1'b0 );
buf ( n6265 , 1'b0 );
buf ( n6266 , n30345 );
buf ( n6267 , n24659 );
buf ( n6268 , 1'b0 );
buf ( n6269 , 1'b0 );
buf ( n6270 , n1 );
buf ( n6271 , n24664 );
buf ( n6272 , 1'b0 );
buf ( n6273 , 1'b0 );
buf ( n6274 , n1 );
buf ( n6275 , n23534 );
buf ( n6276 , 1'b0 );
buf ( n6277 , 1'b0 );
buf ( n6278 , n30355 );
buf ( n6279 , n24670 );
buf ( n6280 , 1'b0 );
buf ( n6281 , 1'b0 );
buf ( n6282 , n30352 );
buf ( n6283 , n24672 );
buf ( n6284 , 1'b0 );
buf ( n6285 , 1'b0 );
buf ( n6286 , n1 );
buf ( n6287 , n27331 );
buf ( n6288 , 1'b0 );
buf ( n6289 , 1'b0 );
buf ( n6290 , n30376 );
buf ( n6291 , n24675 );
buf ( n6292 , 1'b0 );
buf ( n6293 , 1'b0 );
buf ( n6294 , n30355 );
buf ( n6295 , n24680 );
buf ( n6296 , 1'b0 );
buf ( n6297 , 1'b0 );
buf ( n6298 , n30358 );
buf ( n6299 , n24682 );
buf ( n6300 , 1'b0 );
buf ( n6301 , 1'b0 );
buf ( n6302 , n30345 );
buf ( n6303 , n24687 );
buf ( n6304 , 1'b0 );
buf ( n6305 , 1'b0 );
buf ( n6306 , n30345 );
buf ( n6307 , n23098 );
buf ( n6308 , 1'b0 );
buf ( n6309 , 1'b0 );
buf ( n6310 , n30374 );
buf ( n6311 , n24692 );
buf ( n6312 , 1'b0 );
buf ( n6313 , 1'b0 );
buf ( n6314 , n30372 );
buf ( n6315 , n28951 );
buf ( n6316 , 1'b0 );
buf ( n6317 , 1'b0 );
buf ( n6318 , n30374 );
buf ( n6319 , n24703 );
buf ( n6320 , 1'b0 );
buf ( n6321 , 1'b0 );
buf ( n6322 , n30375 );
buf ( n6323 , n24698 );
buf ( n6324 , 1'b0 );
buf ( n6325 , 1'b0 );
buf ( n6326 , n30347 );
buf ( n6327 , n23100 );
buf ( n6328 , 1'b0 );
buf ( n6329 , 1'b0 );
buf ( n6330 , n30358 );
buf ( n6331 , n24708 );
buf ( n6332 , 1'b0 );
buf ( n6333 , 1'b0 );
buf ( n6334 , n30340 );
buf ( n6335 , n24713 );
buf ( n6336 , 1'b0 );
buf ( n6337 , 1'b0 );
buf ( n6338 , n30340 );
buf ( n6339 , n25215 );
buf ( n6340 , 1'b0 );
buf ( n6341 , 1'b0 );
buf ( n6342 , n30340 );
buf ( n6343 , n24715 );
buf ( n6344 , 1'b0 );
buf ( n6345 , 1'b0 );
buf ( n6346 , n30347 );
buf ( n6347 , n23102 );
buf ( n6348 , 1'b0 );
buf ( n6349 , 1'b0 );
buf ( n6350 , n30340 );
buf ( n6351 , n27820 );
buf ( n6352 , 1'b0 );
buf ( n6353 , 1'b0 );
buf ( n6354 , n30372 );
buf ( n6355 , n23104 );
buf ( n6356 , 1'b0 );
buf ( n6357 , 1'b0 );
buf ( n6358 , n30355 );
buf ( n6359 , n26362 );
buf ( n6360 , 1'b0 );
buf ( n6361 , 1'b0 );
buf ( n6362 , n30355 );
buf ( n6363 , n26370 );
buf ( n6364 , 1'b0 );
buf ( n6365 , 1'b0 );
buf ( n6366 , n30357 );
buf ( n6367 , n24720 );
buf ( n6368 , 1'b0 );
buf ( n6369 , 1'b0 );
buf ( n6370 , n30340 );
buf ( n6371 , n24722 );
buf ( n6372 , 1'b0 );
buf ( n6373 , 1'b0 );
buf ( n6374 , n1 );
buf ( n6375 , n24727 );
buf ( n6376 , 1'b0 );
buf ( n6377 , 1'b0 );
buf ( n6378 , n1 );
buf ( n6379 , n24732 );
buf ( n6380 , 1'b0 );
buf ( n6381 , 1'b0 );
buf ( n6382 , n1 );
buf ( n6383 , n25213 );
buf ( n6384 , 1'b0 );
buf ( n6385 , 1'b0 );
buf ( n6386 , n1 );
buf ( n6387 , n24737 );
buf ( n6388 , 1'b0 );
buf ( n6389 , 1'b0 );
buf ( n6390 , n1 );
buf ( n6391 , n24742 );
buf ( n6392 , 1'b0 );
buf ( n6393 , 1'b0 );
buf ( n6394 , n30357 );
buf ( n6395 , n27004 );
buf ( n6396 , 1'b0 );
buf ( n6397 , 1'b0 );
buf ( n6398 , n30357 );
buf ( n6399 , n24747 );
buf ( n6400 , 1'b0 );
buf ( n6401 , 1'b0 );
buf ( n6402 , n30378 );
buf ( n6403 , n15230 );
buf ( n6404 , 1'b0 );
buf ( n6405 , 1'b0 );
buf ( n6406 , n30378 );
buf ( n6407 , n24752 );
buf ( n6408 , 1'b0 );
buf ( n6409 , 1'b0 );
buf ( n6410 , n30375 );
buf ( n6411 , n25208 );
buf ( n6412 , 1'b0 );
buf ( n6413 , 1'b0 );
buf ( n6414 , n30378 );
buf ( n6415 , n24758 );
buf ( n6416 , 1'b0 );
buf ( n6417 , 1'b0 );
buf ( n6418 , n30340 );
buf ( n6419 , n24763 );
buf ( n6420 , 1'b0 );
buf ( n6421 , 1'b0 );
buf ( n6422 , n30357 );
buf ( n6423 , n24768 );
buf ( n6424 , 1'b0 );
buf ( n6425 , 1'b0 );
buf ( n6426 , n30357 );
buf ( n6427 , n25203 );
buf ( n6428 , 1'b0 );
buf ( n6429 , 1'b0 );
buf ( n6430 , n30357 );
buf ( n6431 , n24774 );
buf ( n6432 , 1'b0 );
buf ( n6433 , 1'b0 );
buf ( n6434 , n30349 );
buf ( n6435 , n24779 );
buf ( n6436 , 1'b0 );
buf ( n6437 , 1'b0 );
buf ( n6438 , n30349 );
buf ( n6439 , n24784 );
buf ( n6440 , 1'b0 );
buf ( n6441 , 1'b0 );
buf ( n6442 , n30347 );
buf ( n6443 , n25193 );
buf ( n6444 , 1'b0 );
buf ( n6445 , 1'b0 );
buf ( n6446 , n30349 );
buf ( n6447 , n24789 );
buf ( n6448 , 1'b0 );
buf ( n6449 , 1'b0 );
buf ( n6450 , n30348 );
buf ( n6451 , n24794 );
buf ( n6452 , 1'b0 );
buf ( n6453 , 1'b0 );
buf ( n6454 , n30348 );
buf ( n6455 , n24799 );
buf ( n6456 , 1'b0 );
buf ( n6457 , 1'b0 );
buf ( n6458 , n30340 );
buf ( n6459 , n25198 );
buf ( n6460 , 1'b0 );
buf ( n6461 , 1'b0 );
buf ( n6462 , n30357 );
buf ( n6463 , n24804 );
buf ( n6464 , 1'b0 );
buf ( n6465 , 1'b0 );
buf ( n6466 , n30340 );
buf ( n6467 , n24809 );
buf ( n6468 , 1'b0 );
buf ( n6469 , 1'b0 );
buf ( n6470 , n30347 );
buf ( n6471 , n24814 );
buf ( n6472 , 1'b0 );
buf ( n6473 , 1'b0 );
buf ( n6474 , n30347 );
buf ( n6475 , n25188 );
buf ( n6476 , 1'b0 );
buf ( n6477 , 1'b0 );
buf ( n6478 , n30347 );
buf ( n6479 , n24533 );
buf ( n6480 , 1'b0 );
buf ( n6481 , 1'b0 );
buf ( n6482 , n30348 );
buf ( n6483 , n24507 );
buf ( n6484 , 1'b0 );
buf ( n6485 , 1'b0 );
buf ( n6486 , n30373 );
buf ( n6487 , n24433 );
buf ( n6488 , 1'b0 );
buf ( n6489 , 1'b0 );
buf ( n6490 , n30377 );
buf ( n6491 , n25158 );
buf ( n6492 , 1'b0 );
buf ( n6493 , 1'b0 );
buf ( n6494 , n30377 );
buf ( n6495 , n24383 );
buf ( n6496 , 1'b0 );
buf ( n6497 , 1'b0 );
buf ( n6498 , n30340 );
buf ( n6499 , n25173 );
buf ( n6500 , 1'b0 );
buf ( n6501 , 1'b0 );
buf ( n6502 , n30340 );
buf ( n6503 , n24359 );
buf ( n6504 , 1'b0 );
buf ( n6505 , 1'b0 );
buf ( n6506 , n30373 );
buf ( n6507 , n25183 );
buf ( n6508 , 1'b0 );
buf ( n6509 , 1'b0 );
buf ( n6510 , n30340 );
buf ( n6511 , n24257 );
buf ( n6512 , 1'b0 );
buf ( n6513 , 1'b0 );
buf ( n6514 , n30340 );
buf ( n6515 , n24252 );
buf ( n6516 , 1'b0 );
buf ( n6517 , 1'b0 );
buf ( n6518 , n30340 );
buf ( n6519 , n24218 );
buf ( n6520 , 1'b0 );
buf ( n6521 , 1'b0 );
buf ( n6522 , n30354 );
buf ( n6523 , n25168 );
buf ( n6524 , 1'b0 );
buf ( n6525 , 1'b0 );
buf ( n6526 , n30377 );
buf ( n6527 , n24190 );
buf ( n6528 , 1'b0 );
buf ( n6529 , 1'b0 );
buf ( n6530 , n30357 );
buf ( n6531 , n23575 );
buf ( n6532 , 1'b0 );
buf ( n6533 , 1'b0 );
buf ( n6534 , n30354 );
buf ( n6535 , n23569 );
buf ( n6536 , 1'b0 );
buf ( n6537 , 1'b0 );
buf ( n6538 , n30373 );
buf ( n6539 , n25178 );
buf ( n6540 , 1'b0 );
buf ( n6541 , 1'b0 );
buf ( n6542 , n30373 );
buf ( n6543 , n23563 );
buf ( n6544 , 1'b0 );
buf ( n6545 , 1'b0 );
buf ( n6546 , n30349 );
buf ( n6547 , n23557 );
buf ( n6548 , 1'b0 );
buf ( n6549 , 1'b0 );
buf ( n6550 , n30349 );
buf ( n6551 , n23551 );
buf ( n6552 , 1'b0 );
buf ( n6553 , 1'b0 );
buf ( n6554 , n30348 );
buf ( n6555 , n25153 );
buf ( n6556 , 1'b0 );
buf ( n6557 , 1'b0 );
buf ( n6558 , n30348 );
buf ( n6559 , n23545 );
buf ( n6560 , 1'b0 );
buf ( n6561 , 1'b0 );
buf ( n6562 , n30348 );
buf ( n6563 , n23540 );
buf ( n6564 , 1'b0 );
buf ( n6565 , 1'b0 );
buf ( n6566 , n30373 );
buf ( n6567 , n23521 );
buf ( n6568 , 1'b0 );
buf ( n6569 , 1'b0 );
buf ( n6570 , n30377 );
buf ( n6571 , n25148 );
buf ( n6572 , 1'b0 );
buf ( n6573 , 1'b0 );
buf ( n6574 , n30377 );
buf ( n6575 , n23515 );
buf ( n6576 , 1'b0 );
buf ( n6577 , 1'b0 );
buf ( n6578 , n30354 );
buf ( n6579 , n24838 );
buf ( n6580 , 1'b0 );
buf ( n6581 , 1'b0 );
buf ( n6582 , n30373 );
buf ( n6583 , n24819 );
buf ( n6584 , 1'b0 );
buf ( n6585 , 1'b0 );
buf ( n6586 , n30354 );
buf ( n6587 , n25143 );
buf ( n6588 , 1'b0 );
buf ( n6589 , 1'b0 );
buf ( n6590 , n30354 );
buf ( n6591 , n24824 );
buf ( n6592 , 1'b0 );
buf ( n6593 , 1'b0 );
buf ( n6594 , n30377 );
buf ( n6595 , n24827 );
buf ( n6596 , 1'b0 );
buf ( n6597 , 1'b0 );
buf ( n6598 , n30377 );
buf ( n6599 , n24829 );
buf ( n6600 , 1'b0 );
buf ( n6601 , 1'b0 );
buf ( n6602 , n30349 );
buf ( n6603 , n24831 );
buf ( n6604 , 1'b0 );
buf ( n6605 , 1'b0 );
buf ( n6606 , n30377 );
buf ( n6607 , n24833 );
buf ( n6608 , 1'b0 );
buf ( n6609 , 1'b0 );
buf ( n6610 , n30357 );
buf ( n6611 , n24841 );
buf ( n6612 , 1'b0 );
buf ( n6613 , 1'b0 );
buf ( n6614 , n30372 );
buf ( n6615 , n23107 );
buf ( n6616 , 1'b0 );
buf ( n6617 , 1'b0 );
buf ( n6618 , n30340 );
buf ( n6619 , n23109 );
buf ( n6620 , 1'b0 );
buf ( n6621 , 1'b0 );
buf ( n6622 , n30340 );
buf ( n6623 , n23111 );
buf ( n6624 , 1'b0 );
buf ( n6625 , 1'b0 );
buf ( n6626 , n30373 );
buf ( n6627 , n24843 );
buf ( n6628 , 1'b0 );
buf ( n6629 , 1'b0 );
buf ( n6630 , n30373 );
buf ( n6631 , n23114 );
buf ( n6632 , 1'b0 );
buf ( n6633 , 1'b0 );
buf ( n6634 , n30349 );
buf ( n6635 , n24845 );
buf ( n6636 , 1'b0 );
buf ( n6637 , 1'b0 );
buf ( n6638 , n30373 );
buf ( n6639 , n24847 );
buf ( n6640 , 1'b0 );
buf ( n6641 , 1'b0 );
buf ( n6642 , n30354 );
buf ( n6643 , n24850 );
buf ( n6644 , 1'b0 );
buf ( n6645 , 1'b0 );
buf ( n6646 , n30354 );
buf ( n6647 , n24853 );
buf ( n6648 , 1'b0 );
buf ( n6649 , 1'b0 );
buf ( n6650 , n30372 );
buf ( n6651 , n24855 );
buf ( n6652 , 1'b0 );
buf ( n6653 , 1'b0 );
buf ( n6654 , n30354 );
buf ( n6655 , n23137 );
buf ( n6656 , 1'b0 );
buf ( n6657 , 1'b0 );
buf ( n6658 , n30377 );
buf ( n6659 , n28001 );
buf ( n6660 , 1'b0 );
buf ( n6661 , 1'b0 );
buf ( n6662 , n30354 );
buf ( n6663 , n24857 );
buf ( n6664 , 1'b0 );
buf ( n6665 , 1'b0 );
buf ( n6666 , n30377 );
buf ( n6667 , n24859 );
buf ( n6668 , 1'b0 );
buf ( n6669 , 1'b0 );
buf ( n6670 , n30377 );
buf ( n6671 , n24862 );
buf ( n6672 , 1'b0 );
buf ( n6673 , 1'b0 );
buf ( n6674 , n30349 );
buf ( n6675 , n23140 );
buf ( n6676 , 1'b0 );
buf ( n6677 , 1'b0 );
buf ( n6678 , n30349 );
buf ( n6679 , n24864 );
buf ( n6680 , 1'b0 );
buf ( n6681 , 1'b0 );
buf ( n6682 , n30372 );
buf ( n6683 , n24866 );
buf ( n6684 , 1'b0 );
buf ( n6685 , 1'b0 );
buf ( n6686 , n30349 );
buf ( n6687 , n24870 );
buf ( n6688 , 1'b0 );
buf ( n6689 , 1'b0 );
buf ( n6690 , n30372 );
buf ( n6691 , n24868 );
buf ( n6692 , 1'b0 );
buf ( n6693 , 1'b0 );
buf ( n6694 , n30377 );
buf ( n6695 , n23142 );
buf ( n6696 , 1'b0 );
buf ( n6697 , 1'b0 );
buf ( n6698 , n30372 );
buf ( n6699 , n23145 );
buf ( n6700 , 1'b0 );
buf ( n6701 , 1'b0 );
buf ( n6702 , n30349 );
buf ( n6703 , n23147 );
buf ( n6704 , 1'b0 );
buf ( n6705 , 1'b0 );
buf ( n6706 , n30372 );
buf ( n6707 , n23150 );
buf ( n6708 , 1'b0 );
buf ( n6709 , 1'b0 );
buf ( n6710 , n30372 );
buf ( n6711 , n24873 );
buf ( n6712 , 1'b0 );
buf ( n6713 , 1'b0 );
buf ( n6714 , n30377 );
buf ( n6715 , n23152 );
buf ( n6716 , 1'b0 );
buf ( n6717 , 1'b0 );
buf ( n6718 , n30373 );
buf ( n6719 , n24875 );
buf ( n6720 , 1'b0 );
buf ( n6721 , 1'b0 );
buf ( n6722 , n30354 );
buf ( n6723 , n24879 );
buf ( n6724 , 1'b0 );
buf ( n6725 , 1'b0 );
buf ( n6726 , n30349 );
buf ( n6727 , n24877 );
buf ( n6728 , 1'b0 );
buf ( n6729 , 1'b0 );
buf ( n6730 , n30377 );
buf ( n6731 , n24881 );
buf ( n6732 , 1'b0 );
buf ( n6733 , 1'b0 );
buf ( n6734 , n30372 );
buf ( n6735 , n23165 );
buf ( n6736 , 1'b0 );
buf ( n6737 , 1'b0 );
buf ( n6738 , n30354 );
buf ( n6739 , n23168 );
buf ( n6740 , 1'b0 );
buf ( n6741 , 1'b0 );
buf ( n6742 , n30349 );
buf ( n6743 , n24883 );
buf ( n6744 , 1'b0 );
buf ( n6745 , 1'b0 );
buf ( n6746 , n30348 );
buf ( n6747 , n24886 );
buf ( n6748 , 1'b0 );
buf ( n6749 , 1'b0 );
buf ( n6750 , n30349 );
buf ( n6751 , n24888 );
buf ( n6752 , 1'b0 );
buf ( n6753 , 1'b0 );
buf ( n6754 , n30373 );
buf ( n6755 , n24892 );
buf ( n6756 , 1'b0 );
buf ( n6757 , 1'b0 );
buf ( n6758 , n30354 );
buf ( n6759 , n24890 );
buf ( n6760 , 1'b0 );
buf ( n6761 , 1'b0 );
buf ( n6762 , n30348 );
buf ( n6763 , n24895 );
buf ( n6764 , 1'b0 );
buf ( n6765 , 1'b0 );
buf ( n6766 , n30373 );
buf ( n6767 , n23170 );
buf ( n6768 , 1'b0 );
buf ( n6769 , 1'b0 );
buf ( n6770 , n30349 );
buf ( n6771 , n24897 );
buf ( n6772 , 1'b0 );
buf ( n6773 , 1'b0 );
buf ( n6774 , n30377 );
buf ( n6775 , n23172 );
buf ( n6776 , 1'b0 );
buf ( n6777 , 1'b0 );
buf ( n6778 , n30349 );
buf ( n6779 , n23174 );
buf ( n6780 , 1'b0 );
buf ( n6781 , 1'b0 );
buf ( n6782 , n30357 );
buf ( n6783 , n23176 );
buf ( n6784 , 1'b0 );
buf ( n6785 , 1'b0 );
buf ( n6786 , n30377 );
buf ( n6787 , n23178 );
buf ( n6788 , 1'b0 );
buf ( n6789 , 1'b0 );
buf ( n6790 , n30373 );
buf ( n6791 , n23181 );
buf ( n6792 , 1'b0 );
buf ( n6793 , 1'b0 );
buf ( n6794 , n30373 );
buf ( n6795 , n23184 );
buf ( n6796 , 1'b0 );
buf ( n6797 , 1'b0 );
buf ( n6798 , n30377 );
buf ( n6799 , n24899 );
buf ( n6800 , 1'b0 );
buf ( n6801 , 1'b0 );
buf ( n6802 , n30354 );
buf ( n6803 , n23186 );
buf ( n6804 , 1'b0 );
buf ( n6805 , 1'b0 );
buf ( n6806 , n30354 );
buf ( n6807 , n24901 );
buf ( n6808 , 1'b0 );
buf ( n6809 , 1'b0 );
buf ( n6810 , n30349 );
buf ( n6811 , n24903 );
buf ( n6812 , 1'b0 );
buf ( n6813 , 1'b0 );
buf ( n6814 , n30347 );
buf ( n6815 , n24905 );
buf ( n6816 , 1'b0 );
buf ( n6817 , 1'b0 );
buf ( n6818 , n30348 );
buf ( n6819 , n24907 );
buf ( n6820 , 1'b0 );
buf ( n6821 , 1'b0 );
buf ( n6822 , n30357 );
buf ( n6823 , n23197 );
buf ( n6824 , 1'b0 );
buf ( n6825 , 1'b0 );
buf ( n6826 , n30347 );
buf ( n6827 , n24909 );
buf ( n6828 , 1'b0 );
buf ( n6829 , 1'b0 );
buf ( n6830 , n30354 );
buf ( n6831 , n24912 );
buf ( n6832 , 1'b0 );
buf ( n6833 , 1'b0 );
buf ( n6834 , n30347 );
buf ( n6835 , n24914 );
buf ( n6836 , 1'b0 );
buf ( n6837 , 1'b0 );
buf ( n6838 , n30357 );
buf ( n6839 , n24916 );
buf ( n6840 , 1'b0 );
buf ( n6841 , 1'b0 );
buf ( n6842 , n30348 );
buf ( n6843 , n24919 );
buf ( n6844 , 1'b0 );
buf ( n6845 , 1'b0 );
buf ( n6846 , n30357 );
buf ( n6847 , n24922 );
buf ( n6848 , 1'b0 );
buf ( n6849 , 1'b0 );
buf ( n6850 , n30340 );
buf ( n6851 , n24924 );
buf ( n6852 , 1'b0 );
buf ( n6853 , 1'b0 );
buf ( n6854 , n30354 );
buf ( n6855 , n24926 );
buf ( n6856 , 1'b0 );
buf ( n6857 , 1'b0 );
buf ( n6858 , n30357 );
buf ( n6859 , n24928 );
buf ( n6860 , 1'b0 );
buf ( n6861 , 1'b0 );
buf ( n6862 , n30340 );
buf ( n6863 , n24930 );
buf ( n6864 , 1'b0 );
buf ( n6865 , 1'b0 );
buf ( n6866 , n30343 );
buf ( n6867 , n23199 );
buf ( n6868 , 1'b0 );
buf ( n6869 , 1'b0 );
buf ( n6870 , n30372 );
buf ( n6871 , n24932 );
buf ( n6872 , 1'b0 );
buf ( n6873 , 1'b0 );
buf ( n6874 , n30372 );
buf ( n6875 , n23202 );
buf ( n6876 , 1'b0 );
buf ( n6877 , 1'b0 );
buf ( n6878 , n30372 );
buf ( n6879 , n24934 );
buf ( n6880 , 1'b0 );
buf ( n6881 , 1'b0 );
buf ( n6882 , n30349 );
buf ( n6883 , n24936 );
buf ( n6884 , 1'b0 );
buf ( n6885 , 1'b0 );
buf ( n6886 , n30376 );
buf ( n6887 , n24939 );
buf ( n6888 , 1'b0 );
buf ( n6889 , 1'b0 );
buf ( n6890 , n30375 );
buf ( n6891 , n24941 );
buf ( n6892 , 1'b0 );
buf ( n6893 , 1'b0 );
buf ( n6894 , n30358 );
buf ( n6895 , n24943 );
buf ( n6896 , 1'b0 );
buf ( n6897 , 1'b0 );
buf ( n6898 , n30355 );
buf ( n6899 , n23213 );
buf ( n6900 , 1'b0 );
buf ( n6901 , 1'b0 );
buf ( n6902 , n1 );
buf ( n6903 , n30252 );
buf ( n6904 , 1'b0 );
buf ( n6905 , 1'b0 );
buf ( n6906 , n30375 );
buf ( n6907 , n28856 );
buf ( n6908 , 1'b0 );
buf ( n6909 , 1'b0 );
buf ( n6910 , n30378 );
buf ( n6911 , n28861 );
buf ( n6912 , 1'b0 );
buf ( n6913 , 1'b0 );
buf ( n6914 , n30358 );
buf ( n6915 , n28883 );
buf ( n6916 , 1'b0 );
buf ( n6917 , 1'b0 );
buf ( n6918 , n30378 );
buf ( n6919 , n29055 );
buf ( n6920 , 1'b0 );
buf ( n6921 , 1'b0 );
buf ( n6922 , n30376 );
buf ( n6923 , n29081 );
buf ( n6924 , 1'b0 );
buf ( n6925 , 1'b0 );
buf ( n6926 , n30375 );
buf ( n6927 , n23215 );
buf ( n6928 , 1'b0 );
buf ( n6929 , 1'b0 );
buf ( n6930 , n30374 );
buf ( n6931 , n28948 );
buf ( n6932 , 1'b0 );
buf ( n6933 , 1'b0 );
buf ( n6934 , n30347 );
buf ( n6935 , n22552 );
buf ( n6936 , 1'b0 );
buf ( n6937 , 1'b0 );
buf ( n6938 , n30358 );
buf ( n6939 , n24948 );
buf ( n6940 , 1'b0 );
buf ( n6941 , 1'b0 );
buf ( n6942 , n30372 );
buf ( n6943 , n28851 );
buf ( n6944 , 1'b0 );
buf ( n6945 , 1'b0 );
buf ( n6946 , n30347 );
buf ( n6947 , n24953 );
buf ( n6948 , 1'b0 );
buf ( n6949 , 1'b0 );
buf ( n6950 , n30372 );
buf ( n6951 , n24955 );
buf ( n6952 , 1'b0 );
buf ( n6953 , 1'b0 );
buf ( n6954 , n30351 );
buf ( n6955 , n24957 );
buf ( n6956 , 1'b0 );
buf ( n6957 , 1'b0 );
buf ( n6958 , n30347 );
buf ( n6959 , n24959 );
buf ( n6960 , 1'b0 );
buf ( n6961 , 1'b0 );
buf ( n6962 , n30356 );
buf ( n6963 , n23217 );
buf ( n6964 , 1'b0 );
buf ( n6965 , 1'b0 );
buf ( n6966 , n30345 );
buf ( n6967 , n24964 );
buf ( n6968 , 1'b0 );
buf ( n6969 , 1'b0 );
buf ( n6970 , n30372 );
buf ( n6971 , n23831 );
buf ( n6972 , 1'b0 );
buf ( n6973 , 1'b0 );
buf ( n6974 , n30347 );
buf ( n6975 , n24967 );
buf ( n6976 , 1'b0 );
buf ( n6977 , 1'b0 );
buf ( n6978 , n30355 );
buf ( n6979 , n24969 );
buf ( n6980 , 1'b0 );
buf ( n6981 , 1'b0 );
buf ( n6982 , n30356 );
buf ( n6983 , n24971 );
buf ( n6984 , 1'b0 );
buf ( n6985 , 1'b0 );
buf ( n6986 , n30345 );
buf ( n6987 , n24973 );
buf ( n6988 , 1'b0 );
buf ( n6989 , 1'b0 );
buf ( n6990 , n30378 );
buf ( n6991 , n24975 );
buf ( n6992 , 1'b0 );
buf ( n6993 , 1'b0 );
buf ( n6994 , n30352 );
buf ( n6995 , n23219 );
buf ( n6996 , 1'b0 );
buf ( n6997 , 1'b0 );
buf ( n6998 , n30378 );
buf ( n6999 , n1539 );
buf ( n7000 , 1'b0 );
buf ( n7001 , 1'b0 );
buf ( n7002 , n30343 );
buf ( n7003 , n28516 );
buf ( n7004 , 1'b0 );
buf ( n7005 , 1'b0 );
buf ( n7006 , n30376 );
buf ( n7007 , n24980 );
buf ( n7008 , 1'b0 );
buf ( n7009 , 1'b0 );
buf ( n7010 , n30355 );
buf ( n7011 , n24985 );
buf ( n7012 , 1'b0 );
buf ( n7013 , 1'b0 );
buf ( n7014 , n30376 );
buf ( n7015 , n24987 );
buf ( n7016 , 1'b0 );
buf ( n7017 , 1'b0 );
buf ( n7018 , n30343 );
buf ( n7019 , n24992 );
buf ( n7020 , 1'b0 );
buf ( n7021 , 1'b0 );
buf ( n7022 , n30353 );
buf ( n7023 , n24997 );
buf ( n7024 , 1'b0 );
buf ( n7025 , 1'b0 );
buf ( n7026 , n30374 );
buf ( n7027 , n25002 );
buf ( n7028 , 1'b0 );
buf ( n7029 , 1'b0 );
buf ( n7030 , n30356 );
buf ( n7031 , n25007 );
buf ( n7032 , 1'b0 );
buf ( n7033 , 1'b0 );
buf ( n7034 , n30355 );
buf ( n7035 , n23594 );
buf ( n7036 , 1'b0 );
buf ( n7037 , 1'b0 );
buf ( n7038 , n30353 );
buf ( n7039 , n25022 );
buf ( n7040 , 1'b0 );
buf ( n7041 , 1'b0 );
buf ( n7042 , n30374 );
buf ( n7043 , n25012 );
buf ( n7044 , 1'b0 );
buf ( n7045 , 1'b0 );
buf ( n7046 , n30374 );
buf ( n7047 , n25017 );
buf ( n7048 , 1'b0 );
buf ( n7049 , 1'b0 );
buf ( n7050 , n30345 );
buf ( n7051 , n23582 );
buf ( n7052 , 1'b0 );
buf ( n7053 , 1'b0 );
buf ( n7054 , n30351 );
buf ( n7055 , n23221 );
buf ( n7056 , 1'b0 );
buf ( n7057 , 1'b0 );
buf ( n7058 , n30356 );
buf ( n7059 , n25027 );
buf ( n7060 , 1'b0 );
buf ( n7061 , 1'b0 );
buf ( n7062 , n30376 );
buf ( n7063 , n23223 );
buf ( n7064 , 1'b0 );
buf ( n7065 , 1'b0 );
buf ( n7066 , n30346 );
buf ( n7067 , n25032 );
buf ( n7068 , 1'b0 );
buf ( n7069 , 1'b0 );
buf ( n7070 , n30356 );
buf ( n7071 , n25037 );
buf ( n7072 , 1'b0 );
buf ( n7073 , 1'b0 );
buf ( n7074 , n30371 );
buf ( n7075 , n25039 );
buf ( n7076 , 1'b0 );
buf ( n7077 , 1'b0 );
buf ( n7078 , n30356 );
buf ( n7079 , n25054 );
buf ( n7080 , 1'b0 );
buf ( n7081 , 1'b0 );
buf ( n7082 , n30371 );
buf ( n7083 , n25044 );
buf ( n7084 , 1'b0 );
buf ( n7085 , 1'b0 );
buf ( n7086 , n30352 );
buf ( n7087 , n25049 );
buf ( n7088 , 1'b0 );
buf ( n7089 , 1'b0 );
buf ( n7090 , n30351 );
buf ( n7091 , n25064 );
buf ( n7092 , 1'b0 );
buf ( n7093 , 1'b0 );
buf ( n7094 , n30371 );
buf ( n7095 , n25059 );
buf ( n7096 , 1'b0 );
buf ( n7097 , 1'b0 );
buf ( n7098 , n30343 );
buf ( n7099 , n23225 );
buf ( n7100 , 1'b0 );
buf ( n7101 , 1'b0 );
buf ( n7102 , n30375 );
buf ( n7103 , n23227 );
buf ( n7104 , 1'b0 );
buf ( n7105 , 1'b0 );
buf ( n7106 , n30351 );
buf ( n7107 , n25069 );
buf ( n7108 , 1'b0 );
buf ( n7109 , 1'b0 );
buf ( n7110 , n30375 );
buf ( n7111 , n25072 );
buf ( n7112 , 1'b0 );
buf ( n7113 , 1'b0 );
buf ( n7114 , n30342 );
buf ( n7115 , n25074 );
buf ( n7116 , 1'b0 );
buf ( n7117 , 1'b0 );
buf ( n7118 , n30346 );
buf ( n7119 , n25079 );
buf ( n7120 , 1'b0 );
buf ( n7121 , 1'b0 );
buf ( n7122 , n30346 );
buf ( n7123 , n25081 );
buf ( n7124 , 1'b0 );
buf ( n7125 , 1'b0 );
buf ( n7126 , n30353 );
buf ( n7127 , n25083 );
buf ( n7128 , 1'b0 );
buf ( n7129 , 1'b0 );
buf ( n7130 , n30371 );
buf ( n7131 , n25085 );
buf ( n7132 , 1'b0 );
buf ( n7133 , 1'b0 );
buf ( n7134 , n30356 );
buf ( n7135 , n25087 );
buf ( n7136 , 1'b0 );
buf ( n7137 , 1'b0 );
buf ( n7138 , n30352 );
buf ( n7139 , n28526 );
buf ( n7140 , 1'b0 );
buf ( n7141 , 1'b0 );
buf ( n7142 , n1 );
buf ( n7143 , n27049 );
buf ( n7144 , 1'b0 );
buf ( n7145 , 1'b0 );
buf ( n7146 , n1 );
buf ( n7147 , n27054 );
buf ( n7148 , 1'b0 );
buf ( n7149 , 1'b0 );
buf ( n7150 , n1 );
buf ( n7151 , n26469 );
buf ( n7152 , 1'b0 );
buf ( n7153 , 1'b0 );
buf ( n7154 , n1 );
buf ( n7155 , n27064 );
buf ( n7156 , 1'b0 );
buf ( n7157 , 1'b0 );
buf ( n7158 , n1 );
buf ( n7159 , n27059 );
buf ( n7160 , 1'b0 );
buf ( n7161 , 1'b0 );
buf ( n7162 , n1 );
buf ( n7163 , n26464 );
buf ( n7164 , 1'b0 );
buf ( n7165 , 1'b0 );
buf ( n7166 , n30356 );
buf ( n7167 , n25090 );
buf ( n7168 , 1'b0 );
buf ( n7169 , 1'b0 );
buf ( n7170 , n1 );
buf ( n7171 , n27105 );
buf ( n7172 , 1'b0 );
buf ( n7173 , 1'b0 );
buf ( n7174 , n1 );
buf ( n7175 , n26414 );
buf ( n7176 , 1'b0 );
buf ( n7177 , 1'b0 );
buf ( n7178 , n1 );
buf ( n7179 , n26351 );
buf ( n7180 , 1'b0 );
buf ( n7181 , 1'b0 );
buf ( n7182 , n1 );
buf ( n7183 , n26299 );
buf ( n7184 , 1'b0 );
buf ( n7185 , 1'b0 );
buf ( n7186 , n1 );
buf ( n7187 , n26249 );
buf ( n7188 , 1'b0 );
buf ( n7189 , 1'b0 );
buf ( n7190 , n1 );
buf ( n7191 , n27145 );
buf ( n7192 , 1'b0 );
buf ( n7193 , 1'b0 );
buf ( n7194 , n1 );
buf ( n7195 , n27292 );
buf ( n7196 , 1'b0 );
buf ( n7197 , 1'b0 );
buf ( n7198 , n1 );
buf ( n7199 , n26152 );
buf ( n7200 , 1'b0 );
buf ( n7201 , 1'b0 );
buf ( n7202 , n1 );
buf ( n7203 , n26105 );
buf ( n7204 , 1'b0 );
buf ( n7205 , 1'b0 );
buf ( n7206 , n1 );
buf ( n7207 , n25904 );
buf ( n7208 , 1'b0 );
buf ( n7209 , 1'b0 );
buf ( n7210 , n1 );
buf ( n7211 , n27189 );
buf ( n7212 , 1'b0 );
buf ( n7213 , 1'b0 );
buf ( n7214 , n1 );
buf ( n7215 , n25993 );
buf ( n7216 , 1'b0 );
buf ( n7217 , 1'b0 );
buf ( n7218 , n30346 );
buf ( n7219 , n25092 );
buf ( n7220 , 1'b0 );
buf ( n7221 , 1'b0 );
buf ( n7222 , n30352 );
buf ( n7223 , n18726 );
buf ( n7224 , 1'b0 );
buf ( n7225 , 1'b0 );
buf ( n7226 , n30342 );
buf ( n7227 , n18735 );
buf ( n7228 , 1'b0 );
buf ( n7229 , 1'b0 );
buf ( n7230 , n30352 );
buf ( n7231 , n18744 );
buf ( n7232 , 1'b0 );
buf ( n7233 , 1'b0 );
buf ( n7234 , n30358 );
buf ( n7235 , n18753 );
buf ( n7236 , 1'b0 );
buf ( n7237 , 1'b0 );
buf ( n7238 , n30352 );
buf ( n7239 , n25163 );
buf ( n7240 , 1'b0 );
buf ( n7241 , 1'b0 );
buf ( n7242 , n30371 );
buf ( n7243 , n25095 );
buf ( n7244 , 1'b0 );
buf ( n7245 , 1'b0 );
buf ( n7246 , n30342 );
buf ( n7247 , n25097 );
buf ( n7248 , 1'b0 );
buf ( n7249 , 1'b0 );
buf ( n7250 , n30345 );
buf ( n7251 , n28864 );
buf ( n7252 , 1'b0 );
buf ( n7253 , 1'b0 );
buf ( n7254 , n30378 );
buf ( n7255 , n29900 );
buf ( n7256 , 1'b0 );
buf ( n7257 , 1'b0 );
buf ( n7258 , n1 );
buf ( n7259 , n27807 );
buf ( n7260 , 1'b0 );
buf ( n7261 , 1'b0 );
buf ( n7262 , n30343 );
buf ( n7263 , n25099 );
buf ( n7264 , 1'b0 );
buf ( n7265 , 1'b0 );
buf ( n7266 , n30342 );
buf ( n7267 , n28652 );
buf ( n7268 , 1'b0 );
buf ( n7269 , 1'b0 );
buf ( n7270 , n30345 );
buf ( n7271 , n28867 );
buf ( n7272 , 1'b0 );
buf ( n7273 , 1'b0 );
buf ( n7274 , n1 );
buf ( n7275 , n25813 );
buf ( n7276 , 1'b0 );
buf ( n7277 , 1'b0 );
buf ( n7278 , n1 );
buf ( n7279 , n27194 );
buf ( n7280 , 1'b0 );
buf ( n7281 , 1'b0 );
buf ( n7282 , n1 );
buf ( n7283 , n27199 );
buf ( n7284 , 1'b0 );
buf ( n7285 , 1'b0 );
buf ( n7286 , n1 );
buf ( n7287 , n27214 );
buf ( n7288 , 1'b0 );
buf ( n7289 , 1'b0 );
buf ( n7290 , n1 );
buf ( n7291 , n27204 );
buf ( n7292 , 1'b0 );
buf ( n7293 , 1'b0 );
buf ( n7294 , n1 );
buf ( n7295 , n27209 );
buf ( n7296 , 1'b0 );
buf ( n7297 , 1'b0 );
buf ( n7298 , n1 );
buf ( n7299 , n26567 );
buf ( n7300 , 1'b0 );
buf ( n7301 , 1'b0 );
buf ( n7302 , n1 );
buf ( n7303 , n25634 );
buf ( n7304 , 1'b0 );
buf ( n7305 , 1'b0 );
buf ( n7306 , n1 );
buf ( n7307 , n25629 );
buf ( n7308 , 1'b0 );
buf ( n7309 , 1'b0 );
buf ( n7310 , n1 );
buf ( n7311 , n25257 );
buf ( n7312 , 1'b0 );
buf ( n7313 , 1'b0 );
buf ( n7314 , n1 );
buf ( n7315 , n26562 );
buf ( n7316 , 1'b0 );
buf ( n7317 , 1'b0 );
buf ( n7318 , n1 );
buf ( n7319 , n26557 );
buf ( n7320 , 1'b0 );
buf ( n7321 , 1'b0 );
buf ( n7322 , n30343 );
buf ( n7323 , n23229 );
buf ( n7324 , 1'b0 );
buf ( n7325 , 1'b0 );
buf ( n7326 , n30342 );
buf ( n7327 , n25101 );
buf ( n7328 , 1'b0 );
buf ( n7329 , 1'b0 );
buf ( n7330 , n30351 );
buf ( n7331 , n25103 );
buf ( n7332 , 1'b0 );
buf ( n7333 , 1'b0 );
buf ( n7334 , n30342 );
buf ( n7335 , n28541 );
buf ( n7336 , 1'b0 );
buf ( n7337 , 1'b0 );
buf ( n7338 , n30378 );
buf ( n7339 , n28544 );
buf ( n7340 , 1'b0 );
buf ( n7341 , 1'b0 );
buf ( n7342 , n30346 );
buf ( n7343 , n28547 );
buf ( n7344 , 1'b0 );
buf ( n7345 , 1'b0 );
buf ( n7346 , n30343 );
buf ( n7347 , n28550 );
buf ( n7348 , 1'b0 );
buf ( n7349 , 1'b0 );
buf ( n7350 , n30351 );
buf ( n7351 , n25108 );
buf ( n7352 , 1'b0 );
buf ( n7353 , 1'b0 );
buf ( n7354 , n1 );
buf ( n7355 , n26522 );
buf ( n7356 , 1'b0 );
buf ( n7357 , 1'b0 );
buf ( n7358 , n30346 );
buf ( n7359 , n19229 );
buf ( n7360 , 1'b0 );
buf ( n7361 , 1'b0 );
buf ( n7362 , n30343 );
buf ( n7363 , n19273 );
buf ( n7364 , 1'b0 );
buf ( n7365 , 1'b0 );
buf ( n7366 , n30378 );
buf ( n7367 , n25117 );
buf ( n7368 , 1'b0 );
buf ( n7369 , 1'b0 );
buf ( n7370 , n30346 );
buf ( n7371 , n25110 );
buf ( n7372 , 1'b0 );
buf ( n7373 , 1'b0 );
buf ( n7374 , n30353 );
buf ( n7375 , n25112 );
buf ( n7376 , 1'b0 );
buf ( n7377 , 1'b0 );
buf ( n7378 , n30345 );
buf ( n7379 , n28905 );
buf ( n7380 , 1'b0 );
buf ( n7381 , 1'b0 );
buf ( n7382 , n30346 );
buf ( n7383 , n23231 );
buf ( n7384 , 1'b0 );
buf ( n7385 , 1'b0 );
buf ( n7386 , n30352 );
buf ( n7387 , n23236 );
buf ( n7388 , 1'b0 );
buf ( n7389 , 1'b0 );
buf ( n7390 , n30375 );
buf ( n7391 , n23242 );
buf ( n7392 , 1'b0 );
buf ( n7393 , 1'b0 );
buf ( n7394 , n30376 );
buf ( n7395 , n23248 );
buf ( n7396 , 1'b0 );
buf ( n7397 , 1'b0 );
buf ( n7398 , n30353 );
buf ( n7399 , n23253 );
buf ( n7400 , 1'b0 );
buf ( n7401 , 1'b0 );
buf ( n7402 , n30353 );
buf ( n7403 , n23258 );
buf ( n7404 , 1'b0 );
buf ( n7405 , 1'b0 );
buf ( n7406 , n30342 );
buf ( n7407 , n21757 );
buf ( n7408 , 1'b0 );
buf ( n7409 , 1'b0 );
buf ( n7410 , n30353 );
buf ( n7411 , n23264 );
buf ( n7412 , 1'b0 );
buf ( n7413 , 1'b0 );
buf ( n7414 , n30358 );
buf ( n7415 , n23269 );
buf ( n7416 , 1'b0 );
buf ( n7417 , 1'b0 );
buf ( n7418 , n30356 );
buf ( n7419 , n23274 );
buf ( n7420 , 1'b0 );
buf ( n7421 , 1'b0 );
buf ( n7422 , n30371 );
buf ( n7423 , n21768 );
buf ( n7424 , 1'b0 );
buf ( n7425 , 1'b0 );
buf ( n7426 , n30358 );
buf ( n7427 , n23279 );
buf ( n7428 , 1'b0 );
buf ( n7429 , 1'b0 );
buf ( n7430 , n30351 );
buf ( n7431 , n25275 );
buf ( n7432 , 1'b0 );
buf ( n7433 , 1'b0 );
buf ( n7434 , n30371 );
buf ( n7435 , n23285 );
buf ( n7436 , 1'b0 );
buf ( n7437 , 1'b0 );
buf ( n7438 , n30374 );
buf ( n7439 , n25128 );
buf ( n7440 , 1'b0 );
buf ( n7441 , 1'b0 );
buf ( n7442 , n30345 );
buf ( n7443 , n25123 );
buf ( n7444 , 1'b0 );
buf ( n7445 , 1'b0 );
buf ( n7446 , n30355 );
buf ( n7447 , n23290 );
buf ( n7448 , 1'b0 );
buf ( n7449 , 1'b0 );
buf ( n7450 , n30355 );
buf ( n7451 , n23295 );
buf ( n7452 , 1'b0 );
buf ( n7453 , 1'b0 );
buf ( n7454 , n30374 );
buf ( n7455 , n23300 );
buf ( n7456 , 1'b0 );
buf ( n7457 , 1'b0 );
buf ( n7458 , n1 );
buf ( n7459 , n26517 );
buf ( n7460 , 1'b0 );
buf ( n7461 , 1'b0 );
buf ( n7462 , n1 );
buf ( n7463 , n27568 );
buf ( n7464 , 1'b0 );
buf ( n7465 , 1'b0 );
buf ( n7466 , n1 );
buf ( n7467 , n27591 );
buf ( n7468 , 1'b0 );
buf ( n7469 , 1'b0 );
buf ( n7470 , n1 );
buf ( n7471 , n27252 );
buf ( n7472 , 1'b0 );
buf ( n7473 , 1'b0 );
buf ( n7474 , n30355 );
buf ( n7475 , n25133 );
buf ( n7476 , 1'b0 );
buf ( n7477 , 1'b0 );
buf ( n7478 , n30378 );
buf ( n7479 , n27827 );
buf ( n7480 , 1'b0 );
buf ( n7481 , 1'b0 );
buf ( n7482 , n1 );
buf ( n7483 , n27614 );
buf ( n7484 , 1'b0 );
buf ( n7485 , 1'b0 );
buf ( n7486 , n1 );
buf ( n7487 , n27637 );
buf ( n7488 , 1'b0 );
buf ( n7489 , 1'b0 );
buf ( n7490 , n1 );
buf ( n7491 , n27660 );
buf ( n7492 , 1'b0 );
buf ( n7493 , 1'b0 );
buf ( n7494 , n30355 );
buf ( n7495 , n23308 );
buf ( n7496 , 1'b0 );
buf ( n7497 , 1'b0 );
buf ( n7498 , n30376 );
buf ( n7499 , n23313 );
buf ( n7500 , 1'b0 );
buf ( n7501 , 1'b0 );
buf ( n7502 , n30345 );
buf ( n7503 , n23318 );
buf ( n7504 , 1'b0 );
buf ( n7505 , 1'b0 );
buf ( n7506 , n30358 );
buf ( n7507 , n23324 );
buf ( n7508 , 1'b0 );
buf ( n7509 , 1'b0 );
buf ( n7510 , n30347 );
buf ( n7511 , n23329 );
buf ( n7512 , 1'b0 );
buf ( n7513 , 1'b0 );
buf ( n7514 , n30347 );
buf ( n7515 , n23334 );
buf ( n7516 , 1'b0 );
buf ( n7517 , 1'b0 );
buf ( n7518 , n30372 );
buf ( n7519 , n23489 );
buf ( n7520 , 1'b0 );
buf ( n7521 , 1'b0 );
buf ( n7522 , n30347 );
buf ( n7523 , n23339 );
buf ( n7524 , 1'b0 );
buf ( n7525 , 1'b0 );
buf ( n7526 , n30358 );
buf ( n7527 , n23344 );
buf ( n7528 , 1'b0 );
buf ( n7529 , 1'b0 );
buf ( n7530 , n30378 );
buf ( n7531 , n23349 );
buf ( n7532 , 1'b0 );
buf ( n7533 , 1'b0 );
buf ( n7534 , n30358 );
buf ( n7535 , n23494 );
buf ( n7536 , 1'b0 );
buf ( n7537 , 1'b0 );
buf ( n7538 , n30340 );
buf ( n7539 , n23354 );
buf ( n7540 , 1'b0 );
buf ( n7541 , 1'b0 );
buf ( n7542 , n30347 );
buf ( n7543 , n23359 );
buf ( n7544 , 1'b0 );
buf ( n7545 , 1'b0 );
buf ( n7546 , n30372 );
buf ( n7547 , n23365 );
buf ( n7548 , 1'b0 );
buf ( n7549 , 1'b0 );
buf ( n7550 , n30356 );
buf ( n7551 , n23462 );
buf ( n7552 , 1'b0 );
buf ( n7553 , 1'b0 );
buf ( n7554 , n30340 );
buf ( n7555 , n23370 );
buf ( n7556 , 1'b0 );
buf ( n7557 , 1'b0 );
buf ( n7558 , n30340 );
buf ( n7559 , n23375 );
buf ( n7560 , 1'b0 );
buf ( n7561 , 1'b0 );
buf ( n7562 , n30375 );
buf ( n7563 , n23380 );
buf ( n7564 , 1'b0 );
buf ( n7565 , 1'b0 );
buf ( n7566 , n1 );
buf ( n7567 , n27702 );
buf ( n7568 , 1'b0 );
buf ( n7569 , 1'b0 );
buf ( n7570 , n30378 );
buf ( n7571 , n23385 );
buf ( n7572 , 1'b0 );
buf ( n7573 , 1'b0 );
buf ( n7574 , n30357 );
buf ( n7575 , n23390 );
buf ( n7576 , 1'b0 );
buf ( n7577 , 1'b0 );
buf ( n7578 , n30340 );
buf ( n7579 , n23395 );
buf ( n7580 , 1'b0 );
buf ( n7581 , 1'b0 );
buf ( n7582 , n30347 );
buf ( n7583 , n23400 );
buf ( n7584 , 1'b0 );
buf ( n7585 , 1'b0 );
buf ( n7586 , n30349 );
buf ( n7587 , n23120 );
buf ( n7588 , 1'b0 );
buf ( n7589 , 1'b0 );
buf ( n7590 , n30340 );
buf ( n7591 , n19318 );
buf ( n7592 , 1'b0 );
buf ( n7593 , 1'b0 );
buf ( n7594 , n30357 );
buf ( n7595 , n19361 );
buf ( n7596 , 1'b0 );
buf ( n7597 , 1'b0 );
buf ( n7598 , n30347 );
buf ( n7599 , n23406 );
buf ( n7600 , 1'b0 );
buf ( n7601 , 1'b0 );
buf ( n7602 , n30348 );
buf ( n7603 , n28514 );
buf ( n7604 , 1'b0 );
buf ( n7605 , 1'b0 );
buf ( n7606 , n30373 );
buf ( n7607 , n23411 );
buf ( n7608 , 1'b0 );
buf ( n7609 , 1'b0 );
buf ( n7610 , n30357 );
buf ( n7611 , n23416 );
buf ( n7612 , 1'b0 );
buf ( n7613 , 1'b0 );
buf ( n7614 , n30373 );
buf ( n7615 , n21806 );
buf ( n7616 , 1'b0 );
buf ( n7617 , 1'b0 );
buf ( n7618 , n30340 );
buf ( n7619 , n23421 );
buf ( n7620 , 1'b0 );
buf ( n7621 , 1'b0 );
buf ( n7622 , n30354 );
buf ( n7623 , n23426 );
buf ( n7624 , 1'b0 );
buf ( n7625 , 1'b0 );
buf ( n7626 , n30377 );
buf ( n7627 , n23431 );
buf ( n7628 , 1'b0 );
buf ( n7629 , 1'b0 );
buf ( n7630 , n30354 );
buf ( n7631 , n21811 );
buf ( n7632 , 1'b0 );
buf ( n7633 , 1'b0 );
buf ( n7634 , n30377 );
buf ( n7635 , n1547 );
buf ( n7636 , 1'b0 );
buf ( n7637 , 1'b0 );
buf ( n7638 , n30348 );
buf ( n7639 , n1547 );
buf ( n7640 , 1'b0 );
buf ( n7641 , 1'b0 );
buf ( n7642 , n30348 );
buf ( n7643 , n23436 );
buf ( n7644 , 1'b0 );
buf ( n7645 , 1'b0 );
buf ( n7646 , n30373 );
buf ( n7647 , n23441 );
buf ( n7648 , 1'b0 );
buf ( n7649 , 1'b0 );
buf ( n7650 , n30357 );
buf ( n7651 , n25138 );
buf ( n7652 , 1'b0 );
buf ( n7653 , 1'b0 );
buf ( n7654 , n1 );
buf ( n7655 , n27851 );
buf ( n7656 , 1'b0 );
buf ( n7657 , 1'b0 );
buf ( n7658 , n1 );
buf ( n7659 , n27875 );
buf ( n7660 , 1'b0 );
buf ( n7661 , 1'b0 );
buf ( n7662 , n30373 );
buf ( n7663 , n29325 );
buf ( n7664 , 1'b0 );
buf ( n7665 , 1'b0 );
buf ( n7666 , n30349 );
buf ( n7667 , n29356 );
buf ( n7668 , 1'b0 );
buf ( n7669 , 1'b0 );
buf ( n7670 , n30349 );
buf ( n7671 , n15346 );
buf ( n7672 , 1'b0 );
buf ( n7673 , 1'b0 );
buf ( n7674 , n1 );
buf ( n7675 , n27881 );
buf ( n7676 , 1'b0 );
buf ( n7677 , 1'b0 );
buf ( n7678 , n30377 );
buf ( n7679 , n25247 );
buf ( n7680 , 1'b0 );
buf ( n7681 , 1'b0 );
buf ( n7682 , n1 );
buf ( n7683 , n27892 );
buf ( n7684 , 1'b0 );
buf ( n7685 , 1'b0 );
buf ( n7686 , n30372 );
buf ( n7687 , n28505 );
buf ( n7688 , 1'b0 );
buf ( n7689 , 1'b0 );
buf ( n7690 , n1 );
buf ( n7691 , n27897 );
buf ( n7692 , 1'b0 );
buf ( n7693 , 1'b0 );
buf ( n7694 , n1 );
buf ( n7695 , n28868 );
buf ( n7696 , 1'b0 );
buf ( n7697 , 1'b0 );
buf ( n7698 , n1 );
buf ( n7699 , n27902 );
buf ( n7700 , 1'b0 );
buf ( n7701 , 1'b0 );
buf ( n7702 , n1 );
buf ( n7703 , n27907 );
buf ( n7704 , 1'b0 );
buf ( n7705 , 1'b0 );
buf ( n7706 , n30377 );
buf ( n7707 , n18928 );
buf ( n7708 , 1'b0 );
buf ( n7709 , 1'b0 );
buf ( n7710 , n1 );
buf ( n7711 , n27912 );
buf ( n7712 , 1'b0 );
buf ( n7713 , 1'b0 );
buf ( n7714 , n30349 );
buf ( n7715 , n28510 );
buf ( n7716 , 1'b0 );
buf ( n7717 , 1'b0 );
buf ( n7718 , n30373 );
buf ( n7719 , n20432 );
buf ( n7720 , 1'b0 );
buf ( n7721 , 1'b0 );
buf ( n7722 , n30372 );
buf ( n7723 , n25240 );
buf ( n7724 , 1'b0 );
buf ( n7725 , 1'b0 );
buf ( n7726 , n30354 );
buf ( n7727 , n25234 );
buf ( n7728 , 1'b0 );
buf ( n7729 , 1'b0 );
buf ( n7730 , n30354 );
buf ( n7731 , n25222 );
buf ( n7732 , 1'b0 );
buf ( n7733 , 1'b0 );
buf ( n7734 , n1 );
buf ( n7735 , n27923 );
buf ( n7736 , 1'b0 );
buf ( n7737 , 1'b0 );
buf ( n7738 , n1 );
buf ( n7739 , n28557 );
buf ( n7740 , 1'b0 );
buf ( n7741 , 1'b0 );
buf ( n7742 , n1 );
buf ( n7743 , n28564 );
buf ( n7744 , 1'b0 );
buf ( n7745 , 1'b0 );
buf ( n7746 , n30372 );
buf ( n7747 , n28565 );
buf ( n7748 , 1'b0 );
buf ( n7749 , 1'b0 );
buf ( n7750 , n1 );
buf ( n7751 , n28337 );
buf ( n7752 , 1'b0 );
buf ( n7753 , 1'b0 );
buf ( n7754 , n30372 );
buf ( n7755 , n28567 );
buf ( n7756 , 1'b0 );
buf ( n7757 , 1'b0 );
buf ( n7758 , n30349 );
buf ( n7759 , n28530 );
buf ( n7760 , 1'b0 );
buf ( n7761 , 1'b0 );
buf ( n7762 , n1 );
buf ( n7763 , n28348 );
buf ( n7764 , 1'b0 );
buf ( n7765 , 1'b0 );
buf ( n7766 , n30377 );
buf ( n7767 , n21463 );
buf ( n7768 , 1'b0 );
buf ( n7769 , 1'b0 );
buf ( n7770 , n30349 );
buf ( n7771 , n21470 );
buf ( n7772 , 1'b0 );
buf ( n7773 , 1'b0 );
buf ( n7774 , n30373 );
buf ( n7775 , n21477 );
buf ( n7776 , 1'b0 );
buf ( n7777 , 1'b0 );
buf ( n7778 , n1 );
buf ( n7779 , n28368 );
buf ( n7780 , 1'b0 );
buf ( n7781 , 1'b0 );
buf ( n7782 , n30377 );
buf ( n7783 , n21484 );
buf ( n7784 , 1'b0 );
buf ( n7785 , 1'b0 );
buf ( n7786 , n30377 );
buf ( n7787 , n20427 );
buf ( n7788 , 1'b0 );
buf ( n7789 , 1'b0 );
buf ( n7790 , n1 );
buf ( n7791 , n27988 );
buf ( n7792 , 1'b0 );
buf ( n7793 , 1'b0 );
buf ( n7794 , n1 );
buf ( n7795 , n27934 );
buf ( n7796 , 1'b0 );
buf ( n7797 , 1'b0 );
buf ( n7798 , n30349 );
buf ( n7799 , n27942 );
buf ( n7800 , 1'b0 );
buf ( n7801 , 1'b0 );
buf ( n7802 , n30373 );
buf ( n7803 , n27950 );
buf ( n7804 , 1'b0 );
buf ( n7805 , 1'b0 );
buf ( n7806 , n30354 );
buf ( n7807 , n27958 );
buf ( n7808 , 1'b0 );
buf ( n7809 , 1'b0 );
buf ( n7810 , n30349 );
buf ( n7811 , n27966 );
buf ( n7812 , 1'b0 );
buf ( n7813 , 1'b0 );
buf ( n7814 , n1 );
buf ( n7815 , n28649 );
buf ( n7816 , 1'b0 );
buf ( n7817 , 1'b0 );
buf ( n7818 , n1 );
buf ( n7819 , n28538 );
buf ( n7820 , 1'b0 );
buf ( n7821 , 1'b0 );
buf ( n7822 , n1 );
buf ( n7823 , n28379 );
buf ( n7824 , 1'b0 );
buf ( n7825 , 1'b0 );
buf ( n7826 , n30348 );
buf ( n7827 , n28484 );
buf ( n7828 , 1'b0 );
buf ( n7829 , 1'b0 );
buf ( n7830 , n30357 );
buf ( n7831 , n28571 );
buf ( n7832 , 1'b0 );
buf ( n7833 , 1'b0 );
buf ( n7834 , n30357 );
buf ( n7835 , n20414 );
buf ( n7836 , 1'b0 );
buf ( n7837 , 1'b0 );
buf ( n7838 , n30373 );
buf ( n7839 , n28923 );
buf ( n7840 , 1'b0 );
buf ( n7841 , 1'b0 );
buf ( n7842 , n1 );
buf ( n7843 , n28576 );
buf ( n7844 , 1'b0 );
buf ( n7845 , 1'b0 );
buf ( n7846 , n1 );
buf ( n7847 , n28583 );
buf ( n7848 , 1'b0 );
buf ( n7849 , 1'b0 );
buf ( n7850 , n30373 );
buf ( n7851 , n28326 );
buf ( n7852 , 1'b0 );
buf ( n7853 , 1'b0 );
buf ( n7854 , n30373 );
buf ( n7855 , n29597 );
buf ( n7856 , 1'b0 );
buf ( n7857 , 1'b0 );
buf ( n7858 , n30377 );
buf ( n7859 , n29945 );
buf ( n7860 , 1'b0 );
buf ( n7861 , 1'b0 );
buf ( n7862 , n30347 );
buf ( n7863 , n30369 );
buf ( n7864 , 1'b0 );
buf ( n7865 , 1'b0 );
buf ( n7866 , n1 );
buf ( n7867 , n28590 );
buf ( n7868 , 1'b0 );
buf ( n7869 , 1'b0 );
buf ( n7870 , n1 );
buf ( n7871 , n28596 );
buf ( n7872 , 1'b0 );
buf ( n7873 , 1'b0 );
buf ( n7874 , n1 );
buf ( n7875 , n28317 );
buf ( n7876 , 1'b0 );
buf ( n7877 , 1'b0 );
buf ( n7878 , n30357 );
buf ( n7879 , n29008 );
buf ( n7880 , 1'b0 );
buf ( n7881 , 1'b0 );
buf ( n7882 , n30373 );
buf ( n7883 , n29015 );
buf ( n7884 , 1'b0 );
buf ( n7885 , 1'b0 );
buf ( n7886 , n30357 );
buf ( n7887 , n30402 );
buf ( n7888 , 1'b0 );
buf ( n7889 , 1'b0 );
buf ( n7890 , n30357 );
buf ( n7891 , n28598 );
buf ( n7892 , 1'b0 );
buf ( n7893 , 1'b0 );
buf ( n7894 , n1 );
buf ( n7895 , n28925 );
buf ( n7896 , 1'b0 );
buf ( n7897 , 1'b0 );
buf ( n7898 , n1 );
buf ( n7899 , n28927 );
buf ( n7900 , 1'b0 );
buf ( n7901 , 1'b0 );
buf ( n7902 , n30354 );
buf ( n7903 , n30386 );
buf ( n7904 , 1'b0 );
buf ( n7905 , 1'b0 );
buf ( n7906 , n1 );
buf ( n7907 , n29196 );
buf ( n7908 , 1'b0 );
buf ( n7909 , 1'b0 );
buf ( n7910 , n30376 );
buf ( n7911 , n30394 );
buf ( n7912 , 1'b0 );
buf ( n7913 , 1'b0 );
buf ( n7914 , n30340 );
buf ( n7915 , n29001 );
buf ( n7916 , 1'b0 );
buf ( n7917 , 1'b0 );
buf ( n7918 , n30378 );
buf ( n7919 , n20421 );
buf ( n7920 , 1'b0 );
buf ( n7921 , 1'b0 );
buf ( n7922 , n30358 );
buf ( n7923 , n30116 );
buf ( n7924 , 1'b0 );
buf ( n7925 , 1'b0 );
buf ( n7926 , n1 );
buf ( n7927 , n28996 );
buf ( n7928 , 1'b0 );
buf ( n7929 , 1'b0 );
buf ( n7930 , n1 );
buf ( n7931 , n28603 );
buf ( n7932 , 1'b0 );
buf ( n7933 , 1'b0 );
buf ( n7934 , n1 );
buf ( n7935 , n28608 );
buf ( n7936 , 1'b0 );
buf ( n7937 , 1'b0 );
buf ( n7938 , n1 );
buf ( n7939 , n28708 );
buf ( n7940 , 1'b0 );
buf ( n7941 , 1'b0 );
buf ( n7942 , n1 );
buf ( n7943 , n28875 );
buf ( n7944 , 1'b0 );
buf ( n7945 , 1'b0 );
buf ( n7946 , n1 );
buf ( n7947 , n30366 );
buf ( n7948 , 1'b0 );
buf ( n7949 , 1'b0 );
buf ( n7950 , n1 );
buf ( n7951 , n28993 );
buf ( n7952 , 1'b0 );
buf ( n7953 , 1'b0 );
buf ( n7954 , n1 );
buf ( n7955 , n29882 );
buf ( n7956 , 1'b0 );
buf ( n7957 , 1'b0 );
buf ( n7958 , n1 );
buf ( n7959 , n28929 );
buf ( n7960 , 1'b0 );
buf ( n7961 , 1'b0 );
buf ( n7962 , n1 );
buf ( n7963 , n29309 );
buf ( n7964 , 1'b0 );
buf ( n7965 , 1'b0 );
buf ( n7966 , n1 );
buf ( n7967 , n29199 );
buf ( n7968 , 1'b0 );
buf ( n7969 , 1'b0 );
buf ( n7970 , n30375 );
buf ( n7971 , n28306 );
buf ( n7972 , 1'b0 );
buf ( n7973 , 1'b0 );
buf ( n7974 , n30358 );
buf ( n7975 , n28489 );
buf ( n7976 , 1'b0 );
buf ( n7977 , 1'b0 );
buf ( n7978 , n30376 );
buf ( n7979 , n28901 );
buf ( n7980 , 1'b0 );
buf ( n7981 , 1'b0 );
buf ( n7982 , n30358 );
buf ( n7983 , n1755 );
buf ( n7984 , 1'b0 );
buf ( n7985 , 1'b0 );
buf ( n7986 , n1 );
buf ( n7987 , n29084 );
buf ( n7988 , 1'b0 );
buf ( n7989 , 1'b0 );
buf ( n7990 , n30347 );
buf ( n7991 , n27667 );
buf ( n7992 , 1'b0 );
buf ( n7993 , 1'b0 );
buf ( n7994 , n30347 );
buf ( n7995 , n30387 );
buf ( n7996 , 1'b0 );
buf ( n7997 , 1'b0 );
buf ( n7998 , n30351 );
buf ( n7999 , n30388 );
buf ( n8000 , 1'b0 );
buf ( n8001 , 1'b0 );
buf ( n8002 , n30378 );
buf ( n8003 , n27977 );
buf ( n8004 , 1'b0 );
buf ( n8005 , 1'b0 );
buf ( n8006 , n30372 );
buf ( n8007 , n28931 );
buf ( n8008 , 1'b0 );
buf ( n8009 , 1'b0 );
buf ( n8010 , n1 );
buf ( n8011 , n30334 );
buf ( n8012 , 1'b0 );
buf ( n8013 , 1'b0 );
buf ( n8014 , n1 );
buf ( n8015 , n30359 );
buf ( n8016 , 1'b0 );
buf ( n8017 , 1'b0 );
buf ( n8018 , n1 );
buf ( n8019 , n30365 );
buf ( n8020 , 1'b0 );
buf ( n8021 , 1'b0 );
buf ( n8022 , n30351 );
buf ( n8023 , n30400 );
buf ( n8024 , 1'b0 );
buf ( n8025 , 1'b0 );
buf ( n8026 , n1 );
buf ( n8027 , n28989 );
buf ( n8028 , 1'b0 );
buf ( n8029 , 1'b0 );
buf ( n8030 , n30353 );
buf ( n8031 , n29613 );
buf ( n8032 , 1'b0 );
buf ( n8033 , 1'b0 );
buf ( n8034 , n1 );
buf ( n8035 , n29880 );
buf ( n8036 , 1'b0 );
buf ( n8037 , 1'b0 );
buf ( n8038 , n30352 );
buf ( n8039 , n29014 );
buf ( n8040 , 1'b0 );
buf ( n8041 , 1'b0 );
buf ( n8042 , n30353 );
buf ( n8043 , n29007 );
buf ( n8044 , 1'b0 );
buf ( n8045 , 1'b0 );
buf ( n8046 , n1 );
buf ( n8047 , n28985 );
buf ( n8048 , 1'b0 );
buf ( n8049 , 1'b0 );
buf ( n8050 , n1 );
buf ( n8051 , n28982 );
buf ( n8052 , 1'b0 );
buf ( n8053 , 1'b0 );
buf ( n8054 , n1 );
buf ( n8055 , n28933 );
buf ( n8056 , 1'b0 );
buf ( n8057 , 1'b0 );
buf ( n8058 , n1 );
buf ( n8059 , n28979 );
buf ( n8060 , 1'b0 );
buf ( n8061 , 1'b0 );
buf ( n8062 , n30355 );
buf ( n8063 , n30392 );
buf ( n8064 , 1'b0 );
buf ( n8065 , 1'b0 );
buf ( n8066 , n30343 );
buf ( n8067 , n30360 );
buf ( n8068 , 1'b0 );
buf ( n8069 , 1'b0 );
buf ( n8070 , n30351 );
buf ( n8071 , n29937 );
buf ( n8072 , 1'b0 );
buf ( n8073 , 1'b0 );
buf ( n8074 , n30355 );
buf ( n8075 , n30390 );
buf ( n8076 , 1'b0 );
buf ( n8077 , 1'b0 );
buf ( n8078 , n1 );
buf ( n8079 , n29103 );
buf ( n8080 , 1'b0 );
buf ( n8081 , 1'b0 );
buf ( n8082 , n30343 );
buf ( n8083 , n30396 );
buf ( n8084 , 1'b0 );
buf ( n8085 , 1'b0 );
buf ( n8086 , n30353 );
buf ( n8087 , n27678 );
buf ( n8088 , 1'b0 );
buf ( n8089 , 1'b0 );
buf ( n8090 , n1 );
buf ( n8091 , n29404 );
buf ( n8092 , 1'b0 );
buf ( n8093 , 1'b0 );
buf ( n8094 , n1 );
buf ( n8095 , n28976 );
buf ( n8096 , 1'b0 );
buf ( n8097 , 1'b0 );
buf ( n8098 , n1 );
buf ( n8099 , n28973 );
buf ( n8100 , 1'b0 );
buf ( n8101 , 1'b0 );
buf ( n8102 , n30356 );
buf ( n8103 , n29200 );
buf ( n8104 , 1'b0 );
buf ( n8105 , 1'b0 );
buf ( n8106 , n30346 );
buf ( n8107 , n28938 );
buf ( n8108 , 1'b0 );
buf ( n8109 , 1'b0 );
buf ( n8110 , n30356 );
buf ( n8111 , n28614 );
buf ( n8112 , 1'b0 );
buf ( n8113 , 1'b0 );
buf ( n8114 , n30343 );
buf ( n8115 , n28620 );
buf ( n8116 , 1'b0 );
buf ( n8117 , 1'b0 );
buf ( n8118 , n30351 );
buf ( n8119 , n28626 );
buf ( n8120 , 1'b0 );
buf ( n8121 , 1'b0 );
buf ( n8122 , n30346 );
buf ( n8123 , n28632 );
buf ( n8124 , 1'b0 );
buf ( n8125 , 1'b0 );
buf ( n8126 , n30351 );
buf ( n8127 , n28895 );
buf ( n8128 , 1'b0 );
buf ( n8129 , 1'b0 );
buf ( n8130 , n1 );
buf ( n8131 , n29070 );
buf ( n8132 , 1'b0 );
buf ( n8133 , 1'b0 );
buf ( n8134 , n30342 );
buf ( n8135 , n29331 );
buf ( n8136 , 1'b0 );
buf ( n8137 , 1'b0 );
buf ( n8138 , n1 );
buf ( n8139 , n28970 );
buf ( n8140 , 1'b0 );
buf ( n8141 , 1'b0 );
buf ( n8142 , n1 );
buf ( n8143 , n29884 );
buf ( n8144 , 1'b0 );
buf ( n8145 , 1'b0 );
buf ( n8146 , n1 );
buf ( n8147 , n28966 );
buf ( n8148 , 1'b0 );
buf ( n8149 , 1'b0 );
buf ( n8150 , n1 );
buf ( n8151 , n28941 );
buf ( n8152 , 1'b0 );
buf ( n8153 , 1'b0 );
buf ( n8154 , n1 );
buf ( n8155 , n28878 );
buf ( n8156 , 1'b0 );
buf ( n8157 , 1'b0 );
buf ( n8158 , n1 );
buf ( n8159 , n28944 );
buf ( n8160 , 1'b0 );
buf ( n8161 , 1'b0 );
buf ( n8162 , n1 );
buf ( n8163 , n28947 );
buf ( n8164 , 1'b0 );
buf ( n8165 , 1'b0 );
buf ( n8166 , n30375 );
buf ( n8167 , n1754 );
buf ( n8168 , 1'b0 );
buf ( n8169 , 1'b0 );
buf ( n8170 , n1 );
buf ( n8171 , n1707 );
buf ( n8172 , 1'b0 );
buf ( n8173 , 1'b0 );
buf ( n8174 , n30352 );
buf ( n8175 , n29207 );
buf ( n8176 , 1'b0 );
buf ( n8177 , 1'b0 );
buf ( n8178 , n1 );
buf ( n8179 , n29791 );
buf ( n8180 , 1'b0 );
buf ( n8181 , 1'b0 );
buf ( n8182 , n30352 );
buf ( n8183 , n28300 );
buf ( n8184 , 1'b0 );
buf ( n8185 , 1'b0 );
buf ( n8186 , n30346 );
buf ( n8187 , n28709 );
buf ( n8188 , 1'b0 );
buf ( n8189 , 1'b0 );
buf ( n8190 , n1 );
buf ( n8191 , n1756 );
buf ( n8192 , 1'b0 );
buf ( n8193 , 1'b0 );
buf ( n8194 , n30378 );
buf ( n8195 , n1796 );
buf ( n8196 , 1'b0 );
buf ( n8197 , 1'b0 );
buf ( n8198 , n30358 );
buf ( n8199 , n29362 );
buf ( n8200 , 1'b0 );
buf ( n8201 , 1'b0 );
buf ( n8202 , n1 );
buf ( n8203 , n29878 );
buf ( n8204 , 1'b0 );
buf ( n8205 , 1'b0 );
buf ( n8206 , n30346 );
buf ( n8207 , n28963 );
buf ( n8208 , 1'b0 );
buf ( n8209 , 1'b0 );
buf ( n8210 , n30371 );
buf ( n8211 , n30398 );
buf ( n8212 , 1'b0 );
buf ( n8213 , 1'b0 );
buf ( n8214 , n30343 );
buf ( n8215 , n30397 );
buf ( n8216 , 1'b0 );
buf ( n8217 , 1'b0 );
buf ( n8218 , n30345 );
buf ( n8219 , n28957 );
buf ( n8220 , 1'b0 );
buf ( n8221 , 1'b0 );
buf ( n8222 , n1 );
buf ( n8223 , n29731 );
buf ( n8224 , 1'b0 );
buf ( n8225 , 1'b0 );
buf ( n8226 , n30352 );
buf ( n8227 , n29213 );
buf ( n8228 , 1'b0 );
buf ( n8229 , 1'b0 );
buf ( n8230 , n30351 );
buf ( n8231 , n29219 );
buf ( n8232 , 1'b0 );
buf ( n8233 , 1'b0 );
buf ( n8234 , n30378 );
buf ( n8235 , n29225 );
buf ( n8236 , 1'b0 );
buf ( n8237 , 1'b0 );
buf ( n8238 , n30346 );
buf ( n8239 , n29231 );
buf ( n8240 , 1'b0 );
buf ( n8241 , 1'b0 );
buf ( n8242 , n1 );
buf ( n8243 , n29796 );
buf ( n8244 , 1'b0 );
buf ( n8245 , 1'b0 );
buf ( n8246 , n1 );
buf ( n8247 , n29683 );
buf ( n8248 , 1'b0 );
buf ( n8249 , 1'b0 );
buf ( n8250 , n30343 );
buf ( n8251 , n29475 );
buf ( n8252 , 1'b0 );
buf ( n8253 , 1'b0 );
buf ( n8254 , n30353 );
buf ( n8255 , n29480 );
buf ( n8256 , 1'b0 );
buf ( n8257 , 1'b0 );
buf ( n8258 , n1 );
buf ( n8259 , n30028 );
buf ( n8260 , 1'b0 );
buf ( n8261 , 1'b0 );
buf ( n8262 , n1 );
buf ( n8263 , n30031 );
buf ( n8264 , 1'b0 );
buf ( n8265 , 1'b0 );
buf ( n8266 , n1 );
buf ( n8267 , n30041 );
buf ( n8268 , 1'b0 );
buf ( n8269 , 1'b0 );
buf ( n8270 , n30356 );
buf ( n8271 , n13561 );
buf ( n8272 , 1'b0 );
buf ( n8273 , 1'b0 );
buf ( n8274 , n30352 );
buf ( n8275 , n30032 );
buf ( n8276 , 1'b0 );
buf ( n8277 , 1'b0 );
buf ( n8278 , n30346 );
buf ( n8279 , n28301 );
buf ( n8280 , 1'b0 );
buf ( n8281 , 1'b0 );
buf ( n8282 , n30351 );
buf ( n8283 , n30033 );
buf ( n8284 , 1'b0 );
buf ( n8285 , 1'b0 );
buf ( n8286 , n30351 );
buf ( n8287 , n30037 );
buf ( n8288 , 1'b0 );
buf ( n8289 , 1'b0 );
buf ( n8290 , n30371 );
buf ( n8291 , n29658 );
buf ( n8292 , 1'b0 );
buf ( n8293 , 1'b0 );
buf ( n8294 , n30356 );
buf ( n8295 , n29663 );
buf ( n8296 , 1'b0 );
buf ( n8297 , 1'b0 );
buf ( n8298 , n30374 );
buf ( n8299 , n29485 );
buf ( n8300 , 1'b0 );
buf ( n8301 , 1'b0 );
buf ( n8302 , n30355 );
buf ( n8303 , n29673 );
buf ( n8304 , 1'b0 );
buf ( n8305 , 1'b0 );
buf ( n8306 , n30353 );
buf ( n8307 , n29602 );
buf ( n8308 , 1'b0 );
buf ( n8309 , 1'b0 );
buf ( n8310 , n30352 );
buf ( n8311 , n1083 );
buf ( n8312 , 1'b0 );
buf ( n8313 , 1'b0 );
buf ( n8314 , n30376 );
buf ( n8315 , n26358 );
buf ( n8316 , 1'b0 );
buf ( n8317 , 1'b0 );
buf ( n8318 , n30376 );
buf ( n8319 , n28487 );
buf ( n8320 , 1'b0 );
buf ( n8321 , 1'b0 );
buf ( n8322 , n30347 );
buf ( n8323 , n30325 );
buf ( n8324 , 1'b0 );
buf ( n8325 , 1'b0 );
buf ( n8326 , n30376 );
buf ( n8327 , n29885 );
buf ( n8328 , 1'b0 );
buf ( n8329 , 1'b0 );
buf ( n8330 , n1 );
buf ( n8331 , n29868 );
buf ( n8332 , 1'b0 );
buf ( n8333 , 1'b0 );
buf ( n8334 , n30375 );
buf ( n8335 , n29607 );
buf ( n8336 , 1'b0 );
buf ( n8337 , 1'b0 );
buf ( n8338 , n30372 );
buf ( n8339 , n29490 );
buf ( n8340 , 1'b0 );
buf ( n8341 , 1'b0 );
buf ( n8342 , n30340 );
buf ( n8343 , n29495 );
buf ( n8344 , 1'b0 );
buf ( n8345 , 1'b0 );
buf ( n8346 , n30356 );
buf ( n8347 , n29500 );
buf ( n8348 , 1'b0 );
buf ( n8349 , 1'b0 );
buf ( n8350 , n30340 );
buf ( n8351 , n29505 );
buf ( n8352 , 1'b0 );
buf ( n8353 , 1'b0 );
buf ( n8354 , n30348 );
buf ( n8355 , n29510 );
buf ( n8356 , 1'b0 );
buf ( n8357 , 1'b0 );
buf ( n8358 , n30340 );
buf ( n8359 , n29515 );
buf ( n8360 , 1'b0 );
buf ( n8361 , 1'b0 );
buf ( n8362 , n30340 );
buf ( n8363 , n29520 );
buf ( n8364 , 1'b0 );
buf ( n8365 , 1'b0 );
buf ( n8366 , n30340 );
buf ( n8367 , n29525 );
buf ( n8368 , 1'b0 );
buf ( n8369 , 1'b0 );
buf ( n8370 , n30348 );
buf ( n8371 , n29530 );
buf ( n8372 , 1'b0 );
buf ( n8373 , 1'b0 );
buf ( n8374 , n30357 );
buf ( n8375 , n30005 );
buf ( n8376 , 1'b0 );
buf ( n8377 , 1'b0 );
buf ( n8378 , n30354 );
buf ( n8379 , n29535 );
buf ( n8380 , 1'b0 );
buf ( n8381 , 1'b0 );
buf ( n8382 , n30357 );
buf ( n8383 , n29375 );
buf ( n8384 , 1'b0 );
buf ( n8385 , 1'b0 );
buf ( n8386 , n30377 );
buf ( n8387 , n29540 );
buf ( n8388 , 1'b0 );
buf ( n8389 , 1'b0 );
buf ( n8390 , n30348 );
buf ( n8391 , n29545 );
buf ( n8392 , 1'b0 );
buf ( n8393 , 1'b0 );
buf ( n8394 , n30357 );
buf ( n8395 , n29635 );
buf ( n8396 , 1'b0 );
buf ( n8397 , 1'b0 );
buf ( n8398 , n30349 );
buf ( n8399 , n29550 );
buf ( n8400 , 1'b0 );
buf ( n8401 , 1'b0 );
buf ( n8402 , n30349 );
buf ( n8403 , n29555 );
buf ( n8404 , 1'b0 );
buf ( n8405 , 1'b0 );
buf ( n8406 , n30377 );
buf ( n8407 , n29668 );
buf ( n8408 , 1'b0 );
buf ( n8409 , 1'b0 );
buf ( n8410 , n30373 );
buf ( n8411 , n29560 );
buf ( n8412 , 1'b0 );
buf ( n8413 , 1'b0 );
buf ( n8414 , n1 );
buf ( n8415 , n29873 );
buf ( n8416 , 1'b0 );
buf ( n8417 , 1'b0 );
buf ( n8418 , n30377 );
buf ( n8419 , n29618 );
buf ( n8420 , 1'b0 );
buf ( n8421 , 1'b0 );
buf ( n8422 , n30372 );
buf ( n8423 , n29565 );
buf ( n8424 , 1'b0 );
buf ( n8425 , 1'b0 );
buf ( n8426 , n1 );
buf ( n8427 , n29801 );
buf ( n8428 , 1'b0 );
buf ( n8429 , 1'b0 );
buf ( n8430 , n1 );
buf ( n8431 , n29704 );
buf ( n8432 , 1'b0 );
buf ( n8433 , 1'b0 );
buf ( n8434 , n30372 );
buf ( n8435 , n29570 );
buf ( n8436 , 1'b0 );
buf ( n8437 , 1'b0 );
buf ( n8438 , n30377 );
buf ( n8439 , n29575 );
buf ( n8440 , 1'b0 );
buf ( n8441 , 1'b0 );
buf ( n8442 , n1 );
buf ( n8443 , n29812 );
buf ( n8444 , 1'b0 );
buf ( n8445 , 1'b0 );
buf ( n8446 , n1 );
buf ( n8447 , n29823 );
buf ( n8448 , 1'b0 );
buf ( n8449 , 1'b0 );
buf ( n8450 , n1 );
buf ( n8451 , n29834 );
buf ( n8452 , 1'b0 );
buf ( n8453 , 1'b0 );
buf ( n8454 , n30372 );
buf ( n8455 , n29580 );
buf ( n8456 , 1'b0 );
buf ( n8457 , 1'b0 );
buf ( n8458 , n30372 );
buf ( n8459 , n29585 );
buf ( n8460 , 1'b0 );
buf ( n8461 , 1'b0 );
buf ( n8462 , n1 );
buf ( n8463 , n29726 );
buf ( n8464 , 1'b0 );
buf ( n8465 , 1'b0 );
buf ( n8466 , n1 );
buf ( n8467 , n29715 );
buf ( n8468 , 1'b0 );
buf ( n8469 , 1'b0 );
buf ( n8470 , n1 );
buf ( n8471 , n29699 );
buf ( n8472 , 1'b0 );
buf ( n8473 , 1'b0 );
buf ( n8474 , n1 );
buf ( n8475 , n29845 );
buf ( n8476 , 1'b0 );
buf ( n8477 , 1'b0 );
buf ( n8478 , n1 );
buf ( n8479 , n29856 );
buf ( n8480 , 1'b0 );
buf ( n8481 , 1'b0 );
buf ( n8482 , n30349 );
buf ( n8483 , n29623 );
buf ( n8484 , 1'b0 );
buf ( n8485 , 1'b0 );
buf ( n8486 , n30373 );
buf ( n8487 , n29978 );
buf ( n8488 , 1'b0 );
buf ( n8489 , 1'b0 );
buf ( n8490 , n30377 );
buf ( n8491 , n29947 );
buf ( n8492 , 1'b0 );
buf ( n8493 , 1'b0 );
buf ( n8494 , n30377 );
buf ( n8495 , n29949 );
buf ( n8496 , 1'b0 );
buf ( n8497 , 1'b0 );
buf ( n8498 , n30348 );
buf ( n8499 , n27714 );
buf ( n8500 , 1'b0 );
buf ( n8501 , 1'b0 );
buf ( n8502 , n30348 );
buf ( n8503 , n30361 );
buf ( n8504 , 1'b0 );
buf ( n8505 , 1'b0 );
buf ( n8506 , n30348 );
buf ( n8507 , n30337 );
buf ( n8508 , 1'b0 );
buf ( n8509 , 1'b0 );
buf ( n8510 , n30348 );
buf ( n8511 , n30364 );
buf ( n8512 , 1'b0 );
buf ( n8513 , 1'b0 );
buf ( n8514 , n30340 );
buf ( n8515 , n15647 );
buf ( n8516 , 1'b0 );
buf ( n8517 , 1'b0 );
buf ( n8518 , n30347 );
buf ( n8519 , n29925 );
buf ( n8520 , 1'b0 );
buf ( n8521 , 1'b0 );
buf ( n8522 , n30345 );
buf ( n8523 , n29930 );
buf ( n8524 , 1'b0 );
buf ( n8525 , 1'b0 );
buf ( n8526 , n30358 );
buf ( n8527 , n29236 );
buf ( n8528 , 1'b0 );
buf ( n8529 , 1'b0 );
buf ( n8530 , n30374 );
buf ( n8531 , n29241 );
buf ( n8532 , 1'b0 );
buf ( n8533 , 1'b0 );
buf ( n8534 , n30378 );
buf ( n8535 , n29246 );
buf ( n8536 , 1'b0 );
buf ( n8537 , 1'b0 );
buf ( n8538 , n30351 );
buf ( n8539 , n29251 );
buf ( n8540 , 1'b0 );
buf ( n8541 , 1'b0 );
buf ( n8542 , n30355 );
buf ( n8543 , n29256 );
buf ( n8544 , 1'b0 );
buf ( n8545 , 1'b0 );
buf ( n8546 , n1 );
buf ( n8547 , n30036 );
buf ( n8548 , 1'b0 );
buf ( n8549 , 1'b0 );
buf ( n8550 , n30345 );
buf ( n8551 , n29261 );
buf ( n8552 , 1'b0 );
buf ( n8553 , 1'b0 );
buf ( n8554 , n30351 );
buf ( n8555 , n29266 );
buf ( n8556 , 1'b0 );
buf ( n8557 , 1'b0 );
buf ( n8558 , n30343 );
buf ( n8559 , n29271 );
buf ( n8560 , 1'b0 );
buf ( n8561 , 1'b0 );
buf ( n8562 , n30358 );
buf ( n8563 , n29276 );
buf ( n8564 , 1'b0 );
buf ( n8565 , 1'b0 );
buf ( n8566 , n30356 );
buf ( n8567 , n29101 );
buf ( n8568 , 1'b0 );
buf ( n8569 , 1'b0 );
buf ( n8570 , n30353 );
buf ( n8571 , n29109 );
buf ( n8572 , 1'b0 );
buf ( n8573 , 1'b0 );
buf ( n8574 , n30342 );
buf ( n8575 , n29281 );
buf ( n8576 , 1'b0 );
buf ( n8577 , 1'b0 );
buf ( n8578 , n30375 );
buf ( n8579 , n29286 );
buf ( n8580 , 1'b0 );
buf ( n8581 , 1'b0 );
buf ( n8582 , n30378 );
buf ( n8583 , n29291 );
buf ( n8584 , 1'b0 );
buf ( n8585 , 1'b0 );
buf ( n8586 , n30378 );
buf ( n8587 , n29296 );
buf ( n8588 , 1'b0 );
buf ( n8589 , 1'b0 );
buf ( n8590 , n30346 );
buf ( n8591 , n29301 );
buf ( n8592 , 1'b0 );
buf ( n8593 , 1'b0 );
buf ( n8594 , n30343 );
buf ( n8595 , n29306 );
buf ( n8596 , 1'b0 );
buf ( n8597 , 1'b0 );
buf ( n8598 , n30352 );
buf ( n8599 , n29193 );
buf ( n8600 , 1'b0 );
buf ( n8601 , 1'b0 );
buf ( n8602 , n30352 );
buf ( n8603 , n29188 );
buf ( n8604 , 1'b0 );
buf ( n8605 , 1'b0 );
buf ( n8606 , n30343 );
buf ( n8607 , n29183 );
buf ( n8608 , 1'b0 );
buf ( n8609 , 1'b0 );
buf ( n8610 , n30352 );
buf ( n8611 , n29178 );
buf ( n8612 , 1'b0 );
buf ( n8613 , 1'b0 );
buf ( n8614 , n30375 );
buf ( n8615 , n29166 );
buf ( n8616 , 1'b0 );
buf ( n8617 , 1'b0 );
buf ( n8618 , n30353 );
buf ( n8619 , n29161 );
buf ( n8620 , 1'b0 );
buf ( n8621 , 1'b0 );
buf ( n8622 , n30358 );
buf ( n8623 , n29156 );
buf ( n8624 , 1'b0 );
buf ( n8625 , 1'b0 );
buf ( n8626 , n30356 );
buf ( n8627 , n29151 );
buf ( n8628 , 1'b0 );
buf ( n8629 , 1'b0 );
buf ( n8630 , n30355 );
buf ( n8631 , n29146 );
buf ( n8632 , 1'b0 );
buf ( n8633 , 1'b0 );
buf ( n8634 , n30345 );
buf ( n8635 , n29141 );
buf ( n8636 , 1'b0 );
buf ( n8637 , 1'b0 );
buf ( n8638 , n30358 );
buf ( n8639 , n29136 );
buf ( n8640 , 1'b0 );
buf ( n8641 , 1'b0 );
buf ( n8642 , n30355 );
buf ( n8643 , n29131 );
buf ( n8644 , 1'b0 );
buf ( n8645 , 1'b0 );
buf ( n8646 , n30357 );
buf ( n8647 , n29126 );
buf ( n8648 , 1'b0 );
buf ( n8649 , 1'b0 );
buf ( n8650 , n30348 );
buf ( n8651 , n29120 );
buf ( n8652 , 1'b0 );
buf ( n8653 , 1'b0 );
buf ( n8654 , n30340 );
buf ( n8655 , n29114 );
buf ( n8656 , 1'b0 );
buf ( n8657 , 1'b0 );
buf ( n8658 , n30373 );
buf ( n8659 , n29327 );
buf ( n8660 , 1'b0 );
buf ( n8661 , 1'b0 );
buf ( n8662 , n30354 );
buf ( n8663 , n30303 );
buf ( n8664 , 1'b0 );
buf ( n8665 , 1'b0 );
buf ( n8666 , n30348 );
buf ( n8667 , n30108 );
buf ( n8668 , 1'b0 );
buf ( n8669 , 1'b0 );
buf ( n8670 , n30354 );
buf ( n8671 , n19375 );
buf ( n8672 , 1'b0 );
buf ( n8673 , 1'b0 );
buf ( n8674 , n30349 );
buf ( n8675 , n30038 );
buf ( n8676 , 1'b0 );
buf ( n8677 , 1'b0 );
buf ( n8678 , n30373 );
buf ( n8679 , n29858 );
buf ( n8680 , 1'b0 );
buf ( n8681 , 1'b0 );
buf ( n8682 , n30372 );
buf ( n8683 , n29933 );
buf ( n8684 , 1'b0 );
buf ( n8685 , 1'b0 );
buf ( n8686 , n30377 );
buf ( n8687 , n30363 );
buf ( n8688 , 1'b0 );
buf ( n8689 , 1'b0 );
buf ( n8690 , n30349 );
buf ( n8691 , n29935 );
buf ( n8692 , 1'b0 );
buf ( n8693 , 1'b0 );
buf ( n8694 , n30349 );
buf ( n8695 , n20055 );
buf ( n8696 , 1'b0 );
buf ( n8697 , 1'b0 );
buf ( n8698 , n1 );
buf ( n8699 , n1809 );
buf ( n8700 , 1'b0 );
buf ( n8701 , 1'b0 );
buf ( n8702 , n1 );
buf ( n8703 , n1855 );
buf ( n8704 , 1'b0 );
buf ( n8705 , 1'b0 );
buf ( n8706 , n30349 );
buf ( n8707 , n21342 );
buf ( n8708 , 1'b0 );
buf ( n8709 , 1'b0 );
buf ( n8710 , n1 );
buf ( n8711 , n17011 );
buf ( n8712 , 1'b0 );
buf ( n8713 , 1'b0 );
buf ( n8714 , n30348 );
buf ( n8715 , n1859 );
buf ( n8716 , 1'b0 );
buf ( n8717 , 1'b0 );
buf ( n8718 , n1 );
buf ( n8719 , n1167 );
buf ( n8720 , 1'b0 );
buf ( n8721 , 1'b0 );
buf ( n8722 , n1 );
buf ( n8723 , n1848 );
buf ( n8724 , 1'b0 );
buf ( n8725 , 1'b0 );
buf ( n8726 , n1 );
buf ( n8727 , n1852 );
buf ( n8728 , 1'b0 );
buf ( n8729 , 1'b0 );
buf ( n8730 , n30357 );
buf ( n8731 , n1853 );
buf ( n8732 , 1'b0 );
buf ( n8733 , 1'b0 );
buf ( n8734 , n1 );
buf ( n8735 , n1849 );
buf ( n8736 , 1'b0 );
buf ( n8737 , 1'b0 );
buf ( n8738 , n1 );
buf ( n8739 , n1865 );
buf ( n8740 , 1'b0 );
buf ( n8741 , 1'b0 );
buf ( n8742 , n1 );
buf ( n8743 , n1861 );
buf ( n8744 , 1'b0 );
buf ( n8745 , 1'b0 );
buf ( n8746 , n1 );
buf ( n8747 , n1874 );
buf ( n8748 , 1'b0 );
buf ( n8749 , 1'b0 );
buf ( n8750 , n30347 );
buf ( n8751 , n30338 );
buf ( n8752 , 1'b0 );
buf ( n8753 , 1'b0 );
buf ( n8754 , n1 );
buf ( n8755 , n1859 );
buf ( n8756 , 1'b0 );
buf ( n8757 , 1'b0 );
buf ( n8758 , n30378 );
buf ( n8759 , n1863 );
buf ( n8760 , 1'b0 );
buf ( n8761 , 1'b0 );
buf ( n8762 , n1 );
buf ( n8763 , n1863 );
buf ( n8764 , 1'b0 );
buf ( n8765 , 1'b0 );
buf ( n8766 , n30374 );
buf ( n8767 , n74 );
buf ( n8768 , 1'b0 );
buf ( n8769 , 1'b0 );
buf ( n8770 , n1 );
buf ( n8771 , n1873 );
buf ( n8772 , 1'b0 );
buf ( n8773 , 1'b0 );
buf ( n8774 , n1 );
buf ( n8775 , n1872 );
buf ( n8776 , 1'b0 );
buf ( n8777 , 1'b0 );
buf ( n8778 , n30355 );
buf ( n8779 , n241 );
buf ( n8780 , 1'b0 );
buf ( n8781 , 1'b0 );
buf ( n8782 , n1 );
buf ( n8783 , n1857 );
buf ( n8784 , 1'b0 );
buf ( n8785 , 1'b0 );
buf ( n8786 , n30376 );
buf ( n8787 , n1872 );
buf ( n8788 , 1'b0 );
buf ( n8789 , 1'b0 );
buf ( n8790 , n30358 );
buf ( n8791 , n241 );
buf ( n8792 , 1'b0 );
buf ( n8793 , 1'b0 );
buf ( n8794 , n30353 );
buf ( n8795 , n1857 );
buf ( n8796 , 1'b0 );
buf ( n8797 , 1'b0 );
buf ( n8798 , n1 );
buf ( n8799 , n1850 );
buf ( n8800 , 1'b0 );
buf ( n8801 , 1'b0 );
buf ( n8802 , n1 );
buf ( n8803 , n1167 );
buf ( n8804 , 1'b0 );
buf ( n8805 , 1'b0 );
buf ( n8806 , n1 );
buf ( n8807 , n16941 );
buf ( n8808 , 1'b0 );
buf ( n8809 , 1'b0 );
buf ( n8810 , n1 );
buf ( n8811 , n17081 );
buf ( n8812 , 1'b0 );
buf ( n8813 , 1'b0 );
buf ( n8814 , n1 );
buf ( n8815 , n16868 );
buf ( n8816 , 1'b0 );
buf ( n8817 , 1'b0 );
buf ( n8818 , n30342 );
buf ( n8819 , n29202 );
buf ( n8820 , 1'b0 );
buf ( n8821 , 1'b0 );
buf ( n8822 , n30351 );
buf ( n8823 , n1555 );
buf ( n8824 , 1'b0 );
buf ( n8825 , 1'b0 );
buf ( n8826 , n30343 );
buf ( n8827 , n1557 );
buf ( n8828 , 1'b0 );
buf ( n8829 , 1'b0 );
buf ( n8830 , n30346 );
buf ( n8831 , n1554 );
buf ( n8832 , 1'b0 );
buf ( n8833 , 1'b0 );
buf ( n8834 , n30352 );
buf ( n8835 , n1073 );
buf ( n8836 , 1'b0 );
buf ( n8837 , 1'b0 );
buf ( n8838 , n30371 );
buf ( n8839 , n1548 );
buf ( n8840 , 1'b0 );
buf ( n8841 , 1'b0 );
buf ( n8842 , n30353 );
buf ( n8843 , n1065 );
buf ( n8844 , 1'b0 );
buf ( n8845 , 1'b0 );
buf ( n8846 , n30347 );
buf ( n8847 , n1072 );
buf ( n8848 , 1'b0 );
buf ( n8849 , 1'b0 );
buf ( n8850 , n30374 );
buf ( n8851 , n1061 );
buf ( n8852 , 1'b0 );
buf ( n8853 , 1'b0 );
buf ( n8854 , n30340 );
buf ( n8855 , n1062 );
buf ( n8856 , 1'b0 );
buf ( n8857 , 1'b0 );
buf ( n8858 , n30373 );
buf ( n8859 , n1552 );
buf ( n8860 , 1'b0 );
buf ( n8861 , 1'b0 );
buf ( n8862 , n30348 );
buf ( n8863 , n1060 );
buf ( n8864 , 1'b0 );
buf ( n8865 , 1'b0 );
buf ( n8866 , n30348 );
buf ( n8867 , n1063 );
buf ( n8868 , 1'b0 );
buf ( n8869 , 1'b0 );
buf ( n8870 , n30372 );
buf ( n8871 , n1064 );
buf ( n8872 , 1'b0 );
buf ( n8873 , 1'b0 );
buf ( n8874 , n30357 );
buf ( n8875 , n91 );
buf ( n8876 , 1'b0 );
buf ( n8877 , 1'b0 );
buf ( n8878 , n30348 );
buf ( n8879 , n95 );
buf ( n8880 , 1'b0 );
buf ( n8881 , 1'b0 );
buf ( n8882 , n30340 );
buf ( n8883 , n93 );
buf ( n8884 , 1'b0 );
buf ( n8885 , 1'b0 );
buf ( n8886 , n30378 );
buf ( n8887 , n83 );
buf ( n8888 , 1'b0 );
buf ( n8889 , 1'b0 );
buf ( n8890 , n30378 );
buf ( n8891 , n94 );
buf ( n8892 , 1'b0 );
buf ( n8893 , 1'b0 );
buf ( n8894 , n30351 );
buf ( n8895 , n923 );
buf ( n8896 , 1'b0 );
buf ( n8897 , 1'b0 );
buf ( n8898 , n30342 );
buf ( n8899 , n78 );
buf ( n8900 , 1'b0 );
buf ( n8901 , 1'b0 );
buf ( n8902 , n1 );
buf ( n8903 , n1586 );
buf ( n8904 , 1'b0 );
buf ( n8905 , 1'b0 );
buf ( n8906 , n30378 );
buf ( n8907 , n82 );
buf ( n8908 , 1'b0 );
buf ( n8909 , 1'b0 );
buf ( n8910 , n30371 );
buf ( n8911 , n1691 );
buf ( n8912 , 1'b0 );
buf ( n8913 , 1'b0 );
buf ( n8914 , n30374 );
buf ( n8915 , n1228 );
buf ( n8916 , 1'b0 );
buf ( n8917 , 1'b0 );
buf ( n8918 , n30348 );
buf ( n8919 , n1685 );
buf ( n8920 , 1'b0 );
buf ( n8921 , 1'b0 );
buf ( n8922 , n30348 );
buf ( n8923 , n87 );
buf ( n8924 , 1'b0 );
buf ( n8925 , 1'b0 );
buf ( n8926 , n30348 );
buf ( n8927 , n92 );
buf ( n8928 , 1'b0 );
buf ( n8929 , 1'b0 );
buf ( n8930 , n30354 );
buf ( n8931 , n85 );
buf ( n8932 , 1'b0 );
buf ( n8933 , 1'b0 );
buf ( n8934 , n30340 );
buf ( n8935 , n1690 );
buf ( n8936 , 1'b0 );
buf ( n8937 , 1'b0 );
buf ( n8938 , n30378 );
buf ( n8939 , n80 );
buf ( n8940 , 1'b0 );
buf ( n8941 , 1'b0 );
buf ( n8942 , n30352 );
buf ( n8943 , n89 );
buf ( n8944 , 1'b0 );
buf ( n8945 , 1'b0 );
buf ( n8946 , n30353 );
buf ( n8947 , n86 );
buf ( n8948 , 1'b0 );
buf ( n8949 , 1'b0 );
buf ( n8950 , n30340 );
buf ( n8951 , n79 );
buf ( n8952 , 1'b0 );
buf ( n8953 , 1'b0 );
buf ( n8954 , n30357 );
buf ( n8955 , n87 );
buf ( n8956 , 1'b0 );
buf ( n8957 , 1'b0 );
buf ( n8958 , n30357 );
buf ( n8959 , n81 );
buf ( n8960 , 1'b0 );
buf ( n8961 , 1'b0 );
buf ( n8962 , n30352 );
buf ( n8963 , n84 );
buf ( n8964 , 1'b0 );
buf ( n8965 , 1'b0 );
buf ( n8966 , n30375 );
buf ( n8967 , n86 );
buf ( n8968 , 1'b0 );
buf ( n8969 , 1'b0 );
buf ( n8970 , n30340 );
buf ( n8971 , n1680 );
buf ( n8972 , 1'b0 );
buf ( n8973 , 1'b0 );
buf ( n8974 , n30355 );
buf ( n8975 , n90 );
buf ( n8976 , 1'b0 );
buf ( n8977 , 1'b0 );
buf ( n8978 , n30357 );
buf ( n8979 , n96 );
not ( n12487 , n999 );
not ( n12488 , n1228 );
or ( n12489 , n12487 , n12488 );
not ( n12490 , n994 );
not ( n12491 , n319 );
not ( n12492 , n930 );
nand ( n12493 , n900 , n12492 );
not ( n12494 , n12493 );
not ( n12495 , n900 );
not ( n12496 , n930 );
nand ( n12497 , n12495 , n12496 );
not ( n12498 , n12497 );
nand ( n12499 , n1622 , n12498 );
not ( n12500 , n12499 );
or ( n12501 , n12494 , n12500 );
not ( n12502 , n925 );
nor ( n12503 , n12502 , n12498 );
nand ( n12504 , n12501 , n12503 );
not ( n12505 , n12504 );
not ( n12506 , n12505 );
not ( n12507 , n1587 );
not ( n12508 , n12497 );
not ( n12509 , n12508 );
or ( n12510 , n12507 , n12509 );
not ( n12511 , n900 );
nand ( n12512 , n930 , n12511 );
nand ( n12513 , n12510 , n12512 );
not ( n12514 , n12513 );
buf ( n12515 , n12514 );
not ( n12516 , n12515 );
nand ( n12517 , n12506 , n12516 );
not ( n12518 , n12517 );
buf ( n12519 , n12518 );
not ( n12520 , n12519 );
or ( n12521 , n12491 , n12520 );
not ( n12522 , n993 );
nand ( n12523 , n12521 , n12522 );
not ( n12524 , n12505 );
not ( n12525 , n12524 );
not ( n12526 , n12525 );
not ( n12527 , n318 );
not ( n12528 , n12515 );
not ( n12529 , n12528 );
nor ( n12530 , n12527 , n12529 );
not ( n12531 , n12530 );
buf ( n12532 , n12513 );
not ( n12533 , n12532 );
buf ( n12534 , n12533 );
nand ( n12535 , n365 , n12534 );
nand ( n12536 , n12531 , n12535 );
and ( n12537 , n12526 , n12536 );
not ( n12538 , n1006 );
not ( n12539 , n12525 );
nor ( n12540 , n12538 , n12539 );
nor ( n12541 , n12537 , n12540 );
not ( n12542 , n12541 );
and ( n12543 , n868 , n12542 );
and ( n12544 , n12523 , n12543 );
not ( n12545 , n993 );
nand ( n12546 , n319 , n12519 );
nor ( n12547 , n12545 , n12546 );
nor ( n12548 , n12544 , n12547 );
not ( n12549 , n868 );
nand ( n12550 , n12549 , n12541 );
and ( n12551 , n12523 , n12550 );
not ( n12552 , n1004 );
nand ( n12553 , n264 , n12518 );
not ( n12554 , n12524 );
nand ( n12555 , n888 , n12554 );
not ( n12556 , n12504 );
not ( n12557 , n12556 );
nand ( n12558 , n12533 , n12557 );
not ( n12559 , n12558 );
nand ( n12560 , n372 , n12559 );
nand ( n12561 , n12552 , n12553 , n12555 , n12560 );
not ( n12562 , n12561 );
not ( n12563 , n998 );
nand ( n12564 , n263 , n12518 );
nand ( n12565 , n939 , n12554 );
nand ( n12566 , n353 , n12559 );
and ( n12567 , n12563 , n12564 , n12565 , n12566 );
not ( n12568 , n12567 );
not ( n12569 , n12517 );
nand ( n12570 , n262 , n12569 );
nand ( n12571 , n937 , n12525 );
nand ( n12572 , n370 , n12559 );
nand ( n12573 , n12570 , n12571 , n12572 );
nand ( n12574 , n996 , n12573 );
not ( n12575 , n997 );
not ( n12576 , n12517 );
nand ( n12577 , n12576 , n261 );
nand ( n12578 , n938 , n12525 );
not ( n12579 , n12558 );
nand ( n12580 , n12579 , n371 );
nand ( n12581 , n12575 , n12577 , n12578 , n12580 );
not ( n12582 , n12581 );
or ( n12583 , n12574 , n12582 );
nand ( n12584 , n12577 , n12578 , n12580 );
nand ( n12585 , n997 , n12584 );
nand ( n12586 , n12583 , n12585 );
and ( n12587 , n12568 , n12586 );
nand ( n12588 , n12564 , n12565 , n12566 );
nand ( n12589 , n998 , n12588 );
not ( n12590 , n12589 );
nor ( n12591 , n12587 , n12590 );
or ( n12592 , n12562 , n12591 );
nand ( n12593 , n12553 , n12555 , n12560 );
nand ( n12594 , n1004 , n12593 );
nand ( n12595 , n12592 , n12594 );
nand ( n12596 , n12551 , n12595 );
and ( n12597 , n12548 , n12596 );
not ( n12598 , n903 );
nand ( n12599 , n320 , n12518 );
nand ( n12600 , n12598 , n12599 );
not ( n12601 , n869 );
nand ( n12602 , n321 , n12519 );
nand ( n12603 , n12601 , n12602 );
nand ( n12604 , n12600 , n12603 );
nor ( n12605 , n12597 , n12604 );
not ( n12606 , n12605 );
not ( n12607 , n12599 );
and ( n12608 , n903 , n12607 );
and ( n12609 , n12603 , n12608 );
not ( n12610 , n12602 );
and ( n12611 , n869 , n12610 );
nor ( n12612 , n12609 , n12611 );
not ( n12613 , n12551 );
nor ( n12614 , n12613 , n12604 );
not ( n12615 , n996 );
not ( n12616 , n12573 );
nand ( n12617 , n12615 , n12616 );
not ( n12618 , n12581 );
not ( n12619 , n12618 );
nand ( n12620 , n12617 , n12619 );
not ( n12621 , n12562 );
nand ( n12622 , n12621 , n12568 );
nor ( n12623 , n12620 , n12622 );
not ( n12624 , n12557 );
nand ( n12625 , n936 , n12624 );
not ( n12626 , n12625 );
not ( n12627 , n12532 );
not ( n12628 , n12627 );
nand ( n12629 , n317 , n12628 );
nand ( n12630 , n369 , n12515 );
and ( n12631 , n12629 , n12630 );
not ( n12632 , n12524 );
nor ( n12633 , n12631 , n12632 );
nor ( n12634 , n12626 , n12633 );
not ( n12635 , n12634 );
nand ( n12636 , n871 , n12635 );
not ( n12637 , n12636 );
nand ( n12638 , n280 , n12528 );
not ( n12639 , n12638 );
not ( n12640 , n350 );
not ( n12641 , n12533 );
nor ( n12642 , n12640 , n12641 );
nor ( n12643 , n12639 , n12642 );
or ( n12644 , n12554 , n12643 );
nand ( n12645 , n884 , n12624 );
nand ( n12646 , n12644 , n12645 );
nor ( n12647 , n1074 , n12646 );
not ( n12648 , n12647 );
and ( n12649 , n12637 , n12648 );
and ( n12650 , n1074 , n12646 );
nor ( n12651 , n12649 , n12650 );
not ( n12652 , n871 );
nand ( n12653 , n12652 , n12634 );
not ( n12654 , n12653 );
nor ( n12655 , n12647 , n12654 );
not ( n12656 , n1069 );
not ( n12657 , n12557 );
not ( n12658 , n279 );
or ( n12659 , n12658 , n12514 );
nand ( n12660 , n367 , n12514 );
nand ( n12661 , n12659 , n12660 );
not ( n12662 , n12661 );
or ( n12663 , n12657 , n12662 );
nand ( n12664 , n933 , n12505 );
nand ( n12665 , n12663 , n12664 );
not ( n12666 , n12665 );
nand ( n12667 , n12656 , n12666 );
not ( n12668 , n12556 );
not ( n12669 , n12668 );
not ( n12670 , n277 );
not ( n12671 , n12513 );
or ( n12672 , n12670 , n12671 );
not ( n12673 , n12513 );
nand ( n12674 , n366 , n12673 );
nand ( n12675 , n12672 , n12674 );
not ( n12676 , n12675 );
or ( n12677 , n12669 , n12676 );
nand ( n12678 , n879 , n12556 );
nand ( n12679 , n12677 , n12678 );
nand ( n12680 , n1075 , n12679 );
not ( n12681 , n12504 );
not ( n12682 , n316 );
not ( n12683 , n12513 );
or ( n12684 , n12682 , n12683 );
not ( n12685 , n12513 );
nand ( n12686 , n12685 , n386 );
nand ( n12687 , n12684 , n12686 );
not ( n12688 , n12687 );
or ( n12689 , n12681 , n12688 );
nand ( n12690 , n988 , n12556 );
nand ( n12691 , n12689 , n12690 );
nand ( n12692 , n1024 , n12691 );
not ( n12693 , n12692 );
not ( n12694 , n12679 );
not ( n12695 , n1075 );
nand ( n12696 , n12694 , n12695 );
nand ( n12697 , n12693 , n12696 );
nand ( n12698 , n12680 , n12697 );
and ( n12699 , n12667 , n12698 );
not ( n12700 , n12666 );
nand ( n12701 , n1069 , n12700 );
not ( n12702 , n12701 );
nor ( n12703 , n12699 , n12702 );
not ( n12704 , n12524 );
not ( n12705 , n278 );
or ( n12706 , n12705 , n12533 );
nand ( n12707 , n368 , n12627 );
nand ( n12708 , n12706 , n12707 );
not ( n12709 , n12708 );
or ( n12710 , n12704 , n12709 );
nand ( n12711 , n935 , n12624 );
nand ( n12712 , n12710 , n12711 );
nor ( n12713 , n870 , n12712 );
or ( n12714 , n12703 , n12713 );
nand ( n12715 , n870 , n12712 );
nand ( n12716 , n12714 , n12715 );
nand ( n12717 , n12655 , n12716 );
nand ( n12718 , n12651 , n12717 );
nand ( n12719 , n12623 , n12718 );
not ( n12720 , n12719 );
nand ( n12721 , n12614 , n12720 );
nand ( n12722 , n12606 , n12612 , n12721 );
not ( n12723 , n12722 );
nor ( n12724 , n12490 , n12723 );
or ( n12725 , n994 , n12722 );
not ( n12726 , n1228 );
nand ( n12727 , n12725 , n12726 );
or ( n12728 , n12724 , n12727 );
nand ( n12729 , n12489 , n12728 );
not ( n12730 , n904 );
nand ( n12731 , n994 , n995 );
nor ( n12732 , n12731 , n12604 );
not ( n12733 , n12732 );
not ( n12734 , n12551 );
or ( n12735 , n12589 , n12562 );
nand ( n12736 , n12735 , n12594 );
not ( n12737 , n12736 );
or ( n12738 , n12734 , n12737 );
nand ( n12739 , n12738 , n12548 );
not ( n12740 , n12739 );
or ( n12741 , n12733 , n12740 );
not ( n12742 , n12732 );
not ( n12743 , n12622 );
nand ( n12744 , n12551 , n12743 );
nor ( n12745 , n12742 , n12744 );
not ( n12746 , n12586 );
not ( n12747 , n12651 );
not ( n12748 , n12717 );
or ( n12749 , n12747 , n12748 );
not ( n12750 , n12620 );
nand ( n12751 , n12749 , n12750 );
nand ( n12752 , n12746 , n12751 );
and ( n12753 , n12745 , n12752 );
nor ( n12754 , n12731 , n12612 );
nor ( n12755 , n12753 , n12754 );
nand ( n12756 , n12741 , n12755 );
not ( n12757 , n12756 );
nor ( n12758 , n12730 , n12757 );
or ( n12759 , n904 , n12756 );
nand ( n12760 , n12759 , n12726 );
or ( n12761 , n12758 , n12760 );
not ( n12762 , n946 );
or ( n12763 , n12762 , n12726 );
nand ( n12764 , n12761 , n12763 );
nand ( n12765 , n944 , n1228 );
not ( n12766 , n12611 );
nand ( n12767 , n12766 , n12603 );
nand ( n12768 , n12523 , n12600 );
not ( n12769 , n12768 );
not ( n12770 , n12550 );
not ( n12771 , n12770 );
nand ( n12772 , n12771 , n12561 );
not ( n12773 , n12772 );
not ( n12774 , n12773 );
nor ( n12775 , n12567 , n12618 );
not ( n12776 , n12775 );
not ( n12777 , n12650 );
not ( n12778 , n12617 );
or ( n12779 , n12777 , n12778 );
nand ( n12780 , n12779 , n12574 );
not ( n12781 , n12780 );
or ( n12782 , n12776 , n12781 );
not ( n12783 , n12585 );
and ( n12784 , n12783 , n12568 );
nor ( n12785 , n12784 , n12590 );
nand ( n12786 , n12782 , n12785 );
not ( n12787 , n12786 );
or ( n12788 , n12774 , n12787 );
not ( n12789 , n12770 );
not ( n12790 , n12594 );
and ( n12791 , n12789 , n12790 );
nor ( n12792 , n12791 , n12543 );
nand ( n12793 , n12788 , n12792 );
nand ( n12794 , n12769 , n12793 );
and ( n12795 , n12600 , n12547 );
nor ( n12796 , n12795 , n12608 );
not ( n12797 , n12617 );
not ( n12798 , n12648 );
nor ( n12799 , n12797 , n12798 );
nand ( n12800 , n12799 , n12775 );
not ( n12801 , n12715 );
nand ( n12802 , n12801 , n12653 );
nand ( n12803 , n12636 , n12802 );
nor ( n12804 , n12713 , n12654 );
not ( n12805 , n12680 );
not ( n12806 , n12805 );
not ( n12807 , n12667 );
or ( n12808 , n12806 , n12807 );
nand ( n12809 , n12808 , n12701 );
not ( n12810 , n12809 );
not ( n12811 , n12697 );
nand ( n12812 , n12667 , n12811 );
nand ( n12813 , n12810 , n12812 );
nand ( n12814 , n12804 , n12813 );
not ( n12815 , n12814 );
nor ( n12816 , n12803 , n12815 );
nor ( n12817 , n12800 , n12816 );
nand ( n12818 , n12773 , n12769 , n12817 );
nand ( n12819 , n12794 , n12796 , n12818 );
nand ( n12820 , n12726 , n12767 , n12819 );
not ( n12821 , n12767 );
not ( n12822 , n12819 );
nand ( n12823 , n12726 , n12821 , n12822 );
nand ( n12824 , n12765 , n12820 , n12823 );
not ( n12825 , n138 );
not ( n12826 , n1754 );
or ( n12827 , n12826 , n195 , n1671 );
nand ( n12828 , n184 , n187 , n1821 );
not ( n12829 , n12828 );
buf ( n12830 , n12829 );
not ( n12831 , n190 );
not ( n12832 , n1558 );
nor ( n12833 , n184 , n188 );
and ( n12834 , n12832 , n12833 );
nand ( n12835 , n1551 , n12831 , n12834 );
nor ( n12836 , n1821 , n12835 );
not ( n12837 , n12836 );
not ( n12838 , n1551 );
nand ( n12839 , n12838 , n190 , n12834 );
and ( n12840 , n187 , n1821 );
nor ( n12841 , n225 , n1147 );
nand ( n12842 , n12840 , n12841 );
not ( n12843 , n12842 );
not ( n12844 , n188 );
nor ( n12845 , n190 , n1551 );
and ( n12846 , n12844 , n184 , n12832 , n12845 );
nand ( n12847 , n12843 , n12846 );
nand ( n12848 , n12837 , n12839 , n12847 );
not ( n12849 , n12848 );
buf ( n12850 , n12849 );
nand ( n12851 , n12830 , n12850 );
and ( n12852 , n12827 , n12851 );
buf ( n12853 , n12852 );
buf ( n12854 , n12853 );
not ( n12855 , n12854 );
not ( n12856 , n12855 );
not ( n12857 , n12856 );
nor ( n12858 , n12825 , n12857 );
not ( n12859 , n12858 );
not ( n12860 , n1713 );
not ( n12861 , n322 );
not ( n12862 , n12861 );
not ( n12863 , n1003 );
nand ( n12864 , n12828 , n12863 );
not ( n12865 , n12864 );
not ( n12866 , n12865 );
or ( n12867 , n12862 , n12866 );
nand ( n12868 , n281 , n328 );
nand ( n12869 , n322 , n12868 );
nand ( n12870 , n281 , n328 );
not ( n12871 , n12870 );
nand ( n12872 , n12861 , n12871 );
nand ( n12873 , n12869 , n12872 , n12864 );
nand ( n12874 , n12867 , n12873 );
buf ( n12875 , n12874 );
not ( n12876 , n12875 );
not ( n12877 , n281 );
nand ( n12878 , n328 , n12877 );
not ( n12879 , n328 );
nand ( n12880 , n281 , n12879 );
nand ( n12881 , n12878 , n12880 );
or ( n12882 , n12865 , n12881 );
nand ( n12883 , n12879 , n12865 );
nand ( n12884 , n12882 , n12883 );
not ( n12885 , n12884 );
not ( n12886 , n12877 );
not ( n12887 , n12864 );
or ( n12888 , n12886 , n12887 );
nand ( n12889 , n12865 , n281 );
nand ( n12890 , n12888 , n12889 );
nand ( n12891 , n12876 , n12885 , n12890 );
not ( n12892 , n12891 );
not ( n12893 , n12892 );
or ( n12894 , n12860 , n12893 );
not ( n12895 , n12874 );
not ( n12896 , n12895 );
not ( n12897 , n12890 );
and ( n12898 , n12865 , n12879 );
not ( n12899 , n12865 );
not ( n12900 , n12881 );
and ( n12901 , n12899 , n12900 );
nor ( n12902 , n12898 , n12901 );
not ( n12903 , n12902 );
nand ( n12904 , n12896 , n12897 , n12903 );
not ( n12905 , n12904 );
nand ( n12906 , n12905 , n1761 );
nand ( n12907 , n12894 , n12906 );
not ( n12908 , n1769 );
not ( n12909 , n12890 );
nand ( n12910 , n12909 , n12885 , n12875 );
not ( n12911 , n12910 );
not ( n12912 , n12911 );
or ( n12913 , n12908 , n12912 );
and ( n12914 , n12897 , n12885 , n12895 );
nand ( n12915 , n1720 , n12914 );
nand ( n12916 , n12913 , n12915 );
nor ( n12917 , n12907 , n12916 );
not ( n12918 , n12890 );
not ( n12919 , n12918 );
not ( n12920 , n12895 );
nand ( n12921 , n12919 , n12903 , n12920 );
not ( n12922 , n12921 );
nand ( n12923 , n1770 , n12922 );
not ( n12924 , n1718 );
not ( n12925 , n12875 );
and ( n12926 , n12897 , n12903 , n12925 );
not ( n12927 , n12926 );
or ( n12928 , n12924 , n12927 );
not ( n12929 , n12875 );
nand ( n12930 , n12929 , n12903 , n12890 );
not ( n12931 , n12930 );
nand ( n12932 , n1739 , n12931 );
nand ( n12933 , n12928 , n12932 );
not ( n12934 , n12933 );
not ( n12935 , n12897 );
and ( n12936 , n12935 , n12885 , n12920 );
nand ( n12937 , n1777 , n12936 );
nand ( n12938 , n12917 , n12923 , n12934 , n12937 );
not ( n12939 , n12938 );
not ( n12940 , n1793 );
not ( n12941 , n12921 );
not ( n12942 , n12941 );
or ( n12943 , n12940 , n12942 );
nand ( n12944 , n1774 , n12905 );
nand ( n12945 , n12943 , n12944 );
not ( n12946 , n1773 );
not ( n12947 , n12897 );
not ( n12948 , n12895 );
and ( n12949 , n12947 , n12885 , n12948 );
not ( n12950 , n12949 );
or ( n12951 , n12946 , n12950 );
nand ( n12952 , n1767 , n12911 );
nand ( n12953 , n12951 , n12952 );
nor ( n12954 , n12945 , n12953 );
not ( n12955 , n1715 );
and ( n12956 , n12897 , n12903 , n12925 );
not ( n12957 , n12956 );
or ( n12958 , n12955 , n12957 );
nand ( n12959 , n1743 , n12931 );
nand ( n12960 , n12958 , n12959 );
not ( n12961 , n1692 );
not ( n12962 , n12914 );
or ( n12963 , n12961 , n12962 );
not ( n12964 , n12948 );
not ( n12965 , n12897 );
nand ( n12966 , n12964 , n12965 , n12885 );
not ( n12967 , n12966 );
nand ( n12968 , n1714 , n12967 );
nand ( n12969 , n12963 , n12968 );
nor ( n12970 , n12960 , n12969 );
nand ( n12971 , n12954 , n12970 );
and ( n12972 , n12939 , n12971 );
not ( n12973 , n12939 );
not ( n12974 , n12971 );
and ( n12975 , n12973 , n12974 );
nor ( n12976 , n12972 , n12975 );
not ( n12977 , n12976 );
buf ( n12978 , n12977 );
not ( n12979 , n1789 );
not ( n12980 , n12922 );
or ( n12981 , n12979 , n12980 );
nand ( n12982 , n1775 , n12905 );
nand ( n12983 , n12981 , n12982 );
nand ( n12984 , n1781 , n12936 );
nand ( n12985 , n1783 , n12911 );
nand ( n12986 , n12984 , n12985 );
nor ( n12987 , n12983 , n12986 );
nand ( n12988 , n1744 , n12931 );
nand ( n12989 , n1725 , n12956 );
nand ( n12990 , n1738 , n12967 );
and ( n12991 , n12885 , n12918 , n12925 );
nand ( n12992 , n1706 , n12991 );
nand ( n12993 , n12988 , n12989 , n12990 , n12992 );
not ( n12994 , n12993 );
nand ( n12995 , n12987 , n12994 );
not ( n12996 , n12995 );
not ( n12997 , n1735 );
not ( n12998 , n12956 );
or ( n12999 , n12997 , n12998 );
nand ( n13000 , n1717 , n12931 );
nand ( n13001 , n12999 , n13000 );
not ( n13002 , n1763 );
not ( n13003 , n12936 );
or ( n13004 , n13002 , n13003 );
nand ( n13005 , n1784 , n12911 );
nand ( n13006 , n13004 , n13005 );
nor ( n13007 , n13001 , n13006 );
not ( n13008 , n1791 );
not ( n13009 , n12922 );
or ( n13010 , n13008 , n13009 );
nand ( n13011 , n1771 , n12905 );
nand ( n13012 , n13010 , n13011 );
not ( n13013 , n1727 );
not ( n13014 , n12991 );
or ( n13015 , n13013 , n13014 );
nand ( n13016 , n1721 , n12967 );
nand ( n13017 , n13015 , n13016 );
nor ( n13018 , n13012 , n13017 );
nand ( n13019 , n13007 , n13018 );
not ( n13020 , n13019 );
not ( n13021 , n13020 );
or ( n13022 , n12996 , n13021 );
not ( n13023 , n12983 );
nand ( n13024 , n13023 , n12984 , n12985 );
nor ( n13025 , n13024 , n12993 );
nand ( n13026 , n13019 , n13025 );
nand ( n13027 , n13022 , n13026 );
not ( n13028 , n13027 );
nand ( n13029 , n12978 , n13028 );
not ( n13030 , n13029 );
nor ( n13031 , n12978 , n13028 );
nor ( n13032 , n13030 , n13031 );
not ( n13033 , n13032 );
and ( n13034 , n908 , n1007 );
not ( n13035 , n908 );
not ( n13036 , n1007 );
and ( n13037 , n13035 , n13036 );
or ( n13038 , n13034 , n13037 );
not ( n13039 , n183 );
and ( n13040 , n906 , n13039 );
not ( n13041 , n906 );
and ( n13042 , n13041 , n183 );
nor ( n13043 , n13040 , n13042 );
not ( n13044 , n13043 );
and ( n13045 , n13038 , n13044 );
not ( n13046 , n13038 );
and ( n13047 , n13046 , n13043 );
nor ( n13048 , n13045 , n13047 );
not ( n13049 , n13048 );
not ( n13050 , n154 );
and ( n13051 , n182 , n13050 );
not ( n13052 , n182 );
and ( n13053 , n13052 , n154 );
nor ( n13054 , n13051 , n13053 );
not ( n13055 , n13054 );
and ( n13056 , n907 , n876 );
not ( n13057 , n907 );
not ( n13058 , n876 );
and ( n13059 , n13057 , n13058 );
nor ( n13060 , n13056 , n13059 );
not ( n13061 , n13060 );
and ( n13062 , n13055 , n13061 );
and ( n13063 , n13054 , n13060 );
nor ( n13064 , n13062 , n13063 );
not ( n13065 , n13064 );
or ( n13066 , n13049 , n13065 );
or ( n13067 , n13048 , n13064 );
nand ( n13068 , n13066 , n13067 );
not ( n13069 , n13068 );
not ( n13070 , n1772 );
not ( n13071 , n12949 );
or ( n13072 , n13070 , n13071 );
not ( n13073 , n12904 );
nand ( n13074 , n13073 , n1764 );
nand ( n13075 , n13072 , n13074 );
not ( n13076 , n1728 );
not ( n13077 , n12991 );
or ( n13078 , n13076 , n13077 );
nand ( n13079 , n1703 , n12892 );
nand ( n13080 , n13078 , n13079 );
nor ( n13081 , n13075 , n13080 );
not ( n13082 , n1722 );
not ( n13083 , n12931 );
or ( n13084 , n13082 , n13083 );
nand ( n13085 , n1778 , n12941 );
nand ( n13086 , n13084 , n13085 );
not ( n13087 , n1724 );
not ( n13088 , n12926 );
or ( n13089 , n13087 , n13088 );
nand ( n13090 , n1788 , n12911 );
nand ( n13091 , n13089 , n13090 );
nor ( n13092 , n13086 , n13091 );
nand ( n13093 , n13081 , n13092 );
not ( n13094 , n1704 );
not ( n13095 , n12956 );
or ( n13096 , n13094 , n13095 );
nand ( n13097 , n1729 , n12931 );
nand ( n13098 , n13096 , n13097 );
not ( n13099 , n1792 );
not ( n13100 , n12941 );
or ( n13101 , n13099 , n13100 );
nand ( n13102 , n1765 , n12911 );
nand ( n13103 , n13101 , n13102 );
nor ( n13104 , n13098 , n13103 );
not ( n13105 , n1762 );
not ( n13106 , n12936 );
or ( n13107 , n13105 , n13106 );
nand ( n13108 , n1787 , n12905 );
nand ( n13109 , n13107 , n13108 );
not ( n13110 , n1730 );
not ( n13111 , n12991 );
or ( n13112 , n13110 , n13111 );
nand ( n13113 , n1702 , n12967 );
nand ( n13114 , n13112 , n13113 );
nor ( n13115 , n13109 , n13114 );
nand ( n13116 , n13104 , n13115 );
xor ( n13117 , n13093 , n13116 );
not ( n13118 , n13117 );
not ( n13119 , n13118 );
or ( n13120 , n13069 , n13119 );
not ( n13121 , n13117 );
or ( n13122 , n13121 , n13068 );
nand ( n13123 , n13120 , n13122 );
not ( n13124 , n13123 );
not ( n13125 , n13124 );
not ( n13126 , n1782 );
not ( n13127 , n12941 );
or ( n13128 , n13126 , n13127 );
nand ( n13129 , n13073 , n1780 );
nand ( n13130 , n13128 , n13129 );
not ( n13131 , n1790 );
not ( n13132 , n12949 );
or ( n13133 , n13131 , n13132 );
nand ( n13134 , n1786 , n12911 );
nand ( n13135 , n13133 , n13134 );
nor ( n13136 , n13130 , n13135 );
not ( n13137 , n1693 );
not ( n13138 , n12926 );
or ( n13139 , n13137 , n13138 );
not ( n13140 , n12891 );
nand ( n13141 , n1731 , n13140 );
nand ( n13142 , n13139 , n13141 );
not ( n13143 , n1726 );
not ( n13144 , n12931 );
or ( n13145 , n13143 , n13144 );
nand ( n13146 , n1732 , n12914 );
nand ( n13147 , n13145 , n13146 );
nor ( n13148 , n13142 , n13147 );
nand ( n13149 , n13136 , n13148 );
not ( n13150 , n13149 );
not ( n13151 , n13150 );
not ( n13152 , n1716 );
not ( n13153 , n12926 );
or ( n13154 , n13152 , n13153 );
nand ( n13155 , n1719 , n12931 );
nand ( n13156 , n13154 , n13155 );
not ( n13157 , n13156 );
not ( n13158 , n1768 );
not ( n13159 , n12949 );
or ( n13160 , n13158 , n13159 );
nand ( n13161 , n12911 , n1785 );
nand ( n13162 , n13160 , n13161 );
not ( n13163 , n13162 );
and ( n13164 , n1734 , n12991 );
and ( n13165 , n1779 , n13073 );
nor ( n13166 , n13164 , n13165 );
and ( n13167 , n1776 , n12922 );
not ( n13168 , n1705 );
nor ( n13169 , n13168 , n12891 );
nor ( n13170 , n13167 , n13169 );
nand ( n13171 , n13157 , n13163 , n13166 , n13170 );
not ( n13172 , n13171 );
not ( n13173 , n13172 );
or ( n13174 , n13151 , n13173 );
not ( n13175 , n13171 );
not ( n13176 , n13149 );
or ( n13177 , n13175 , n13176 );
nand ( n13178 , n13174 , n13177 );
not ( n13179 , n13178 );
not ( n13180 , n13179 );
not ( n13181 , n138 );
and ( n13182 , n13180 , n13181 );
and ( n13183 , n138 , n13179 );
nor ( n13184 , n13182 , n13183 );
not ( n13185 , n13184 );
not ( n13186 , n13185 );
or ( n13187 , n13125 , n13186 );
nand ( n13188 , n13184 , n13123 );
nand ( n13189 , n13187 , n13188 );
not ( n13190 , n13189 );
or ( n13191 , n13033 , n13190 );
or ( n13192 , n13032 , n13189 );
nand ( n13193 , n13191 , n13192 );
not ( n13194 , n12856 );
nand ( n13195 , n13193 , n13194 );
not ( n13196 , n12841 );
buf ( n13197 , n13196 );
buf ( n13198 , n13197 );
and ( n13199 , n12826 , n13198 );
not ( n13200 , n13199 );
nand ( n13201 , n12859 , n13195 , n13200 );
not ( n13202 , n891 );
not ( n13203 , n1587 );
not ( n13204 , n12508 );
or ( n13205 , n13203 , n13204 );
nor ( n13206 , n896 , n1599 );
not ( n13207 , n13206 );
not ( n13208 , n13207 );
nor ( n13209 , n1600 , n13208 );
not ( n13210 , n925 );
not ( n13211 , n900 );
not ( n13212 , n930 );
nand ( n13213 , n13211 , n13212 );
nand ( n13214 , n13209 , n13210 , n13213 );
nand ( n13215 , n13205 , n13214 );
not ( n13216 , n13215 );
not ( n13217 , n13216 );
not ( n13218 , n13217 );
not ( n13219 , n13218 );
or ( n13220 , n13202 , n13219 );
not ( n13221 , n13217 );
not ( n13222 , n13221 );
nand ( n13223 , n878 , n13222 );
nand ( n13224 , n13220 , n13223 );
or ( n13225 , n1129 , n13224 );
not ( n13226 , n1130 );
not ( n13227 , n897 );
or ( n13228 , n13227 , n13219 );
not ( n13229 , n13221 );
nand ( n13230 , n981 , n13229 );
nand ( n13231 , n13228 , n13230 );
not ( n13232 , n13231 );
nand ( n13233 , n13226 , n13232 );
and ( n13234 , n13225 , n13233 );
not ( n13235 , n1141 );
not ( n13236 , n955 );
not ( n13237 , n13218 );
or ( n13238 , n13236 , n13237 );
nand ( n13239 , n978 , n13217 );
nand ( n13240 , n13238 , n13239 );
not ( n13241 , n13240 );
nor ( n13242 , n13235 , n13241 );
not ( n13243 , n13242 );
not ( n13244 , n1142 );
not ( n13245 , n13218 );
and ( n13246 , n13245 , n979 );
not ( n13247 , n13245 );
and ( n13248 , n13247 , n956 );
nor ( n13249 , n13246 , n13248 );
nand ( n13250 , n13244 , n13249 );
not ( n13251 , n13250 );
or ( n13252 , n13243 , n13251 );
not ( n13253 , n13249 );
nand ( n13254 , n1142 , n13253 );
nand ( n13255 , n13252 , n13254 );
and ( n13256 , n13234 , n13255 );
nand ( n13257 , n1129 , n13224 );
not ( n13258 , n13233 );
nor ( n13259 , n13257 , n13258 );
nor ( n13260 , n13256 , n13259 );
nand ( n13261 , n1130 , n13231 );
nand ( n13262 , n13235 , n13241 );
and ( n13263 , n13262 , n13250 );
and ( n13264 , n13234 , n13263 );
not ( n13265 , n901 );
not ( n13266 , n1587 );
not ( n13267 , n13213 );
not ( n13268 , n13267 );
or ( n13269 , n13266 , n13268 );
not ( n13270 , n925 );
not ( n13271 , n1600 );
nand ( n13272 , n13270 , n13213 , n13271 , n13207 );
nand ( n13273 , n13269 , n13272 );
buf ( n13274 , n13273 );
or ( n13275 , n13265 , n13274 );
nand ( n13276 , n877 , n13274 );
nand ( n13277 , n13275 , n13276 );
not ( n13278 , n13277 );
not ( n13279 , n13278 );
nor ( n13280 , n1139 , n13279 );
not ( n13281 , n13280 );
not ( n13282 , n1140 );
buf ( n13283 , n13215 );
or ( n13284 , n954 , n13283 );
not ( n13285 , n977 );
nand ( n13286 , n13285 , n13283 );
nand ( n13287 , n13284 , n13286 );
not ( n13288 , n13287 );
not ( n13289 , n13288 );
not ( n13290 , n13289 );
not ( n13291 , n13290 );
nand ( n13292 , n13282 , n13291 );
and ( n13293 , n13281 , n13292 );
not ( n13294 , n13293 );
not ( n13295 , n1138 );
not ( n13296 , n953 );
or ( n13297 , n13296 , n13283 );
nand ( n13298 , n976 , n13283 );
nand ( n13299 , n13297 , n13298 );
not ( n13300 , n13299 );
buf ( n13301 , n13300 );
nand ( n13302 , n13295 , n13301 );
not ( n13303 , n1137 );
or ( n13304 , n952 , n13283 );
not ( n13305 , n13273 );
not ( n13306 , n13305 );
not ( n13307 , n975 );
nand ( n13308 , n13306 , n13307 );
nand ( n13309 , n13304 , n13308 );
nand ( n13310 , n13303 , n13309 );
and ( n13311 , n13302 , n13310 );
not ( n13312 , n880 );
not ( n13313 , n13274 );
or ( n13314 , n13312 , n13313 );
not ( n13315 , n13273 );
nand ( n13316 , n899 , n13315 );
nand ( n13317 , n13314 , n13316 );
nand ( n13318 , n1135 , n13317 );
or ( n13319 , n974 , n13216 );
not ( n13320 , n951 );
nand ( n13321 , n13320 , n13305 );
nand ( n13322 , n13319 , n13321 );
buf ( n13323 , n13322 );
not ( n13324 , n13323 );
nor ( n13325 , n1136 , n13324 );
or ( n13326 , n13318 , n13325 );
not ( n13327 , n13323 );
nand ( n13328 , n1136 , n13327 );
nand ( n13329 , n13326 , n13328 );
not ( n13330 , n13329 );
not ( n13331 , n1134 );
not ( n13332 , n973 );
not ( n13333 , n13283 );
or ( n13334 , n13332 , n13333 );
nand ( n13335 , n950 , n13305 );
nand ( n13336 , n13334 , n13335 );
buf ( n13337 , n13336 );
not ( n13338 , n13337 );
nor ( n13339 , n13331 , n13338 );
not ( n13340 , n13339 );
not ( n13341 , n13340 );
not ( n13342 , n971 );
not ( n13343 , n13274 );
or ( n13344 , n13342 , n13343 );
nand ( n13345 , n948 , n13305 );
nand ( n13346 , n13344 , n13345 );
not ( n13347 , n13346 );
not ( n13348 , n13347 );
nand ( n13349 , n1128 , n13348 );
not ( n13350 , n13349 );
not ( n13351 , n1128 );
nand ( n13352 , n13351 , n13347 );
not ( n13353 , n1127 );
not ( n13354 , n1000 );
not ( n13355 , n13315 );
or ( n13356 , n13354 , n13355 );
nand ( n13357 , n883 , n13274 );
nand ( n13358 , n13356 , n13357 );
not ( n13359 , n13358 );
nand ( n13360 , n13353 , n13359 );
not ( n13361 , n13360 );
not ( n13362 , n1126 );
and ( n13363 , n13216 , n947 );
not ( n13364 , n13216 );
and ( n13365 , n13364 , n970 );
nor ( n13366 , n13363 , n13365 );
nor ( n13367 , n13362 , n13366 );
not ( n13368 , n13367 );
or ( n13369 , n13361 , n13368 );
nand ( n13370 , n1127 , n13358 );
nand ( n13371 , n13369 , n13370 );
nand ( n13372 , n13352 , n13371 );
not ( n13373 , n13372 );
or ( n13374 , n13350 , n13373 );
not ( n13375 , n1134 );
not ( n13376 , n13337 );
nand ( n13377 , n13375 , n13376 );
nand ( n13378 , n13374 , n13377 );
not ( n13379 , n13378 );
or ( n13380 , n13341 , n13379 );
or ( n13381 , n1135 , n13317 );
not ( n13382 , n13381 );
nor ( n13383 , n13382 , n13325 );
nand ( n13384 , n13380 , n13383 );
nand ( n13385 , n13330 , n13384 );
and ( n13386 , n13311 , n13385 );
not ( n13387 , n13301 );
nand ( n13388 , n1138 , n13387 );
not ( n13389 , n13309 );
nand ( n13390 , n1137 , n13389 );
not ( n13391 , n13390 );
nand ( n13392 , n13391 , n13302 );
nand ( n13393 , n13388 , n13392 );
nor ( n13394 , n13386 , n13393 );
or ( n13395 , n13294 , n13394 );
not ( n13396 , n13278 );
not ( n13397 , n13396 );
not ( n13398 , n13397 );
and ( n13399 , n1139 , n13398 );
and ( n13400 , n13399 , n13292 );
nor ( n13401 , n13282 , n13289 );
nor ( n13402 , n13400 , n13401 );
nand ( n13403 , n13395 , n13402 );
nand ( n13404 , n13264 , n13403 );
nand ( n13405 , n13260 , n13261 , n13404 );
and ( n13406 , n13405 , n1131 );
not ( n13407 , n13405 );
not ( n13408 , n1131 );
and ( n13409 , n13407 , n13408 );
nor ( n13410 , n13406 , n13409 );
not ( n13411 , n995 );
nand ( n13412 , n994 , n12603 );
not ( n13413 , n13412 );
not ( n13414 , n12796 );
and ( n13415 , n13413 , n13414 );
and ( n13416 , n994 , n12611 );
nor ( n13417 , n13415 , n13416 );
nor ( n13418 , n13412 , n12768 );
not ( n13419 , n12773 );
not ( n13420 , n12785 );
not ( n13421 , n13420 );
or ( n13422 , n13419 , n13421 );
nand ( n13423 , n13422 , n12792 );
nand ( n13424 , n13418 , n13423 );
not ( n13425 , n12775 );
nor ( n13426 , n12772 , n13425 );
not ( n13427 , n12780 );
not ( n13428 , n12803 );
not ( n13429 , n13428 );
not ( n13430 , n12814 );
or ( n13431 , n13429 , n13430 );
nand ( n13432 , n13431 , n12799 );
nand ( n13433 , n13427 , n13432 );
nand ( n13434 , n13418 , n13426 , n13433 );
nand ( n13435 , n13417 , n13424 , n13434 );
not ( n13436 , n13435 );
nor ( n13437 , n13411 , n13436 );
or ( n13438 , n995 , n13435 );
nand ( n13439 , n13438 , n12726 );
or ( n13440 , n13437 , n13439 );
not ( n13441 , n945 );
or ( n13442 , n13441 , n12726 );
nand ( n13443 , n13440 , n13442 );
not ( n13444 , n12600 );
nor ( n13445 , n13444 , n12608 );
not ( n13446 , n12744 );
not ( n13447 , n13446 );
not ( n13448 , n12752 );
or ( n13449 , n13447 , n13448 );
not ( n13450 , n12739 );
nand ( n13451 , n13449 , n13450 );
nor ( n13452 , n13445 , n13451 );
not ( n13453 , n13445 );
not ( n13454 , n13451 );
or ( n13455 , n13453 , n13454 );
nand ( n13456 , n13455 , n12726 );
or ( n13457 , n13452 , n13456 );
not ( n13458 , n943 );
or ( n13459 , n13458 , n12726 );
nand ( n13460 , n13457 , n13459 );
not ( n13461 , n142 );
nor ( n13462 , n13461 , n12855 );
not ( n13463 , n13462 );
and ( n13464 , n12939 , n12971 );
not ( n13465 , n12939 );
and ( n13466 , n13465 , n12974 );
nor ( n13467 , n13464 , n13466 );
and ( n13468 , n13178 , n13467 );
not ( n13469 , n13178 );
and ( n13470 , n13469 , n12977 );
or ( n13471 , n13468 , n13470 );
and ( n13472 , n183 , n13050 );
not ( n13473 , n183 );
and ( n13474 , n13473 , n154 );
nor ( n13475 , n13472 , n13474 );
not ( n13476 , n906 );
and ( n13477 , n1007 , n13476 );
not ( n13478 , n1007 );
and ( n13479 , n13478 , n906 );
nor ( n13480 , n13477 , n13479 );
not ( n13481 , n13480 );
or ( n13482 , n13475 , n13481 );
not ( n13483 , n13475 );
or ( n13484 , n13480 , n13483 );
nand ( n13485 , n13482 , n13484 );
not ( n13486 , n13485 );
and ( n13487 , n876 , n12825 );
not ( n13488 , n876 );
and ( n13489 , n13488 , n138 );
nor ( n13490 , n13487 , n13489 );
xnor ( n13491 , n908 , n907 );
not ( n13492 , n13491 );
and ( n13493 , n13490 , n13492 );
not ( n13494 , n13490 );
and ( n13495 , n13494 , n13491 );
nor ( n13496 , n13493 , n13495 );
not ( n13497 , n13496 );
or ( n13498 , n13486 , n13497 );
or ( n13499 , n13496 , n13485 );
nand ( n13500 , n13498 , n13499 );
not ( n13501 , n13500 );
not ( n13502 , n13117 );
not ( n13503 , n13502 );
or ( n13504 , n13501 , n13503 );
not ( n13505 , n13500 );
nand ( n13506 , n13505 , n13117 );
nand ( n13507 , n13504 , n13506 );
not ( n13508 , n13028 );
and ( n13509 , n13507 , n13508 );
not ( n13510 , n13507 );
and ( n13511 , n13510 , n13028 );
nor ( n13512 , n13509 , n13511 );
xnor ( n13513 , n13471 , n13512 );
nand ( n13514 , n13194 , n13513 );
nand ( n13515 , n13463 , n13200 , n13514 );
buf ( n13516 , n12498 );
not ( n13517 , n13516 );
not ( n13518 , n1357 );
nand ( n13519 , n1356 , n13518 );
not ( n13520 , n13519 );
not ( n13521 , n1365 );
nor ( n13522 , n13521 , n1358 );
nand ( n13523 , n13520 , n13522 );
not ( n13524 , n13523 );
not ( n13525 , n13524 );
or ( n13526 , n13517 , n13525 );
nand ( n13527 , n13526 , n12512 );
not ( n13528 , n13527 );
nor ( n13529 , n217 , n238 );
nor ( n13530 , n218 , n237 );
not ( n13531 , n239 );
not ( n13532 , n224 );
nor ( n13533 , n240 , n241 );
nand ( n13534 , n13531 , n13532 , n13533 );
nor ( n13535 , n221 , n13534 );
and ( n13536 , n13529 , n13530 , n13535 );
not ( n13537 , n909 );
nor ( n13538 , n13537 , n927 );
not ( n13539 , n1608 );
not ( n13540 , n1365 );
nand ( n13541 , n13540 , n1358 );
not ( n13542 , n13541 );
nor ( n13543 , n1356 , n1357 );
nand ( n13544 , n13542 , n13543 );
nor ( n13545 , n13539 , n13544 );
nor ( n13546 , n13538 , n13545 );
not ( n13547 , n927 );
nor ( n13548 , n13547 , n909 );
not ( n13549 , n13541 );
nand ( n13550 , n13520 , n13549 );
nand ( n13551 , n481 , n13550 );
or ( n13552 , n13548 , n13551 );
not ( n13553 , n1599 );
not ( n13554 , n1600 );
or ( n13555 , n13553 , n13554 );
not ( n13556 , n13516 );
not ( n13557 , n13556 );
not ( n13558 , n1599 );
nor ( n13559 , n1358 , n1365 );
nand ( n13560 , n13520 , n13559 );
not ( n13561 , n13560 );
not ( n13562 , n13561 );
or ( n13563 , n13558 , n13562 );
not ( n13564 , n13523 );
nand ( n13565 , n13564 , n1600 );
nand ( n13566 , n13563 , n13565 );
and ( n13567 , n13557 , n13566 );
or ( n13568 , n254 , n12493 );
or ( n13569 , n514 , n12512 );
nand ( n13570 , n13568 , n13569 );
not ( n13571 , n13570 );
not ( n13572 , n12503 );
nor ( n13573 , n13571 , n13572 );
nor ( n13574 , n13567 , n13573 );
nand ( n13575 , n13555 , n13574 );
nor ( n13576 , n13552 , n13575 );
nand ( n13577 , n13536 , n13546 , n13576 );
nor ( n13578 , n13528 , n13577 );
or ( n13579 , n250 , n13578 );
nand ( n13580 , n1220 , n1230 );
nor ( n13581 , n198 , n203 );
not ( n13582 , n13581 );
nor ( n13583 , n13582 , n204 , n199 );
nor ( n13584 , n209 , n210 );
nor ( n13585 , n211 , n212 );
nand ( n13586 , n13584 , n13585 );
nor ( n13587 , n202 , n205 );
not ( n13588 , n207 );
not ( n13589 , n206 );
nor ( n13590 , n200 , n208 );
and ( n13591 , n13588 , n13589 , n13590 );
nand ( n13592 , n13587 , n13591 );
nor ( n13593 , n13586 , n13592 );
nand ( n13594 , n13583 , n13593 );
nand ( n13595 , n12829 , n13594 );
nand ( n13596 , n13580 , n13595 );
not ( n13597 , n13596 );
and ( n13598 , n212 , n13597 );
not ( n13599 , n211 );
not ( n13600 , n200 );
nand ( n13601 , n13589 , n13587 );
nor ( n13602 , n207 , n13601 );
nand ( n13603 , n13600 , n13602 );
nor ( n13604 , n208 , n13603 );
and ( n13605 , n13599 , n13584 , n13604 );
and ( n13606 , n212 , n13605 );
nor ( n13607 , n212 , n13605 );
nor ( n13608 , n13606 , n13607 , n13597 );
nor ( n13609 , n13598 , n13608 );
nor ( n13610 , n13579 , n13609 );
not ( n13611 , n13610 );
not ( n13612 , n13290 );
nor ( n13613 , n13224 , n13231 );
not ( n13614 , n13287 );
nand ( n13615 , n13614 , n13279 );
or ( n13616 , n939 , n13615 );
not ( n13617 , n13288 );
or ( n13618 , n888 , n13617 );
nand ( n13619 , n13616 , n13618 );
nor ( n13620 , n888 , n939 );
and ( n13621 , n13620 , n13396 );
not ( n13622 , n13621 );
not ( n13623 , n937 );
not ( n13624 , n13299 );
and ( n13625 , n938 , n13624 );
nor ( n13626 , n13625 , n13309 );
and ( n13627 , n888 , n13287 );
not ( n13628 , n939 );
nor ( n13629 , n13628 , n13277 );
nor ( n13630 , n13627 , n13629 );
nand ( n13631 , n13623 , n13626 , n13630 );
not ( n13632 , n13300 );
not ( n13633 , n938 );
nand ( n13634 , n13632 , n13633 , n13630 );
nand ( n13635 , n13622 , n13631 , n13634 );
or ( n13636 , n13619 , n13635 );
or ( n13637 , n12538 , n13240 );
nand ( n13638 , n13636 , n13637 );
nand ( n13639 , n13613 , n13638 );
not ( n13640 , n13639 );
nor ( n13641 , n879 , n988 );
not ( n13642 , n13641 );
nand ( n13643 , n879 , n988 );
not ( n13644 , n13643 );
not ( n13645 , n13644 );
and ( n13646 , n13283 , n970 );
not ( n13647 , n13283 );
and ( n13648 , n13647 , n947 );
nor ( n13649 , n13646 , n13648 );
not ( n13650 , n13649 );
or ( n13651 , n13645 , n13650 );
or ( n13652 , n879 , n13366 );
nand ( n13653 , n13652 , n13359 );
nand ( n13654 , n13651 , n13653 );
nand ( n13655 , n13642 , n13654 );
and ( n13656 , n884 , n13323 );
not ( n13657 , n13317 );
and ( n13658 , n13657 , n936 );
nor ( n13659 , n13656 , n13658 );
not ( n13660 , n935 );
not ( n13661 , n13660 );
not ( n13662 , n13346 );
or ( n13663 , n13661 , n13662 );
not ( n13664 , n933 );
nand ( n13665 , n13664 , n13336 );
nand ( n13666 , n13663 , n13665 );
not ( n13667 , n13666 );
nand ( n13668 , n13664 , n13660 );
nand ( n13669 , n13346 , n13336 );
nand ( n13670 , n13667 , n13668 , n13669 );
nand ( n13671 , n13655 , n13659 , n13670 );
and ( n13672 , n13660 , n13337 , n13659 );
nor ( n13673 , n884 , n13323 );
nor ( n13674 , n13672 , n13673 );
not ( n13675 , n936 );
nor ( n13676 , n13657 , n13323 );
nand ( n13677 , n13675 , n13676 );
not ( n13678 , n13347 );
not ( n13679 , n13336 );
and ( n13680 , n935 , n13679 );
nor ( n13681 , n13680 , n933 );
and ( n13682 , n13678 , n13681 , n13659 );
or ( n13683 , n884 , n936 );
nor ( n13684 , n13683 , n13657 );
nor ( n13685 , n13682 , n13684 );
nand ( n13686 , n13671 , n13674 , n13677 , n13685 );
or ( n13687 , n937 , n13624 );
not ( n13688 , n13626 );
nor ( n13689 , n937 , n938 );
not ( n13690 , n13689 );
nand ( n13691 , n13687 , n13688 , n13690 );
and ( n13692 , n13637 , n13630 );
nand ( n13693 , n13686 , n13691 , n13692 );
not ( n13694 , n1006 );
not ( n13695 , n13249 );
or ( n13696 , n13694 , n13695 );
nand ( n13697 , n13241 , n13249 );
nand ( n13698 , n13696 , n13697 );
nand ( n13699 , n13640 , n13693 , n13698 );
buf ( n13700 , n13699 );
or ( n13701 , n13612 , n13700 );
nand ( n13702 , n888 , n13700 );
nand ( n13703 , n13701 , n13702 );
nand ( n13704 , n13579 , n13703 );
nand ( n13705 , n13611 , n2 , n13704 );
not ( n13706 , n13250 );
and ( n13707 , n13262 , n13401 );
nor ( n13708 , n13707 , n13242 );
or ( n13709 , n13706 , n13708 );
nand ( n13710 , n13709 , n13254 );
nand ( n13711 , n13225 , n13710 );
and ( n13712 , n13262 , n13292 );
and ( n13713 , n13250 , n13712 );
not ( n13714 , n13302 );
or ( n13715 , n13280 , n13714 );
not ( n13716 , n13325 );
and ( n13717 , n13716 , n13310 );
not ( n13718 , n13339 );
not ( n13719 , n13381 );
or ( n13720 , n13718 , n13719 );
nand ( n13721 , n13720 , n13318 );
not ( n13722 , n13721 );
and ( n13723 , n13381 , n13377 );
nand ( n13724 , n13349 , n13372 );
nand ( n13725 , n13723 , n13724 );
nand ( n13726 , n13722 , n13725 );
and ( n13727 , n13717 , n13726 );
not ( n13728 , n13328 );
nand ( n13729 , n13310 , n13728 );
nand ( n13730 , n13390 , n13729 );
nor ( n13731 , n13727 , n13730 );
or ( n13732 , n13715 , n13731 );
not ( n13733 , n13388 );
not ( n13734 , n13280 );
and ( n13735 , n13733 , n13734 );
nor ( n13736 , n13735 , n13399 );
nand ( n13737 , n13732 , n13736 );
nand ( n13738 , n13713 , n13225 , n13737 );
nand ( n13739 , n13711 , n13257 , n13738 );
nand ( n13740 , n13261 , n13233 );
not ( n13741 , n13740 );
and ( n13742 , n13739 , n13741 );
not ( n13743 , n13739 );
and ( n13744 , n13743 , n13740 );
nor ( n13745 , n13742 , n13744 );
not ( n13746 , n12526 );
not ( n13747 , n13746 );
not ( n13748 , n13747 );
buf ( n13749 , n12534 );
buf ( n13750 , n13749 );
buf ( n13751 , n13750 );
not ( n13752 , n13751 );
not ( n13753 , n988 );
not ( n13754 , n13700 );
or ( n13755 , n13753 , n13754 );
not ( n13756 , n13649 );
not ( n13757 , n13756 );
not ( n13758 , n13757 );
not ( n13759 , n13639 );
and ( n13760 , n13759 , n13698 , n13693 );
nand ( n13761 , n13758 , n13760 );
nand ( n13762 , n13755 , n13761 );
and ( n13763 , n13752 , n13762 );
not ( n13764 , n12686 );
nor ( n13765 , n13763 , n13764 );
or ( n13766 , n13748 , n13765 );
nand ( n13767 , n13766 , n12690 );
not ( n13768 , n13751 );
not ( n13769 , n879 );
not ( n13770 , n13700 );
or ( n13771 , n13769 , n13770 );
or ( n13772 , n13359 , n13700 );
nand ( n13773 , n13771 , n13772 );
and ( n13774 , n13768 , n13773 );
not ( n13775 , n12674 );
nor ( n13776 , n13774 , n13775 );
or ( n13777 , n13748 , n13776 );
nand ( n13778 , n13777 , n12678 );
not ( n13779 , n935 );
not ( n13780 , n13700 );
or ( n13781 , n13779 , n13780 );
buf ( n13782 , n13376 );
not ( n13783 , n13782 );
buf ( n13784 , n13783 );
not ( n13785 , n13784 );
buf ( n13786 , n13785 );
or ( n13787 , n13786 , n13700 );
nand ( n13788 , n13781 , n13787 );
and ( n13789 , n13768 , n13788 );
not ( n13790 , n12707 );
nor ( n13791 , n13789 , n13790 );
or ( n13792 , n13748 , n13791 );
nand ( n13793 , n13792 , n12711 );
not ( n13794 , n884 );
not ( n13795 , n13700 );
or ( n13796 , n13794 , n13795 );
not ( n13797 , n13327 );
or ( n13798 , n13797 , n13700 );
nand ( n13799 , n13796 , n13798 );
and ( n13800 , n13752 , n13799 );
nor ( n13801 , n13800 , n12642 );
or ( n13802 , n13748 , n13801 );
nand ( n13803 , n13802 , n12645 );
not ( n13804 , n936 );
not ( n13805 , n13700 );
or ( n13806 , n13804 , n13805 );
or ( n13807 , n13657 , n13700 );
nand ( n13808 , n13806 , n13807 );
and ( n13809 , n13752 , n13808 );
not ( n13810 , n12630 );
nor ( n13811 , n13809 , n13810 );
or ( n13812 , n13748 , n13811 );
nand ( n13813 , n13812 , n12625 );
not ( n13814 , n13747 );
not ( n13815 , n1006 );
not ( n13816 , n13700 );
or ( n13817 , n13815 , n13816 );
or ( n13818 , n13241 , n13700 );
nand ( n13819 , n13817 , n13818 );
and ( n13820 , n13752 , n13819 );
not ( n13821 , n12535 );
nor ( n13822 , n13820 , n13821 );
or ( n13823 , n13814 , n13822 );
not ( n13824 , n12540 );
nand ( n13825 , n13823 , n13824 );
and ( n13826 , n13579 , n13762 );
not ( n13827 , n13579 );
not ( n13828 , n202 );
and ( n13829 , n13828 , n13597 );
and ( n13830 , n202 , n13596 );
nor ( n13831 , n13829 , n13830 );
and ( n13832 , n13827 , n13831 );
nor ( n13833 , n13826 , n13832 );
nand ( n13834 , n2 , n13833 );
not ( n13835 , n139 );
nor ( n13836 , n13835 , n12855 );
not ( n13837 , n13836 );
xor ( n13838 , n13496 , n13471 );
or ( n13839 , n13039 , n13481 );
or ( n13840 , n183 , n13480 );
nand ( n13841 , n13839 , n13840 );
nand ( n13842 , n13092 , n13081 );
xor ( n13843 , n13841 , n13842 );
not ( n13844 , n13843 );
not ( n13845 , n13027 );
or ( n13846 , n13844 , n13845 );
or ( n13847 , n13843 , n13027 );
nand ( n13848 , n13846 , n13847 );
xnor ( n13849 , n13838 , n13848 );
nand ( n13850 , n13849 , n13194 );
nand ( n13851 , n13837 , n13850 , n13200 );
and ( n13852 , n13828 , n13596 );
not ( n13853 , n205 );
nor ( n13854 , n13852 , n13853 );
or ( n13855 , n13587 , n13854 );
or ( n13856 , n205 , n13596 );
not ( n13857 , n13579 );
nand ( n13858 , n13855 , n13856 , n13857 );
nand ( n13859 , n13579 , n13773 );
nand ( n13860 , n13858 , n2 , n13859 );
not ( n13861 , n937 );
not ( n13862 , n13700 );
or ( n13863 , n13861 , n13862 );
not ( n13864 , n13309 );
not ( n13865 , n13864 );
or ( n13866 , n13865 , n13700 );
nand ( n13867 , n13863 , n13866 );
or ( n13868 , n13857 , n13867 );
and ( n13869 , n209 , n13597 );
not ( n13870 , n13592 );
or ( n13871 , n209 , n13870 );
and ( n13872 , n209 , n13870 );
nor ( n13873 , n13872 , n13597 );
nand ( n13874 , n13871 , n13873 );
nand ( n13875 , n13874 , n13857 );
or ( n13876 , n13869 , n13875 );
nand ( n13877 , n13868 , n13876 );
nand ( n13878 , n2 , n13877 );
not ( n13879 , n13747 );
buf ( n13880 , n13750 );
not ( n13881 , n13347 );
not ( n13882 , n13881 );
not ( n13883 , n13882 );
not ( n13884 , n13760 );
or ( n13885 , n13883 , n13884 );
or ( n13886 , n933 , n13760 );
nand ( n13887 , n13885 , n13886 );
or ( n13888 , n13880 , n13887 );
nand ( n13889 , n13888 , n12660 );
not ( n13890 , n13889 );
or ( n13891 , n13879 , n13890 );
nand ( n13892 , n13891 , n12664 );
not ( n13893 , n938 );
not ( n13894 , n13700 );
or ( n13895 , n13893 , n13894 );
not ( n13896 , n13387 );
or ( n13897 , n13896 , n13700 );
nand ( n13898 , n13895 , n13897 );
or ( n13899 , n13857 , n13898 );
and ( n13900 , n210 , n13597 );
not ( n13901 , n209 );
and ( n13902 , n13901 , n13590 , n13602 );
or ( n13903 , n210 , n13902 );
and ( n13904 , n210 , n13902 );
nor ( n13905 , n13904 , n13597 );
nand ( n13906 , n13903 , n13905 );
nand ( n13907 , n13906 , n13857 );
or ( n13908 , n13900 , n13907 );
nand ( n13909 , n13899 , n13908 );
nand ( n13910 , n2 , n13909 );
nor ( n13911 , n12543 , n12770 );
not ( n13912 , n12595 );
nand ( n13913 , n13912 , n12719 );
nor ( n13914 , n13911 , n13913 );
not ( n13915 , n13911 );
not ( n13916 , n13913 );
or ( n13917 , n13915 , n13916 );
nand ( n13918 , n13917 , n12726 );
or ( n13919 , n13914 , n13918 );
not ( n13920 , n941 );
or ( n13921 , n13920 , n12726 );
nand ( n13922 , n13919 , n13921 );
not ( n13923 , n12523 );
nor ( n13924 , n13923 , n12547 );
not ( n13925 , n13423 );
nand ( n13926 , n13426 , n13433 );
nand ( n13927 , n13925 , n13926 );
nor ( n13928 , n13924 , n13927 );
not ( n13929 , n13924 );
not ( n13930 , n13927 );
or ( n13931 , n13929 , n13930 );
nand ( n13932 , n13931 , n12726 );
or ( n13933 , n13928 , n13932 );
not ( n13934 , n942 );
or ( n13935 , n13934 , n12726 );
nand ( n13936 , n13933 , n13935 );
not ( n13937 , n12519 );
not ( n13938 , n13937 );
not ( n13939 , n13938 );
not ( n13940 , n13703 );
or ( n13941 , n13939 , n13940 );
and ( n13942 , n12555 , n12560 );
nand ( n13943 , n13941 , n13942 );
not ( n13944 , n13579 );
not ( n13945 , n939 );
not ( n13946 , n13700 );
or ( n13947 , n13945 , n13946 );
not ( n13948 , n13398 );
or ( n13949 , n13948 , n13700 );
nand ( n13950 , n13947 , n13949 );
not ( n13951 , n13950 );
or ( n13952 , n13944 , n13951 );
nand ( n13953 , n13590 , n13584 , n13602 );
and ( n13954 , n13953 , n211 );
not ( n13955 , n13953 );
and ( n13956 , n13955 , n13599 );
nor ( n13957 , n13954 , n13956 );
or ( n13958 , n13957 , n13597 );
or ( n13959 , n13599 , n13596 );
nand ( n13960 , n13958 , n13959 );
and ( n13961 , n13857 , n13960 );
not ( n13962 , n2 );
nor ( n13963 , n13961 , n13962 );
nand ( n13964 , n13952 , n13963 );
not ( n13965 , n12594 );
nor ( n13966 , n13965 , n12562 );
not ( n13967 , n12786 );
not ( n13968 , n12817 );
nand ( n13969 , n13967 , n13968 );
nor ( n13970 , n13966 , n13969 );
not ( n13971 , n13966 );
not ( n13972 , n13969 );
or ( n13973 , n13971 , n13972 );
nand ( n13974 , n13973 , n12726 );
or ( n13975 , n13970 , n13974 );
not ( n13976 , n963 );
or ( n13977 , n13976 , n12726 );
nand ( n13978 , n13975 , n13977 );
or ( n13979 , n13050 , n12855 );
and ( n13980 , n142 , n13058 );
not ( n13981 , n142 );
and ( n13982 , n13981 , n876 );
nor ( n13983 , n13980 , n13982 );
not ( n13984 , n13983 );
not ( n13985 , n13984 );
buf ( n13986 , n13184 );
not ( n13987 , n13986 );
or ( n13988 , n13985 , n13987 );
not ( n13989 , n13986 );
and ( n13990 , n13983 , n13989 );
nor ( n13991 , n13990 , n12854 );
nand ( n13992 , n13988 , n13991 );
nand ( n13993 , n13979 , n13200 , n13992 );
and ( n13994 , n12589 , n12568 );
nor ( n13995 , n13994 , n12752 );
not ( n13996 , n13994 );
not ( n13997 , n12752 );
or ( n13998 , n13996 , n13997 );
nand ( n13999 , n13998 , n12726 );
or ( n14000 , n13995 , n13999 );
not ( n14001 , n962 );
or ( n14002 , n14001 , n12726 );
nand ( n14003 , n14000 , n14002 );
not ( n14004 , n13579 );
not ( n14005 , n13819 );
or ( n14006 , n14004 , n14005 );
not ( n14007 , n198 );
not ( n14008 , n13597 );
or ( n14009 , n14007 , n14008 );
xnor ( n14010 , n13593 , n198 );
or ( n14011 , n13597 , n14010 );
nand ( n14012 , n14009 , n14011 );
and ( n14013 , n13857 , n14012 );
not ( n14014 , n2 );
nor ( n14015 , n14013 , n14014 );
nand ( n14016 , n14006 , n14015 );
not ( n14017 , n13579 );
not ( n14018 , n13808 );
or ( n14019 , n14017 , n14018 );
not ( n14020 , n200 );
nand ( n14021 , n14020 , n13597 );
not ( n14022 , n13602 );
or ( n14023 , n14022 , n13597 );
nand ( n14024 , n14023 , n200 );
nand ( n14025 , n13603 , n14024 );
and ( n14026 , n14021 , n14025 , n13857 );
not ( n14027 , n2 );
nor ( n14028 , n14026 , n14027 );
nand ( n14029 , n14019 , n14028 );
not ( n14030 , n13579 );
nand ( n14031 , n13253 , n13760 );
not ( n14032 , n14031 );
or ( n14033 , n14030 , n14032 );
nand ( n14034 , n203 , n13597 );
not ( n14035 , n13902 );
or ( n14036 , n198 , n212 );
nor ( n14037 , n14035 , n210 , n211 , n14036 );
or ( n14038 , n203 , n14037 );
and ( n14039 , n203 , n14037 );
nor ( n14040 , n14039 , n13597 );
nand ( n14041 , n14038 , n14040 );
nand ( n14042 , n14034 , n14041 , n13857 );
nand ( n14043 , n14033 , n14042 );
nand ( n14044 , n2 , n14043 );
not ( n14045 , n13579 );
nand ( n14046 , n13231 , n13760 );
not ( n14047 , n14046 );
or ( n14048 , n14045 , n14047 );
nand ( n14049 , n204 , n13597 );
not ( n14050 , n13605 );
nor ( n14051 , n14050 , n199 , n203 , n14036 );
or ( n14052 , n204 , n14051 );
and ( n14053 , n204 , n14051 );
nor ( n14054 , n14053 , n13597 );
nand ( n14055 , n14052 , n14054 );
nand ( n14056 , n14049 , n14055 , n13857 );
nand ( n14057 , n14048 , n14056 );
nand ( n14058 , n2 , n14057 );
not ( n14059 , n13579 );
not ( n14060 , n13788 );
or ( n14061 , n14059 , n14060 );
not ( n14062 , n207 );
not ( n14063 , n13596 );
and ( n14064 , n14062 , n14063 );
or ( n14065 , n13601 , n13597 );
nand ( n14066 , n14065 , n207 );
and ( n14067 , n14022 , n14066 );
nor ( n14068 , n14064 , n14067 );
and ( n14069 , n14068 , n13857 );
not ( n14070 , n2 );
nor ( n14071 , n14069 , n14070 );
nand ( n14072 , n14061 , n14071 );
not ( n14073 , n13579 );
not ( n14074 , n13799 );
or ( n14075 , n14073 , n14074 );
not ( n14076 , n208 );
not ( n14077 , n13596 );
and ( n14078 , n14076 , n14077 );
not ( n14079 , n13604 );
or ( n14080 , n13603 , n13597 );
nand ( n14081 , n14080 , n208 );
and ( n14082 , n14079 , n14081 );
nor ( n14083 , n14078 , n14082 );
and ( n14084 , n14083 , n13857 );
not ( n14085 , n2 );
nor ( n14086 , n14084 , n14085 );
nand ( n14087 , n14075 , n14086 );
not ( n14088 , n13938 );
not ( n14089 , n13950 );
or ( n14090 , n14088 , n14089 );
and ( n14091 , n12565 , n12566 );
nand ( n14092 , n14090 , n14091 );
not ( n14093 , n13242 );
nand ( n14094 , n14093 , n13262 );
not ( n14095 , n13403 );
and ( n14096 , n14094 , n14095 );
not ( n14097 , n14094 );
and ( n14098 , n14097 , n13403 );
nor ( n14099 , n14096 , n14098 );
not ( n14100 , n13938 );
not ( n14101 , n13867 );
or ( n14102 , n14100 , n14101 );
and ( n14103 , n12571 , n12572 );
nand ( n14104 , n14102 , n14103 );
not ( n14105 , n13938 );
not ( n14106 , n13898 );
or ( n14107 , n14105 , n14106 );
and ( n14108 , n12578 , n12580 );
nand ( n14109 , n14107 , n14108 );
and ( n14110 , n13717 , n13721 );
nor ( n14111 , n14110 , n13730 );
or ( n14112 , n13715 , n14111 );
nand ( n14113 , n14112 , n13736 );
nand ( n14114 , n13712 , n14113 );
not ( n14115 , n13715 );
not ( n14116 , n13725 );
nand ( n14117 , n13717 , n14116 );
not ( n14118 , n14117 );
nand ( n14119 , n13712 , n14115 , n14118 );
nand ( n14120 , n14114 , n13708 , n14119 );
nand ( n14121 , n13254 , n13250 );
not ( n14122 , n14121 );
and ( n14123 , n14120 , n14122 );
not ( n14124 , n14120 );
and ( n14125 , n14124 , n14121 );
nor ( n14126 , n14123 , n14125 );
or ( n14127 , n13857 , n13887 );
not ( n14128 , n206 );
not ( n14129 , n13596 );
and ( n14130 , n14128 , n14129 );
not ( n14131 , n13587 );
not ( n14132 , n13596 );
or ( n14133 , n14131 , n14132 );
nand ( n14134 , n14133 , n206 );
and ( n14135 , n13601 , n14134 );
nor ( n14136 , n14130 , n14135 );
and ( n14137 , n14136 , n13857 );
not ( n14138 , n2 );
nor ( n14139 , n14137 , n14138 );
nand ( n14140 , n14127 , n14139 );
nand ( n14141 , n177 , n12854 );
not ( n14142 , n13492 );
buf ( n14143 , n12978 );
not ( n14144 , n14143 );
or ( n14145 , n14142 , n14144 );
not ( n14146 , n14143 );
and ( n14147 , n13491 , n14146 );
nor ( n14148 , n14147 , n12853 );
nand ( n14149 , n14145 , n14148 );
nand ( n14150 , n14141 , n13200 , n14149 );
nand ( n14151 , n13224 , n13760 );
or ( n14152 , n13857 , n14151 );
not ( n14153 , n13579 );
not ( n14154 , n199 );
not ( n14155 , n13953 );
nand ( n14156 , n14155 , n13581 , n13585 );
not ( n14157 , n14156 );
or ( n14158 , n14154 , n14157 );
or ( n14159 , n199 , n14156 );
nand ( n14160 , n14158 , n14159 );
and ( n14161 , n13596 , n14160 );
and ( n14162 , n199 , n13597 );
nor ( n14163 , n14161 , n14162 );
not ( n14164 , n14163 );
and ( n14165 , n14153 , n14164 );
not ( n14166 , n2 );
nor ( n14167 , n14165 , n14166 );
nand ( n14168 , n14152 , n14167 );
not ( n14169 , n13292 );
nor ( n14170 , n14169 , n13401 );
and ( n14171 , n14170 , n13737 );
not ( n14172 , n14170 );
not ( n14173 , n13737 );
and ( n14174 , n14172 , n14173 );
nor ( n14175 , n14171 , n14174 );
not ( n14176 , n1708 );
nand ( n14177 , n1230 , n14176 );
not ( n14178 , n14177 );
xor ( n14179 , n173 , n167 );
and ( n14180 , n14178 , n14179 );
not ( n14181 , n14178 );
and ( n14182 , n14181 , n173 );
nor ( n14183 , n14180 , n14182 );
or ( n14184 , n226 , n250 );
not ( n14185 , n162 );
nand ( n14186 , n160 , n171 );
nand ( n14187 , n166 , n174 );
not ( n14188 , n14187 );
nand ( n14189 , n164 , n165 );
not ( n14190 , n168 );
nand ( n14191 , n169 , n167 , n173 );
nor ( n14192 , n14190 , n14191 );
and ( n14193 , n170 , n14192 );
nand ( n14194 , n163 , n14193 );
nor ( n14195 , n14189 , n14194 );
nand ( n14196 , n14188 , n14195 );
nor ( n14197 , n14186 , n14196 );
and ( n14198 , n161 , n172 , n14197 );
not ( n14199 , n14198 );
nand ( n14200 , n14185 , n14199 );
and ( n14201 , n162 , n14198 );
not ( n14202 , n14178 );
not ( n14203 , n14202 );
not ( n14204 , n14203 );
buf ( n14205 , n14204 );
not ( n14206 , n14205 );
not ( n14207 , n14206 );
not ( n14208 , n14207 );
not ( n14209 , n14208 );
nor ( n14210 , n14201 , n14209 );
and ( n14211 , n14200 , n14210 );
and ( n14212 , n162 , n14209 );
nor ( n14213 , n14211 , n14212 );
nor ( n14214 , n220 , n14213 );
not ( n14215 , n14214 );
not ( n14216 , n172 );
not ( n14217 , n14208 );
not ( n14218 , n14217 );
or ( n14219 , n14216 , n14218 );
nor ( n14220 , n172 , n14197 );
not ( n14221 , n14220 );
nand ( n14222 , n172 , n14197 );
nand ( n14223 , n14221 , n14208 , n14222 );
nand ( n14224 , n14219 , n14223 );
xor ( n14225 , n14224 , n242 );
not ( n14226 , n219 );
not ( n14227 , n161 );
not ( n14228 , n14186 );
nand ( n14229 , n165 , n166 );
and ( n14230 , n163 , n164 );
nand ( n14231 , n14230 , n14193 );
nor ( n14232 , n14229 , n14231 );
nand ( n14233 , n174 , n14232 );
not ( n14234 , n14233 );
nand ( n14235 , n14228 , n172 , n14234 );
nand ( n14236 , n14227 , n14235 );
not ( n14237 , n14235 );
and ( n14238 , n161 , n14237 );
nor ( n14239 , n14238 , n14207 );
and ( n14240 , n14236 , n14239 );
and ( n14241 , n161 , n14207 );
nor ( n14242 , n14240 , n14241 );
not ( n14243 , n14242 );
or ( n14244 , n14226 , n14243 );
or ( n14245 , n219 , n14242 );
nand ( n14246 , n14244 , n14245 );
nor ( n14247 , n14225 , n14246 );
not ( n14248 , n171 );
nand ( n14249 , n14248 , n14196 );
not ( n14250 , n14196 );
and ( n14251 , n171 , n14250 );
buf ( n14252 , n14205 );
nor ( n14253 , n14251 , n14252 );
and ( n14254 , n14249 , n14253 );
and ( n14255 , n171 , n14252 );
nor ( n14256 , n14254 , n14255 );
not ( n14257 , n231 );
and ( n14258 , n14256 , n14257 );
not ( n14259 , n14256 );
and ( n14260 , n14259 , n231 );
nor ( n14261 , n14258 , n14260 );
not ( n14262 , n14192 );
or ( n14263 , n14202 , n14191 );
nand ( n14264 , n14263 , n14190 );
and ( n14265 , n14262 , n14264 );
and ( n14266 , n168 , n14202 );
nor ( n14267 , n14265 , n14266 );
xor ( n14268 , n14267 , n411 );
not ( n14269 , n14193 );
or ( n14270 , n14202 , n14262 );
not ( n14271 , n170 );
nand ( n14272 , n14270 , n14271 );
and ( n14273 , n14269 , n14272 );
and ( n14274 , n170 , n14202 );
nor ( n14275 , n14273 , n14274 );
xor ( n14276 , n14275 , n344 );
or ( n14277 , n14202 , n14269 );
not ( n14278 , n163 );
nand ( n14279 , n14277 , n14278 );
and ( n14280 , n14194 , n14279 );
and ( n14281 , n163 , n14204 );
nor ( n14282 , n14280 , n14281 );
xor ( n14283 , n14282 , n345 );
not ( n14284 , n13572 );
not ( n14285 , n830 );
not ( n14286 , n167 );
not ( n14287 , n14177 );
or ( n14288 , n14286 , n14287 );
or ( n14289 , n167 , n14177 );
nand ( n14290 , n14288 , n14289 );
not ( n14291 , n14290 );
or ( n14292 , n14285 , n14291 );
or ( n14293 , n830 , n14290 );
nand ( n14294 , n14292 , n14293 );
xor ( n14295 , n490 , n14183 );
nand ( n14296 , n169 , n14177 );
nand ( n14297 , n167 , n173 );
or ( n14298 , n14297 , n14177 );
not ( n14299 , n169 );
nand ( n14300 , n14298 , n14299 );
nand ( n14301 , n14191 , n14300 );
and ( n14302 , n14296 , n14301 );
xor ( n14303 , n14302 , n389 );
and ( n14304 , n14284 , n14294 , n14295 , n14303 );
nand ( n14305 , n14268 , n14276 , n14283 , n14304 );
nor ( n14306 , n14261 , n14305 );
not ( n14307 , n171 );
not ( n14308 , n14234 );
or ( n14309 , n14307 , n14308 );
not ( n14310 , n160 );
nand ( n14311 , n14309 , n14310 );
and ( n14312 , n160 , n171 , n14234 );
nor ( n14313 , n14312 , n14252 );
and ( n14314 , n14311 , n14313 );
and ( n14315 , n160 , n14207 );
nor ( n14316 , n14314 , n14315 );
xor ( n14317 , n251 , n14316 );
not ( n14318 , n165 );
nand ( n14319 , n14318 , n14231 );
not ( n14320 , n14231 );
and ( n14321 , n165 , n14320 );
not ( n14322 , n14203 );
nor ( n14323 , n14321 , n14322 );
and ( n14324 , n14319 , n14323 );
and ( n14325 , n165 , n14205 );
nor ( n14326 , n14324 , n14325 );
not ( n14327 , n14326 );
and ( n14328 , n374 , n14327 );
not ( n14329 , n374 );
and ( n14330 , n14329 , n14326 );
nor ( n14331 , n14328 , n14330 );
not ( n14332 , n268 );
not ( n14333 , n166 );
not ( n14334 , n14195 );
nand ( n14335 , n14333 , n14334 );
not ( n14336 , n14335 );
and ( n14337 , n166 , n14195 );
nor ( n14338 , n14337 , n14322 );
not ( n14339 , n14338 );
or ( n14340 , n14336 , n14339 );
nand ( n14341 , n166 , n14322 );
nand ( n14342 , n14340 , n14341 );
not ( n14343 , n14342 );
and ( n14344 , n14332 , n14343 );
and ( n14345 , n268 , n14342 );
nor ( n14346 , n14344 , n14345 );
nor ( n14347 , n14331 , n14346 );
not ( n14348 , n269 );
not ( n14349 , n164 );
not ( n14350 , n14322 );
or ( n14351 , n14349 , n14350 );
not ( n14352 , n164 );
not ( n14353 , n14352 );
not ( n14354 , n14194 );
or ( n14355 , n14353 , n14354 );
not ( n14356 , n14194 );
and ( n14357 , n164 , n14356 );
nor ( n14358 , n14357 , n14322 );
nand ( n14359 , n14355 , n14358 );
nand ( n14360 , n14351 , n14359 );
not ( n14361 , n14360 );
or ( n14362 , n14348 , n14361 );
or ( n14363 , n269 , n14360 );
nand ( n14364 , n14362 , n14363 );
not ( n14365 , n249 );
not ( n14366 , n174 );
not ( n14367 , n14252 );
or ( n14368 , n14366 , n14367 );
nor ( n14369 , n174 , n14232 );
not ( n14370 , n14369 );
nand ( n14371 , n14370 , n14206 , n14233 );
nand ( n14372 , n14368 , n14371 );
not ( n14373 , n14372 );
or ( n14374 , n14365 , n14373 );
or ( n14375 , n249 , n14372 );
nand ( n14376 , n14374 , n14375 );
and ( n14377 , n14347 , n14364 , n14376 );
and ( n14378 , n14306 , n14317 , n14377 );
nand ( n14379 , n220 , n14213 );
nand ( n14380 , n14215 , n14247 , n14378 , n14379 );
not ( n14381 , n14380 );
or ( n14382 , n14183 , n14184 , n14381 );
nand ( n14383 , n1134 , n14184 );
nand ( n14384 , n14382 , n14383 );
and ( n14385 , n12574 , n12617 );
nor ( n14386 , n14385 , n12718 );
not ( n14387 , n14385 );
not ( n14388 , n12718 );
or ( n14389 , n14387 , n14388 );
nand ( n14390 , n14389 , n12726 );
or ( n14391 , n14386 , n14390 );
not ( n14392 , n961 );
or ( n14393 , n14392 , n12726 );
nand ( n14394 , n14391 , n14393 );
not ( n14395 , n12619 );
nor ( n14396 , n12783 , n14395 );
nor ( n14397 , n14396 , n13433 );
not ( n14398 , n14396 );
not ( n14399 , n13433 );
or ( n14400 , n14398 , n14399 );
nand ( n14401 , n14400 , n12726 );
or ( n14402 , n14397 , n14401 );
not ( n14403 , n886 );
or ( n14404 , n14403 , n12726 );
nand ( n14405 , n14402 , n14404 );
or ( n14406 , n14282 , n14184 , n14381 );
nand ( n14407 , n1138 , n14184 );
nand ( n14408 , n14406 , n14407 );
or ( n14409 , n14302 , n14184 , n14381 );
nand ( n14410 , n1135 , n14184 );
nand ( n14411 , n14409 , n14410 );
or ( n14412 , n14275 , n14184 , n14381 );
nand ( n14413 , n1137 , n14184 );
nand ( n14414 , n14412 , n14413 );
not ( n14415 , n14380 );
or ( n14416 , n14267 , n14184 , n14415 );
nand ( n14417 , n1136 , n14184 );
nand ( n14418 , n14416 , n14417 );
nand ( n14419 , n179 , n12854 );
not ( n14420 , n13483 );
not ( n14421 , n13121 );
not ( n14422 , n14421 );
or ( n14423 , n14420 , n14422 );
and ( n14424 , n13475 , n13121 );
nor ( n14425 , n14424 , n12853 );
nand ( n14426 , n14423 , n14425 );
nand ( n14427 , n14419 , n13200 , n14426 );
nand ( n14428 , n182 , n12853 );
not ( n14429 , n12939 );
not ( n14430 , n14429 );
not ( n14431 , n13176 );
not ( n14432 , n14431 );
and ( n14433 , n13060 , n14432 );
not ( n14434 , n13060 );
and ( n14435 , n14434 , n14431 );
nor ( n14436 , n14433 , n14435 );
not ( n14437 , n14436 );
not ( n14438 , n14437 );
or ( n14439 , n14430 , n14438 );
not ( n14440 , n14429 );
and ( n14441 , n14440 , n14436 );
nor ( n14442 , n14441 , n12853 );
nand ( n14443 , n14439 , n14442 );
nand ( n14444 , n14428 , n13200 , n14443 );
not ( n14445 , n13224 );
nand ( n14446 , n256 , n14445 );
nand ( n14447 , n255 , n13249 );
nand ( n14448 , n14446 , n14447 );
nand ( n14449 , n248 , n13241 );
nor ( n14450 , n230 , n13289 );
and ( n14451 , n14449 , n14450 );
nor ( n14452 , n248 , n13241 );
nor ( n14453 , n14451 , n14452 );
or ( n14454 , n14448 , n14453 );
not ( n14455 , n14446 );
not ( n14456 , n255 );
nand ( n14457 , n14456 , n13253 );
or ( n14458 , n14455 , n14457 );
nand ( n14459 , n14454 , n14458 );
nand ( n14460 , n230 , n13289 );
nand ( n14461 , n14449 , n14460 );
nor ( n14462 , n14448 , n14461 );
not ( n14463 , n14462 );
not ( n14464 , n13396 );
nand ( n14465 , n229 , n14464 );
not ( n14466 , n14465 );
nand ( n14467 , n228 , n13624 );
not ( n14468 , n14467 );
nor ( n14469 , n14466 , n14468 );
nand ( n14470 , n236 , n13323 );
nand ( n14471 , n227 , n13309 );
and ( n14472 , n14470 , n14471 );
and ( n14473 , n14469 , n14472 );
not ( n14474 , n14473 );
nand ( n14475 , n246 , n13657 );
not ( n14476 , n14475 );
not ( n14477 , n235 );
nand ( n14478 , n14477 , n13783 );
or ( n14479 , n14476 , n14478 );
nor ( n14480 , n246 , n13657 );
not ( n14481 , n14480 );
nand ( n14482 , n14479 , n14481 );
not ( n14483 , n14482 );
nand ( n14484 , n235 , n13782 );
and ( n14485 , n14475 , n14484 );
nand ( n14486 , n234 , n13347 );
not ( n14487 , n14486 );
nand ( n14488 , n233 , n13359 );
not ( n14489 , n14488 );
nand ( n14490 , n232 , n13649 );
not ( n14491 , n14490 );
or ( n14492 , n14489 , n14491 );
not ( n14493 , n233 );
nand ( n14494 , n14493 , n13358 );
nand ( n14495 , n14492 , n14494 );
not ( n14496 , n14495 );
or ( n14497 , n14487 , n14496 );
not ( n14498 , n234 );
and ( n14499 , n14498 , n13346 );
not ( n14500 , n14499 );
nand ( n14501 , n14497 , n14500 );
nand ( n14502 , n14485 , n14501 );
nand ( n14503 , n14483 , n14502 );
not ( n14504 , n14503 );
or ( n14505 , n14474 , n14504 );
or ( n14506 , n228 , n13301 );
not ( n14507 , n14506 );
and ( n14508 , n14465 , n14507 );
nor ( n14509 , n229 , n13397 );
nor ( n14510 , n14508 , n14509 );
nor ( n14511 , n227 , n13309 );
not ( n14512 , n14511 );
nor ( n14513 , n236 , n13323 );
nand ( n14514 , n14471 , n14513 );
nand ( n14515 , n14512 , n14514 );
nand ( n14516 , n14469 , n14515 );
and ( n14517 , n14510 , n14516 );
nand ( n14518 , n14505 , n14517 );
not ( n14519 , n14518 );
or ( n14520 , n14463 , n14519 );
not ( n14521 , n256 );
nand ( n14522 , n14521 , n13224 );
nand ( n14523 , n14520 , n14522 );
nor ( n14524 , n14459 , n14523 );
not ( n14525 , n252 );
not ( n14526 , n13231 );
and ( n14527 , n14525 , n14526 );
and ( n14528 , n252 , n13231 );
nor ( n14529 , n14527 , n14528 );
and ( n14530 , n14524 , n14529 );
not ( n14531 , n14524 );
not ( n14532 , n14529 );
and ( n14533 , n14531 , n14532 );
nor ( n14534 , n14530 , n14533 );
nor ( n14535 , n13937 , n14046 );
nor ( n14536 , n13937 , n14031 );
nor ( n14537 , n13937 , n14151 );
nand ( n14538 , n365 , n13249 );
and ( n14539 , n14538 , n13697 );
not ( n14540 , n1103 );
nor ( n14541 , n14539 , n14540 );
nand ( n14542 , n365 , n13241 );
not ( n14543 , n371 );
not ( n14544 , n13615 );
not ( n14545 , n14544 );
not ( n14546 , n353 );
not ( n14547 , n13617 );
and ( n14548 , n14546 , n14547 );
not ( n14549 , n372 );
and ( n14550 , n14549 , n13279 );
nor ( n14551 , n14548 , n14550 );
not ( n14552 , n353 );
nand ( n14553 , n14552 , n14549 );
nand ( n14554 , n14545 , n14551 , n14553 );
nand ( n14555 , n14543 , n13387 , n14554 );
not ( n14556 , n14553 );
not ( n14557 , n13948 );
and ( n14558 , n14556 , n14557 );
nor ( n14559 , n372 , n13612 );
nor ( n14560 , n14558 , n14559 );
nand ( n14561 , n13632 , n13864 );
or ( n14562 , n370 , n14561 );
nor ( n14563 , n370 , n371 );
nand ( n14564 , n14563 , n13864 );
nand ( n14565 , n14562 , n14564 );
and ( n14566 , n14565 , n14554 );
and ( n14567 , n14552 , n14544 );
nor ( n14568 , n14566 , n14567 );
nand ( n14569 , n14555 , n14560 , n14568 );
nand ( n14570 , n14542 , n14569 );
nand ( n14571 , n14541 , n13613 , n14570 );
nand ( n14572 , n366 , n386 );
and ( n14573 , n14572 , n13358 );
nor ( n14574 , n366 , n386 );
and ( n14575 , n366 , n13359 );
nor ( n14576 , n14575 , n13757 );
nor ( n14577 , n14573 , n14574 , n14576 );
or ( n14578 , n367 , n13785 );
or ( n14579 , n368 , n13882 );
nand ( n14580 , n14578 , n14579 );
nor ( n14581 , n367 , n368 );
not ( n14582 , n13669 );
nor ( n14583 , n14580 , n14581 , n14582 );
not ( n14584 , n13327 );
or ( n14585 , n369 , n14584 );
or ( n14586 , n350 , n13657 );
nand ( n14587 , n14585 , n14586 );
nor ( n14588 , n350 , n369 );
nor ( n14589 , n14587 , n14588 , n13676 );
nor ( n14590 , n14577 , n14583 , n14589 );
not ( n14591 , n368 );
and ( n14592 , n14591 , n13784 );
not ( n14593 , n367 );
and ( n14594 , n14593 , n14582 );
and ( n14595 , n14581 , n13881 );
nor ( n14596 , n14592 , n14594 , n14595 );
or ( n14597 , n14596 , n14589 );
not ( n14598 , n13676 );
or ( n14599 , n369 , n14598 );
not ( n14600 , n350 );
not ( n14601 , n13797 );
and ( n14602 , n14600 , n14601 );
and ( n14603 , n14588 , n13317 );
nor ( n14604 , n14602 , n14603 );
nand ( n14605 , n14597 , n14599 , n14604 );
or ( n14606 , n14571 , n14590 , n14605 );
or ( n14607 , n371 , n13865 );
or ( n14608 , n370 , n13896 );
not ( n14609 , n14561 );
nor ( n14610 , n14563 , n14609 );
nand ( n14611 , n14607 , n14608 , n14610 );
and ( n14612 , n14611 , n14542 , n14554 );
or ( n14613 , n14612 , n14571 );
nand ( n14614 , n14606 , n14613 );
not ( n14615 , n13887 );
nor ( n14616 , n12650 , n12798 );
not ( n14617 , n12816 );
nor ( n14618 , n14616 , n14617 );
not ( n14619 , n14616 );
not ( n14620 , n14617 );
or ( n14621 , n14619 , n14620 );
nand ( n14622 , n14621 , n12726 );
or ( n14623 , n14618 , n14622 );
not ( n14624 , n960 );
or ( n14625 , n14624 , n12726 );
nand ( n14626 , n14623 , n14625 );
not ( n14627 , n14316 );
not ( n14628 , n14184 );
nand ( n14629 , n14627 , n14628 );
not ( n14630 , n14380 );
or ( n14631 , n14629 , n14630 );
or ( n14632 , n13226 , n14628 );
nand ( n14633 , n14631 , n14632 );
not ( n14634 , n14242 );
nand ( n14635 , n14628 , n14634 );
or ( n14636 , n14635 , n14630 );
not ( n14637 , n1132 );
or ( n14638 , n14637 , n14628 );
nand ( n14639 , n14636 , n14638 );
not ( n14640 , n14213 );
nand ( n14641 , n14628 , n14640 );
or ( n14642 , n14641 , n14630 );
not ( n14643 , n1133 );
or ( n14644 , n14643 , n14628 );
nand ( n14645 , n14642 , n14644 );
nand ( n14646 , n14628 , n14360 );
or ( n14647 , n14646 , n14630 );
not ( n14648 , n1139 );
or ( n14649 , n14648 , n14628 );
nand ( n14650 , n14647 , n14649 );
nand ( n14651 , n14628 , n14327 );
or ( n14652 , n14651 , n14630 );
or ( n14653 , n13282 , n14628 );
nand ( n14654 , n14652 , n14653 );
nand ( n14655 , n14628 , n14342 );
or ( n14656 , n14655 , n14630 );
or ( n14657 , n13235 , n14628 );
nand ( n14658 , n14656 , n14657 );
nand ( n14659 , n14628 , n14290 );
or ( n14660 , n14659 , n14415 );
nand ( n14661 , n1128 , n14184 );
nand ( n14662 , n14660 , n14661 );
not ( n14663 , n14256 );
nand ( n14664 , n14663 , n14628 );
or ( n14665 , n14664 , n14630 );
not ( n14666 , n1129 );
or ( n14667 , n14666 , n14628 );
nand ( n14668 , n14665 , n14667 );
nand ( n14669 , n14628 , n14224 );
or ( n14670 , n14669 , n14415 );
or ( n14671 , n13408 , n14628 );
nand ( n14672 , n14670 , n14671 );
nand ( n14673 , n14628 , n14372 );
or ( n14674 , n14673 , n14415 );
or ( n14675 , n13244 , n14628 );
nand ( n14676 , n14674 , n14675 );
nand ( n14677 , n181 , n12854 );
not ( n14678 , n13481 );
not ( n14679 , n13028 );
not ( n14680 , n14679 );
or ( n14681 , n14678 , n14680 );
not ( n14682 , n13481 );
not ( n14683 , n14679 );
and ( n14684 , n14682 , n14683 );
nor ( n14685 , n14684 , n12853 );
nand ( n14686 , n14681 , n14685 );
nand ( n14687 , n14677 , n13200 , n14686 );
nand ( n14688 , n189 , n12853 );
not ( n14689 , n12971 );
not ( n14690 , n14689 );
not ( n14691 , n13038 );
not ( n14692 , n13019 );
not ( n14693 , n14692 );
and ( n14694 , n14691 , n14693 );
and ( n14695 , n13038 , n14692 );
nor ( n14696 , n14694 , n14695 );
not ( n14697 , n14696 );
not ( n14698 , n14697 );
or ( n14699 , n14690 , n14698 );
not ( n14700 , n14689 );
and ( n14701 , n14700 , n14696 );
nor ( n14702 , n14701 , n12853 );
nand ( n14703 , n14699 , n14702 );
nand ( n14704 , n14688 , n13200 , n14703 );
nand ( n14705 , n14467 , n14471 );
not ( n14706 , n14705 );
and ( n14707 , n14465 , n14460 );
and ( n14708 , n14706 , n14707 );
not ( n14709 , n14708 );
and ( n14710 , n14475 , n14470 );
not ( n14711 , n14710 );
nand ( n14712 , n14495 , n14486 , n14484 );
nor ( n14713 , n14711 , n14712 );
not ( n14714 , n14713 );
or ( n14715 , n14709 , n14714 );
not ( n14716 , n14706 );
not ( n14717 , n14710 );
nand ( n14718 , n14484 , n14499 );
nand ( n14719 , n14478 , n14718 );
not ( n14720 , n14719 );
or ( n14721 , n14717 , n14720 );
and ( n14722 , n14480 , n14470 );
nor ( n14723 , n14722 , n14513 );
nand ( n14724 , n14721 , n14723 );
not ( n14725 , n14724 );
or ( n14726 , n14716 , n14725 );
nand ( n14727 , n14467 , n14511 );
and ( n14728 , n14506 , n14727 );
nand ( n14729 , n14726 , n14728 );
and ( n14730 , n14707 , n14729 );
and ( n14731 , n14509 , n14460 );
nor ( n14732 , n14731 , n14450 );
not ( n14733 , n14732 );
nor ( n14734 , n14730 , n14733 );
nand ( n14735 , n14715 , n14734 );
not ( n14736 , n14452 );
nand ( n14737 , n14736 , n14449 );
not ( n14738 , n14737 );
and ( n14739 , n14735 , n14738 );
not ( n14740 , n14735 );
and ( n14741 , n14740 , n14737 );
nor ( n14742 , n14739 , n14741 );
not ( n14743 , n14151 );
not ( n14744 , n14031 );
not ( n14745 , n14046 );
not ( n14746 , n14461 );
not ( n14747 , n14502 );
nand ( n14748 , n14746 , n14473 , n14747 );
not ( n14749 , n14469 );
not ( n14750 , n14472 );
not ( n14751 , n14482 );
or ( n14752 , n14750 , n14751 );
not ( n14753 , n14515 );
nand ( n14754 , n14752 , n14753 );
not ( n14755 , n14754 );
or ( n14756 , n14749 , n14755 );
nand ( n14757 , n14756 , n14510 );
nand ( n14758 , n14746 , n14757 );
nand ( n14759 , n14748 , n14453 , n14758 );
nand ( n14760 , n14457 , n14447 );
not ( n14761 , n14760 );
and ( n14762 , n14759 , n14761 );
not ( n14763 , n14759 );
and ( n14764 , n14763 , n14760 );
nor ( n14765 , n14762 , n14764 );
nand ( n14766 , n13257 , n13225 );
not ( n14767 , n14766 );
not ( n14768 , n13402 );
and ( n14769 , n13311 , n13329 );
nor ( n14770 , n14769 , n13393 );
not ( n14771 , n14770 );
nand ( n14772 , n14771 , n13293 );
not ( n14773 , n14772 );
or ( n14774 , n14768 , n14773 );
nand ( n14775 , n14774 , n13263 );
not ( n14776 , n13255 );
and ( n14777 , n13383 , n13311 );
nand ( n14778 , n13340 , n13378 );
nand ( n14779 , n13263 , n13293 , n14777 , n14778 );
nand ( n14780 , n14775 , n14776 , n14779 );
not ( n14781 , n14780 );
or ( n14782 , n14767 , n14781 );
or ( n14783 , n14766 , n14780 );
nand ( n14784 , n14782 , n14783 );
nor ( n14785 , n222 , n13197 );
nor ( n14786 , n197 , n14785 );
nor ( n14787 , n74 , n14786 );
not ( n14788 , n14787 );
nor ( n14789 , n1796 , n14788 );
nand ( n14790 , n149 , n14789 );
nor ( n14791 , n194 , n222 );
nor ( n14792 , n14791 , n14787 );
not ( n14793 , n14792 );
nand ( n14794 , n1558 , n12833 , n12845 );
nand ( n14795 , n14794 , n12835 );
nand ( n14796 , n12839 , n12847 );
not ( n14797 , n13197 );
not ( n14798 , n184 );
and ( n14799 , n12832 , n12845 );
and ( n14800 , n188 , n14798 , n14799 );
not ( n14801 , n14800 );
or ( n14802 , n14797 , n14801 );
and ( n14803 , n223 , n13196 );
nand ( n14804 , n14803 , n14800 );
nand ( n14805 , n14802 , n14804 );
or ( n14806 , n14795 , n14796 , n14805 );
or ( n14807 , n14806 , n14432 );
not ( n14808 , n14806 );
buf ( n14809 , n12850 );
not ( n14810 , n14809 );
and ( n14811 , n13058 , n14810 );
not ( n14812 , n14809 );
nor ( n14813 , n177 , n14812 );
nor ( n14814 , n14811 , n14813 );
or ( n14815 , n14808 , n14814 );
nand ( n14816 , n1551 , n1821 );
and ( n14817 , n14816 , n14794 , n12849 );
not ( n14818 , n14817 );
not ( n14819 , n14818 );
nand ( n14820 , n14819 , n14806 );
nand ( n14821 , n14807 , n14815 , n14820 );
nand ( n14822 , n14788 , n14821 );
nand ( n14823 , n14790 , n14793 , n14822 );
nand ( n14824 , n180 , n12853 );
not ( n14825 , n13842 );
not ( n14826 , n14825 );
and ( n14827 , n12995 , n13044 );
not ( n14828 , n12995 );
and ( n14829 , n14828 , n13043 );
nor ( n14830 , n14827 , n14829 );
not ( n14831 , n14830 );
not ( n14832 , n14831 );
or ( n14833 , n14826 , n14832 );
and ( n14834 , n13842 , n14830 );
nor ( n14835 , n14834 , n12853 );
nand ( n14836 , n14833 , n14835 );
nand ( n14837 , n14824 , n13200 , n14836 );
not ( n14838 , n12853 );
or ( n14839 , n13039 , n14838 );
not ( n14840 , n138 );
not ( n14841 , n139 );
buf ( n14842 , n13175 );
not ( n14843 , n14842 );
and ( n14844 , n14841 , n14843 );
and ( n14845 , n139 , n14842 );
nor ( n14846 , n14844 , n14845 );
not ( n14847 , n14846 );
not ( n14848 , n14847 );
or ( n14849 , n14840 , n14848 );
and ( n14850 , n12825 , n14846 );
nor ( n14851 , n14850 , n12853 );
nand ( n14852 , n14849 , n14851 );
nand ( n14853 , n14839 , n13200 , n14852 );
not ( n14854 , n129 );
not ( n14855 , n14789 );
or ( n14856 , n14854 , n14855 );
not ( n14857 , n133 );
not ( n14858 , n134 );
and ( n14859 , n14857 , n14858 );
and ( n14860 , n133 , n134 );
nor ( n14861 , n14859 , n14860 );
or ( n14862 , n14791 , n14861 );
not ( n14863 , n14808 );
not ( n14864 , n14689 );
or ( n14865 , n14863 , n14864 );
nand ( n14866 , n1111 , n14819 );
not ( n14867 , n908 );
not ( n14868 , n14809 );
not ( n14869 , n14868 );
or ( n14870 , n14867 , n14869 );
and ( n14871 , n181 , n12850 );
nor ( n14872 , n14871 , n14817 );
nand ( n14873 , n14870 , n14872 );
nand ( n14874 , n14866 , n14806 , n14873 );
nand ( n14875 , n14865 , n14874 );
nand ( n14876 , n14791 , n14875 );
nand ( n14877 , n14862 , n14788 , n14876 );
nand ( n14878 , n14856 , n14877 );
not ( n14879 , n131 );
not ( n14880 , n14789 );
or ( n14881 , n14879 , n14880 );
or ( n14882 , n134 , n14791 );
nand ( n14883 , n14882 , n14788 );
not ( n14884 , n14808 );
not ( n14885 , n14819 );
or ( n14886 , n189 , n14810 );
or ( n14887 , n907 , n14809 );
nand ( n14888 , n14886 , n14887 );
and ( n14889 , n14885 , n14888 );
and ( n14890 , n1145 , n14819 );
nor ( n14891 , n14889 , n14890 );
not ( n14892 , n14891 );
and ( n14893 , n14884 , n14892 );
not ( n14894 , n14808 );
not ( n14895 , n14429 );
or ( n14896 , n14894 , n14895 );
nand ( n14897 , n14896 , n14791 );
nor ( n14898 , n14893 , n14897 );
or ( n14899 , n14883 , n14898 );
nand ( n14900 , n14881 , n14899 );
not ( n14901 , n132 );
not ( n14902 , n14789 );
or ( n14903 , n14901 , n14902 );
not ( n14904 , n14791 );
nand ( n14905 , n134 , n14904 );
and ( n14906 , n12850 , n139 );
not ( n14907 , n12850 );
and ( n14908 , n14907 , n183 );
nor ( n14909 , n14906 , n14908 );
and ( n14910 , n14818 , n14909 );
not ( n14911 , n1145 );
and ( n14912 , n14911 , n14817 );
nor ( n14913 , n14910 , n14912 );
nor ( n14914 , n14808 , n14913 );
not ( n14915 , n14914 );
nand ( n14916 , n14808 , n13842 );
nand ( n14917 , n14915 , n14791 , n14916 );
nand ( n14918 , n14905 , n14788 , n14917 );
nand ( n14919 , n14903 , n14918 );
not ( n14920 , n959 );
not ( n14921 , n1228 );
or ( n14922 , n14920 , n14921 );
nor ( n14923 , n12637 , n12654 );
not ( n14924 , n14923 );
not ( n14925 , n14924 );
not ( n14926 , n12716 );
not ( n14927 , n14926 );
or ( n14928 , n14925 , n14927 );
and ( n14929 , n14923 , n12716 );
nor ( n14930 , n14929 , n1228 );
nand ( n14931 , n14928 , n14930 );
nand ( n14932 , n14922 , n14931 );
or ( n14933 , n13399 , n13280 );
not ( n14934 , n14933 );
nand ( n14935 , n14777 , n14778 );
nand ( n14936 , n14770 , n14935 );
not ( n14937 , n14936 );
or ( n14938 , n14934 , n14937 );
or ( n14939 , n14933 , n14936 );
nand ( n14940 , n14938 , n14939 );
nand ( n14941 , n14111 , n14117 );
nand ( n14942 , n13388 , n13302 );
not ( n14943 , n14942 );
and ( n14944 , n14941 , n14943 );
not ( n14945 , n14941 );
and ( n14946 , n14945 , n14942 );
nor ( n14947 , n14944 , n14946 );
not ( n14948 , n14522 );
nor ( n14949 , n14948 , n14455 );
not ( n14950 , n14949 );
and ( n14951 , n14447 , n14449 , n14707 );
nor ( n14952 , n14711 , n14705 );
not ( n14953 , n14952 );
not ( n14954 , n14719 );
nand ( n14955 , n14954 , n14712 );
not ( n14956 , n14955 );
or ( n14957 , n14953 , n14956 );
not ( n14958 , n14723 );
nand ( n14959 , n14958 , n14706 );
and ( n14960 , n14728 , n14959 );
nand ( n14961 , n14957 , n14960 );
and ( n14962 , n14951 , n14961 );
not ( n14963 , n14449 );
or ( n14964 , n14963 , n14732 );
nand ( n14965 , n14964 , n14736 );
nand ( n14966 , n14447 , n14965 );
nand ( n14967 , n14457 , n14966 );
nor ( n14968 , n14962 , n14967 );
not ( n14969 , n14968 );
or ( n14970 , n14950 , n14969 );
or ( n14971 , n14949 , n14968 );
nand ( n14972 , n14970 , n14971 );
not ( n14973 , n1251 );
not ( n14974 , n1819 );
not ( n14975 , n508 );
nand ( n14976 , n1559 , n1700 );
nand ( n14977 , n1176 , n1559 );
nand ( n14978 , n1559 , n1655 );
and ( n14979 , n14976 , n14977 , n14978 );
not ( n14980 , n14979 );
not ( n14981 , n14980 );
not ( n14982 , n14981 );
not ( n14983 , n14982 );
not ( n14984 , n14983 );
or ( n14985 , n14975 , n14984 );
not ( n14986 , n508 );
not ( n14987 , n14986 );
not ( n14988 , n515 );
nand ( n14989 , n14988 , n1396 );
not ( n14990 , n595 );
nand ( n14991 , n1248 , n14990 );
and ( n14992 , n14989 , n14991 );
not ( n14993 , n1399 );
nor ( n14994 , n14993 , n516 );
not ( n14995 , n14994 );
not ( n14996 , n609 );
nand ( n14997 , n1403 , n14996 );
and ( n14998 , n14995 , n14997 );
nand ( n14999 , n14992 , n14998 );
not ( n15000 , n613 );
nand ( n15001 , n15000 , n1250 );
not ( n15002 , n638 );
nand ( n15003 , n1401 , n15002 );
and ( n15004 , n15001 , n15003 );
not ( n15005 , n637 );
nand ( n15006 , n1152 , n15005 );
not ( n15007 , n537 );
nand ( n15008 , n1151 , n15007 );
not ( n15009 , n15008 );
not ( n15010 , n636 );
nand ( n15011 , n15010 , n1406 );
not ( n15012 , n15011 );
nor ( n15013 , n15009 , n15012 );
nand ( n15014 , n15006 , n15013 );
not ( n15015 , n15014 );
nand ( n15016 , n15004 , n15015 );
nor ( n15017 , n14999 , n15016 );
not ( n15018 , n14992 );
not ( n15019 , n14998 );
not ( n15020 , n1250 );
nand ( n15021 , n15020 , n613 );
not ( n15022 , n1401 );
nand ( n15023 , n15022 , n638 );
nand ( n15024 , n15021 , n15023 );
not ( n15025 , n15024 );
not ( n15026 , n15006 );
not ( n15027 , n636 );
nor ( n15028 , n15027 , n1406 );
not ( n15029 , n15028 );
or ( n15030 , n15026 , n15029 );
not ( n15031 , n1152 );
nand ( n15032 , n15031 , n637 );
nand ( n15033 , n15030 , n15032 );
not ( n15034 , n15033 );
nand ( n15035 , n15025 , n15034 );
not ( n15036 , n15001 );
nand ( n15037 , n15021 , n15036 );
not ( n15038 , n15037 );
nand ( n15039 , n15038 , n15034 );
not ( n15040 , n15004 );
nand ( n15041 , n15024 , n15037 );
nand ( n15042 , n15040 , n15041 );
nand ( n15043 , n15035 , n15039 , n15042 );
not ( n15044 , n15043 );
not ( n15045 , n15044 );
or ( n15046 , n15019 , n15045 );
not ( n15047 , n14994 );
not ( n15048 , n1403 );
nand ( n15049 , n15048 , n609 );
not ( n15050 , n15049 );
and ( n15051 , n15047 , n15050 );
not ( n15052 , n516 );
nor ( n15053 , n15052 , n1399 );
nor ( n15054 , n15051 , n15053 );
nand ( n15055 , n15046 , n15054 );
not ( n15056 , n15055 );
or ( n15057 , n15018 , n15056 );
not ( n15058 , n515 );
nor ( n15059 , n15058 , n1396 );
and ( n15060 , n14991 , n15059 );
nor ( n15061 , n14990 , n1248 );
nor ( n15062 , n15060 , n15061 );
nand ( n15063 , n15057 , n15062 );
nor ( n15064 , n15017 , n15063 );
not ( n15065 , n15064 );
not ( n15066 , n15065 );
or ( n15067 , n14987 , n15066 );
and ( n15068 , n508 , n15064 );
nor ( n15069 , n15068 , n14983 );
nand ( n15070 , n15067 , n15069 );
nand ( n15071 , n14985 , n15070 );
and ( n15072 , n14974 , n15071 );
nand ( n15073 , n515 , n516 );
not ( n15074 , n15073 );
nand ( n15075 , n537 , n636 );
not ( n15076 , n15075 );
nand ( n15077 , n637 , n638 );
not ( n15078 , n15077 );
nand ( n15079 , n613 , n15076 , n15078 );
not ( n15080 , n15079 );
nand ( n15081 , n595 , n609 , n15074 , n15080 );
and ( n15082 , n15081 , n14986 );
not ( n15083 , n15081 );
and ( n15084 , n15083 , n508 );
nor ( n15085 , n15082 , n15084 );
and ( n15086 , n1819 , n15085 );
nor ( n15087 , n15072 , n15086 );
nor ( n15088 , n14973 , n15087 );
not ( n15089 , n1272 );
not ( n15090 , n1826 );
not ( n15091 , n487 );
or ( n15092 , n1655 , n1698 );
nand ( n15093 , n15092 , n1588 );
nand ( n15094 , n1176 , n1588 );
nand ( n15095 , n15093 , n15094 );
not ( n15096 , n15095 );
not ( n15097 , n15096 );
not ( n15098 , n15097 );
not ( n15099 , n15098 );
not ( n15100 , n15099 );
not ( n15101 , n15100 );
or ( n15102 , n15091 , n15101 );
not ( n15103 , n487 );
not ( n15104 , n15103 );
not ( n15105 , n695 );
nand ( n15106 , n15105 , n1163 );
not ( n15107 , n752 );
nand ( n15108 , n1268 , n15107 );
and ( n15109 , n15106 , n15108 );
not ( n15110 , n1394 );
nor ( n15111 , n15110 , n698 );
not ( n15112 , n15111 );
not ( n15113 , n777 );
nand ( n15114 , n1271 , n15113 );
and ( n15115 , n15112 , n15114 );
nand ( n15116 , n15109 , n15115 );
not ( n15117 , n779 );
nand ( n15118 , n15117 , n1162 );
not ( n15119 , n783 );
nand ( n15120 , n1387 , n15119 );
and ( n15121 , n15118 , n15120 );
not ( n15122 , n782 );
nand ( n15123 , n1270 , n15122 );
not ( n15124 , n715 );
nand ( n15125 , n1161 , n15124 );
not ( n15126 , n791 );
nand ( n15127 , n1471 , n15126 );
nand ( n15128 , n15125 , n15127 );
not ( n15129 , n15128 );
nand ( n15130 , n15123 , n15129 );
not ( n15131 , n15130 );
nand ( n15132 , n15121 , n15131 );
nor ( n15133 , n15116 , n15132 );
not ( n15134 , n15109 );
not ( n15135 , n15115 );
not ( n15136 , n1162 );
nand ( n15137 , n15136 , n779 );
not ( n15138 , n1387 );
nand ( n15139 , n15138 , n783 );
nand ( n15140 , n15137 , n15139 );
not ( n15141 , n15140 );
not ( n15142 , n15123 );
not ( n15143 , n791 );
nor ( n15144 , n15143 , n1471 );
not ( n15145 , n15144 );
or ( n15146 , n15142 , n15145 );
not ( n15147 , n1270 );
nand ( n15148 , n15147 , n782 );
nand ( n15149 , n15146 , n15148 );
not ( n15150 , n15149 );
nand ( n15151 , n15141 , n15150 );
not ( n15152 , n15118 );
nand ( n15153 , n15137 , n15152 );
not ( n15154 , n15153 );
nand ( n15155 , n15154 , n15150 );
not ( n15156 , n15121 );
nand ( n15157 , n15140 , n15153 );
nand ( n15158 , n15156 , n15157 );
nand ( n15159 , n15151 , n15155 , n15158 );
not ( n15160 , n15159 );
not ( n15161 , n15160 );
or ( n15162 , n15135 , n15161 );
not ( n15163 , n15111 );
not ( n15164 , n1271 );
nand ( n15165 , n15164 , n777 );
not ( n15166 , n15165 );
and ( n15167 , n15163 , n15166 );
not ( n15168 , n698 );
nor ( n15169 , n15168 , n1394 );
nor ( n15170 , n15167 , n15169 );
nand ( n15171 , n15162 , n15170 );
not ( n15172 , n15171 );
or ( n15173 , n15134 , n15172 );
not ( n15174 , n695 );
nor ( n15175 , n15174 , n1163 );
and ( n15176 , n15108 , n15175 );
nor ( n15177 , n15107 , n1268 );
nor ( n15178 , n15176 , n15177 );
nand ( n15179 , n15173 , n15178 );
nor ( n15180 , n15133 , n15179 );
not ( n15181 , n15180 );
not ( n15182 , n15181 );
or ( n15183 , n15104 , n15182 );
and ( n15184 , n487 , n15180 );
nor ( n15185 , n15184 , n15100 );
nand ( n15186 , n15183 , n15185 );
nand ( n15187 , n15102 , n15186 );
and ( n15188 , n15090 , n15187 );
nand ( n15189 , n695 , n698 );
not ( n15190 , n15189 );
not ( n15191 , n779 );
nand ( n15192 , n782 , n783 );
nand ( n15193 , n715 , n791 );
nor ( n15194 , n15191 , n15192 , n15193 );
nand ( n15195 , n752 , n777 , n15190 , n15194 );
and ( n15196 , n15195 , n15103 );
not ( n15197 , n15195 );
and ( n15198 , n15197 , n487 );
nor ( n15199 , n15196 , n15198 );
and ( n15200 , n1826 , n15199 );
nor ( n15201 , n15188 , n15200 );
nor ( n15202 , n15089 , n15201 );
not ( n15203 , n1230 );
not ( n15204 , n15203 );
not ( n15205 , n438 );
not ( n15206 , n465 );
not ( n15207 , n1499 );
not ( n15208 , n1220 );
nor ( n15209 , n538 , n1217 );
nand ( n15210 , n15207 , n15208 , n15209 );
nor ( n15211 , n789 , n15210 );
nand ( n15212 , n1219 , n15205 , n15206 , n15211 );
nor ( n15213 , n15208 , n1499 );
nor ( n15214 , n465 , n789 );
nor ( n15215 , n438 , n1219 );
and ( n15216 , n15213 , n15209 , n15214 , n15215 );
not ( n15217 , n1217 );
nor ( n15218 , n15217 , n1499 );
not ( n15219 , n538 );
and ( n15220 , n15208 , n15214 , n15215 );
and ( n15221 , n15218 , n15219 , n15220 );
nor ( n15222 , n15216 , n15221 );
and ( n15223 , n15212 , n15222 );
not ( n15224 , n15212 );
and ( n15225 , n15224 , n267 );
nor ( n15226 , n15223 , n15225 );
not ( n15227 , n15226 );
or ( n15228 , n15204 , n15227 );
not ( n15229 , n325 );
nand ( n15230 , n15228 , n15229 );
not ( n15231 , n15230 );
not ( n15232 , n15231 );
not ( n15233 , n15230 );
nand ( n15234 , n15233 , n775 );
not ( n15235 , n15234 );
not ( n15236 , n15235 );
not ( n15237 , n15236 );
not ( n15238 , n1817 );
nor ( n15239 , n15238 , n53 );
nand ( n15240 , n3 , n15239 );
not ( n15241 , n15240 );
not ( n15242 , n3 );
nand ( n15243 , n53 , n1817 );
nor ( n15244 , n15242 , n15243 );
nor ( n15245 , n15241 , n15244 );
not ( n15246 , n831 );
not ( n15247 , n845 );
not ( n15248 , n1530 );
nor ( n15249 , n763 , n806 );
nand ( n15250 , n15248 , n15249 );
not ( n15251 , n15250 );
and ( n15252 , n15247 , n15251 );
nand ( n15253 , n15246 , n748 , n15252 );
nor ( n15254 , n15245 , n15253 );
not ( n15255 , n15254 );
nor ( n15256 , n748 , n831 );
nand ( n15257 , n845 , n15256 , n15251 );
not ( n15258 , n15257 );
nand ( n15259 , n15258 , n15234 );
not ( n15260 , n748 );
nand ( n15261 , n831 , n15260 , n15252 );
not ( n15262 , n15261 );
nand ( n15263 , n15262 , n15234 );
nand ( n15264 , n15255 , n15259 , n15263 );
not ( n15265 , n15264 );
not ( n15266 , n15265 );
or ( n15267 , n15237 , n15266 );
nand ( n15268 , n15267 , n15231 );
buf ( n15269 , n15268 );
nand ( n15270 , n15232 , n1798 , n15269 );
nor ( n15271 , n831 , n845 );
not ( n15272 , n15271 );
nor ( n15273 , n15272 , n15250 );
not ( n15274 , n15273 );
nand ( n15275 , n831 , n15236 );
and ( n15276 , n15274 , n15275 );
and ( n15277 , n15246 , n15244 );
nor ( n15278 , n15277 , n15274 );
nor ( n15279 , n15276 , n15265 , n15278 );
not ( n15280 , n15236 );
not ( n15281 , n15265 );
or ( n15282 , n15280 , n15281 );
nand ( n15283 , n15282 , n15231 );
buf ( n15284 , n15283 );
not ( n15285 , n15284 );
nand ( n15286 , n15279 , n15285 );
nand ( n15287 , n15270 , n15286 );
not ( n15288 , n150 );
not ( n15289 , n14789 );
or ( n15290 , n15288 , n15289 );
not ( n15291 , n14820 );
not ( n15292 , n14842 );
and ( n15293 , n14808 , n15292 );
not ( n15294 , n14808 );
and ( n15295 , n182 , n14809 );
and ( n15296 , n138 , n14810 );
nor ( n15297 , n15295 , n15296 );
and ( n15298 , n15294 , n15297 );
nor ( n15299 , n15293 , n15298 );
not ( n15300 , n15299 );
or ( n15301 , n15291 , n15300 );
nor ( n15302 , n14904 , n14787 );
nand ( n15303 , n15301 , n15302 );
nand ( n15304 , n15290 , n15303 );
not ( n15305 , n196 );
nor ( n15306 , n15305 , n217 );
not ( n15307 , n237 );
not ( n15308 , n238 );
not ( n15309 , n218 );
not ( n15310 , n221 );
and ( n15311 , n15309 , n15310 );
nand ( n15312 , n15307 , n15308 , n15311 );
nor ( n15313 , n15312 , n13534 );
and ( n15314 , n15306 , n15313 );
nand ( n15315 , n13552 , n15314 );
not ( n15316 , n15315 );
and ( n15317 , n196 , n15316 );
not ( n15318 , n1362 );
not ( n15319 , n1356 );
and ( n15320 , n1357 , n15319 );
nand ( n15321 , n15320 , n13559 );
nor ( n15322 , n15318 , n15321 );
or ( n15323 , n15305 , n15322 );
not ( n15324 , n1546 );
nand ( n15325 , n15323 , n15324 );
not ( n15326 , n217 );
and ( n15327 , n15305 , n15326 );
and ( n15328 , n15308 , n237 , n15327 );
not ( n15329 , n15328 );
not ( n15330 , n13534 );
nand ( n15331 , n15311 , n15330 );
nor ( n15332 , n15329 , n15331 );
and ( n15333 , n15325 , n15332 );
nor ( n15334 , n15317 , n15333 );
nand ( n15335 , n15307 , n15327 );
nor ( n15336 , n238 , n15335 );
and ( n15337 , n15336 , n15330 );
and ( n15338 , n15310 , n218 , n15337 );
not ( n15339 , n196 );
not ( n15340 , n1756 );
and ( n15341 , n1755 , n15340 );
not ( n15342 , n825 );
nor ( n15343 , n511 , n824 );
nand ( n15344 , n15342 , n776 , n15343 );
or ( n15345 , n15341 , n15344 );
not ( n15346 , n15345 );
not ( n15347 , n15346 );
not ( n15348 , n15347 );
not ( n15349 , n15348 );
not ( n15350 , n15349 );
or ( n15351 , n15339 , n15350 );
nand ( n15352 , n858 , n862 , n856 , n875 );
nor ( n15353 , n860 , n866 );
nor ( n15354 , n859 , n867 );
nand ( n15355 , n15353 , n15354 );
nor ( n15356 , n15352 , n15355 );
nor ( n15357 , n852 , n861 );
nor ( n15358 , n864 , n873 );
nand ( n15359 , n15357 , n15358 );
nor ( n15360 , n851 , n865 );
nor ( n15361 , n863 , n874 );
nand ( n15362 , n15360 , n15361 );
nor ( n15363 , n15359 , n15362 );
and ( n15364 , n15356 , n15363 );
nor ( n15365 , n15345 , n15364 );
nor ( n15366 , n1545 , n267 , n15365 );
nand ( n15367 , n15351 , n15366 );
and ( n15368 , n15338 , n15367 );
not ( n15369 , n240 );
nand ( n15370 , n13532 , n15327 );
nor ( n15371 , n239 , n15370 , n15312 );
and ( n15372 , n241 , n15369 , n15371 );
nor ( n15373 , n15308 , n15335 , n15331 );
and ( n15374 , n267 , n15373 );
nor ( n15375 , n15372 , n15374 );
not ( n15376 , n754 );
not ( n15377 , n267 );
nor ( n15378 , n854 , n872 );
nand ( n15379 , n15376 , n15377 , n15378 );
not ( n15380 , n15312 );
nand ( n15381 , n15380 , n13533 );
nor ( n15382 , n13531 , n15370 , n15381 );
and ( n15383 , n15379 , n15382 );
not ( n15384 , n15313 );
nor ( n15385 , n196 , n15384 );
and ( n15386 , n217 , n15385 );
nor ( n15387 , n15383 , n15386 );
nand ( n15388 , n15375 , n15387 );
nor ( n15389 , n15368 , n15388 );
not ( n15390 , n13557 );
not ( n15391 , n15390 );
nand ( n15392 , n1358 , n1365 );
not ( n15393 , n15392 );
nand ( n15394 , n15393 , n13520 );
and ( n15395 , n15394 , n13560 );
not ( n15396 , n15395 );
and ( n15397 , n15391 , n15396 );
not ( n15398 , n12493 );
nor ( n15399 , n15397 , n15398 );
nand ( n15400 , n13528 , n15399 );
not ( n15401 , n13576 );
nor ( n15402 , n15400 , n15401 );
nand ( n15403 , n13546 , n15314 , n196 , n15402 );
not ( n15404 , n15321 );
not ( n15405 , n1168 );
and ( n15406 , n1223 , n15405 );
not ( n15407 , n1223 );
and ( n15408 , n15407 , n1168 );
nor ( n15409 , n15406 , n15408 );
not ( n15410 , n1169 );
and ( n15411 , n1224 , n15410 );
not ( n15412 , n1224 );
and ( n15413 , n15412 , n1169 );
nor ( n15414 , n15411 , n15413 );
not ( n15415 , n1170 );
and ( n15416 , n1198 , n15415 );
not ( n15417 , n1198 );
and ( n15418 , n15417 , n1170 );
nor ( n15419 , n15416 , n15418 );
not ( n15420 , n1178 );
and ( n15421 , n1225 , n15420 );
not ( n15422 , n1225 );
and ( n15423 , n15422 , n1178 );
nor ( n15424 , n15421 , n15423 );
nand ( n15425 , n15409 , n15414 , n15419 , n15424 );
or ( n15426 , n1608 , n13544 );
nand ( n15427 , n15426 , n1363 );
nor ( n15428 , n15404 , n15425 , n15427 , n15318 );
and ( n15429 , n15393 , n13543 );
and ( n15430 , n15320 , n13542 );
nor ( n15431 , n15429 , n15430 );
not ( n15432 , n1171 );
and ( n15433 , n1226 , n15432 );
not ( n15434 , n1226 );
and ( n15435 , n15434 , n1171 );
nor ( n15436 , n15433 , n15435 );
not ( n15437 , n1146 );
and ( n15438 , n1227 , n15437 );
not ( n15439 , n1227 );
and ( n15440 , n15439 , n1146 );
nor ( n15441 , n15438 , n15440 );
nand ( n15442 , n15431 , n15436 , n15441 );
and ( n15443 , n13522 , n13543 );
and ( n15444 , n1197 , n1172 );
not ( n15445 , n1197 );
not ( n15446 , n1172 );
and ( n15447 , n15445 , n15446 );
nor ( n15448 , n15444 , n15447 );
nor ( n15449 , n15443 , n15448 );
not ( n15450 , n15392 );
not ( n15451 , n13522 );
not ( n15452 , n15451 );
or ( n15453 , n15450 , n15452 );
nand ( n15454 , n15453 , n15320 );
not ( n15455 , n1173 );
not ( n15456 , n1466 );
or ( n15457 , n15455 , n15456 );
or ( n15458 , n1173 , n1466 );
nand ( n15459 , n15457 , n15458 );
not ( n15460 , n15459 );
xor ( n15461 , n1168 , n1169 );
not ( n15462 , n15461 );
or ( n15463 , n15460 , n15462 );
or ( n15464 , n15461 , n15459 );
nand ( n15465 , n15463 , n15464 );
xnor ( n15466 , n1171 , n1172 );
not ( n15467 , n1447 );
and ( n15468 , n15466 , n15467 );
not ( n15469 , n15466 );
and ( n15470 , n15469 , n1447 );
nor ( n15471 , n15468 , n15470 );
xor ( n15472 , n15465 , n15471 );
and ( n15473 , n1173 , n1465 );
not ( n15474 , n1173 );
not ( n15475 , n1465 );
and ( n15476 , n15474 , n15475 );
or ( n15477 , n15473 , n15476 );
xor ( n15478 , n15477 , n15461 );
not ( n15479 , n1442 );
not ( n15480 , n1170 );
not ( n15481 , n1178 );
and ( n15482 , n15480 , n15481 );
and ( n15483 , n1170 , n1178 );
nor ( n15484 , n15482 , n15483 );
not ( n15485 , n15484 );
or ( n15486 , n15479 , n15485 );
or ( n15487 , n1442 , n15484 );
nand ( n15488 , n15486 , n15487 );
and ( n15489 , n1171 , n1447 );
not ( n15490 , n1171 );
and ( n15491 , n15490 , n15467 );
nor ( n15492 , n15489 , n15491 );
not ( n15493 , n15492 );
and ( n15494 , n15488 , n15493 );
not ( n15495 , n15488 );
and ( n15496 , n15495 , n15492 );
nor ( n15497 , n15494 , n15496 );
not ( n15498 , n15497 );
and ( n15499 , n15478 , n15498 );
not ( n15500 , n15478 );
and ( n15501 , n15500 , n15497 );
nor ( n15502 , n15499 , n15501 );
nor ( n15503 , n15472 , n15502 );
not ( n15504 , n15503 );
xor ( n15505 , n1146 , n1446 );
not ( n15506 , n15505 );
not ( n15507 , n15461 );
or ( n15508 , n15506 , n15507 );
or ( n15509 , n15461 , n15505 );
nand ( n15510 , n15508 , n15509 );
xor ( n15511 , n1173 , n1464 );
not ( n15512 , n15511 );
not ( n15513 , n15484 );
or ( n15514 , n15512 , n15513 );
or ( n15515 , n15484 , n15511 );
nand ( n15516 , n15514 , n15515 );
xnor ( n15517 , n15510 , n15516 );
and ( n15518 , n1463 , n1178 );
not ( n15519 , n1463 );
and ( n15520 , n15519 , n15420 );
nor ( n15521 , n15518 , n15520 );
not ( n15522 , n1442 );
and ( n15523 , n15521 , n15522 );
not ( n15524 , n15521 );
and ( n15525 , n15524 , n1442 );
nor ( n15526 , n15523 , n15525 );
not ( n15527 , n15526 );
not ( n15528 , n15461 );
xor ( n15529 , n1146 , n1172 );
not ( n15530 , n15529 );
and ( n15531 , n15528 , n15530 );
and ( n15532 , n15529 , n15461 );
nor ( n15533 , n15531 , n15532 );
not ( n15534 , n15533 );
or ( n15535 , n15527 , n15534 );
not ( n15536 , n15526 );
not ( n15537 , n15533 );
and ( n15538 , n15536 , n15537 );
not ( n15539 , n15505 );
not ( n15540 , n15539 );
xor ( n15541 , n1171 , n1414 );
and ( n15542 , n1170 , n1168 );
not ( n15543 , n1170 );
and ( n15544 , n15543 , n15405 );
nor ( n15545 , n15542 , n15544 );
xor ( n15546 , n15541 , n15545 );
not ( n15547 , n15546 );
or ( n15548 , n15540 , n15547 );
or ( n15549 , n15539 , n15546 );
nand ( n15550 , n15548 , n15549 );
nor ( n15551 , n15538 , n15550 );
nand ( n15552 , n15535 , n15551 );
nor ( n15553 , n15517 , n15552 );
not ( n15554 , n15553 );
or ( n15555 , n15504 , n15554 );
nand ( n15556 , n15555 , n1362 );
nand ( n15557 , n15449 , n15454 , n15556 );
nor ( n15558 , n15442 , n15557 );
nand ( n15559 , n15428 , n15558 );
nand ( n15560 , n2 , n15559 );
not ( n15561 , n15560 );
nand ( n15562 , n15334 , n15389 , n15403 , n15561 );
not ( n15563 , n481 );
not ( n15564 , n854 );
or ( n15565 , n15563 , n15564 );
nand ( n15566 , n15306 , n13530 , n15308 , n13535 );
not ( n15567 , n15559 );
and ( n15568 , n15566 , n15567 );
nor ( n15569 , n15568 , n373 );
nand ( n15570 , n15565 , n15569 );
nand ( n15571 , n13310 , n13390 );
not ( n15572 , n15571 );
not ( n15573 , n13385 );
or ( n15574 , n15572 , n15573 );
or ( n15575 , n15571 , n13385 );
nand ( n15576 , n15574 , n15575 );
not ( n15577 , n431 );
nand ( n15578 , n429 , n430 );
nand ( n15579 , n15577 , n15578 );
nor ( n15580 , n1113 , n1174 );
nor ( n15581 , n1100 , n1124 );
nor ( n15582 , n1095 , n1148 );
nand ( n15583 , n15581 , n15582 );
not ( n15584 , n15583 );
not ( n15585 , n1806 );
nor ( n15586 , n1045 , n1175 );
nand ( n15587 , n15585 , n15586 );
nor ( n15588 , n902 , n1066 );
nor ( n15589 , n889 , n1150 );
nand ( n15590 , n15588 , n15589 );
nor ( n15591 , n15587 , n15590 );
nand ( n15592 , n15580 , n15584 , n15591 );
not ( n15593 , n15592 );
not ( n15594 , n1179 );
nand ( n15595 , n15593 , n15594 , n1083 );
not ( n15596 , n15595 );
not ( n15597 , n15596 );
not ( n15598 , n1124 );
and ( n15599 , n15598 , n15582 );
not ( n15600 , n15599 );
nor ( n15601 , n1083 , n1179 );
nand ( n15602 , n15580 , n15601 );
not ( n15603 , n15602 );
nand ( n15604 , n15603 , n15591 );
nor ( n15605 , n15600 , n15604 );
nand ( n15606 , n1100 , n15605 );
nor ( n15607 , n15583 , n15590 );
nand ( n15608 , n15603 , n15607 );
not ( n15609 , n15608 );
not ( n15610 , n1175 );
nor ( n15611 , n15610 , n1045 );
nand ( n15612 , n15609 , n15585 , n15611 );
nand ( n15613 , n15597 , n15606 , n15612 );
not ( n15614 , n15613 );
not ( n15615 , n15614 );
nand ( n15616 , n914 , n1608 );
nand ( n15617 , n914 , n13539 );
not ( n15618 , n15617 );
nor ( n15619 , n15616 , n15618 );
not ( n15620 , n15619 );
nor ( n15621 , n1474 , n1608 );
nand ( n15622 , n15621 , n853 , n1089 );
nand ( n15623 , n15620 , n15622 );
and ( n15624 , n1045 , n15610 );
not ( n15625 , n15624 );
nor ( n15626 , n15625 , n15608 );
nand ( n15627 , n15585 , n15626 );
not ( n15628 , n15604 );
not ( n15629 , n1148 );
nor ( n15630 , n15629 , n1095 );
not ( n15631 , n1100 );
and ( n15632 , n15631 , n15598 );
nand ( n15633 , n15628 , n15630 , n15632 );
not ( n15634 , n15604 );
nand ( n15635 , n1100 , n15599 , n15634 );
nand ( n15636 , n15627 , n15633 , n15635 );
not ( n15637 , n15604 );
and ( n15638 , n1095 , n15629 );
nand ( n15639 , n15637 , n15638 , n15632 );
and ( n15640 , n15595 , n15633 , n15639 );
and ( n15641 , n15636 , n15640 );
and ( n15642 , n15623 , n15641 );
not ( n15643 , n15640 );
and ( n15644 , n391 , n15643 , n15636 );
nor ( n15645 , n15642 , n15644 );
or ( n15646 , n15615 , n15645 );
nor ( n15647 , n1866 , n1868 );
nand ( n15648 , n1758 , n15647 );
not ( n15649 , n15648 );
nand ( n15650 , n853 , n15649 );
not ( n15651 , n15650 );
not ( n15652 , n15636 );
not ( n15653 , n15652 );
nand ( n15654 , n15651 , n15640 , n15615 , n15653 );
nand ( n15655 , n15646 , n15654 );
not ( n15656 , n15655 );
not ( n15657 , n406 );
not ( n15658 , n15636 );
and ( n15659 , n15613 , n15658 );
not ( n15660 , n15659 );
or ( n15661 , n15657 , n15660 );
not ( n15662 , n15613 );
nand ( n15663 , n15647 , n15662 , n15652 );
nand ( n15664 , n15661 , n15663 );
and ( n15665 , n15643 , n15664 );
not ( n15666 , n15648 );
and ( n15667 , n405 , n15666 );
not ( n15668 , n15667 );
nor ( n15669 , n15668 , n15643 );
and ( n15670 , n15669 , n15615 , n15652 );
nor ( n15671 , n15665 , n15670 );
nand ( n15672 , n15643 , n15652 );
not ( n15673 , n15641 );
nand ( n15674 , n1806 , n15586 );
nor ( n15675 , n15674 , n15608 );
not ( n15676 , n15612 );
nor ( n15677 , n15675 , n15676 );
not ( n15678 , n15596 );
nand ( n15679 , n15677 , n15639 , n15678 , n15658 );
not ( n15680 , n15614 );
not ( n15681 , n15680 );
not ( n15682 , n15636 );
or ( n15683 , n15681 , n15682 );
nand ( n15684 , n15662 , n15658 );
nand ( n15685 , n15683 , n15684 );
nand ( n15686 , n15672 , n15673 , n15679 , n15685 );
nand ( n15687 , n15656 , n15671 , n15686 );
not ( n15688 , n15687 );
nand ( n15689 , n432 , n15579 , n15688 );
not ( n15690 , n413 );
not ( n15691 , n435 );
nand ( n15692 , n15690 , n15691 );
or ( n15693 , n434 , n433 , n15692 );
nand ( n15694 , n15693 , n15688 );
nand ( n15695 , n15689 , n15694 );
not ( n15696 , n14460 );
nor ( n15697 , n15696 , n14450 );
and ( n15698 , n15697 , n14518 );
not ( n15699 , n15697 );
not ( n15700 , n14518 );
and ( n15701 , n15699 , n15700 );
nor ( n15702 , n15698 , n15701 );
not ( n15703 , n1260 );
not ( n15704 , n1808 );
not ( n15705 , n597 );
nand ( n15706 , n1576 , n1701 );
nand ( n15707 , n1176 , n1576 );
nand ( n15708 , n1576 , n1655 );
nand ( n15709 , n15706 , n15707 , n15708 );
buf ( n15710 , n15709 );
not ( n15711 , n15710 );
not ( n15712 , n15711 );
not ( n15713 , n15712 );
not ( n15714 , n15713 );
or ( n15715 , n15705 , n15714 );
not ( n15716 , n597 );
not ( n15717 , n15716 );
not ( n15718 , n509 );
not ( n15719 , n662 );
nand ( n15720 , n1256 , n15719 );
not ( n15721 , n612 );
nor ( n15722 , n15721 , n1158 );
and ( n15723 , n15720 , n15722 );
nor ( n15724 , n15719 , n1256 );
nor ( n15725 , n15723 , n15724 );
and ( n15726 , n15718 , n15725 );
not ( n15727 , n691 );
nand ( n15728 , n1158 , n15721 );
and ( n15729 , n15728 , n15720 );
not ( n15730 , n1212 );
nand ( n15731 , n15730 , n696 );
not ( n15732 , n15731 );
not ( n15733 , n696 );
nand ( n15734 , n1212 , n15733 );
or ( n15735 , n15732 , n15734 );
not ( n15736 , n1157 );
nand ( n15737 , n751 , n15736 );
nand ( n15738 , n15737 , n15731 );
not ( n15739 , n614 );
nand ( n15740 , n1205 , n15739 );
not ( n15741 , n678 );
nand ( n15742 , n1259 , n15741 );
and ( n15743 , n15740 , n15742 );
nand ( n15744 , n15735 , n15738 , n15743 );
not ( n15745 , n751 );
nand ( n15746 , n15745 , n1157 );
nand ( n15747 , n15734 , n15746 );
not ( n15748 , n15747 );
and ( n15749 , n15743 , n15748 );
not ( n15750 , n716 );
nand ( n15751 , n1258 , n15750 );
not ( n15752 , n635 );
nand ( n15753 , n1156 , n15752 );
not ( n15754 , n747 );
nand ( n15755 , n1439 , n15754 );
nand ( n15756 , n15753 , n15755 );
not ( n15757 , n15756 );
nand ( n15758 , n15751 , n15757 );
not ( n15759 , n15751 );
nor ( n15760 , n15754 , n1439 );
not ( n15761 , n15760 );
or ( n15762 , n15759 , n15761 );
nor ( n15763 , n15750 , n1258 );
not ( n15764 , n15763 );
nand ( n15765 , n15762 , n15764 );
not ( n15766 , n15765 );
nand ( n15767 , n15758 , n15766 );
and ( n15768 , n15749 , n15767 );
not ( n15769 , n1205 );
nand ( n15770 , n15769 , n614 );
nor ( n15771 , n15741 , n1259 );
nand ( n15772 , n15740 , n15771 );
nand ( n15773 , n15770 , n15772 );
nor ( n15774 , n15768 , n15773 );
nand ( n15775 , n15744 , n15774 );
nand ( n15776 , n15729 , n15775 );
nand ( n15777 , n15726 , n15727 , n15776 );
not ( n15778 , n15777 );
or ( n15779 , n15717 , n15778 );
not ( n15780 , n15777 );
and ( n15781 , n597 , n15780 );
not ( n15782 , n15712 );
nor ( n15783 , n15781 , n15782 );
nand ( n15784 , n15779 , n15783 );
nand ( n15785 , n15715 , n15784 );
and ( n15786 , n15704 , n15785 );
not ( n15787 , n597 );
nand ( n15788 , n509 , n662 );
not ( n15789 , n15788 );
not ( n15790 , n15789 );
not ( n15791 , n15790 );
nand ( n15792 , n678 , n696 );
nand ( n15793 , n635 , n747 );
nor ( n15794 , n15750 , n15793 );
nand ( n15795 , n751 , n15794 );
nor ( n15796 , n15792 , n15795 );
nand ( n15797 , n614 , n15796 );
not ( n15798 , n15797 );
and ( n15799 , n612 , n15798 );
nand ( n15800 , n691 , n15791 , n15799 );
not ( n15801 , n15800 );
or ( n15802 , n15787 , n15801 );
or ( n15803 , n597 , n15800 );
nand ( n15804 , n15802 , n15803 );
and ( n15805 , n1808 , n15804 );
nor ( n15806 , n15786 , n15805 );
nor ( n15807 , n15703 , n15806 );
not ( n15808 , n750 );
not ( n15809 , n15100 );
or ( n15810 , n15808 , n15809 );
not ( n15811 , n750 );
not ( n15812 , n15811 );
and ( n15813 , n15103 , n15178 );
not ( n15814 , n774 );
not ( n15815 , n15157 );
nand ( n15816 , n15115 , n15815 );
and ( n15817 , n15115 , n15121 );
not ( n15818 , n15149 );
nand ( n15819 , n15818 , n15130 );
nand ( n15820 , n15817 , n15819 );
nand ( n15821 , n15816 , n15170 , n15820 );
nand ( n15822 , n15109 , n15821 );
nand ( n15823 , n15813 , n15814 , n15822 );
not ( n15824 , n15823 );
or ( n15825 , n15812 , n15824 );
not ( n15826 , n15823 );
and ( n15827 , n750 , n15826 );
buf ( n15828 , n15095 );
not ( n15829 , n15828 );
not ( n15830 , n15829 );
not ( n15831 , n15830 );
nor ( n15832 , n15827 , n15831 );
nand ( n15833 , n15825 , n15832 );
nand ( n15834 , n15810 , n15833 );
and ( n15835 , n15090 , n15834 );
not ( n15836 , n750 );
nand ( n15837 , n487 , n752 );
not ( n15838 , n15837 );
nand ( n15839 , n777 , n779 );
nor ( n15840 , n15122 , n15193 );
nand ( n15841 , n783 , n15840 );
nor ( n15842 , n15839 , n15841 );
nand ( n15843 , n698 , n15842 );
not ( n15844 , n15843 );
and ( n15845 , n695 , n15844 );
nand ( n15846 , n774 , n15838 , n15845 );
not ( n15847 , n15846 );
or ( n15848 , n15836 , n15847 );
or ( n15849 , n750 , n15846 );
nand ( n15850 , n15848 , n15849 );
and ( n15851 , n1826 , n15850 );
nor ( n15852 , n15835 , n15851 );
nor ( n15853 , n15089 , n15852 );
not ( n15854 , n510 );
not ( n15855 , n14983 );
or ( n15856 , n15854 , n15855 );
not ( n15857 , n510 );
not ( n15858 , n15857 );
and ( n15859 , n14986 , n15062 );
not ( n15860 , n599 );
not ( n15861 , n15041 );
nand ( n15862 , n14998 , n15861 );
and ( n15863 , n14998 , n15004 );
not ( n15864 , n15033 );
nand ( n15865 , n15864 , n15014 );
nand ( n15866 , n15863 , n15865 );
nand ( n15867 , n15862 , n15054 , n15866 );
nand ( n15868 , n14992 , n15867 );
nand ( n15869 , n15859 , n15860 , n15868 );
not ( n15870 , n15869 );
or ( n15871 , n15858 , n15870 );
not ( n15872 , n15869 );
and ( n15873 , n510 , n15872 );
not ( n15874 , n14979 );
buf ( n15875 , n15874 );
not ( n15876 , n15875 );
nor ( n15877 , n15873 , n15876 );
nand ( n15878 , n15871 , n15877 );
nand ( n15879 , n15856 , n15878 );
and ( n15880 , n14974 , n15879 );
not ( n15881 , n510 );
nand ( n15882 , n508 , n595 );
not ( n15883 , n15882 );
not ( n15884 , n15883 );
not ( n15885 , n15884 );
nand ( n15886 , n609 , n613 );
nor ( n15887 , n15005 , n15075 );
nand ( n15888 , n638 , n15887 );
nor ( n15889 , n15886 , n15888 );
nand ( n15890 , n516 , n15889 );
not ( n15891 , n15890 );
and ( n15892 , n515 , n15891 );
nand ( n15893 , n599 , n15885 , n15892 );
not ( n15894 , n15893 );
or ( n15895 , n15881 , n15894 );
or ( n15896 , n510 , n15893 );
nand ( n15897 , n15895 , n15896 );
and ( n15898 , n1819 , n15897 );
nor ( n15899 , n15880 , n15898 );
nor ( n15900 , n14973 , n15899 );
not ( n15901 , n46 );
or ( n15902 , n15901 , n15284 );
nand ( n15903 , n308 , n15269 );
nand ( n15904 , n15902 , n15903 );
not ( n15905 , n5 );
or ( n15906 , n15905 , n15284 );
nand ( n15907 , n161 , n15269 );
nand ( n15908 , n15906 , n15907 );
not ( n15909 , n6 );
or ( n15910 , n15909 , n15284 );
buf ( n15911 , n15268 );
nand ( n15912 , n172 , n15911 );
nand ( n15913 , n15910 , n15912 );
not ( n15914 , n7 );
or ( n15915 , n15914 , n15284 );
nand ( n15916 , n160 , n15911 );
nand ( n15917 , n15915 , n15916 );
not ( n15918 , n8 );
or ( n15919 , n15918 , n15284 );
buf ( n15920 , n15268 );
nand ( n15921 , n171 , n15920 );
nand ( n15922 , n15919 , n15921 );
not ( n15923 , n9 );
or ( n15924 , n15923 , n15284 );
nand ( n15925 , n174 , n15269 );
nand ( n15926 , n15924 , n15925 );
not ( n15927 , n10 );
or ( n15928 , n15927 , n15284 );
nand ( n15929 , n166 , n15920 );
nand ( n15930 , n15928 , n15929 );
not ( n15931 , n11 );
or ( n15932 , n15931 , n15284 );
nand ( n15933 , n165 , n15269 );
nand ( n15934 , n15932 , n15933 );
not ( n15935 , n12 );
or ( n15936 , n15935 , n15284 );
nand ( n15937 , n164 , n15269 );
nand ( n15938 , n15936 , n15937 );
not ( n15939 , n13 );
or ( n15940 , n15939 , n15284 );
nand ( n15941 , n163 , n15911 );
nand ( n15942 , n15940 , n15941 );
not ( n15943 , n14 );
or ( n15944 , n15943 , n15284 );
nand ( n15945 , n170 , n15911 );
nand ( n15946 , n15944 , n15945 );
not ( n15947 , n15 );
or ( n15948 , n15947 , n15284 );
nand ( n15949 , n168 , n15911 );
nand ( n15950 , n15948 , n15949 );
not ( n15951 , n16 );
not ( n15952 , n15951 );
not ( n15953 , n15952 );
or ( n15954 , n15953 , n15284 );
nand ( n15955 , n169 , n15920 );
nand ( n15956 , n15954 , n15955 );
not ( n15957 , n17 );
or ( n15958 , n15957 , n15284 );
nand ( n15959 , n173 , n15920 );
nand ( n15960 , n15958 , n15959 );
not ( n15961 , n18 );
or ( n15962 , n15961 , n15284 );
nand ( n15963 , n167 , n15911 );
nand ( n15964 , n15962 , n15963 );
not ( n15965 , n21 );
or ( n15966 , n15965 , n15284 );
nand ( n15967 , n305 , n15269 );
nand ( n15968 , n15966 , n15967 );
not ( n15969 , n22 );
or ( n15970 , n15969 , n15284 );
nand ( n15971 , n270 , n15920 );
nand ( n15972 , n15970 , n15971 );
not ( n15973 , n23 );
or ( n15974 , n15973 , n15284 );
nand ( n15975 , n303 , n15920 );
nand ( n15976 , n15974 , n15975 );
not ( n15977 , n25 );
or ( n15978 , n15977 , n15284 );
nand ( n15979 , n274 , n15269 );
nand ( n15980 , n15978 , n15979 );
not ( n15981 , n26 );
or ( n15982 , n15981 , n15284 );
nand ( n15983 , n301 , n15911 );
nand ( n15984 , n15982 , n15983 );
not ( n15985 , n27 );
or ( n15986 , n15985 , n15284 );
nand ( n15987 , n300 , n15920 );
nand ( n15988 , n15986 , n15987 );
not ( n15989 , n28 );
or ( n15990 , n15989 , n15284 );
nand ( n15991 , n299 , n15920 );
nand ( n15992 , n15990 , n15991 );
not ( n15993 , n29 );
or ( n15994 , n15993 , n15284 );
nand ( n15995 , n298 , n15920 );
nand ( n15996 , n15994 , n15995 );
not ( n15997 , n30 );
or ( n15998 , n15997 , n15284 );
nand ( n15999 , n297 , n15269 );
nand ( n16000 , n15998 , n15999 );
not ( n16001 , n31 );
or ( n16002 , n16001 , n15284 );
nand ( n16003 , n296 , n15920 );
nand ( n16004 , n16002 , n16003 );
not ( n16005 , n32 );
or ( n16006 , n16005 , n15284 );
nand ( n16007 , n295 , n15911 );
nand ( n16008 , n16006 , n16007 );
not ( n16009 , n33 );
or ( n16010 , n16009 , n15284 );
nand ( n16011 , n294 , n15911 );
nand ( n16012 , n16010 , n16011 );
not ( n16013 , n34 );
or ( n16014 , n16013 , n15284 );
nand ( n16015 , n293 , n15911 );
nand ( n16016 , n16014 , n16015 );
not ( n16017 , n35 );
or ( n16018 , n16017 , n15284 );
nand ( n16019 , n292 , n15911 );
nand ( n16020 , n16018 , n16019 );
not ( n16021 , n36 );
or ( n16022 , n16021 , n15284 );
nand ( n16023 , n276 , n15911 );
nand ( n16024 , n16022 , n16023 );
not ( n16025 , n37 );
or ( n16026 , n16025 , n15284 );
nand ( n16027 , n291 , n15911 );
nand ( n16028 , n16026 , n16027 );
not ( n16029 , n38 );
or ( n16030 , n16029 , n15284 );
nand ( n16031 , n290 , n15269 );
nand ( n16032 , n16030 , n16031 );
not ( n16033 , n39 );
or ( n16034 , n16033 , n15284 );
nand ( n16035 , n289 , n15911 );
nand ( n16036 , n16034 , n16035 );
not ( n16037 , n4 );
or ( n16038 , n16037 , n15284 );
nand ( n16039 , n162 , n15269 );
nand ( n16040 , n16038 , n16039 );
not ( n16041 , n41 );
or ( n16042 , n16041 , n15284 );
nand ( n16043 , n288 , n15920 );
nand ( n16044 , n16042 , n16043 );
not ( n16045 , n42 );
or ( n16046 , n16045 , n15284 );
nand ( n16047 , n286 , n15920 );
nand ( n16048 , n16046 , n16047 );
not ( n16049 , n43 );
or ( n16050 , n16049 , n15284 );
nand ( n16051 , n311 , n15920 );
nand ( n16052 , n16050 , n16051 );
not ( n16053 , n44 );
or ( n16054 , n16053 , n15284 );
nand ( n16055 , n310 , n15920 );
nand ( n16056 , n16054 , n16055 );
not ( n16057 , n45 );
or ( n16058 , n16057 , n15284 );
nand ( n16059 , n309 , n15269 );
nand ( n16060 , n16058 , n16059 );
not ( n16061 , n47 );
or ( n16062 , n16061 , n15284 );
nand ( n16063 , n273 , n15269 );
nand ( n16064 , n16062 , n16063 );
not ( n16065 , n24 );
or ( n16066 , n16065 , n15284 );
nand ( n16067 , n302 , n15920 );
nand ( n16068 , n16066 , n16067 );
not ( n16069 , n49 );
or ( n16070 , n16069 , n15284 );
nand ( n16071 , n306 , n15920 );
nand ( n16072 , n16070 , n16071 );
not ( n16073 , n50 );
or ( n16074 , n16073 , n15284 );
nand ( n16075 , n304 , n15911 );
nand ( n16076 , n16074 , n16075 );
not ( n16077 , n51 );
or ( n16078 , n16077 , n15284 );
nand ( n16079 , n275 , n15269 );
nand ( n16080 , n16078 , n16079 );
not ( n16081 , n40 );
or ( n16082 , n16081 , n15284 );
nand ( n16083 , n287 , n15269 );
nand ( n16084 , n16082 , n16083 );
not ( n16085 , n48 );
or ( n16086 , n16085 , n15284 );
nand ( n16087 , n307 , n15269 );
nand ( n16088 , n16086 , n16087 );
not ( n16089 , n52 );
or ( n16090 , n16089 , n15284 );
nand ( n16091 , n285 , n15911 );
nand ( n16092 , n16090 , n16091 );
not ( n16093 , n14904 );
xor ( n16094 , n133 , n134 );
not ( n16095 , n16094 );
or ( n16096 , n16093 , n16095 );
and ( n16097 , n14808 , n13104 , n13115 );
not ( n16098 , n1111 );
and ( n16099 , n16098 , n14817 );
not ( n16100 , n12850 );
and ( n16101 , n154 , n16100 );
and ( n16102 , n142 , n12849 );
nor ( n16103 , n16101 , n16102 , n14817 );
nor ( n16104 , n16099 , n14808 , n16103 );
nor ( n16105 , n16097 , n16104 );
or ( n16106 , n14904 , n16105 );
nand ( n16107 , n16096 , n16106 );
or ( n16108 , n14787 , n16107 );
not ( n16109 , n130 );
not ( n16110 , n14789 );
or ( n16111 , n16109 , n16110 );
nand ( n16112 , n16108 , n16111 );
not ( n16113 , n1380 );
and ( n16114 , n221 , n15309 , n15337 );
nand ( n16115 , n16113 , n16114 );
and ( n16116 , n221 , n15399 );
nor ( n16117 , n16116 , n13527 );
not ( n16118 , n13546 );
nor ( n16119 , n16117 , n16118 , n15401 );
or ( n16120 , n13552 , n16119 );
nand ( n16121 , n16120 , n15314 );
and ( n16122 , n16115 , n16121 );
and ( n16123 , n15314 , n16119 );
nor ( n16124 , n16123 , n221 );
nor ( n16125 , n16122 , n16124 , n15560 );
xnor ( n16126 , n408 , n423 );
not ( n16127 , n1750 );
not ( n16128 , n15687 );
nand ( n16129 , n16127 , n16128 );
nor ( n16130 , n16126 , n16129 );
not ( n16131 , n412 );
nor ( n16132 , n421 , n422 );
and ( n16133 , n16131 , n16132 );
not ( n16134 , n420 );
nor ( n16135 , n416 , n417 );
not ( n16136 , n16135 );
or ( n16137 , n418 , n16136 );
nand ( n16138 , n16137 , n419 );
nand ( n16139 , n16134 , n16132 , n16138 );
nand ( n16140 , n16139 , n15688 );
nor ( n16141 , n16133 , n16140 );
not ( n16142 , n418 );
nand ( n16143 , n416 , n417 );
nor ( n16144 , n16142 , n16143 );
nand ( n16145 , n419 , n16144 );
nor ( n16146 , n16134 , n16145 );
not ( n16147 , n16146 );
nand ( n16148 , n16147 , n16131 );
nand ( n16149 , n412 , n16146 );
and ( n16150 , n16148 , n1750 , n16149 );
and ( n16151 , n412 , n16127 );
nor ( n16152 , n16150 , n16151 );
not ( n16153 , n1663 );
nand ( n16154 , n16153 , n16128 );
nor ( n16155 , n16152 , n16154 );
and ( n16156 , n416 , n16127 );
not ( n16157 , n416 );
and ( n16158 , n16157 , n1750 );
nor ( n16159 , n16156 , n16158 );
nor ( n16160 , n16159 , n16154 );
and ( n16161 , n16143 , n1750 , n16136 );
and ( n16162 , n417 , n16127 );
nor ( n16163 , n16161 , n16162 );
nor ( n16164 , n16163 , n16154 );
and ( n16165 , n418 , n16127 );
and ( n16166 , n16142 , n16143 );
nor ( n16167 , n16166 , n16127 , n16144 );
nor ( n16168 , n16165 , n16167 );
nor ( n16169 , n16168 , n16154 );
or ( n16170 , n419 , n16144 );
and ( n16171 , n16170 , n1750 , n16145 );
and ( n16172 , n419 , n16127 );
nor ( n16173 , n16171 , n16172 );
nor ( n16174 , n16173 , n16154 );
and ( n16175 , n420 , n16127 );
and ( n16176 , n16134 , n16145 );
nor ( n16177 , n16176 , n16127 , n16146 );
nor ( n16178 , n16175 , n16177 );
nor ( n16179 , n16178 , n16154 );
and ( n16180 , n421 , n16127 );
not ( n16181 , n421 );
and ( n16182 , n16181 , n16149 );
nor ( n16183 , n16181 , n16149 );
nor ( n16184 , n16182 , n16127 , n16183 );
nor ( n16185 , n16180 , n16184 );
nor ( n16186 , n16185 , n16154 );
and ( n16187 , n422 , n16127 );
and ( n16188 , n422 , n16183 );
nor ( n16189 , n422 , n16183 );
nor ( n16190 , n16188 , n16189 , n16127 );
nor ( n16191 , n16187 , n16190 );
nor ( n16192 , n16191 , n16154 );
nor ( n16193 , n423 , n16129 );
not ( n16194 , n424 );
nand ( n16195 , n408 , n423 );
not ( n16196 , n16195 );
and ( n16197 , n16194 , n16196 );
and ( n16198 , n424 , n16195 );
nor ( n16199 , n16197 , n16198 );
nor ( n16200 , n16199 , n16129 );
not ( n16201 , n425 );
not ( n16202 , n16195 );
nand ( n16203 , n16202 , n424 );
not ( n16204 , n16203 );
nand ( n16205 , n436 , n16204 );
not ( n16206 , n16205 );
and ( n16207 , n16201 , n16206 );
and ( n16208 , n425 , n16205 );
nor ( n16209 , n16207 , n16208 );
nor ( n16210 , n16209 , n16129 );
not ( n16211 , n426 );
not ( n16212 , n16205 );
nand ( n16213 , n16212 , n425 );
not ( n16214 , n16213 );
and ( n16215 , n16211 , n16214 );
and ( n16216 , n426 , n16213 );
nor ( n16217 , n16215 , n16216 );
nor ( n16218 , n16217 , n16129 );
not ( n16219 , n427 );
not ( n16220 , n16213 );
nand ( n16221 , n16220 , n426 );
not ( n16222 , n16221 );
and ( n16223 , n16219 , n16222 );
and ( n16224 , n427 , n16221 );
nor ( n16225 , n16223 , n16224 );
nor ( n16226 , n16225 , n16129 );
not ( n16227 , n436 );
not ( n16228 , n16203 );
and ( n16229 , n16227 , n16228 );
and ( n16230 , n436 , n16203 );
nor ( n16231 , n16229 , n16230 );
nor ( n16232 , n16231 , n16129 );
not ( n16233 , n437 );
not ( n16234 , n16221 );
nand ( n16235 , n16234 , n427 );
not ( n16236 , n16235 );
and ( n16237 , n16233 , n16236 );
and ( n16238 , n437 , n16235 );
nor ( n16239 , n16237 , n16238 );
nor ( n16240 , n16239 , n16129 );
not ( n16241 , n14465 );
nor ( n16242 , n16241 , n14509 );
not ( n16243 , n16242 );
not ( n16244 , n14961 );
not ( n16245 , n16244 );
or ( n16246 , n16243 , n16245 );
or ( n16247 , n16242 , n16244 );
nand ( n16248 , n16246 , n16247 );
nand ( n16249 , n14506 , n14467 );
and ( n16250 , n14472 , n14747 );
nor ( n16251 , n16250 , n14754 );
and ( n16252 , n16249 , n16251 );
not ( n16253 , n16249 );
not ( n16254 , n16251 );
and ( n16255 , n16253 , n16254 );
nor ( n16256 , n16252 , n16255 );
not ( n16257 , n1240 );
not ( n16258 , n1828 );
not ( n16259 , n488 );
nand ( n16260 , n1609 , n1723 );
nand ( n16261 , n1176 , n1609 );
not ( n16262 , n16261 );
not ( n16263 , n16262 );
nand ( n16264 , n1609 , n1655 );
and ( n16265 , n16260 , n16263 , n16264 );
not ( n16266 , n16265 );
not ( n16267 , n16266 );
not ( n16268 , n16267 );
buf ( n16269 , n16268 );
not ( n16270 , n16269 );
not ( n16271 , n16270 );
or ( n16272 , n16259 , n16271 );
not ( n16273 , n1237 );
nor ( n16274 , n16273 , n846 );
not ( n16275 , n16274 );
not ( n16276 , n16275 );
not ( n16277 , n837 );
nand ( n16278 , n1236 , n16277 );
not ( n16279 , n16278 );
nor ( n16280 , n16276 , n16279 );
not ( n16281 , n848 );
nand ( n16282 , n1235 , n16281 );
not ( n16283 , n826 );
nand ( n16284 , n1234 , n16283 );
not ( n16285 , n847 );
nand ( n16286 , n1467 , n16285 );
nand ( n16287 , n16284 , n16286 );
not ( n16288 , n16287 );
nand ( n16289 , n16282 , n16288 );
not ( n16290 , n16289 );
and ( n16291 , n16280 , n16290 );
not ( n16292 , n804 );
nand ( n16293 , n1239 , n16292 );
not ( n16294 , n841 );
nand ( n16295 , n1231 , n16294 );
and ( n16296 , n16293 , n16295 );
not ( n16297 , n843 );
nand ( n16298 , n1210 , n16297 );
not ( n16299 , n16298 );
not ( n16300 , n1238 );
nor ( n16301 , n16300 , n807 );
nor ( n16302 , n16299 , n16301 );
and ( n16303 , n16291 , n16296 , n16302 );
not ( n16304 , n16296 );
not ( n16305 , n16302 );
not ( n16306 , n1236 );
nand ( n16307 , n16306 , n837 );
nand ( n16308 , n846 , n16273 );
nand ( n16309 , n16307 , n16308 );
nand ( n16310 , n16308 , n16274 );
nand ( n16311 , n16309 , n16310 );
not ( n16312 , n16309 );
not ( n16313 , n16312 );
nor ( n16314 , n16285 , n1467 );
and ( n16315 , n16282 , n16314 );
nor ( n16316 , n16281 , n1235 );
nor ( n16317 , n16315 , n16316 );
not ( n16318 , n16317 );
or ( n16319 , n16313 , n16318 );
nand ( n16320 , n16319 , n16280 );
and ( n16321 , n16311 , n16320 );
not ( n16322 , n16310 );
and ( n16323 , n16322 , n16317 );
nor ( n16324 , n16321 , n16323 );
not ( n16325 , n16324 );
or ( n16326 , n16305 , n16325 );
not ( n16327 , n16301 );
not ( n16328 , n1210 );
nand ( n16329 , n16328 , n843 );
not ( n16330 , n16329 );
and ( n16331 , n16327 , n16330 );
not ( n16332 , n807 );
nor ( n16333 , n16332 , n1238 );
nor ( n16334 , n16331 , n16333 );
nand ( n16335 , n16326 , n16334 );
not ( n16336 , n16335 );
or ( n16337 , n16304 , n16336 );
not ( n16338 , n1239 );
and ( n16339 , n804 , n16338 );
and ( n16340 , n16295 , n16339 );
nor ( n16341 , n16294 , n1231 );
nor ( n16342 , n16340 , n16341 );
nand ( n16343 , n16337 , n16342 );
nor ( n16344 , n16303 , n16343 );
or ( n16345 , n488 , n16344 );
and ( n16346 , n488 , n16344 );
buf ( n16347 , n16265 );
not ( n16348 , n16347 );
not ( n16349 , n16348 );
nor ( n16350 , n16346 , n16349 );
nand ( n16351 , n16345 , n16350 );
nand ( n16352 , n16272 , n16351 );
and ( n16353 , n16258 , n16352 );
not ( n16354 , n488 );
nand ( n16355 , n804 , n807 );
not ( n16356 , n16355 );
not ( n16357 , n846 );
nand ( n16358 , n826 , n847 );
nand ( n16359 , n837 , n848 );
not ( n16360 , n16359 );
not ( n16361 , n16360 );
nor ( n16362 , n16357 , n16358 , n16361 );
nand ( n16363 , n841 , n843 , n16356 , n16362 );
not ( n16364 , n16363 );
or ( n16365 , n16354 , n16364 );
or ( n16366 , n488 , n16363 );
nand ( n16367 , n16365 , n16366 );
and ( n16368 , n1828 , n16367 );
nor ( n16369 , n16353 , n16368 );
nor ( n16370 , n16257 , n16369 );
not ( n16371 , n509 );
not ( n16372 , n15713 );
or ( n16373 , n16371 , n16372 );
nor ( n16374 , n15747 , n15758 );
and ( n16375 , n16374 , n15729 , n15743 );
not ( n16376 , n15729 );
not ( n16377 , n15743 );
not ( n16378 , n15748 );
not ( n16379 , n15765 );
or ( n16380 , n16378 , n16379 );
nand ( n16381 , n15738 , n15735 );
nand ( n16382 , n16380 , n16381 );
not ( n16383 , n16382 );
or ( n16384 , n16377 , n16383 );
not ( n16385 , n15773 );
nand ( n16386 , n16384 , n16385 );
not ( n16387 , n16386 );
or ( n16388 , n16376 , n16387 );
nand ( n16389 , n16388 , n15725 );
nor ( n16390 , n16375 , n16389 );
or ( n16391 , n509 , n16390 );
and ( n16392 , n509 , n16390 );
not ( n16393 , n15710 );
buf ( n16394 , n16393 );
nor ( n16395 , n16392 , n16394 );
nand ( n16396 , n16391 , n16395 );
nand ( n16397 , n16373 , n16396 );
and ( n16398 , n15704 , n16397 );
not ( n16399 , n509 );
nand ( n16400 , n612 , n614 );
not ( n16401 , n16400 );
nand ( n16402 , n716 , n751 );
nor ( n16403 , n15733 , n15793 , n16402 );
nand ( n16404 , n662 , n678 , n16401 , n16403 );
not ( n16405 , n16404 );
or ( n16406 , n16399 , n16405 );
or ( n16407 , n509 , n16404 );
nand ( n16408 , n16406 , n16407 );
and ( n16409 , n1808 , n16408 );
nor ( n16410 , n16398 , n16409 );
nor ( n16411 , n15703 , n16410 );
not ( n16412 , n794 );
not ( n16413 , n16270 );
or ( n16414 , n16412 , n16413 );
not ( n16415 , n488 );
nand ( n16416 , n16415 , n16342 );
not ( n16417 , n16296 );
not ( n16418 , n16311 );
nand ( n16419 , n16418 , n16302 );
and ( n16420 , n16302 , n16280 );
nand ( n16421 , n16289 , n16317 );
nand ( n16422 , n16420 , n16421 );
nand ( n16423 , n16419 , n16334 , n16422 );
not ( n16424 , n16423 );
or ( n16425 , n16417 , n16424 );
not ( n16426 , n793 );
nand ( n16427 , n16425 , n16426 );
nor ( n16428 , n16416 , n16427 );
or ( n16429 , n794 , n16428 );
and ( n16430 , n794 , n16428 );
not ( n16431 , n16269 );
nor ( n16432 , n16430 , n16431 );
nand ( n16433 , n16429 , n16432 );
nand ( n16434 , n16414 , n16433 );
and ( n16435 , n16258 , n16434 );
not ( n16436 , n794 );
nand ( n16437 , n488 , n841 );
not ( n16438 , n16437 );
nand ( n16439 , n843 , n846 );
nor ( n16440 , n16281 , n16358 );
nand ( n16441 , n837 , n16440 );
nor ( n16442 , n16439 , n16441 );
nand ( n16443 , n807 , n16442 );
not ( n16444 , n16443 );
and ( n16445 , n804 , n16444 );
nand ( n16446 , n793 , n16438 , n16445 );
not ( n16447 , n16446 );
or ( n16448 , n16436 , n16447 );
or ( n16449 , n794 , n16446 );
nand ( n16450 , n16448 , n16449 );
and ( n16451 , n1828 , n16450 );
nor ( n16452 , n16435 , n16451 );
nor ( n16453 , n16257 , n16452 );
or ( n16454 , n432 , n15579 );
nand ( n16455 , n16454 , n16128 );
nand ( n16456 , n16455 , n15694 );
not ( n16457 , n1546 );
not ( n16458 , n15322 );
nand ( n16459 , n16457 , n16458 , n15332 , n237 );
and ( n16460 , n237 , n15316 );
not ( n16461 , n929 );
and ( n16462 , n928 , n16461 );
and ( n16463 , n1380 , n16462 );
or ( n16464 , n237 , n1380 );
nand ( n16465 , n16464 , n16114 );
nor ( n16466 , n16463 , n16465 );
nor ( n16467 , n16460 , n16466 );
and ( n16468 , n16459 , n16467 );
nor ( n16469 , n16468 , n15560 );
and ( n16470 , n146 , n14789 );
nor ( n16471 , n16470 , n14792 );
not ( n16472 , n14808 );
not ( n16473 , n13019 );
or ( n16474 , n16472 , n16473 );
and ( n16475 , n14809 , n180 );
not ( n16476 , n14809 );
and ( n16477 , n16476 , n1007 );
nor ( n16478 , n16475 , n16477 );
nor ( n16479 , n14819 , n14808 );
nand ( n16480 , n16478 , n16479 );
nand ( n16481 , n16474 , n16480 );
nand ( n16482 , n14788 , n16481 );
nand ( n16483 , n16471 , n16482 );
not ( n16484 , n155 );
not ( n16485 , n14789 );
or ( n16486 , n16484 , n16485 );
not ( n16487 , n14808 );
not ( n16488 , n12995 );
or ( n16489 , n16487 , n16488 );
and ( n16490 , n14809 , n179 );
not ( n16491 , n14809 );
and ( n16492 , n16491 , n906 );
nor ( n16493 , n16490 , n16492 );
nand ( n16494 , n16493 , n16479 );
nand ( n16495 , n16489 , n16494 );
nand ( n16496 , n15302 , n16495 );
nand ( n16497 , n16486 , n16496 );
and ( n16498 , n1112 , n12726 );
and ( n16499 , n885 , n1228 );
nor ( n16500 , n16498 , n16499 );
not ( n16501 , n141 );
buf ( n16502 , n14284 );
not ( n16503 , n16502 );
or ( n16504 , n16501 , n16503 );
nand ( n16505 , n16504 , n224 );
not ( n16506 , n16505 );
or ( n16507 , n16500 , n16506 );
not ( n16508 , n12715 );
nor ( n16509 , n16508 , n12713 );
not ( n16510 , n16509 );
not ( n16511 , n16510 );
not ( n16512 , n12813 );
not ( n16513 , n16512 );
or ( n16514 , n16511 , n16513 );
and ( n16515 , n16509 , n12813 );
nor ( n16516 , n16515 , n16505 );
nand ( n16517 , n16514 , n16516 );
nand ( n16518 , n16507 , n16517 );
not ( n16519 , n15400 );
and ( n16520 , n217 , n16519 );
nor ( n16521 , n16520 , n16118 );
or ( n16522 , n13552 , n16521 );
not ( n16523 , n13575 );
nor ( n16524 , n13552 , n16523 );
not ( n16525 , n16524 );
nand ( n16526 , n16522 , n16525 );
and ( n16527 , n15314 , n16526 );
not ( n16528 , n16115 );
and ( n16529 , n217 , n16528 );
nor ( n16530 , n16527 , n16529 );
nor ( n16531 , n16530 , n15560 );
not ( n16532 , n15349 );
not ( n16533 , n16532 );
nand ( n16534 , n15338 , n15366 );
not ( n16535 , n16534 );
nand ( n16536 , n218 , n16533 , n16535 );
not ( n16537 , n13552 );
or ( n16538 , n218 , n16537 );
not ( n16539 , n15309 );
not ( n16540 , n15399 );
or ( n16541 , n16539 , n16540 );
nand ( n16542 , n16541 , n16523 );
nor ( n16543 , n16542 , n16118 , n13527 );
or ( n16544 , n13552 , n16543 );
nand ( n16545 , n16538 , n16544 , n15314 );
and ( n16546 , n16536 , n16545 );
nor ( n16547 , n16546 , n15560 );
and ( n16548 , n224 , n15316 );
not ( n16549 , n15379 );
and ( n16550 , n16549 , n15382 );
nor ( n16551 , n16548 , n16550 );
or ( n16552 , n224 , n15322 );
nand ( n16553 , n16552 , n15324 , n15332 );
not ( n16554 , n241 );
and ( n16555 , n16554 , n240 , n15371 );
not ( n16556 , n16462 );
and ( n16557 , n1380 , n16556 );
or ( n16558 , n224 , n1380 );
nand ( n16559 , n16558 , n16114 );
nor ( n16560 , n16557 , n16559 );
nor ( n16561 , n16555 , n16560 );
and ( n16562 , n16551 , n16553 , n16561 );
nor ( n16563 , n16562 , n15560 );
or ( n16564 , n16153 , n312 );
and ( n16565 , n433 , n16564 );
not ( n16566 , n433 );
not ( n16567 , n431 );
nor ( n16568 , n16567 , n15578 );
nand ( n16569 , n432 , n16568 );
or ( n16570 , n15690 , n16569 );
or ( n16571 , n15691 , n16570 );
and ( n16572 , n16566 , n16571 );
nor ( n16573 , n16566 , n16571 );
nor ( n16574 , n16572 , n16564 , n16573 );
nor ( n16575 , n16565 , n16574 );
not ( n16576 , n16128 );
nor ( n16577 , n16575 , n16576 );
and ( n16578 , n239 , n15316 );
and ( n16579 , n15377 , n15373 );
nor ( n16580 , n16578 , n16579 );
nor ( n16581 , n16580 , n15560 );
nand ( n16582 , n16115 , n15315 );
and ( n16583 , n240 , n16582 );
and ( n16584 , n15369 , n15349 );
nor ( n16585 , n16462 , n15347 );
nor ( n16586 , n16584 , n16585 , n16534 );
nor ( n16587 , n16583 , n16586 );
nor ( n16588 , n16587 , n15560 );
and ( n16589 , n241 , n15316 );
not ( n16590 , n15327 );
nor ( n16591 , n16590 , n13532 , n239 , n15381 );
nor ( n16592 , n16589 , n16591 );
nor ( n16593 , n16592 , n15560 );
or ( n16594 , n15308 , n16532 );
not ( n16595 , n16585 );
nand ( n16596 , n16594 , n16595 );
and ( n16597 , n16596 , n16535 );
and ( n16598 , n238 , n16582 );
nor ( n16599 , n16597 , n16598 );
nor ( n16600 , n16599 , n15560 );
not ( n16601 , n16564 );
nor ( n16602 , n429 , n430 );
not ( n16603 , n16602 );
and ( n16604 , n15578 , n16601 , n16603 );
and ( n16605 , n430 , n16564 );
nor ( n16606 , n16604 , n16605 );
not ( n16607 , n16128 );
nor ( n16608 , n16606 , n16607 );
not ( n16609 , n431 );
nand ( n16610 , n16609 , n434 , n16602 );
not ( n16611 , n432 );
or ( n16612 , n15692 , n16610 , n16611 , n16566 );
nor ( n16613 , n16612 , n16607 );
not ( n16614 , n13325 );
nand ( n16615 , n16614 , n13328 );
not ( n16616 , n16615 );
and ( n16617 , n13726 , n16616 );
not ( n16618 , n13726 );
and ( n16619 , n16618 , n16615 );
nor ( n16620 , n16617 , n16619 );
not ( n16621 , n13524 );
nand ( n16622 , n16621 , n15395 );
not ( n16623 , n16622 );
nor ( n16624 , n15318 , n16623 , n15567 );
or ( n16625 , n16564 , n16569 );
nand ( n16626 , n16625 , n15690 );
and ( n16627 , n16570 , n16626 );
and ( n16628 , n413 , n16564 );
nor ( n16629 , n16627 , n16628 );
nor ( n16630 , n16629 , n16576 );
and ( n16631 , n429 , n16564 );
not ( n16632 , n429 );
and ( n16633 , n16632 , n16601 );
nor ( n16634 , n16631 , n16633 );
nor ( n16635 , n16634 , n16607 );
not ( n16636 , n16568 );
and ( n16637 , n16601 , n15579 , n16636 );
and ( n16638 , n431 , n16564 );
nor ( n16639 , n16637 , n16638 );
nor ( n16640 , n16639 , n16576 );
or ( n16641 , n16564 , n16570 );
nand ( n16642 , n16641 , n15691 );
and ( n16643 , n16571 , n16642 );
and ( n16644 , n435 , n16564 );
nor ( n16645 , n16643 , n16644 );
nor ( n16646 , n16645 , n16576 );
or ( n16647 , n16564 , n16636 );
nand ( n16648 , n16647 , n16611 );
and ( n16649 , n16569 , n16648 );
and ( n16650 , n432 , n16564 );
nor ( n16651 , n16649 , n16650 );
nor ( n16652 , n16651 , n16576 );
not ( n16653 , n595 );
not ( n16654 , n15876 );
or ( n16655 , n16653 , n16654 );
not ( n16656 , n14991 );
nor ( n16657 , n16656 , n15061 );
not ( n16658 , n16657 );
not ( n16659 , n16658 );
not ( n16660 , n14989 );
nor ( n16661 , n16660 , n14994 );
not ( n16662 , n16661 );
and ( n16663 , n14997 , n15001 );
not ( n16664 , n16663 );
not ( n16665 , n15003 );
not ( n16666 , n15032 );
not ( n16667 , n16666 );
or ( n16668 , n16665 , n16667 );
nand ( n16669 , n16668 , n15023 );
not ( n16670 , n16669 );
and ( n16671 , n15006 , n15003 );
not ( n16672 , n15028 );
not ( n16673 , n15013 );
nand ( n16674 , n16672 , n16673 );
nand ( n16675 , n16671 , n16674 );
nand ( n16676 , n16670 , n16675 );
not ( n16677 , n16676 );
or ( n16678 , n16664 , n16677 );
not ( n16679 , n15021 );
and ( n16680 , n14997 , n16679 );
not ( n16681 , n15049 );
nor ( n16682 , n16680 , n16681 );
nand ( n16683 , n16678 , n16682 );
not ( n16684 , n16683 );
or ( n16685 , n16662 , n16684 );
and ( n16686 , n14989 , n15053 );
nor ( n16687 , n16686 , n15059 );
nand ( n16688 , n16685 , n16687 );
not ( n16689 , n16688 );
not ( n16690 , n16689 );
or ( n16691 , n16659 , n16690 );
and ( n16692 , n16657 , n16688 );
not ( n16693 , n15875 );
nor ( n16694 , n16692 , n16693 );
nand ( n16695 , n16691 , n16694 );
nand ( n16696 , n16655 , n16695 );
and ( n16697 , n14974 , n16696 );
not ( n16698 , n595 );
nand ( n16699 , n15074 , n15889 );
not ( n16700 , n16699 );
or ( n16701 , n16698 , n16700 );
or ( n16702 , n595 , n16699 );
nand ( n16703 , n16701 , n16702 );
and ( n16704 , n1819 , n16703 );
nor ( n16705 , n16697 , n16704 );
nor ( n16706 , n14973 , n16705 );
and ( n16707 , n434 , n16564 );
and ( n16708 , n434 , n16573 );
nor ( n16709 , n434 , n16573 );
nor ( n16710 , n16708 , n16709 , n16564 );
nor ( n16711 , n16707 , n16710 );
nor ( n16712 , n16711 , n16576 );
not ( n16713 , n841 );
not ( n16714 , n16270 );
or ( n16715 , n16713 , n16714 );
not ( n16716 , n16295 );
nor ( n16717 , n16716 , n16341 );
not ( n16718 , n16717 );
not ( n16719 , n16718 );
not ( n16720 , n16301 );
nand ( n16721 , n16720 , n16293 );
nand ( n16722 , n16298 , n16275 );
not ( n16723 , n16722 );
and ( n16724 , n16278 , n16316 );
not ( n16725 , n16307 );
nor ( n16726 , n16724 , n16725 );
not ( n16727 , n16314 );
nand ( n16728 , n16727 , n16287 );
nand ( n16729 , n16282 , n16278 , n16728 );
nand ( n16730 , n16726 , n16729 );
and ( n16731 , n16723 , n16730 );
not ( n16732 , n16298 );
not ( n16733 , n16308 );
not ( n16734 , n16733 );
or ( n16735 , n16732 , n16734 );
nand ( n16736 , n16735 , n16329 );
nor ( n16737 , n16731 , n16736 );
or ( n16738 , n16721 , n16737 );
and ( n16739 , n16293 , n16333 );
nor ( n16740 , n16739 , n16339 );
nand ( n16741 , n16738 , n16740 );
not ( n16742 , n16741 );
not ( n16743 , n16742 );
or ( n16744 , n16719 , n16743 );
and ( n16745 , n16717 , n16741 );
not ( n16746 , n16265 );
not ( n16747 , n16746 );
buf ( n16748 , n16747 );
nor ( n16749 , n16745 , n16748 );
nand ( n16750 , n16744 , n16749 );
nand ( n16751 , n16715 , n16750 );
and ( n16752 , n16258 , n16751 );
not ( n16753 , n841 );
nand ( n16754 , n16356 , n16442 );
not ( n16755 , n16754 );
or ( n16756 , n16753 , n16755 );
or ( n16757 , n841 , n16754 );
nand ( n16758 , n16756 , n16757 );
and ( n16759 , n1828 , n16758 );
nor ( n16760 , n16752 , n16759 );
nor ( n16761 , n16257 , n16760 );
nand ( n16762 , n13318 , n13381 );
not ( n16763 , n16762 );
not ( n16764 , n14778 );
or ( n16765 , n16763 , n16764 );
or ( n16766 , n16762 , n14778 );
nand ( n16767 , n16765 , n16766 );
and ( n16768 , n14471 , n14512 );
not ( n16769 , n16768 );
nor ( n16770 , n14713 , n14724 );
not ( n16771 , n16770 );
or ( n16772 , n16769 , n16771 );
or ( n16773 , n16768 , n16770 );
nand ( n16774 , n16772 , n16773 );
not ( n16775 , n752 );
not ( n16776 , n15831 );
or ( n16777 , n16775 , n16776 );
not ( n16778 , n15108 );
nor ( n16779 , n16778 , n15177 );
not ( n16780 , n16779 );
not ( n16781 , n16780 );
not ( n16782 , n15106 );
nor ( n16783 , n16782 , n15111 );
not ( n16784 , n16783 );
and ( n16785 , n15114 , n15118 );
not ( n16786 , n16785 );
not ( n16787 , n15120 );
not ( n16788 , n15148 );
not ( n16789 , n16788 );
or ( n16790 , n16787 , n16789 );
nand ( n16791 , n16790 , n15139 );
not ( n16792 , n16791 );
not ( n16793 , n15144 );
nand ( n16794 , n16793 , n15128 );
nand ( n16795 , n15123 , n15120 , n16794 );
nand ( n16796 , n16792 , n16795 );
not ( n16797 , n16796 );
or ( n16798 , n16786 , n16797 );
not ( n16799 , n15137 );
and ( n16800 , n15114 , n16799 );
not ( n16801 , n15165 );
nor ( n16802 , n16800 , n16801 );
nand ( n16803 , n16798 , n16802 );
not ( n16804 , n16803 );
or ( n16805 , n16784 , n16804 );
and ( n16806 , n15106 , n15169 );
nor ( n16807 , n16806 , n15175 );
nand ( n16808 , n16805 , n16807 );
not ( n16809 , n16808 );
not ( n16810 , n16809 );
or ( n16811 , n16781 , n16810 );
and ( n16812 , n16779 , n16808 );
nor ( n16813 , n16812 , n15831 );
nand ( n16814 , n16811 , n16813 );
nand ( n16815 , n16777 , n16814 );
and ( n16816 , n15090 , n16815 );
not ( n16817 , n752 );
nand ( n16818 , n15190 , n15842 );
not ( n16819 , n16818 );
or ( n16820 , n16817 , n16819 );
or ( n16821 , n752 , n16818 );
nand ( n16822 , n16820 , n16821 );
and ( n16823 , n1826 , n16822 );
nor ( n16824 , n16816 , n16823 );
nor ( n16825 , n15089 , n16824 );
not ( n16826 , n844 );
nand ( n16827 , n1398 , n16826 );
not ( n16828 , n1398 );
nand ( n16829 , n844 , n16828 );
nand ( n16830 , n16827 , n16829 );
not ( n16831 , n16830 );
not ( n16832 , n1475 );
nor ( n16833 , n16832 , n838 );
nand ( n16834 , n838 , n16832 );
not ( n16835 , n16834 );
not ( n16836 , n1287 );
and ( n16837 , n849 , n16836 );
not ( n16838 , n16837 );
not ( n16839 , n1404 );
nor ( n16840 , n16839 , n808 );
not ( n16841 , n16840 );
not ( n16842 , n16841 );
and ( n16843 , n16838 , n16842 );
nor ( n16844 , n16836 , n849 );
nor ( n16845 , n16843 , n16844 );
nor ( n16846 , n16835 , n16845 );
or ( n16847 , n16833 , n16846 );
not ( n16848 , n1288 );
nand ( n16849 , n792 , n16848 );
nand ( n16850 , n16847 , n16849 );
not ( n16851 , n792 );
nand ( n16852 , n1288 , n16851 );
not ( n16853 , n1286 );
nand ( n16854 , n836 , n16853 );
not ( n16855 , n1285 );
nand ( n16856 , n839 , n16855 );
not ( n16857 , n16856 );
not ( n16858 , n1284 );
nand ( n16859 , n798 , n16858 );
not ( n16860 , n16859 );
not ( n16861 , n1283 );
nand ( n16862 , n828 , n16861 );
not ( n16863 , n16862 );
not ( n16864 , n1412 );
nor ( n16865 , n16864 , n827 );
not ( n16866 , n16865 );
nand ( n16867 , n827 , n16864 );
not ( n16868 , n1460 );
nand ( n16869 , n829 , n16868 );
nand ( n16870 , n16867 , n16869 );
nand ( n16871 , n16866 , n16870 );
not ( n16872 , n16871 );
or ( n16873 , n16863 , n16872 );
not ( n16874 , n828 );
nand ( n16875 , n1283 , n16874 );
nand ( n16876 , n16873 , n16875 );
not ( n16877 , n16876 );
or ( n16878 , n16860 , n16877 );
not ( n16879 , n798 );
nand ( n16880 , n16879 , n1284 );
nand ( n16881 , n16878 , n16880 );
not ( n16882 , n16881 );
or ( n16883 , n16857 , n16882 );
not ( n16884 , n839 );
nand ( n16885 , n1285 , n16884 );
nand ( n16886 , n16883 , n16885 );
and ( n16887 , n16854 , n16886 );
nor ( n16888 , n16853 , n836 );
nor ( n16889 , n16887 , n16888 );
nand ( n16890 , n808 , n16839 );
not ( n16891 , n16890 );
nor ( n16892 , n16889 , n16837 , n16891 );
nand ( n16893 , n16849 , n16834 , n16892 );
nand ( n16894 , n16850 , n16852 , n16893 );
not ( n16895 , n16894 );
or ( n16896 , n16831 , n16895 );
or ( n16897 , n16830 , n16894 );
nand ( n16898 , n16896 , n16897 );
not ( n16899 , n610 );
nand ( n16900 , n1306 , n16899 );
not ( n16901 , n1306 );
nand ( n16902 , n610 , n16901 );
nand ( n16903 , n16900 , n16902 );
not ( n16904 , n16903 );
not ( n16905 , n1211 );
nand ( n16906 , n513 , n16905 );
not ( n16907 , n16906 );
not ( n16908 , n1305 );
nand ( n16909 , n570 , n16908 );
not ( n16910 , n1218 );
nand ( n16911 , n611 , n16910 );
not ( n16912 , n1304 );
nor ( n16913 , n16912 , n517 );
and ( n16914 , n16911 , n16913 );
nor ( n16915 , n16910 , n611 );
nor ( n16916 , n16914 , n16915 );
not ( n16917 , n16916 );
and ( n16918 , n16909 , n16917 );
nor ( n16919 , n16908 , n570 );
nor ( n16920 , n16918 , n16919 );
or ( n16921 , n16907 , n16920 );
not ( n16922 , n513 );
nand ( n16923 , n1211 , n16922 );
nand ( n16924 , n517 , n16912 );
nand ( n16925 , n16911 , n16924 );
not ( n16926 , n1222 );
nand ( n16927 , n639 , n16926 );
not ( n16928 , n1303 );
nand ( n16929 , n571 , n16928 );
not ( n16930 , n16929 );
not ( n16931 , n1216 );
nand ( n16932 , n542 , n16931 );
not ( n16933 , n16932 );
not ( n16934 , n1302 );
nand ( n16935 , n541 , n16934 );
not ( n16936 , n16935 );
not ( n16937 , n1206 );
nor ( n16938 , n16937 , n540 );
not ( n16939 , n16938 );
nand ( n16940 , n540 , n16937 );
not ( n16941 , n1370 );
nand ( n16942 , n539 , n16941 );
nand ( n16943 , n16940 , n16942 );
nand ( n16944 , n16939 , n16943 );
not ( n16945 , n16944 );
or ( n16946 , n16936 , n16945 );
not ( n16947 , n541 );
nand ( n16948 , n1302 , n16947 );
nand ( n16949 , n16946 , n16948 );
not ( n16950 , n16949 );
or ( n16951 , n16933 , n16950 );
nor ( n16952 , n16931 , n542 );
not ( n16953 , n16952 );
nand ( n16954 , n16951 , n16953 );
not ( n16955 , n16954 );
or ( n16956 , n16930 , n16955 );
not ( n16957 , n571 );
nand ( n16958 , n1303 , n16957 );
nand ( n16959 , n16956 , n16958 );
and ( n16960 , n16927 , n16959 );
nor ( n16961 , n16926 , n639 );
nor ( n16962 , n16960 , n16961 );
nor ( n16963 , n16925 , n16962 );
nand ( n16964 , n16909 , n16906 , n16963 );
nand ( n16965 , n16921 , n16923 , n16964 );
not ( n16966 , n16965 );
or ( n16967 , n16904 , n16966 );
or ( n16968 , n16903 , n16965 );
nand ( n16969 , n16967 , n16968 );
not ( n16970 , n693 );
nand ( n16971 , n1330 , n16970 );
not ( n16972 , n1330 );
nand ( n16973 , n693 , n16972 );
nand ( n16974 , n16971 , n16973 );
not ( n16975 , n16974 );
not ( n16976 , n1378 );
nand ( n16977 , n601 , n16976 );
not ( n16978 , n16977 );
not ( n16979 , n1328 );
nand ( n16980 , n689 , n16979 );
not ( n16981 , n1327 );
nand ( n16982 , n694 , n16981 );
not ( n16983 , n1326 );
nor ( n16984 , n16983 , n615 );
and ( n16985 , n16982 , n16984 );
nor ( n16986 , n16981 , n694 );
nor ( n16987 , n16985 , n16986 );
not ( n16988 , n16987 );
and ( n16989 , n16980 , n16988 );
nor ( n16990 , n16979 , n689 );
nor ( n16991 , n16989 , n16990 );
or ( n16992 , n16978 , n16991 );
not ( n16993 , n601 );
nand ( n16994 , n1378 , n16993 );
nand ( n16995 , n615 , n16983 );
nand ( n16996 , n16995 , n16982 );
not ( n16997 , n1393 );
nand ( n16998 , n717 , n16997 );
not ( n16999 , n1325 );
nand ( n17000 , n670 , n16999 );
not ( n17001 , n17000 );
not ( n17002 , n1324 );
nand ( n17003 , n643 , n17002 );
not ( n17004 , n17003 );
not ( n17005 , n1323 );
nand ( n17006 , n642 , n17005 );
not ( n17007 , n17006 );
not ( n17008 , n1405 );
nor ( n17009 , n17008 , n641 );
not ( n17010 , n17009 );
not ( n17011 , n1321 );
nand ( n17012 , n640 , n17011 );
nand ( n17013 , n641 , n17008 );
nand ( n17014 , n17012 , n17013 );
nand ( n17015 , n17010 , n17014 );
not ( n17016 , n17015 );
or ( n17017 , n17007 , n17016 );
not ( n17018 , n642 );
nand ( n17019 , n1323 , n17018 );
nand ( n17020 , n17017 , n17019 );
not ( n17021 , n17020 );
or ( n17022 , n17004 , n17021 );
nor ( n17023 , n17002 , n643 );
not ( n17024 , n17023 );
nand ( n17025 , n17022 , n17024 );
not ( n17026 , n17025 );
or ( n17027 , n17001 , n17026 );
not ( n17028 , n670 );
nand ( n17029 , n1325 , n17028 );
nand ( n17030 , n17027 , n17029 );
and ( n17031 , n16998 , n17030 );
nor ( n17032 , n16997 , n717 );
nor ( n17033 , n17031 , n17032 );
nor ( n17034 , n16996 , n17033 );
nand ( n17035 , n16980 , n16977 , n17034 );
nand ( n17036 , n16992 , n16994 , n17035 );
not ( n17037 , n17036 );
or ( n17038 , n16975 , n17037 );
or ( n17039 , n16974 , n17036 );
nand ( n17040 , n17038 , n17039 );
not ( n17041 , n778 );
nand ( n17042 , n1361 , n17041 );
not ( n17043 , n1361 );
nand ( n17044 , n778 , n17043 );
nand ( n17045 , n17042 , n17044 );
not ( n17046 , n17045 );
not ( n17047 , n1185 );
nor ( n17048 , n17047 , n771 );
nand ( n17049 , n771 , n17047 );
not ( n17050 , n17049 );
not ( n17051 , n1348 );
nand ( n17052 , n760 , n17051 );
not ( n17053 , n1347 );
nor ( n17054 , n17053 , n697 );
and ( n17055 , n17052 , n17054 );
nor ( n17056 , n17051 , n760 );
nor ( n17057 , n17055 , n17056 );
nor ( n17058 , n17050 , n17057 );
or ( n17059 , n17048 , n17058 );
not ( n17060 , n1186 );
nand ( n17061 , n681 , n17060 );
nand ( n17062 , n17059 , n17061 );
not ( n17063 , n681 );
nand ( n17064 , n1186 , n17063 );
nand ( n17065 , n697 , n17053 );
nand ( n17066 , n17065 , n17052 );
not ( n17067 , n1346 );
nand ( n17068 , n784 , n17067 );
not ( n17069 , n1195 );
nand ( n17070 , n17069 , n756 );
not ( n17071 , n17070 );
not ( n17072 , n1345 );
nand ( n17073 , n720 , n17072 );
not ( n17074 , n17073 );
not ( n17075 , n1344 );
nand ( n17076 , n719 , n17075 );
not ( n17077 , n17076 );
not ( n17078 , n1343 );
nor ( n17079 , n17078 , n718 );
not ( n17080 , n17079 );
not ( n17081 , n1342 );
nand ( n17082 , n723 , n17081 );
nand ( n17083 , n718 , n17078 );
nand ( n17084 , n17082 , n17083 );
nand ( n17085 , n17080 , n17084 );
not ( n17086 , n17085 );
or ( n17087 , n17077 , n17086 );
not ( n17088 , n719 );
nand ( n17089 , n1344 , n17088 );
nand ( n17090 , n17087 , n17089 );
not ( n17091 , n17090 );
or ( n17092 , n17074 , n17091 );
nor ( n17093 , n17072 , n720 );
not ( n17094 , n17093 );
nand ( n17095 , n17092 , n17094 );
not ( n17096 , n17095 );
or ( n17097 , n17071 , n17096 );
not ( n17098 , n1195 );
or ( n17099 , n17098 , n756 );
nand ( n17100 , n17097 , n17099 );
and ( n17101 , n17068 , n17100 );
nor ( n17102 , n17067 , n784 );
nor ( n17103 , n17101 , n17102 );
nor ( n17104 , n17066 , n17103 );
nand ( n17105 , n17061 , n17049 , n17104 );
nand ( n17106 , n17062 , n17064 , n17105 );
not ( n17107 , n17106 );
or ( n17108 , n17046 , n17107 );
or ( n17109 , n17045 , n17106 );
nand ( n17110 , n17108 , n17109 );
not ( n17111 , n2 );
not ( n17112 , n776 );
and ( n17113 , n825 , n17112 , n15343 );
nand ( n17114 , n511 , n1755 );
not ( n17115 , n17114 );
nand ( n17116 , n1356 , n1357 );
not ( n17117 , n17116 );
nand ( n17118 , n17117 , n13542 );
nor ( n17119 , n17116 , n15392 );
not ( n17120 , n17119 );
nand ( n17121 , n17117 , n13522 );
nand ( n17122 , n17117 , n13559 );
and ( n17123 , n17118 , n17120 , n17121 , n17122 );
nand ( n17124 , n13550 , n13544 );
nor ( n17125 , n17124 , n16622 );
nand ( n17126 , n1757 , n17123 , n17125 );
nand ( n17127 , n15341 , n17126 );
not ( n17128 , n17127 );
or ( n17129 , n17115 , n17128 );
or ( n17130 , n511 , n17127 );
nand ( n17131 , n17129 , n17130 );
nor ( n17132 , n1756 , n15321 );
nand ( n17133 , n1755 , n1757 );
nor ( n17134 , n1756 , n17133 );
not ( n17135 , n17123 );
and ( n17136 , n17134 , n17135 );
or ( n17137 , n17131 , n17132 , n17136 );
not ( n17138 , n17134 );
nor ( n17139 , n17138 , n17125 );
not ( n17140 , n17139 );
or ( n17141 , n17132 , n17140 );
nand ( n17142 , n17137 , n17141 );
and ( n17143 , n17113 , n17142 );
not ( n17144 , n17114 );
and ( n17145 , n17113 , n17132 );
and ( n17146 , n17144 , n17145 );
not ( n17147 , n15341 );
not ( n17148 , n17147 );
or ( n17149 , n17114 , n17148 );
not ( n17150 , n511 );
not ( n17151 , n17148 );
or ( n17152 , n17150 , n17151 );
nand ( n17153 , n17149 , n17152 );
not ( n17154 , n824 );
nor ( n17155 , n776 , n825 );
nand ( n17156 , n17154 , n511 , n17155 );
or ( n17157 , n17134 , n17156 );
nand ( n17158 , n17157 , n15344 );
and ( n17159 , n17153 , n17158 );
nor ( n17160 , n17143 , n17146 , n17159 );
nor ( n17161 , n17111 , n17160 );
not ( n17162 , n691 );
not ( n17163 , n15713 );
or ( n17164 , n17162 , n17163 );
and ( n17165 , n15742 , n15734 );
not ( n17166 , n17165 );
and ( n17167 , n15751 , n15746 );
not ( n17168 , n15760 );
nand ( n17169 , n17168 , n15756 );
nand ( n17170 , n17167 , n17169 );
nor ( n17171 , n17166 , n17170 );
and ( n17172 , n15728 , n15740 );
nand ( n17173 , n17171 , n15720 , n17172 );
nor ( n17174 , n509 , n15724 );
not ( n17175 , n17172 );
not ( n17176 , n17165 );
not ( n17177 , n15746 );
not ( n17178 , n15763 );
or ( n17179 , n17177 , n17178 );
nand ( n17180 , n17179 , n15737 );
not ( n17181 , n17180 );
or ( n17182 , n17176 , n17181 );
and ( n17183 , n15742 , n15732 );
nor ( n17184 , n17183 , n15771 );
nand ( n17185 , n17182 , n17184 );
not ( n17186 , n17185 );
or ( n17187 , n17175 , n17186 );
not ( n17188 , n15770 );
and ( n17189 , n15728 , n17188 );
nor ( n17190 , n17189 , n15722 );
nand ( n17191 , n17187 , n17190 );
nand ( n17192 , n15720 , n17191 );
and ( n17193 , n17173 , n17174 , n17192 );
or ( n17194 , n691 , n17193 );
and ( n17195 , n691 , n17193 );
not ( n17196 , n15709 );
not ( n17197 , n17196 );
not ( n17198 , n17197 );
nor ( n17199 , n17195 , n17198 );
nand ( n17200 , n17194 , n17199 );
nand ( n17201 , n17164 , n17200 );
and ( n17202 , n15704 , n17201 );
nand ( n17203 , n16401 , n15796 );
nor ( n17204 , n15790 , n17203 );
and ( n17205 , n17204 , n691 );
not ( n17206 , n17204 );
and ( n17207 , n17206 , n15727 );
nor ( n17208 , n17205 , n17207 );
and ( n17209 , n1808 , n17208 );
nor ( n17210 , n17202 , n17209 );
nor ( n17211 , n15703 , n17210 );
not ( n17212 , n662 );
not ( n17213 , n16394 );
or ( n17214 , n17212 , n17213 );
not ( n17215 , n15720 );
nor ( n17216 , n17215 , n15724 );
not ( n17217 , n17216 );
not ( n17218 , n17217 );
not ( n17219 , n17172 );
not ( n17220 , n17165 );
not ( n17221 , n17180 );
nand ( n17222 , n17221 , n17170 );
not ( n17223 , n17222 );
or ( n17224 , n17220 , n17223 );
nand ( n17225 , n17224 , n17184 );
not ( n17226 , n17225 );
or ( n17227 , n17219 , n17226 );
nand ( n17228 , n17227 , n17190 );
not ( n17229 , n17228 );
not ( n17230 , n17229 );
or ( n17231 , n17218 , n17230 );
and ( n17232 , n17216 , n17228 );
nor ( n17233 , n17232 , n17198 );
nand ( n17234 , n17231 , n17233 );
nand ( n17235 , n17214 , n17234 );
and ( n17236 , n15704 , n17235 );
not ( n17237 , n662 );
not ( n17238 , n17203 );
or ( n17239 , n17237 , n17238 );
or ( n17240 , n662 , n17203 );
nand ( n17241 , n17239 , n17240 );
and ( n17242 , n1808 , n17241 );
nor ( n17243 , n17236 , n17242 );
nor ( n17244 , n15703 , n17243 );
and ( n17245 , n1023 , n12726 );
and ( n17246 , n957 , n1228 );
nor ( n17247 , n17245 , n17246 );
or ( n17248 , n17247 , n16506 );
not ( n17249 , n12667 );
nor ( n17250 , n17249 , n12702 );
or ( n17251 , n17250 , n12698 );
and ( n17252 , n17250 , n12698 );
nor ( n17253 , n17252 , n16505 );
nand ( n17254 , n17251 , n17253 );
nand ( n17255 , n17248 , n17254 );
not ( n17256 , n14513 );
nand ( n17257 , n17256 , n14470 );
not ( n17258 , n17257 );
not ( n17259 , n14503 );
or ( n17260 , n17258 , n17259 );
or ( n17261 , n17257 , n14503 );
nand ( n17262 , n17260 , n17261 );
not ( n17263 , n512 );
not ( n17264 , n15876 );
or ( n17265 , n17263 , n17264 );
not ( n17266 , n512 );
nor ( n17267 , n570 , n1248 );
nor ( n17268 , n611 , n1396 );
nor ( n17269 , n17267 , n17268 );
not ( n17270 , n17269 );
not ( n17271 , n1250 );
nand ( n17272 , n17271 , n16957 );
not ( n17273 , n17272 );
nor ( n17274 , n542 , n1401 );
nor ( n17275 , n17273 , n17274 );
nor ( n17276 , n517 , n1399 );
nor ( n17277 , n639 , n1403 );
nor ( n17278 , n17276 , n17277 );
and ( n17279 , n17275 , n17278 );
not ( n17280 , n17279 );
nand ( n17281 , n540 , n1406 );
nor ( n17282 , n541 , n1152 );
or ( n17283 , n17281 , n17282 );
nand ( n17284 , n541 , n1152 );
nand ( n17285 , n17283 , n17284 );
not ( n17286 , n17285 );
not ( n17287 , n17282 );
nand ( n17288 , n539 , n1151 );
nor ( n17289 , n540 , n1406 );
nor ( n17290 , n17288 , n17289 );
nand ( n17291 , n17287 , n17290 );
nand ( n17292 , n17286 , n17291 );
not ( n17293 , n17292 );
or ( n17294 , n17280 , n17293 );
nand ( n17295 , n542 , n1401 );
not ( n17296 , n17295 );
not ( n17297 , n17296 );
not ( n17298 , n17272 );
or ( n17299 , n17297 , n17298 );
nand ( n17300 , n571 , n1250 );
nand ( n17301 , n17299 , n17300 );
and ( n17302 , n17278 , n17301 );
nand ( n17303 , n639 , n1403 );
or ( n17304 , n17303 , n17276 );
nand ( n17305 , n517 , n1399 );
nand ( n17306 , n17304 , n17305 );
nor ( n17307 , n17302 , n17306 );
nand ( n17308 , n17294 , n17307 );
not ( n17309 , n17308 );
or ( n17310 , n17270 , n17309 );
nand ( n17311 , n611 , n1396 );
or ( n17312 , n17311 , n17267 );
nand ( n17313 , n570 , n1248 );
nand ( n17314 , n17312 , n17313 );
not ( n17315 , n17314 );
nand ( n17316 , n17310 , n17315 );
nand ( n17317 , n610 , n513 , n17316 );
not ( n17318 , n17317 );
not ( n17319 , n17318 );
or ( n17320 , n17266 , n17319 );
not ( n17321 , n512 );
and ( n17322 , n17321 , n17317 );
nor ( n17323 , n17322 , n16693 );
nand ( n17324 , n17320 , n17323 );
nand ( n17325 , n17265 , n17324 );
and ( n17326 , n14974 , n17325 );
not ( n17327 , n512 );
nor ( n17328 , n513 , n570 );
not ( n17329 , n517 );
nor ( n17330 , n571 , n639 );
nor ( n17331 , n539 , n540 );
nand ( n17332 , n16947 , n17331 );
nor ( n17333 , n542 , n17332 );
nand ( n17334 , n17329 , n17330 , n17333 );
nor ( n17335 , n611 , n17334 );
nand ( n17336 , n16899 , n17328 , n17335 );
not ( n17337 , n17336 );
or ( n17338 , n17327 , n17337 );
or ( n17339 , n512 , n17336 );
nand ( n17340 , n17338 , n17339 );
and ( n17341 , n1819 , n17340 );
nor ( n17342 , n17326 , n17341 );
nor ( n17343 , n14973 , n17342 );
not ( n17344 , n600 );
not ( n17345 , n16394 );
or ( n17346 , n17344 , n17345 );
not ( n17347 , n600 );
nor ( n17348 , n694 , n1158 );
nor ( n17349 , n689 , n1256 );
nor ( n17350 , n17348 , n17349 );
not ( n17351 , n17350 );
not ( n17352 , n1212 );
nand ( n17353 , n17352 , n17028 );
not ( n17354 , n17353 );
nor ( n17355 , n643 , n1157 );
nor ( n17356 , n17354 , n17355 );
nor ( n17357 , n615 , n1205 );
nor ( n17358 , n717 , n1259 );
nor ( n17359 , n17357 , n17358 );
and ( n17360 , n17356 , n17359 );
not ( n17361 , n17360 );
nand ( n17362 , n641 , n1439 );
nor ( n17363 , n642 , n1258 );
or ( n17364 , n17362 , n17363 );
nand ( n17365 , n642 , n1258 );
nand ( n17366 , n17364 , n17365 );
not ( n17367 , n17366 );
not ( n17368 , n17363 );
nand ( n17369 , n640 , n1156 );
nor ( n17370 , n641 , n1439 );
nor ( n17371 , n17369 , n17370 );
nand ( n17372 , n17368 , n17371 );
nand ( n17373 , n17367 , n17372 );
not ( n17374 , n17373 );
or ( n17375 , n17361 , n17374 );
nand ( n17376 , n643 , n1157 );
not ( n17377 , n17376 );
not ( n17378 , n17377 );
not ( n17379 , n17353 );
or ( n17380 , n17378 , n17379 );
nand ( n17381 , n670 , n1212 );
nand ( n17382 , n17380 , n17381 );
and ( n17383 , n17359 , n17382 );
nand ( n17384 , n717 , n1259 );
or ( n17385 , n17384 , n17357 );
nand ( n17386 , n615 , n1205 );
nand ( n17387 , n17385 , n17386 );
nor ( n17388 , n17383 , n17387 );
nand ( n17389 , n17375 , n17388 );
not ( n17390 , n17389 );
or ( n17391 , n17351 , n17390 );
nand ( n17392 , n694 , n1158 );
or ( n17393 , n17392 , n17349 );
nand ( n17394 , n689 , n1256 );
nand ( n17395 , n17393 , n17394 );
not ( n17396 , n17395 );
nand ( n17397 , n17391 , n17396 );
nand ( n17398 , n693 , n601 , n17397 );
not ( n17399 , n17398 );
not ( n17400 , n17399 );
or ( n17401 , n17347 , n17400 );
not ( n17402 , n600 );
and ( n17403 , n17402 , n17398 );
nor ( n17404 , n17403 , n16394 );
nand ( n17405 , n17401 , n17404 );
nand ( n17406 , n17346 , n17405 );
and ( n17407 , n15704 , n17406 );
not ( n17408 , n600 );
nor ( n17409 , n601 , n689 );
not ( n17410 , n615 );
nor ( n17411 , n670 , n717 );
nor ( n17412 , n640 , n641 );
nand ( n17413 , n17018 , n17412 );
nor ( n17414 , n643 , n17413 );
nand ( n17415 , n17410 , n17411 , n17414 );
nor ( n17416 , n694 , n17415 );
nand ( n17417 , n16970 , n17409 , n17416 );
not ( n17418 , n17417 );
or ( n17419 , n17408 , n17418 );
or ( n17420 , n600 , n17417 );
nand ( n17421 , n17419 , n17420 );
and ( n17422 , n1808 , n17421 );
nor ( n17423 , n17407 , n17422 );
nor ( n17424 , n15703 , n17423 );
not ( n17425 , n599 );
not ( n17426 , n14983 );
or ( n17427 , n17425 , n17426 );
not ( n17428 , n16663 );
nor ( n17429 , n17428 , n16675 );
and ( n17430 , n17429 , n14991 , n16661 );
not ( n17431 , n14991 );
not ( n17432 , n16661 );
not ( n17433 , n16663 );
not ( n17434 , n16669 );
or ( n17435 , n17433 , n17434 );
nand ( n17436 , n17435 , n16682 );
not ( n17437 , n17436 );
or ( n17438 , n17432 , n17437 );
nand ( n17439 , n17438 , n16687 );
not ( n17440 , n17439 );
or ( n17441 , n17431 , n17440 );
nor ( n17442 , n508 , n15061 );
nand ( n17443 , n17441 , n17442 );
nor ( n17444 , n17430 , n17443 );
or ( n17445 , n599 , n17444 );
and ( n17446 , n599 , n17444 );
nor ( n17447 , n17446 , n16693 );
nand ( n17448 , n17445 , n17447 );
nand ( n17449 , n17427 , n17448 );
and ( n17450 , n14974 , n17449 );
nor ( n17451 , n15884 , n16699 );
and ( n17452 , n17451 , n599 );
not ( n17453 , n17451 );
and ( n17454 , n17453 , n15860 );
nor ( n17455 , n17452 , n17454 );
and ( n17456 , n1819 , n17455 );
nor ( n17457 , n17450 , n17456 );
nor ( n17458 , n14973 , n17457 );
not ( n17459 , n774 );
not ( n17460 , n15100 );
or ( n17461 , n17459 , n17460 );
nand ( n17462 , n15108 , n16783 );
not ( n17463 , n16795 );
nand ( n17464 , n17463 , n16785 );
nor ( n17465 , n17462 , n17464 );
not ( n17466 , n15108 );
not ( n17467 , n16783 );
not ( n17468 , n16785 );
not ( n17469 , n16791 );
or ( n17470 , n17468 , n17469 );
nand ( n17471 , n17470 , n16802 );
not ( n17472 , n17471 );
or ( n17473 , n17467 , n17472 );
nand ( n17474 , n17473 , n16807 );
not ( n17475 , n17474 );
or ( n17476 , n17466 , n17475 );
nor ( n17477 , n487 , n15177 );
nand ( n17478 , n17476 , n17477 );
nor ( n17479 , n17465 , n17478 );
or ( n17480 , n774 , n17479 );
and ( n17481 , n774 , n17479 );
nor ( n17482 , n17481 , n15098 );
nand ( n17483 , n17480 , n17482 );
nand ( n17484 , n17461 , n17483 );
and ( n17485 , n15090 , n17484 );
nor ( n17486 , n15837 , n16818 );
and ( n17487 , n17486 , n774 );
not ( n17488 , n17486 );
and ( n17489 , n17488 , n15814 );
nor ( n17490 , n17487 , n17489 );
and ( n17491 , n1826 , n17490 );
nor ( n17492 , n17485 , n17491 );
nor ( n17493 , n15089 , n17492 );
or ( n17494 , n16426 , n16269 );
not ( n17495 , n16426 );
nor ( n17496 , n16716 , n16721 );
not ( n17497 , n17496 );
not ( n17498 , n16723 );
nor ( n17499 , n17498 , n16729 );
not ( n17500 , n17499 );
or ( n17501 , n17497 , n17500 );
nor ( n17502 , n488 , n16341 );
nand ( n17503 , n17501 , n17502 );
not ( n17504 , n16721 );
or ( n17505 , n16722 , n16726 );
not ( n17506 , n16736 );
nand ( n17507 , n17505 , n17506 );
nand ( n17508 , n17504 , n17507 );
and ( n17509 , n16740 , n17508 );
nor ( n17510 , n17509 , n16716 );
nor ( n17511 , n17503 , n17510 );
not ( n17512 , n17511 );
not ( n17513 , n17512 );
or ( n17514 , n17495 , n17513 );
and ( n17515 , n793 , n17511 );
nor ( n17516 , n17515 , n16748 );
nand ( n17517 , n17514 , n17516 );
nand ( n17518 , n17494 , n17517 );
and ( n17519 , n16258 , n17518 );
nor ( n17520 , n16437 , n16754 );
and ( n17521 , n17520 , n793 );
not ( n17522 , n17520 );
and ( n17523 , n17522 , n16426 );
nor ( n17524 , n17521 , n17523 );
and ( n17525 , n1828 , n17524 );
nor ( n17526 , n17519 , n17525 );
nor ( n17527 , n16257 , n17526 );
not ( n17528 , n803 );
not ( n17529 , n16270 );
or ( n17530 , n17528 , n17529 );
not ( n17531 , n803 );
nor ( n17532 , n838 , n1231 );
nor ( n17533 , n849 , n1239 );
nor ( n17534 , n17532 , n17533 );
not ( n17535 , n17534 );
not ( n17536 , n1237 );
nand ( n17537 , n17536 , n16884 );
not ( n17538 , n17537 );
nor ( n17539 , n798 , n1236 );
nor ( n17540 , n17538 , n17539 );
nor ( n17541 , n836 , n1210 );
nor ( n17542 , n808 , n1238 );
nor ( n17543 , n17541 , n17542 );
and ( n17544 , n17540 , n17543 );
not ( n17545 , n17544 );
nand ( n17546 , n827 , n1467 );
nor ( n17547 , n828 , n1235 );
or ( n17548 , n17546 , n17547 );
nand ( n17549 , n828 , n1235 );
nand ( n17550 , n17548 , n17549 );
not ( n17551 , n17550 );
not ( n17552 , n17547 );
nand ( n17553 , n829 , n1234 );
nor ( n17554 , n827 , n1467 );
nor ( n17555 , n17553 , n17554 );
nand ( n17556 , n17552 , n17555 );
nand ( n17557 , n17551 , n17556 );
not ( n17558 , n17557 );
or ( n17559 , n17545 , n17558 );
nand ( n17560 , n798 , n1236 );
not ( n17561 , n17560 );
not ( n17562 , n17561 );
not ( n17563 , n17537 );
or ( n17564 , n17562 , n17563 );
nand ( n17565 , n839 , n1237 );
nand ( n17566 , n17564 , n17565 );
and ( n17567 , n17543 , n17566 );
nand ( n17568 , n836 , n1210 );
or ( n17569 , n17568 , n17542 );
nand ( n17570 , n808 , n1238 );
nand ( n17571 , n17569 , n17570 );
nor ( n17572 , n17567 , n17571 );
nand ( n17573 , n17559 , n17572 );
not ( n17574 , n17573 );
or ( n17575 , n17535 , n17574 );
nand ( n17576 , n849 , n1239 );
or ( n17577 , n17576 , n17532 );
nand ( n17578 , n838 , n1231 );
nand ( n17579 , n17577 , n17578 );
not ( n17580 , n17579 );
nand ( n17581 , n17575 , n17580 );
nand ( n17582 , n844 , n792 , n17581 );
not ( n17583 , n17582 );
not ( n17584 , n17583 );
or ( n17585 , n17531 , n17584 );
not ( n17586 , n803 );
and ( n17587 , n17586 , n17582 );
nor ( n17588 , n17587 , n16748 );
nand ( n17589 , n17585 , n17588 );
nand ( n17590 , n17530 , n17589 );
and ( n17591 , n16258 , n17590 );
nor ( n17592 , n792 , n838 );
not ( n17593 , n808 );
not ( n17594 , n836 );
and ( n17595 , n17594 , n16884 );
nor ( n17596 , n827 , n829 );
nand ( n17597 , n16874 , n17596 );
nor ( n17598 , n798 , n17597 );
nand ( n17599 , n17593 , n17595 , n17598 );
nor ( n17600 , n849 , n17599 );
nand ( n17601 , n16826 , n17592 , n17600 );
xnor ( n17602 , n803 , n17601 );
and ( n17603 , n1828 , n17602 );
nor ( n17604 , n17591 , n17603 );
nor ( n17605 , n16257 , n17604 );
not ( n17606 , n692 );
not ( n17607 , n15831 );
or ( n17608 , n17606 , n17607 );
not ( n17609 , n692 );
nor ( n17610 , n760 , n1163 );
nor ( n17611 , n771 , n1268 );
nor ( n17612 , n17610 , n17611 );
not ( n17613 , n17612 );
not ( n17614 , n1162 );
not ( n17615 , n756 );
nand ( n17616 , n17614 , n17615 );
not ( n17617 , n17616 );
nor ( n17618 , n720 , n1387 );
nor ( n17619 , n17617 , n17618 );
nor ( n17620 , n784 , n1271 );
nor ( n17621 , n697 , n1394 );
nor ( n17622 , n17620 , n17621 );
and ( n17623 , n17619 , n17622 );
not ( n17624 , n17623 );
nand ( n17625 , n718 , n1471 );
nor ( n17626 , n719 , n1270 );
or ( n17627 , n17625 , n17626 );
nand ( n17628 , n719 , n1270 );
nand ( n17629 , n17627 , n17628 );
not ( n17630 , n17629 );
not ( n17631 , n17626 );
nand ( n17632 , n723 , n1161 );
nor ( n17633 , n718 , n1471 );
nor ( n17634 , n17632 , n17633 );
nand ( n17635 , n17631 , n17634 );
nand ( n17636 , n17630 , n17635 );
not ( n17637 , n17636 );
or ( n17638 , n17624 , n17637 );
nand ( n17639 , n720 , n1387 );
not ( n17640 , n17639 );
not ( n17641 , n17640 );
not ( n17642 , n17616 );
or ( n17643 , n17641 , n17642 );
nand ( n17644 , n756 , n1162 );
nand ( n17645 , n17643 , n17644 );
and ( n17646 , n17622 , n17645 );
nand ( n17647 , n784 , n1271 );
or ( n17648 , n17647 , n17621 );
nand ( n17649 , n697 , n1394 );
nand ( n17650 , n17648 , n17649 );
nor ( n17651 , n17646 , n17650 );
nand ( n17652 , n17638 , n17651 );
not ( n17653 , n17652 );
or ( n17654 , n17613 , n17653 );
nand ( n17655 , n760 , n1163 );
or ( n17656 , n17655 , n17611 );
nand ( n17657 , n771 , n1268 );
nand ( n17658 , n17656 , n17657 );
not ( n17659 , n17658 );
nand ( n17660 , n17654 , n17659 );
nand ( n17661 , n778 , n681 , n17660 );
not ( n17662 , n17661 );
not ( n17663 , n17662 );
or ( n17664 , n17609 , n17663 );
not ( n17665 , n692 );
and ( n17666 , n17665 , n17661 );
not ( n17667 , n15830 );
nor ( n17668 , n17666 , n17667 );
nand ( n17669 , n17664 , n17668 );
nand ( n17670 , n17608 , n17669 );
and ( n17671 , n15090 , n17670 );
not ( n17672 , n692 );
nor ( n17673 , n681 , n771 );
not ( n17674 , n697 );
nor ( n17675 , n756 , n784 );
nor ( n17676 , n718 , n723 );
nand ( n17677 , n17088 , n17676 );
nor ( n17678 , n720 , n17677 );
nand ( n17679 , n17674 , n17675 , n17678 );
nor ( n17680 , n760 , n17679 );
nand ( n17681 , n17041 , n17673 , n17680 );
not ( n17682 , n17681 );
or ( n17683 , n17672 , n17682 );
or ( n17684 , n692 , n17681 );
nand ( n17685 , n17683 , n17684 );
and ( n17686 , n1826 , n17685 );
nor ( n17687 , n17671 , n17686 );
nor ( n17688 , n15089 , n17687 );
not ( n17689 , n838 );
not ( n17690 , n16270 );
or ( n17691 , n17689 , n17690 );
not ( n17692 , n17578 );
or ( n17693 , n17692 , n17532 );
nor ( n17694 , n17542 , n17533 );
not ( n17695 , n17537 );
nor ( n17696 , n17541 , n17695 );
not ( n17697 , n17696 );
or ( n17698 , n17549 , n17539 );
nand ( n17699 , n17698 , n17560 );
not ( n17700 , n17699 );
nor ( n17701 , n17547 , n17539 );
not ( n17702 , n17555 );
nand ( n17703 , n17546 , n17702 );
nand ( n17704 , n17701 , n17703 );
nand ( n17705 , n17700 , n17704 );
not ( n17706 , n17705 );
or ( n17707 , n17697 , n17706 );
or ( n17708 , n17565 , n17541 );
nand ( n17709 , n17708 , n17568 );
not ( n17710 , n17709 );
nand ( n17711 , n17707 , n17710 );
and ( n17712 , n17694 , n17711 );
or ( n17713 , n17570 , n17533 );
nand ( n17714 , n17713 , n17576 );
nor ( n17715 , n17712 , n17714 );
or ( n17716 , n17693 , n17715 );
nand ( n17717 , n17693 , n17715 );
nand ( n17718 , n17716 , n17717 , n16269 );
nand ( n17719 , n17691 , n17718 );
and ( n17720 , n16258 , n17719 );
not ( n17721 , n838 );
not ( n17722 , n17721 );
nor ( n17723 , n808 , n849 );
nand ( n17724 , n17595 , n17723 );
not ( n17725 , n17598 );
nor ( n17726 , n17724 , n17725 );
not ( n17727 , n17726 );
or ( n17728 , n17722 , n17727 );
or ( n17729 , n17721 , n17726 );
nand ( n17730 , n17728 , n17729 );
and ( n17731 , n1828 , n17730 );
nor ( n17732 , n17720 , n17731 );
nor ( n17733 , n16257 , n17732 );
not ( n17734 , n2 );
nand ( n17735 , n776 , n1755 );
not ( n17736 , n17127 );
or ( n17737 , n17735 , n17736 );
and ( n17738 , n776 , n17736 );
nor ( n17739 , n17738 , n17136 );
nand ( n17740 , n17737 , n17739 );
not ( n17741 , n17113 );
nor ( n17742 , n17741 , n17132 );
and ( n17743 , n17740 , n17742 , n17140 );
and ( n17744 , n17151 , n17735 );
not ( n17745 , n17151 );
and ( n17746 , n17745 , n17112 );
nor ( n17747 , n17744 , n17746 );
and ( n17748 , n17747 , n17158 );
nor ( n17749 , n17743 , n17748 );
nor ( n17750 , n17734 , n17749 );
not ( n17751 , n771 );
not ( n17752 , n15831 );
or ( n17753 , n17751 , n17752 );
not ( n17754 , n17657 );
or ( n17755 , n17754 , n17611 );
nor ( n17756 , n17610 , n17621 );
not ( n17757 , n17616 );
nor ( n17758 , n17757 , n17620 );
not ( n17759 , n17758 );
or ( n17760 , n17628 , n17618 );
nand ( n17761 , n17760 , n17639 );
not ( n17762 , n17761 );
nor ( n17763 , n17626 , n17618 );
not ( n17764 , n17634 );
nand ( n17765 , n17625 , n17764 );
nand ( n17766 , n17763 , n17765 );
nand ( n17767 , n17762 , n17766 );
not ( n17768 , n17767 );
or ( n17769 , n17759 , n17768 );
or ( n17770 , n17644 , n17620 );
nand ( n17771 , n17770 , n17647 );
not ( n17772 , n17771 );
nand ( n17773 , n17769 , n17772 );
and ( n17774 , n17756 , n17773 );
or ( n17775 , n17649 , n17610 );
nand ( n17776 , n17775 , n17655 );
nor ( n17777 , n17774 , n17776 );
or ( n17778 , n17755 , n17777 );
nand ( n17779 , n17755 , n17777 );
nand ( n17780 , n17778 , n17779 , n15099 );
nand ( n17781 , n17753 , n17780 );
and ( n17782 , n15090 , n17781 );
nor ( n17783 , n697 , n760 );
nand ( n17784 , n17783 , n17675 );
not ( n17785 , n17784 );
nand ( n17786 , n17785 , n17678 );
not ( n17787 , n771 );
xor ( n17788 , n17786 , n17787 );
and ( n17789 , n1826 , n17788 );
nor ( n17790 , n17782 , n17789 );
nor ( n17791 , n15089 , n17790 );
not ( n17792 , n402 );
not ( n17793 , n1146 );
or ( n17794 , n17792 , n17793 );
or ( n17795 , n402 , n1146 );
nand ( n17796 , n17794 , n17795 );
not ( n17797 , n1173 );
and ( n17798 , n381 , n17797 );
not ( n17799 , n381 );
and ( n17800 , n17799 , n1173 );
nor ( n17801 , n17798 , n17800 );
and ( n17802 , n400 , n15410 );
not ( n17803 , n400 );
and ( n17804 , n17803 , n1169 );
nor ( n17805 , n17802 , n17804 );
and ( n17806 , n392 , n15446 );
not ( n17807 , n392 );
and ( n17808 , n17807 , n1172 );
nor ( n17809 , n17806 , n17808 );
nand ( n17810 , n17796 , n17801 , n17805 , n17809 );
not ( n17811 , n1446 );
and ( n17812 , n384 , n17811 );
and ( n17813 , n379 , n1447 );
not ( n17814 , n379 );
and ( n17815 , n17814 , n15467 );
nor ( n17816 , n17813 , n17815 );
nor ( n17817 , n17811 , n384 );
nor ( n17818 , n17812 , n17816 , n17817 );
not ( n17819 , n382 );
not ( n17820 , n1442 );
or ( n17821 , n17819 , n17820 );
or ( n17822 , n382 , n1442 );
nand ( n17823 , n17821 , n17822 );
and ( n17824 , n398 , n15405 );
not ( n17825 , n399 );
not ( n17826 , n1170 );
and ( n17827 , n17825 , n17826 );
and ( n17828 , n399 , n1170 );
nor ( n17829 , n17827 , n17828 );
nor ( n17830 , n15405 , n398 );
nor ( n17831 , n17824 , n17829 , n17830 );
and ( n17832 , n401 , n15420 );
not ( n17833 , n380 );
not ( n17834 , n1171 );
and ( n17835 , n17833 , n17834 );
and ( n17836 , n380 , n1171 );
nor ( n17837 , n17835 , n17836 );
nor ( n17838 , n15420 , n401 );
nor ( n17839 , n17832 , n17837 , n17838 );
nand ( n17840 , n17818 , n17823 , n17831 , n17839 );
not ( n17841 , n15556 );
nor ( n17842 , n15318 , n13550 , n17841 );
not ( n17843 , n17842 );
nor ( n17844 , n17810 , n17840 , n17843 );
not ( n17845 , n570 );
not ( n17846 , n15876 );
or ( n17847 , n17845 , n17846 );
not ( n17848 , n17313 );
or ( n17849 , n17848 , n17267 );
nor ( n17850 , n17268 , n17276 );
not ( n17851 , n17272 );
nor ( n17852 , n17851 , n17277 );
not ( n17853 , n17852 );
or ( n17854 , n17284 , n17274 );
nand ( n17855 , n17854 , n17295 );
not ( n17856 , n17855 );
nor ( n17857 , n17282 , n17274 );
not ( n17858 , n17290 );
nand ( n17859 , n17281 , n17858 );
nand ( n17860 , n17857 , n17859 );
nand ( n17861 , n17856 , n17860 );
not ( n17862 , n17861 );
or ( n17863 , n17853 , n17862 );
or ( n17864 , n17300 , n17277 );
nand ( n17865 , n17864 , n17303 );
not ( n17866 , n17865 );
nand ( n17867 , n17863 , n17866 );
and ( n17868 , n17850 , n17867 );
or ( n17869 , n17305 , n17268 );
nand ( n17870 , n17869 , n17311 );
nor ( n17871 , n17868 , n17870 );
or ( n17872 , n17849 , n17871 );
nand ( n17873 , n17849 , n17871 );
nand ( n17874 , n17872 , n17873 , n14982 );
nand ( n17875 , n17847 , n17874 );
and ( n17876 , n14974 , n17875 );
not ( n17877 , n570 );
not ( n17878 , n17877 );
nor ( n17879 , n517 , n611 );
nand ( n17880 , n17879 , n17330 );
not ( n17881 , n17333 );
nor ( n17882 , n17880 , n17881 );
not ( n17883 , n17882 );
or ( n17884 , n17878 , n17883 );
or ( n17885 , n17877 , n17882 );
nand ( n17886 , n17884 , n17885 );
and ( n17887 , n1819 , n17886 );
nor ( n17888 , n17876 , n17887 );
nor ( n17889 , n14973 , n17888 );
nand ( n17890 , n14481 , n14475 );
not ( n17891 , n17890 );
not ( n17892 , n14955 );
or ( n17893 , n17891 , n17892 );
or ( n17894 , n17890 , n14955 );
nand ( n17895 , n17893 , n17894 );
not ( n17896 , n689 );
not ( n17897 , n15713 );
or ( n17898 , n17896 , n17897 );
not ( n17899 , n17394 );
or ( n17900 , n17899 , n17349 );
nor ( n17901 , n17348 , n17357 );
not ( n17902 , n17353 );
nor ( n17903 , n17902 , n17358 );
not ( n17904 , n17903 );
or ( n17905 , n17365 , n17355 );
nand ( n17906 , n17905 , n17376 );
not ( n17907 , n17906 );
nor ( n17908 , n17355 , n17363 );
not ( n17909 , n17371 );
nand ( n17910 , n17362 , n17909 );
nand ( n17911 , n17908 , n17910 );
nand ( n17912 , n17907 , n17911 );
not ( n17913 , n17912 );
or ( n17914 , n17904 , n17913 );
or ( n17915 , n17381 , n17358 );
nand ( n17916 , n17915 , n17384 );
not ( n17917 , n17916 );
nand ( n17918 , n17914 , n17917 );
and ( n17919 , n17901 , n17918 );
or ( n17920 , n17386 , n17348 );
nand ( n17921 , n17920 , n17392 );
nor ( n17922 , n17919 , n17921 );
or ( n17923 , n17900 , n17922 );
nand ( n17924 , n17900 , n17922 );
nand ( n17925 , n17923 , n17924 , n15712 );
nand ( n17926 , n17898 , n17925 );
and ( n17927 , n15704 , n17926 );
nor ( n17928 , n615 , n694 );
nand ( n17929 , n17928 , n17411 );
not ( n17930 , n17929 );
nand ( n17931 , n17930 , n17414 );
not ( n17932 , n689 );
xor ( n17933 , n17931 , n17932 );
and ( n17934 , n1808 , n17933 );
nor ( n17935 , n17927 , n17934 );
nor ( n17936 , n15703 , n17935 );
not ( n17937 , n17742 );
nor ( n17938 , n17937 , n17139 );
and ( n17939 , n17136 , n17938 );
nor ( n17940 , n17138 , n15344 );
nor ( n17941 , n17939 , n17940 );
buf ( n17942 , n17941 );
buf ( n17943 , n17942 );
nand ( n17944 , n874 , n17943 );
not ( n17945 , n1755 );
nor ( n17946 , n17945 , n1625 );
not ( n17947 , n17946 );
not ( n17948 , n17942 );
not ( n17949 , n860 );
and ( n17950 , n873 , n17949 );
not ( n17951 , n873 );
and ( n17952 , n17951 , n860 );
nor ( n17953 , n17950 , n17952 );
not ( n17954 , n1851 );
and ( n17955 , n1856 , n17954 );
not ( n17956 , n1856 );
and ( n17957 , n17956 , n1851 );
nor ( n17958 , n17955 , n17957 );
xor ( n17959 , n17953 , n17958 );
nand ( n17960 , n17948 , n17959 );
nand ( n17961 , n17944 , n17947 , n17960 );
not ( n17962 , n867 );
not ( n17963 , n17942 );
or ( n17964 , n17962 , n17963 );
and ( n17965 , n851 , n1862 );
not ( n17966 , n851 );
not ( n17967 , n1862 );
and ( n17968 , n17966 , n17967 );
nor ( n17969 , n17965 , n17968 );
or ( n17970 , n856 , n17969 );
nand ( n17971 , n856 , n17969 );
not ( n17972 , n17942 );
nand ( n17973 , n17970 , n17971 , n17972 );
nand ( n17974 , n17964 , n17947 , n17973 );
not ( n17975 , n866 );
not ( n17976 , n17942 );
or ( n17977 , n17975 , n17976 );
not ( n17978 , n861 );
and ( n17979 , n858 , n17978 );
not ( n17980 , n858 );
and ( n17981 , n17980 , n861 );
nor ( n17982 , n17979 , n17981 );
and ( n17983 , n1862 , n1870 );
not ( n17984 , n1862 );
not ( n17985 , n1870 );
and ( n17986 , n17984 , n17985 );
or ( n17987 , n17983 , n17986 );
and ( n17988 , n17987 , n856 );
not ( n17989 , n17987 );
not ( n17990 , n856 );
and ( n17991 , n17989 , n17990 );
nor ( n17992 , n17988 , n17991 );
or ( n17993 , n17982 , n17992 );
and ( n17994 , n17982 , n17992 );
nor ( n17995 , n17994 , n17942 );
nand ( n17996 , n17993 , n17995 );
nand ( n17997 , n17977 , n17947 , n17996 );
not ( n17998 , n12680 );
not ( n17999 , n12696 );
nor ( n18000 , n17998 , n17999 );
xor ( n18001 , n18000 , n12692 );
or ( n18002 , n16505 , n18001 );
and ( n18003 , n1228 , n949 , n16505 );
not ( n18004 , n141 );
and ( n18005 , n934 , n18004 );
and ( n18006 , n896 , n934 );
nor ( n18007 , n896 , n934 );
nor ( n18008 , n18006 , n18004 , n18007 );
nor ( n18009 , n18005 , n18008 );
not ( n18010 , n16502 );
nand ( n18011 , n12726 , n18010 );
nor ( n18012 , n18009 , n18011 , n16506 );
nor ( n18013 , n18003 , n18012 );
nand ( n18014 , n18002 , n18013 );
nand ( n18015 , n865 , n17943 );
and ( n18016 , n873 , n17978 );
not ( n18017 , n873 );
and ( n18018 , n18017 , n861 );
nor ( n18019 , n18016 , n18018 );
and ( n18020 , n1851 , n17985 );
and ( n18021 , n1870 , n17954 );
nor ( n18022 , n18020 , n18021 );
or ( n18023 , n18019 , n18022 );
and ( n18024 , n18019 , n18022 );
nor ( n18025 , n18024 , n17942 );
nand ( n18026 , n18023 , n18025 );
nand ( n18027 , n18015 , n17947 , n18026 );
nand ( n18028 , n13340 , n13377 );
not ( n18029 , n18028 );
not ( n18030 , n13724 );
or ( n18031 , n18029 , n18030 );
or ( n18032 , n18028 , n13724 );
nand ( n18033 , n18031 , n18032 );
not ( n18034 , n513 );
not ( n18035 , n14983 );
or ( n18036 , n18034 , n18035 );
not ( n18037 , n17314 );
not ( n18038 , n17291 );
nand ( n18039 , n17275 , n18038 );
not ( n18040 , n18039 );
nand ( n18041 , n18040 , n17269 , n17278 );
not ( n18042 , n17278 );
and ( n18043 , n17275 , n17285 );
nor ( n18044 , n18043 , n17301 );
or ( n18045 , n18042 , n18044 );
not ( n18046 , n17306 );
nand ( n18047 , n18045 , n18046 );
nand ( n18048 , n17269 , n18047 );
nand ( n18049 , n18037 , n18041 , n18048 );
or ( n18050 , n513 , n18049 );
nand ( n18051 , n513 , n18049 );
nand ( n18052 , n18050 , n18051 , n14982 );
nand ( n18053 , n18036 , n18052 );
and ( n18054 , n14974 , n18053 );
not ( n18055 , n513 );
not ( n18056 , n639 );
not ( n18057 , n540 );
nor ( n18058 , n541 , n542 );
nand ( n18059 , n18057 , n18058 );
nor ( n18060 , n571 , n539 , n18059 );
nand ( n18061 , n18056 , n18060 );
not ( n18062 , n18061 );
nand ( n18063 , n17877 , n17879 , n18062 );
not ( n18064 , n18063 );
or ( n18065 , n18055 , n18064 );
or ( n18066 , n513 , n18063 );
nand ( n18067 , n18065 , n18066 );
and ( n18068 , n1819 , n18067 );
nor ( n18069 , n18054 , n18068 );
nor ( n18070 , n14973 , n18069 );
not ( n18071 , n515 );
not ( n18072 , n16693 );
or ( n18073 , n18071 , n18072 );
not ( n18074 , n14989 );
nor ( n18075 , n18074 , n15059 );
or ( n18076 , n18075 , n15867 );
and ( n18077 , n18075 , n15867 );
not ( n18078 , n14980 );
nor ( n18079 , n18077 , n18078 );
nand ( n18080 , n18076 , n18079 );
nand ( n18081 , n18073 , n18080 );
and ( n18082 , n14974 , n18081 );
xor ( n18083 , n515 , n15891 );
and ( n18084 , n1819 , n18083 );
nor ( n18085 , n18082 , n18084 );
nor ( n18086 , n14973 , n18085 );
not ( n18087 , n601 );
not ( n18088 , n15713 );
or ( n18089 , n18087 , n18088 );
not ( n18090 , n17395 );
not ( n18091 , n17372 );
nand ( n18092 , n17356 , n18091 );
not ( n18093 , n18092 );
nand ( n18094 , n18093 , n17350 , n17359 );
not ( n18095 , n17359 );
and ( n18096 , n17356 , n17366 );
nor ( n18097 , n18096 , n17382 );
or ( n18098 , n18095 , n18097 );
not ( n18099 , n17387 );
nand ( n18100 , n18098 , n18099 );
nand ( n18101 , n17350 , n18100 );
nand ( n18102 , n18090 , n18094 , n18101 );
or ( n18103 , n601 , n18102 );
nand ( n18104 , n601 , n18102 );
nand ( n18105 , n18103 , n18104 , n15712 );
nand ( n18106 , n18089 , n18105 );
and ( n18107 , n15704 , n18106 );
not ( n18108 , n601 );
not ( n18109 , n717 );
not ( n18110 , n641 );
nor ( n18111 , n642 , n643 );
nand ( n18112 , n18110 , n18111 );
nor ( n18113 , n670 , n640 , n18112 );
nand ( n18114 , n18109 , n18113 );
not ( n18115 , n18114 );
nand ( n18116 , n17932 , n17928 , n18115 );
not ( n18117 , n18116 );
or ( n18118 , n18108 , n18117 );
or ( n18119 , n601 , n18116 );
nand ( n18120 , n18118 , n18119 );
and ( n18121 , n1808 , n18120 );
nor ( n18122 , n18107 , n18121 );
nor ( n18123 , n15703 , n18122 );
not ( n18124 , n610 );
not ( n18125 , n15876 );
or ( n18126 , n18124 , n18125 );
nor ( n18127 , n16922 , n17267 );
and ( n18128 , n18127 , n17870 );
and ( n18129 , n513 , n17848 );
nor ( n18130 , n18128 , n18129 );
nand ( n18131 , n18127 , n17850 );
not ( n18132 , n18131 );
not ( n18133 , n17852 );
nor ( n18134 , n18133 , n17860 );
nand ( n18135 , n18132 , n18134 );
and ( n18136 , n17852 , n17855 );
nor ( n18137 , n18136 , n17865 );
or ( n18138 , n18131 , n18137 );
nand ( n18139 , n18130 , n18135 , n18138 );
or ( n18140 , n610 , n18139 );
nand ( n18141 , n610 , n18139 );
nand ( n18142 , n18140 , n18141 , n14982 );
nand ( n18143 , n18126 , n18142 );
and ( n18144 , n14974 , n18143 );
nand ( n18145 , n17330 , n17331 , n18058 );
not ( n18146 , n18145 );
nand ( n18147 , n18146 , n17328 , n17879 );
and ( n18148 , n18147 , n16899 );
not ( n18149 , n18147 );
and ( n18150 , n18149 , n610 );
nor ( n18151 , n18148 , n18150 );
and ( n18152 , n1819 , n18151 );
nor ( n18153 , n18144 , n18152 );
nor ( n18154 , n14973 , n18153 );
not ( n18155 , n612 );
not ( n18156 , n17198 );
or ( n18157 , n18155 , n18156 );
not ( n18158 , n15728 );
nor ( n18159 , n18158 , n15722 );
or ( n18160 , n18159 , n15775 );
and ( n18161 , n18159 , n15775 );
not ( n18162 , n15709 );
nor ( n18163 , n18161 , n18162 );
nand ( n18164 , n18160 , n18163 );
nand ( n18165 , n18157 , n18164 );
and ( n18166 , n15704 , n18165 );
xor ( n18167 , n612 , n15798 );
and ( n18168 , n1808 , n18167 );
nor ( n18169 , n18166 , n18168 );
nor ( n18170 , n15703 , n18169 );
not ( n18171 , n681 );
not ( n18172 , n15100 );
or ( n18173 , n18171 , n18172 );
not ( n18174 , n17658 );
not ( n18175 , n17635 );
nand ( n18176 , n17619 , n18175 );
not ( n18177 , n18176 );
nand ( n18178 , n18177 , n17612 , n17622 );
not ( n18179 , n17622 );
and ( n18180 , n17619 , n17629 );
nor ( n18181 , n18180 , n17645 );
or ( n18182 , n18179 , n18181 );
not ( n18183 , n17650 );
nand ( n18184 , n18182 , n18183 );
nand ( n18185 , n17612 , n18184 );
nand ( n18186 , n18174 , n18178 , n18185 );
or ( n18187 , n681 , n18186 );
nand ( n18188 , n681 , n18186 );
nand ( n18189 , n18187 , n18188 , n15099 );
nand ( n18190 , n18173 , n18189 );
and ( n18191 , n15090 , n18190 );
not ( n18192 , n681 );
not ( n18193 , n784 );
not ( n18194 , n718 );
nor ( n18195 , n719 , n720 );
nand ( n18196 , n18194 , n18195 );
nor ( n18197 , n756 , n723 , n18196 );
nand ( n18198 , n18193 , n18197 );
not ( n18199 , n18198 );
nand ( n18200 , n17787 , n17783 , n18199 );
not ( n18201 , n18200 );
or ( n18202 , n18192 , n18201 );
or ( n18203 , n681 , n18200 );
nand ( n18204 , n18202 , n18203 );
and ( n18205 , n1826 , n18204 );
nor ( n18206 , n18191 , n18205 );
nor ( n18207 , n15089 , n18206 );
not ( n18208 , n693 );
not ( n18209 , n16394 );
or ( n18210 , n18208 , n18209 );
nor ( n18211 , n16993 , n17349 );
and ( n18212 , n18211 , n17921 );
and ( n18213 , n601 , n17899 );
nor ( n18214 , n18212 , n18213 );
nand ( n18215 , n18211 , n17901 );
not ( n18216 , n18215 );
not ( n18217 , n17903 );
nor ( n18218 , n18217 , n17911 );
nand ( n18219 , n18216 , n18218 );
and ( n18220 , n17903 , n17906 );
nor ( n18221 , n18220 , n17916 );
or ( n18222 , n18215 , n18221 );
nand ( n18223 , n18214 , n18219 , n18222 );
or ( n18224 , n693 , n18223 );
nand ( n18225 , n693 , n18223 );
nand ( n18226 , n18224 , n18225 , n15712 );
nand ( n18227 , n18210 , n18226 );
and ( n18228 , n15704 , n18227 );
nand ( n18229 , n17412 , n18111 , n17411 );
not ( n18230 , n18229 );
nand ( n18231 , n18230 , n17409 , n17928 );
and ( n18232 , n18231 , n16970 );
not ( n18233 , n18231 );
and ( n18234 , n18233 , n693 );
nor ( n18235 , n18232 , n18234 );
and ( n18236 , n1808 , n18235 );
nor ( n18237 , n18228 , n18236 );
nor ( n18238 , n15703 , n18237 );
not ( n18239 , n695 );
not ( n18240 , n17667 );
or ( n18241 , n18239 , n18240 );
not ( n18242 , n15106 );
nor ( n18243 , n18242 , n15175 );
or ( n18244 , n18243 , n15821 );
and ( n18245 , n18243 , n15821 );
nor ( n18246 , n18245 , n15829 );
nand ( n18247 , n18244 , n18246 );
nand ( n18248 , n18241 , n18247 );
and ( n18249 , n15090 , n18248 );
xor ( n18250 , n695 , n15844 );
and ( n18251 , n1826 , n18250 );
nor ( n18252 , n18249 , n18251 );
nor ( n18253 , n15089 , n18252 );
not ( n18254 , n778 );
not ( n18255 , n15831 );
or ( n18256 , n18254 , n18255 );
nor ( n18257 , n17063 , n17611 );
and ( n18258 , n18257 , n17776 );
and ( n18259 , n681 , n17754 );
nor ( n18260 , n18258 , n18259 );
nand ( n18261 , n18257 , n17756 );
not ( n18262 , n18261 );
not ( n18263 , n17758 );
nor ( n18264 , n18263 , n17766 );
nand ( n18265 , n18262 , n18264 );
and ( n18266 , n17758 , n17761 );
nor ( n18267 , n18266 , n17771 );
or ( n18268 , n18261 , n18267 );
nand ( n18269 , n18260 , n18265 , n18268 );
or ( n18270 , n778 , n18269 );
nand ( n18271 , n778 , n18269 );
nand ( n18272 , n18270 , n18271 , n15830 );
nand ( n18273 , n18256 , n18272 );
and ( n18274 , n15090 , n18273 );
nand ( n18275 , n17676 , n18195 , n17675 );
not ( n18276 , n18275 );
nand ( n18277 , n18276 , n17783 , n17673 );
and ( n18278 , n18277 , n17041 );
not ( n18279 , n18277 );
and ( n18280 , n18279 , n778 );
nor ( n18281 , n18278 , n18280 );
and ( n18282 , n1826 , n18281 );
nor ( n18283 , n18274 , n18282 );
nor ( n18284 , n15089 , n18283 );
not ( n18285 , n792 );
not ( n18286 , n16270 );
or ( n18287 , n18285 , n18286 );
not ( n18288 , n17579 );
not ( n18289 , n17556 );
nand ( n18290 , n17540 , n18289 );
not ( n18291 , n18290 );
nand ( n18292 , n18291 , n17543 , n17534 );
not ( n18293 , n17543 );
and ( n18294 , n17540 , n17550 );
nor ( n18295 , n18294 , n17566 );
or ( n18296 , n18293 , n18295 );
not ( n18297 , n17571 );
nand ( n18298 , n18296 , n18297 );
nand ( n18299 , n17534 , n18298 );
nand ( n18300 , n18288 , n18292 , n18299 );
or ( n18301 , n792 , n18300 );
nand ( n18302 , n792 , n18300 );
nand ( n18303 , n18301 , n18302 , n16269 );
nand ( n18304 , n18287 , n18303 );
and ( n18305 , n16258 , n18304 );
not ( n18306 , n792 );
not ( n18307 , n827 );
nor ( n18308 , n798 , n828 );
nand ( n18309 , n18307 , n18308 );
nor ( n18310 , n839 , n829 , n18309 );
nand ( n18311 , n17594 , n18310 );
not ( n18312 , n18311 );
nand ( n18313 , n17721 , n17723 , n18312 );
not ( n18314 , n18313 );
or ( n18315 , n18306 , n18314 );
or ( n18316 , n792 , n18313 );
nand ( n18317 , n18315 , n18316 );
and ( n18318 , n1828 , n18317 );
nor ( n18319 , n18305 , n18318 );
nor ( n18320 , n16257 , n18319 );
not ( n18321 , n804 );
not ( n18322 , n16748 );
or ( n18323 , n18321 , n18322 );
not ( n18324 , n16293 );
nor ( n18325 , n18324 , n16339 );
or ( n18326 , n18325 , n16423 );
and ( n18327 , n18325 , n16423 );
nor ( n18328 , n18327 , n16747 );
nand ( n18329 , n18326 , n18328 );
nand ( n18330 , n18323 , n18329 );
and ( n18331 , n16258 , n18330 );
xor ( n18332 , n804 , n16444 );
and ( n18333 , n1828 , n18332 );
nor ( n18334 , n18331 , n18333 );
nor ( n18335 , n16257 , n18334 );
not ( n18336 , n844 );
not ( n18337 , n16349 );
or ( n18338 , n18336 , n18337 );
nor ( n18339 , n16851 , n17532 );
and ( n18340 , n18339 , n17714 );
and ( n18341 , n792 , n17692 );
nor ( n18342 , n18340 , n18341 );
nand ( n18343 , n18339 , n17694 );
not ( n18344 , n18343 );
not ( n18345 , n17696 );
nor ( n18346 , n18345 , n17704 );
nand ( n18347 , n18344 , n18346 );
and ( n18348 , n17696 , n17699 );
nor ( n18349 , n18348 , n17709 );
or ( n18350 , n18343 , n18349 );
nand ( n18351 , n18342 , n18347 , n18350 );
or ( n18352 , n844 , n18351 );
nand ( n18353 , n844 , n18351 );
nand ( n18354 , n18352 , n18353 , n16348 );
nand ( n18355 , n18338 , n18354 );
and ( n18356 , n16258 , n18355 );
nand ( n18357 , n17596 , n18308 , n17595 );
not ( n18358 , n18357 );
nand ( n18359 , n18358 , n17592 , n17723 );
and ( n18360 , n18359 , n16826 );
not ( n18361 , n18359 );
and ( n18362 , n18361 , n844 );
nor ( n18363 , n18360 , n18362 );
and ( n18364 , n1828 , n18363 );
nor ( n18365 , n18356 , n18364 );
nor ( n18366 , n16257 , n18365 );
nand ( n18367 , n851 , n17943 );
not ( n18368 , n852 );
not ( n18369 , n18368 );
not ( n18370 , n859 );
and ( n18371 , n18369 , n18370 );
and ( n18372 , n859 , n18368 );
nor ( n18373 , n18371 , n18372 );
and ( n18374 , n18373 , n17962 );
not ( n18375 , n18373 );
and ( n18376 , n18375 , n867 );
nor ( n18377 , n18374 , n18376 );
and ( n18378 , n1864 , n1869 );
not ( n18379 , n1864 );
not ( n18380 , n1869 );
and ( n18381 , n18379 , n18380 );
nor ( n18382 , n18378 , n18381 );
not ( n18383 , n18382 );
and ( n18384 , n1867 , n18383 );
not ( n18385 , n1867 );
and ( n18386 , n18385 , n18382 );
nor ( n18387 , n18384 , n18386 );
and ( n18388 , n18377 , n18387 );
nor ( n18389 , n18387 , n18377 );
nor ( n18390 , n18388 , n18389 );
not ( n18391 , n17958 );
and ( n18392 , n17987 , n18391 );
not ( n18393 , n17987 );
and ( n18394 , n18393 , n17958 );
nor ( n18395 , n18392 , n18394 );
not ( n18396 , n18395 );
or ( n18397 , n17990 , n861 );
or ( n18398 , n17978 , n856 );
nand ( n18399 , n18397 , n18398 );
not ( n18400 , n18399 );
not ( n18401 , n17953 );
or ( n18402 , n18400 , n18401 );
or ( n18403 , n17953 , n18399 );
nand ( n18404 , n18402 , n18403 );
not ( n18405 , n18404 );
and ( n18406 , n18396 , n18405 );
and ( n18407 , n18404 , n18395 );
nor ( n18408 , n18406 , n18407 );
or ( n18409 , n18390 , n18408 );
and ( n18410 , n18390 , n18408 );
nor ( n18411 , n17942 , n18410 );
nand ( n18412 , n18409 , n18411 );
nand ( n18413 , n18367 , n17947 , n18412 );
or ( n18414 , n17990 , n17963 );
and ( n18415 , n865 , n866 );
not ( n18416 , n865 );
and ( n18417 , n18416 , n17975 );
nor ( n18418 , n18415 , n18417 );
and ( n18419 , n1854 , n1867 );
not ( n18420 , n1854 );
and ( n18421 , n18420 , n18385 );
nor ( n18422 , n18419 , n18421 );
xor ( n18423 , n18418 , n18422 );
and ( n18424 , n18383 , n18391 );
not ( n18425 , n18383 );
and ( n18426 , n18425 , n17958 );
nor ( n18427 , n18424 , n18426 );
and ( n18428 , n18423 , n18427 );
nor ( n18429 , n18427 , n18423 );
nor ( n18430 , n18428 , n18429 );
and ( n18431 , n859 , n867 );
not ( n18432 , n859 );
and ( n18433 , n18432 , n17962 );
or ( n18434 , n18431 , n18433 );
and ( n18435 , n860 , n18368 );
not ( n18436 , n860 );
and ( n18437 , n18436 , n852 );
nor ( n18438 , n18435 , n18437 );
xnor ( n18439 , n18434 , n18438 );
not ( n18440 , n18439 );
xor ( n18441 , n17992 , n18019 );
not ( n18442 , n18441 );
and ( n18443 , n18440 , n18442 );
and ( n18444 , n18439 , n18441 );
nor ( n18445 , n18443 , n18444 );
or ( n18446 , n18430 , n18445 );
and ( n18447 , n18430 , n18445 );
nor ( n18448 , n17942 , n18447 );
nand ( n18449 , n18446 , n18448 );
nand ( n18450 , n18414 , n17947 , n18449 );
nand ( n18451 , n858 , n17943 );
not ( n18452 , n18373 );
not ( n18453 , n18382 );
and ( n18454 , n18452 , n18453 );
and ( n18455 , n18382 , n18373 );
nor ( n18456 , n18454 , n18455 );
and ( n18457 , n866 , n17962 );
and ( n18458 , n867 , n17975 );
nor ( n18459 , n18457 , n18458 );
not ( n18460 , n18459 );
not ( n18461 , n18422 );
and ( n18462 , n18460 , n18461 );
and ( n18463 , n18422 , n18459 );
nor ( n18464 , n18462 , n18463 );
xnor ( n18465 , n18456 , n18464 );
or ( n18466 , n18465 , n18408 );
and ( n18467 , n18465 , n18408 );
nor ( n18468 , n17942 , n18467 );
nand ( n18469 , n18466 , n18468 );
nand ( n18470 , n18451 , n17947 , n18469 );
nand ( n18471 , n862 , n17943 );
and ( n18472 , n1864 , n18385 );
not ( n18473 , n1864 );
and ( n18474 , n1867 , n18473 );
nor ( n18475 , n18472 , n18474 );
or ( n18476 , n18434 , n18475 );
and ( n18477 , n18434 , n18475 );
nor ( n18478 , n18477 , n17942 );
nand ( n18479 , n18476 , n18478 );
nand ( n18480 , n18471 , n17947 , n18479 );
nand ( n18481 , n864 , n17943 );
and ( n18482 , n1856 , n18380 );
not ( n18483 , n1856 );
and ( n18484 , n1869 , n18483 );
nor ( n18485 , n18482 , n18484 );
or ( n18486 , n18438 , n18485 );
and ( n18487 , n18438 , n18485 );
nor ( n18488 , n18487 , n17942 );
nand ( n18489 , n18486 , n18488 );
nand ( n18490 , n18481 , n17947 , n18489 );
not ( n18491 , n17963 );
or ( n18492 , n18385 , n18491 );
not ( n18493 , n17972 );
nand ( n18494 , n1052 , n18493 );
nand ( n18495 , n18492 , n18494 );
or ( n18496 , n516 , n15889 );
nand ( n18497 , n18496 , n1819 , n15890 );
nor ( n18498 , n15052 , n15875 );
or ( n18499 , n14994 , n15053 );
nor ( n18500 , n17429 , n17436 );
and ( n18501 , n18499 , n18500 );
or ( n18502 , n18499 , n18500 );
nand ( n18503 , n18502 , n15874 );
nor ( n18504 , n18501 , n18503 );
or ( n18505 , n18498 , n18504 );
nand ( n18506 , n18505 , n14974 );
and ( n18507 , n18497 , n18506 );
nor ( n18508 , n18507 , n14973 );
not ( n18509 , n517 );
not ( n18510 , n16693 );
or ( n18511 , n18509 , n18510 );
not ( n18512 , n17305 );
nor ( n18513 , n18512 , n17276 );
not ( n18514 , n18134 );
nand ( n18515 , n18514 , n18137 );
or ( n18516 , n18513 , n18515 );
and ( n18517 , n18513 , n18515 );
nor ( n18518 , n18517 , n18078 );
nand ( n18519 , n18516 , n18518 );
nand ( n18520 , n18511 , n18519 );
and ( n18521 , n14974 , n18520 );
and ( n18522 , n18145 , n17329 );
not ( n18523 , n18145 );
and ( n18524 , n18523 , n517 );
nor ( n18525 , n18522 , n18524 );
and ( n18526 , n1819 , n18525 );
nor ( n18527 , n18521 , n18526 );
nor ( n18528 , n14973 , n18527 );
not ( n18529 , n609 );
not ( n18530 , n15876 );
or ( n18531 , n18529 , n18530 );
and ( n18532 , n14997 , n15049 );
nand ( n18533 , n15016 , n15043 );
or ( n18534 , n18532 , n18533 );
and ( n18535 , n18532 , n18533 );
not ( n18536 , n15874 );
nor ( n18537 , n18535 , n18536 );
nand ( n18538 , n18534 , n18537 );
nand ( n18539 , n18531 , n18538 );
and ( n18540 , n14974 , n18539 );
not ( n18541 , n609 );
not ( n18542 , n15079 );
or ( n18543 , n18541 , n18542 );
or ( n18544 , n609 , n15079 );
nand ( n18545 , n18543 , n18544 );
and ( n18546 , n1819 , n18545 );
nor ( n18547 , n18540 , n18546 );
nor ( n18548 , n14973 , n18547 );
not ( n18549 , n615 );
not ( n18550 , n17198 );
or ( n18551 , n18549 , n18550 );
not ( n18552 , n17386 );
nor ( n18553 , n18552 , n17357 );
not ( n18554 , n18218 );
nand ( n18555 , n18554 , n18221 );
or ( n18556 , n18553 , n18555 );
and ( n18557 , n18553 , n18555 );
nor ( n18558 , n18557 , n18162 );
nand ( n18559 , n18556 , n18558 );
nand ( n18560 , n18551 , n18559 );
and ( n18561 , n15704 , n18560 );
and ( n18562 , n18229 , n17410 );
not ( n18563 , n18229 );
and ( n18564 , n18563 , n615 );
nor ( n18565 , n18562 , n18564 );
and ( n18566 , n1808 , n18565 );
nor ( n18567 , n18561 , n18566 );
nor ( n18568 , n15703 , n18567 );
not ( n18569 , n678 );
not ( n18570 , n16394 );
or ( n18571 , n18569 , n18570 );
not ( n18572 , n15771 );
and ( n18573 , n15742 , n18572 );
or ( n18574 , n16374 , n16382 );
or ( n18575 , n18573 , n18574 );
and ( n18576 , n18573 , n18574 );
nor ( n18577 , n18576 , n18162 );
nand ( n18578 , n18575 , n18577 );
nand ( n18579 , n18571 , n18578 );
and ( n18580 , n15704 , n18579 );
xor ( n18581 , n678 , n16403 );
and ( n18582 , n1808 , n18581 );
nor ( n18583 , n18580 , n18582 );
nor ( n18584 , n15703 , n18583 );
not ( n18585 , n697 );
not ( n18586 , n17667 );
or ( n18587 , n18585 , n18586 );
not ( n18588 , n17649 );
nor ( n18589 , n18588 , n17621 );
not ( n18590 , n18264 );
nand ( n18591 , n18590 , n18267 );
or ( n18592 , n18589 , n18591 );
and ( n18593 , n18589 , n18591 );
nor ( n18594 , n18593 , n15829 );
nand ( n18595 , n18592 , n18594 );
nand ( n18596 , n18587 , n18595 );
and ( n18597 , n15090 , n18596 );
and ( n18598 , n18275 , n17674 );
not ( n18599 , n18275 );
and ( n18600 , n18599 , n697 );
nor ( n18601 , n18598 , n18600 );
and ( n18602 , n1826 , n18601 );
nor ( n18603 , n18597 , n18602 );
nor ( n18604 , n15089 , n18603 );
or ( n18605 , n698 , n15842 );
nand ( n18606 , n18605 , n1826 , n15843 );
nor ( n18607 , n15168 , n15099 );
or ( n18608 , n15111 , n15169 );
not ( n18609 , n17464 );
nor ( n18610 , n18609 , n17471 );
and ( n18611 , n18608 , n18610 );
or ( n18612 , n18608 , n18610 );
nand ( n18613 , n18612 , n15830 );
nor ( n18614 , n18611 , n18613 );
or ( n18615 , n18607 , n18614 );
nand ( n18616 , n18615 , n15090 );
and ( n18617 , n18606 , n18616 );
nor ( n18618 , n18617 , n15089 );
and ( n18619 , n2 , n15231 , n15236 , n15264 );
not ( n18620 , n777 );
not ( n18621 , n17667 );
or ( n18622 , n18620 , n18621 );
and ( n18623 , n15114 , n15165 );
nand ( n18624 , n15132 , n15159 );
or ( n18625 , n18623 , n18624 );
and ( n18626 , n18623 , n18624 );
not ( n18627 , n15828 );
nor ( n18628 , n18626 , n18627 );
nand ( n18629 , n18625 , n18628 );
nand ( n18630 , n18622 , n18629 );
and ( n18631 , n15090 , n18630 );
xor ( n18632 , n777 , n15194 );
and ( n18633 , n1826 , n18632 );
nor ( n18634 , n18631 , n18633 );
nor ( n18635 , n15089 , n18634 );
not ( n18636 , n808 );
not ( n18637 , n16748 );
or ( n18638 , n18636 , n18637 );
not ( n18639 , n17570 );
nor ( n18640 , n18639 , n17542 );
not ( n18641 , n18346 );
nand ( n18642 , n18641 , n18349 );
or ( n18643 , n18640 , n18642 );
and ( n18644 , n18640 , n18642 );
nor ( n18645 , n18644 , n16267 );
nand ( n18646 , n18643 , n18645 );
nand ( n18647 , n18638 , n18646 );
and ( n18648 , n16258 , n18647 );
and ( n18649 , n18357 , n17593 );
not ( n18650 , n18357 );
and ( n18651 , n18650 , n808 );
nor ( n18652 , n18649 , n18651 );
and ( n18653 , n1828 , n18652 );
nor ( n18654 , n18648 , n18653 );
nor ( n18655 , n16257 , n18654 );
nor ( n18656 , n15342 , n17945 );
and ( n18657 , n18656 , n17145 );
not ( n18658 , n18656 );
not ( n18659 , n17148 );
and ( n18660 , n18658 , n18659 );
or ( n18661 , n825 , n17147 );
nand ( n18662 , n18661 , n17158 );
nor ( n18663 , n18660 , n18662 );
nor ( n18664 , n18657 , n18663 );
not ( n18665 , n15342 );
not ( n18666 , n17133 );
or ( n18667 , n18665 , n18666 );
not ( n18668 , n17155 );
nor ( n18669 , n17154 , n511 , n18668 );
nand ( n18670 , n18667 , n18669 );
or ( n18671 , n18656 , n17736 );
or ( n18672 , n825 , n17127 );
not ( n18673 , n17938 );
nor ( n18674 , n17136 , n18673 );
nand ( n18675 , n18671 , n18672 , n18674 );
and ( n18676 , n18664 , n18670 , n18675 );
not ( n18677 , n2 );
nor ( n18678 , n18676 , n18677 );
not ( n18679 , n2 );
or ( n18680 , n15247 , n15244 );
nand ( n18681 , n18680 , n15240 );
nor ( n18682 , n3 , n15243 );
not ( n18683 , n18682 );
not ( n18684 , n15239 );
nor ( n18685 , n3 , n18684 );
nor ( n18686 , n18685 , n15253 );
and ( n18687 , n18681 , n18683 , n18686 );
not ( n18688 , n15259 );
and ( n18689 , n845 , n18688 );
nor ( n18690 , n18687 , n18689 );
nor ( n18691 , n18679 , n18690 );
not ( n18692 , n2 );
not ( n18693 , n17942 );
and ( n18694 , n1046 , n18693 );
and ( n18695 , n918 , n16533 );
nor ( n18696 , n18694 , n18695 );
nor ( n18697 , n18692 , n18696 );
or ( n18698 , n18380 , n18491 );
not ( n18699 , n17972 );
nand ( n18700 , n1016 , n18699 );
nand ( n18701 , n18698 , n18700 );
or ( n18702 , n17985 , n18491 );
nand ( n18703 , n1018 , n18493 );
nand ( n18704 , n18702 , n18703 );
not ( n18705 , n17963 );
or ( n18706 , n18483 , n18705 );
nand ( n18707 , n1019 , n18699 );
nand ( n18708 , n18706 , n18707 );
or ( n18709 , n17967 , n18705 );
nand ( n18710 , n1047 , n18699 );
nand ( n18711 , n18709 , n18710 );
or ( n18712 , n17954 , n18705 );
nand ( n18713 , n1049 , n18699 );
nand ( n18714 , n18712 , n18713 );
or ( n18715 , n18473 , n18705 );
nand ( n18716 , n1051 , n18493 );
nand ( n18717 , n18715 , n18716 );
not ( n18718 , n16833 );
nand ( n18719 , n18718 , n16834 );
not ( n18720 , n18719 );
not ( n18721 , n16892 );
nand ( n18722 , n18721 , n16845 );
not ( n18723 , n18722 );
or ( n18724 , n18720 , n18723 );
or ( n18725 , n18719 , n18722 );
nand ( n18726 , n18724 , n18725 );
not ( n18727 , n16919 );
nand ( n18728 , n18727 , n16909 );
not ( n18729 , n18728 );
not ( n18730 , n16963 );
nand ( n18731 , n18730 , n16916 );
not ( n18732 , n18731 );
or ( n18733 , n18729 , n18732 );
or ( n18734 , n18728 , n18731 );
nand ( n18735 , n18733 , n18734 );
not ( n18736 , n16990 );
nand ( n18737 , n18736 , n16980 );
not ( n18738 , n18737 );
not ( n18739 , n17034 );
nand ( n18740 , n18739 , n16987 );
not ( n18741 , n18740 );
or ( n18742 , n18738 , n18741 );
or ( n18743 , n18737 , n18740 );
nand ( n18744 , n18742 , n18743 );
not ( n18745 , n17048 );
nand ( n18746 , n18745 , n17049 );
not ( n18747 , n18746 );
not ( n18748 , n17104 );
nand ( n18749 , n18748 , n17057 );
not ( n18750 , n18749 );
or ( n18751 , n18747 , n18750 );
or ( n18752 , n18746 , n18749 );
nand ( n18753 , n18751 , n18752 );
not ( n18754 , n1854 );
or ( n18755 , n18754 , n18491 );
nand ( n18756 , n1053 , n18493 );
nand ( n18757 , n18755 , n18756 );
not ( n18758 , n1051 );
not ( n18759 , n17942 );
not ( n18760 , n18759 );
or ( n18761 , n18758 , n18760 );
buf ( n18762 , n17942 );
nand ( n18763 , n1057 , n18762 );
nand ( n18764 , n18761 , n18763 );
not ( n18765 , n1019 );
not ( n18766 , n18759 );
or ( n18767 , n18765 , n18766 );
nand ( n18768 , n1056 , n18762 );
nand ( n18769 , n18767 , n18768 );
not ( n18770 , n1049 );
not ( n18771 , n18759 );
or ( n18772 , n18770 , n18771 );
buf ( n18773 , n17942 );
nand ( n18774 , n1055 , n18773 );
nand ( n18775 , n18772 , n18774 );
not ( n18776 , n1018 );
not ( n18777 , n17976 );
or ( n18778 , n18776 , n18777 );
nand ( n18779 , n1054 , n18773 );
nand ( n18780 , n18778 , n18779 );
nand ( n18781 , n1046 , n16533 );
and ( n18782 , n18781 , n18491 );
not ( n18783 , n2 );
nor ( n18784 , n18782 , n18783 );
not ( n18785 , n1016 );
not ( n18786 , n17976 );
or ( n18787 , n18785 , n18786 );
nand ( n18788 , n1013 , n18773 );
nand ( n18789 , n18787 , n18788 );
not ( n18790 , n1047 );
not ( n18791 , n17976 );
or ( n18792 , n18790 , n18791 );
nand ( n18793 , n1010 , n18773 );
nand ( n18794 , n18792 , n18793 );
and ( n18795 , n560 , n13633 );
and ( n18796 , n484 , n13623 );
nor ( n18797 , n18795 , n18796 );
nand ( n18798 , n484 , n560 );
and ( n18799 , n18797 , n18798 , n13690 );
not ( n18800 , n347 );
nand ( n18801 , n18800 , n1006 );
not ( n18802 , n888 );
nand ( n18803 , n18802 , n482 );
not ( n18804 , n939 );
nand ( n18805 , n18804 , n409 );
nand ( n18806 , n409 , n482 );
not ( n18807 , n13620 );
nand ( n18808 , n18803 , n18805 , n18806 , n18807 );
nand ( n18809 , n18801 , n18808 );
nor ( n18810 , n18799 , n18809 );
not ( n18811 , n329 );
not ( n18812 , n939 );
not ( n18813 , n18806 );
and ( n18814 , n18812 , n18813 );
not ( n18815 , n888 );
and ( n18816 , n409 , n18815 );
nor ( n18817 , n18814 , n18816 );
nand ( n18818 , n13633 , n484 , n18808 );
not ( n18819 , n560 );
or ( n18820 , n18819 , n13690 );
or ( n18821 , n937 , n18798 );
nand ( n18822 , n18820 , n18821 );
and ( n18823 , n18822 , n18808 );
and ( n18824 , n482 , n13620 );
nor ( n18825 , n18823 , n18824 );
nand ( n18826 , n18817 , n18818 , n18825 );
and ( n18827 , n18801 , n18826 );
and ( n18828 , n347 , n12538 );
nor ( n18829 , n18827 , n18828 );
nor ( n18830 , n215 , n410 );
nand ( n18831 , n18811 , n18829 , n18830 );
or ( n18832 , n18810 , n18831 );
not ( n18833 , n13683 );
and ( n18834 , n749 , n18833 );
not ( n18835 , n884 );
and ( n18836 , n462 , n18835 );
nor ( n18837 , n18834 , n18836 );
nand ( n18838 , n462 , n749 );
not ( n18839 , n18838 );
and ( n18840 , n13675 , n18839 );
and ( n18841 , n462 , n13675 );
and ( n18842 , n749 , n18835 );
nor ( n18843 , n18841 , n18842 );
and ( n18844 , n18843 , n18838 , n13683 );
not ( n18845 , n802 );
or ( n18846 , n18845 , n13668 );
nand ( n18847 , n674 , n802 );
or ( n18848 , n933 , n18847 );
not ( n18849 , n674 );
or ( n18850 , n18849 , n935 );
nand ( n18851 , n18846 , n18848 , n18850 );
and ( n18852 , n802 , n13660 );
and ( n18853 , n674 , n13664 );
nor ( n18854 , n18852 , n18853 );
and ( n18855 , n18854 , n18847 , n13668 );
not ( n18856 , n855 );
nand ( n18857 , n18856 , n879 );
and ( n18858 , n1487 , n18857 );
and ( n18859 , n855 , n13643 );
nor ( n18860 , n18858 , n18859 , n13641 );
nor ( n18861 , n18855 , n18860 );
nor ( n18862 , n18851 , n18861 );
nor ( n18863 , n18844 , n18862 );
nor ( n18864 , n18840 , n18863 , n18831 );
nand ( n18865 , n18837 , n18864 );
nand ( n18866 , n18832 , n18865 );
or ( n18867 , n18464 , n18705 );
and ( n18868 , n875 , n17942 );
nor ( n18869 , n18868 , n17946 );
nand ( n18870 , n18867 , n18869 );
not ( n18871 , n613 );
not ( n18872 , n18536 );
or ( n18873 , n18871 , n18872 );
nor ( n18874 , n15036 , n16679 );
or ( n18875 , n18874 , n16676 );
and ( n18876 , n18874 , n16676 );
nor ( n18877 , n18876 , n14979 );
nand ( n18878 , n18875 , n18877 );
nand ( n18879 , n18873 , n18878 );
and ( n18880 , n14974 , n18879 );
not ( n18881 , n613 );
not ( n18882 , n15888 );
or ( n18883 , n18881 , n18882 );
or ( n18884 , n613 , n15888 );
nand ( n18885 , n18883 , n18884 );
and ( n18886 , n1819 , n18885 );
nor ( n18887 , n18880 , n18886 );
nor ( n18888 , n14973 , n18887 );
nand ( n18889 , n14478 , n14484 );
not ( n18890 , n18889 );
not ( n18891 , n14501 );
or ( n18892 , n18890 , n18891 );
or ( n18893 , n18889 , n14501 );
nand ( n18894 , n18892 , n18893 );
and ( n18895 , n15247 , n15256 );
nand ( n18896 , n1530 , n15249 , n18895 );
not ( n18897 , n15257 );
not ( n18898 , n15261 );
or ( n18899 , n18897 , n18898 );
or ( n18900 , n806 , n15235 );
nand ( n18901 , n18899 , n18900 );
and ( n18902 , n18896 , n18901 );
not ( n18903 , n2 );
nor ( n18904 , n18902 , n18903 );
or ( n18905 , n807 , n16442 );
nand ( n18906 , n18905 , n1828 , n16443 );
nor ( n18907 , n16332 , n16269 );
or ( n18908 , n16301 , n16333 );
nor ( n18909 , n17499 , n17507 );
and ( n18910 , n18908 , n18909 );
or ( n18911 , n18908 , n18909 );
nand ( n18912 , n18911 , n16268 );
nor ( n18913 , n18910 , n18912 );
or ( n18914 , n18907 , n18913 );
nand ( n18915 , n18914 , n16258 );
and ( n18916 , n18906 , n18915 );
nor ( n18917 , n18916 , n16257 );
and ( n18918 , n824 , n17133 , n18669 );
and ( n18919 , n15344 , n17156 );
and ( n18920 , n17154 , n17148 );
nand ( n18921 , n1755 , n17154 );
not ( n18922 , n18921 );
and ( n18923 , n17147 , n18922 );
nor ( n18924 , n18919 , n18920 , n18923 );
nor ( n18925 , n18918 , n18924 );
not ( n18926 , n2 );
not ( n18927 , n17156 );
and ( n18928 , n17134 , n18927 );
nor ( n18929 , n18926 , n18928 );
nand ( n18930 , n18921 , n17145 );
or ( n18931 , n18921 , n17736 );
or ( n18932 , n824 , n17127 );
nand ( n18933 , n18931 , n18932 , n18674 );
nand ( n18934 , n18925 , n18929 , n18930 , n18933 );
not ( n18935 , n843 );
not ( n18936 , n16349 );
or ( n18937 , n18935 , n18936 );
nand ( n18938 , n16298 , n16329 );
nor ( n18939 , n16291 , n16324 );
or ( n18940 , n18938 , n18939 );
nand ( n18941 , n18938 , n18939 );
nand ( n18942 , n18940 , n18941 , n16348 );
nand ( n18943 , n18937 , n18942 );
and ( n18944 , n16258 , n18943 );
xor ( n18945 , n843 , n16362 );
and ( n18946 , n1828 , n18945 );
nor ( n18947 , n18944 , n18946 );
nor ( n18948 , n16257 , n18947 );
not ( n18949 , n1395 );
and ( n18950 , n774 , n18949 );
and ( n18951 , n750 , n17043 );
nor ( n18952 , n18950 , n18951 );
nand ( n18953 , n750 , n774 );
nand ( n18954 , n17043 , n18949 );
nand ( n18955 , n18952 , n18953 , n18954 );
or ( n18956 , n15107 , n1186 );
and ( n18957 , n487 , n17047 );
nor ( n18958 , n1185 , n1186 );
nor ( n18959 , n18957 , n18958 );
nand ( n18960 , n18956 , n15837 , n18959 );
nand ( n18961 , n18955 , n18960 );
and ( n18962 , n695 , n17051 );
not ( n18963 , n698 );
not ( n18964 , n17051 );
or ( n18965 , n18963 , n18964 );
nand ( n18966 , n18965 , n15189 );
and ( n18967 , n17053 , n18966 );
not ( n18968 , n695 );
nand ( n18969 , n18968 , n1348 );
nand ( n18970 , n17053 , n18969 );
not ( n18971 , n18966 );
nand ( n18972 , n18970 , n18971 );
nand ( n18973 , n17067 , n777 , n18972 );
and ( n18974 , n777 , n17098 );
nor ( n18975 , n1195 , n1346 );
nor ( n18976 , n18974 , n18975 );
not ( n18977 , n18976 );
nand ( n18978 , n779 , n18977 , n18972 );
nand ( n18979 , n18973 , n18978 );
nor ( n18980 , n18962 , n18967 , n18979 );
or ( n18981 , n18961 , n18980 );
not ( n18982 , n1273 );
nor ( n18983 , n18982 , n1388 );
not ( n18984 , n18961 );
or ( n18985 , n1344 , n15192 );
nor ( n18986 , n1344 , n1345 );
and ( n18987 , n782 , n18986 );
and ( n18988 , n783 , n17072 );
nor ( n18989 , n18987 , n18988 );
or ( n18990 , n17078 , n791 );
and ( n18991 , n782 , n17072 );
and ( n18992 , n783 , n17075 );
nor ( n18993 , n18991 , n18992 );
not ( n18994 , n18986 );
and ( n18995 , n18993 , n15192 , n18994 );
and ( n18996 , n791 , n17078 );
nand ( n18997 , n1342 , n15124 );
nor ( n18998 , n18996 , n18997 );
nor ( n18999 , n18995 , n18998 );
nand ( n19000 , n18990 , n18999 );
nand ( n19001 , n18985 , n18989 , n19000 );
or ( n19002 , n15191 , n1346 );
nand ( n19003 , n19002 , n15839 , n18976 );
nand ( n19004 , n18984 , n19001 , n19003 , n18972 );
nand ( n19005 , n18981 , n18983 , n19004 );
or ( n19006 , n1361 , n18953 );
or ( n19007 , n15811 , n1395 );
not ( n19008 , n18959 );
and ( n19009 , n752 , n19008 , n18955 );
not ( n19010 , n18955 );
or ( n19011 , n1186 , n15103 , n19010 );
or ( n19012 , n15814 , n18954 );
nand ( n19013 , n19011 , n19012 );
nor ( n19014 , n19009 , n19013 );
nand ( n19015 , n19006 , n19007 , n19014 );
or ( n19016 , n19005 , n15089 , n19015 );
nand ( n19017 , n1388 , n18982 );
not ( n19018 , n17784 );
nand ( n19019 , n19018 , n17665 , n17041 , n17673 );
nor ( n19020 , n723 , n18196 , n19019 );
or ( n19021 , n15089 , n19017 , n19020 );
nand ( n19022 , n19016 , n19021 );
not ( n19023 , n19022 );
nor ( n19024 , n19023 , n1826 , n1872 , n1712 );
nor ( n19025 , n1289 , n1398 );
not ( n19026 , n19025 );
not ( n19027 , n794 );
not ( n19028 , n19027 );
not ( n19029 , n1398 );
and ( n19030 , n19028 , n19029 );
not ( n19031 , n1289 );
and ( n19032 , n793 , n19031 );
nor ( n19033 , n19030 , n19032 );
nand ( n19034 , n793 , n794 );
nand ( n19035 , n19026 , n19033 , n19034 );
or ( n19036 , n16294 , n1288 );
and ( n19037 , n488 , n16832 );
nor ( n19038 , n1288 , n1475 );
nor ( n19039 , n19037 , n19038 );
nand ( n19040 , n19036 , n16437 , n19039 );
nand ( n19041 , n19035 , n19040 );
and ( n19042 , n804 , n16836 );
not ( n19043 , n807 );
not ( n19044 , n16836 );
or ( n19045 , n19043 , n19044 );
nand ( n19046 , n19045 , n16355 );
and ( n19047 , n16839 , n19046 );
not ( n19048 , n804 );
nand ( n19049 , n19048 , n1287 );
nand ( n19050 , n16839 , n19049 );
not ( n19051 , n19046 );
nand ( n19052 , n19050 , n19051 );
nand ( n19053 , n16853 , n843 , n19052 );
and ( n19054 , n843 , n16855 );
nor ( n19055 , n1285 , n1286 );
nor ( n19056 , n19054 , n19055 );
not ( n19057 , n19056 );
nand ( n19058 , n846 , n19057 , n19052 );
nand ( n19059 , n19053 , n19058 );
nor ( n19060 , n19042 , n19047 , n19059 );
or ( n19061 , n19041 , n19060 );
not ( n19062 , n1242 );
and ( n19063 , n1241 , n19062 );
not ( n19064 , n19041 );
or ( n19065 , n1283 , n16361 );
or ( n19066 , n16277 , n1284 );
nand ( n19067 , n1412 , n16285 );
and ( n19068 , n848 , n16858 );
and ( n19069 , n837 , n16861 );
nor ( n19070 , n19068 , n19069 );
nor ( n19071 , n1283 , n1284 );
nor ( n19072 , n16360 , n19071 );
and ( n19073 , n19070 , n19072 );
nand ( n19074 , n847 , n16864 );
nor ( n19075 , n16868 , n826 );
and ( n19076 , n19074 , n19075 );
nor ( n19077 , n19073 , n19076 );
and ( n19078 , n19067 , n19077 );
and ( n19079 , n848 , n19071 );
nor ( n19080 , n19078 , n19079 );
nand ( n19081 , n19065 , n19066 , n19080 );
or ( n19082 , n16357 , n1286 );
nand ( n19083 , n19082 , n16439 , n19056 );
nand ( n19084 , n19064 , n19081 , n19083 , n19052 );
nand ( n19085 , n19061 , n19063 , n19084 );
not ( n19086 , n1398 );
not ( n19087 , n19034 );
and ( n19088 , n19086 , n19087 );
and ( n19089 , n794 , n19031 );
nor ( n19090 , n19088 , n19089 );
not ( n19091 , n19039 );
nand ( n19092 , n841 , n19091 , n19035 );
and ( n19093 , n16848 , n488 , n19035 );
and ( n19094 , n793 , n19025 );
nor ( n19095 , n19093 , n19094 );
nand ( n19096 , n19090 , n19092 , n19095 );
or ( n19097 , n19085 , n16257 , n19096 );
not ( n19098 , n1241 );
nand ( n19099 , n1242 , n19098 );
not ( n19100 , n17724 );
nand ( n19101 , n19100 , n17586 , n16826 , n17592 );
nor ( n19102 , n829 , n18309 , n19101 );
or ( n19103 , n16257 , n19099 , n19102 );
nand ( n19104 , n19097 , n19103 );
not ( n19105 , n19104 );
nor ( n19106 , n19105 , n1828 , n1857 , n1733 );
not ( n19107 , n862 );
not ( n19108 , n17976 );
or ( n19109 , n19107 , n19108 );
and ( n19110 , n852 , n17942 );
nor ( n19111 , n19110 , n17946 );
nand ( n19112 , n19109 , n19111 );
not ( n19113 , n875 );
not ( n19114 , n17976 );
or ( n19115 , n19113 , n19114 );
and ( n19116 , n859 , n17942 );
nor ( n19117 , n19116 , n17946 );
nand ( n19118 , n19115 , n19117 );
not ( n19119 , n863 );
not ( n19120 , n17976 );
or ( n19121 , n19119 , n19120 );
and ( n19122 , n860 , n17942 );
nor ( n19123 , n19122 , n17946 );
nand ( n19124 , n19121 , n19123 );
not ( n19125 , n874 );
not ( n19126 , n17976 );
or ( n19127 , n19125 , n19126 );
and ( n19128 , n861 , n17942 );
nor ( n19129 , n19128 , n17946 );
nand ( n19130 , n19127 , n19129 );
or ( n19131 , n18456 , n18705 );
and ( n19132 , n863 , n17942 );
nor ( n19133 , n19132 , n17946 );
nand ( n19134 , n19131 , n19133 );
not ( n19135 , n864 );
not ( n19136 , n17976 );
or ( n19137 , n19135 , n19136 );
and ( n19138 , n873 , n17942 );
nor ( n19139 , n19138 , n17946 );
nand ( n19140 , n19137 , n19139 );
not ( n19141 , n1053 );
not ( n19142 , n17976 );
or ( n19143 , n19141 , n19142 );
nand ( n19144 , n1059 , n18762 );
nand ( n19145 , n19143 , n19144 );
not ( n19146 , n1054 );
not ( n19147 , n17976 );
or ( n19148 , n19146 , n19147 );
nand ( n19149 , n1060 , n18773 );
nand ( n19150 , n19148 , n19149 );
not ( n19151 , n1056 );
not ( n19152 , n18759 );
or ( n19153 , n19151 , n19152 );
nand ( n19154 , n1062 , n18762 );
nand ( n19155 , n19153 , n19154 );
not ( n19156 , n1057 );
not ( n19157 , n18759 );
or ( n19158 , n19156 , n19157 );
nand ( n19159 , n1063 , n18773 );
nand ( n19160 , n19158 , n19159 );
not ( n19161 , n1058 );
not ( n19162 , n18759 );
or ( n19163 , n19161 , n19162 );
nand ( n19164 , n1064 , n18762 );
nand ( n19165 , n19163 , n19164 );
not ( n19166 , n1059 );
not ( n19167 , n17976 );
or ( n19168 , n19166 , n19167 );
nand ( n19169 , n1065 , n18762 );
nand ( n19170 , n19168 , n19169 );
not ( n19171 , n1055 );
not ( n19172 , n17976 );
or ( n19173 , n19171 , n19172 );
nand ( n19174 , n1061 , n18773 );
nand ( n19175 , n19173 , n19174 );
not ( n19176 , n1010 );
not ( n19177 , n18759 );
or ( n19178 , n19176 , n19177 );
nand ( n19179 , n1072 , n18773 );
nand ( n19180 , n19178 , n19179 );
not ( n19181 , n1013 );
not ( n19182 , n17976 );
or ( n19183 , n19181 , n19182 );
nand ( n19184 , n1073 , n18762 );
nand ( n19185 , n19183 , n19184 );
not ( n19186 , n1308 );
and ( n19187 , n512 , n19186 );
and ( n19188 , n1308 , n17321 );
nor ( n19189 , n19187 , n19188 );
not ( n19190 , n19189 );
not ( n19191 , n16906 );
not ( n19192 , n16919 );
nand ( n19193 , n16909 , n16915 );
nand ( n19194 , n19192 , n19193 );
not ( n19195 , n19194 );
or ( n19196 , n19191 , n19195 );
nand ( n19197 , n19196 , n16923 );
nand ( n19198 , n16902 , n19197 );
and ( n19199 , n16911 , n16909 );
and ( n19200 , n16927 , n16924 );
not ( n19201 , n19200 );
not ( n19202 , n16932 );
not ( n19203 , n16929 );
nor ( n19204 , n19202 , n19203 );
not ( n19205 , n19204 );
not ( n19206 , n16943 );
nand ( n19207 , n16935 , n19206 );
not ( n19208 , n16935 );
not ( n19209 , n16938 );
or ( n19210 , n19208 , n19209 );
nand ( n19211 , n19210 , n16948 );
not ( n19212 , n19211 );
nand ( n19213 , n19207 , n19212 );
not ( n19214 , n19213 );
or ( n19215 , n19205 , n19214 );
nand ( n19216 , n16929 , n16952 );
and ( n19217 , n16958 , n19216 );
nand ( n19218 , n19215 , n19217 );
not ( n19219 , n19218 );
or ( n19220 , n19201 , n19219 );
and ( n19221 , n16924 , n16961 );
nor ( n19222 , n19221 , n16913 );
nand ( n19223 , n19220 , n19222 );
nand ( n19224 , n16906 , n19199 , n16902 , n19223 );
and ( n19225 , n19198 , n16900 , n19224 );
not ( n19226 , n19225 );
or ( n19227 , n19190 , n19226 );
or ( n19228 , n19189 , n19225 );
nand ( n19229 , n19227 , n19228 );
not ( n19230 , n1165 );
and ( n19231 , n600 , n19230 );
and ( n19232 , n1165 , n17402 );
nor ( n19233 , n19231 , n19232 );
not ( n19234 , n19233 );
not ( n19235 , n16977 );
not ( n19236 , n16990 );
nand ( n19237 , n16980 , n16986 );
nand ( n19238 , n19236 , n19237 );
not ( n19239 , n19238 );
or ( n19240 , n19235 , n19239 );
nand ( n19241 , n19240 , n16994 );
nand ( n19242 , n16973 , n19241 );
and ( n19243 , n16982 , n16980 );
and ( n19244 , n16995 , n16998 );
not ( n19245 , n19244 );
not ( n19246 , n17003 );
not ( n19247 , n17000 );
nor ( n19248 , n19246 , n19247 );
not ( n19249 , n19248 );
not ( n19250 , n17014 );
nand ( n19251 , n17006 , n19250 );
not ( n19252 , n17006 );
not ( n19253 , n17009 );
or ( n19254 , n19252 , n19253 );
nand ( n19255 , n19254 , n17019 );
not ( n19256 , n19255 );
nand ( n19257 , n19251 , n19256 );
not ( n19258 , n19257 );
or ( n19259 , n19249 , n19258 );
nand ( n19260 , n17000 , n17023 );
and ( n19261 , n17029 , n19260 );
nand ( n19262 , n19259 , n19261 );
not ( n19263 , n19262 );
or ( n19264 , n19245 , n19263 );
and ( n19265 , n16995 , n17032 );
nor ( n19266 , n19265 , n16984 );
nand ( n19267 , n19264 , n19266 );
nand ( n19268 , n16977 , n19243 , n16973 , n19267 );
and ( n19269 , n19242 , n16971 , n19268 );
not ( n19270 , n19269 );
or ( n19271 , n19234 , n19270 );
or ( n19272 , n19233 , n19269 );
nand ( n19273 , n19271 , n19272 );
and ( n19274 , n803 , n19031 );
and ( n19275 , n1289 , n17586 );
nor ( n19276 , n19274 , n19275 );
not ( n19277 , n19276 );
not ( n19278 , n16849 );
not ( n19279 , n16833 );
nand ( n19280 , n16834 , n16844 );
nand ( n19281 , n19279 , n19280 );
not ( n19282 , n19281 );
or ( n19283 , n19278 , n19282 );
nand ( n19284 , n19283 , n16852 );
nand ( n19285 , n16829 , n19284 );
not ( n19286 , n16834 );
nor ( n19287 , n16837 , n19286 );
and ( n19288 , n16854 , n16890 );
not ( n19289 , n19288 );
not ( n19290 , n16859 );
not ( n19291 , n16856 );
nor ( n19292 , n19290 , n19291 );
not ( n19293 , n19292 );
not ( n19294 , n16870 );
nand ( n19295 , n16862 , n19294 );
not ( n19296 , n16862 );
not ( n19297 , n16865 );
or ( n19298 , n19296 , n19297 );
nand ( n19299 , n19298 , n16875 );
not ( n19300 , n19299 );
nand ( n19301 , n19295 , n19300 );
not ( n19302 , n19301 );
or ( n19303 , n19293 , n19302 );
not ( n19304 , n16880 );
nand ( n19305 , n19304 , n16856 );
and ( n19306 , n16885 , n19305 );
nand ( n19307 , n19303 , n19306 );
not ( n19308 , n19307 );
or ( n19309 , n19289 , n19308 );
and ( n19310 , n16890 , n16888 );
nor ( n19311 , n19310 , n16840 );
nand ( n19312 , n19309 , n19311 );
nand ( n19313 , n16849 , n19287 , n16829 , n19312 );
and ( n19314 , n19285 , n16827 , n19313 );
not ( n19315 , n19314 );
or ( n19316 , n19277 , n19315 );
or ( n19317 , n19276 , n19314 );
nand ( n19318 , n19316 , n19317 );
and ( n19319 , n692 , n18949 );
and ( n19320 , n1395 , n17665 );
nor ( n19321 , n19319 , n19320 );
not ( n19322 , n19321 );
not ( n19323 , n17061 );
not ( n19324 , n17048 );
nand ( n19325 , n17049 , n17056 );
nand ( n19326 , n19324 , n19325 );
not ( n19327 , n19326 );
or ( n19328 , n19323 , n19327 );
nand ( n19329 , n19328 , n17064 );
nand ( n19330 , n17044 , n19329 );
and ( n19331 , n17049 , n17052 );
and ( n19332 , n17068 , n17065 );
not ( n19333 , n19332 );
not ( n19334 , n17073 );
not ( n19335 , n17070 );
nor ( n19336 , n19334 , n19335 );
not ( n19337 , n19336 );
not ( n19338 , n17084 );
nand ( n19339 , n17076 , n19338 );
not ( n19340 , n17076 );
not ( n19341 , n17079 );
or ( n19342 , n19340 , n19341 );
nand ( n19343 , n19342 , n17089 );
not ( n19344 , n19343 );
nand ( n19345 , n19339 , n19344 );
not ( n19346 , n19345 );
or ( n19347 , n19337 , n19346 );
nand ( n19348 , n17070 , n17093 );
and ( n19349 , n17099 , n19348 );
nand ( n19350 , n19347 , n19349 );
not ( n19351 , n19350 );
or ( n19352 , n19333 , n19351 );
and ( n19353 , n17065 , n17102 );
nor ( n19354 , n19353 , n17054 );
nand ( n19355 , n19352 , n19354 );
nand ( n19356 , n17061 , n19331 , n17044 , n19355 );
and ( n19357 , n19330 , n17042 , n19356 );
not ( n19358 , n19357 );
or ( n19359 , n19322 , n19358 );
or ( n19360 , n19321 , n19357 );
nand ( n19361 , n19359 , n19360 );
not ( n19362 , n1052 );
not ( n19363 , n18759 );
or ( n19364 , n19362 , n19363 );
nand ( n19365 , n1058 , n18762 );
nand ( n19366 , n19364 , n19365 );
not ( n19367 , n1794 );
or ( n19368 , n19367 , n1001 );
not ( n19369 , n19368 );
and ( n19370 , n1834 , n19369 );
and ( n19371 , n916 , n19368 );
nor ( n19372 , n19370 , n19371 );
not ( n19373 , n1673 );
not ( n19374 , n1868 );
nor ( n19375 , n19374 , n1866 );
nand ( n19376 , n1797 , n19375 );
not ( n19377 , n19376 );
nand ( n19378 , n405 , n19377 );
nor ( n19379 , n19378 , n15667 );
not ( n19380 , n15608 );
nand ( n19381 , n19380 , n15585 , n15624 );
nand ( n19382 , n19379 , n19381 , n15676 );
not ( n19383 , n15622 );
nor ( n19384 , n15617 , n19383 );
nor ( n19385 , n15676 , n15627 );
nand ( n19386 , n19384 , n19385 );
not ( n19387 , n19385 );
nand ( n19388 , n19381 , n15676 );
not ( n19389 , n1083 );
not ( n19390 , n15592 );
and ( n19391 , n1179 , n19389 , n19390 );
nand ( n19392 , n19387 , n19388 , n19391 );
and ( n19393 , n19382 , n19386 , n19392 );
nand ( n19394 , n19373 , n1474 , n19393 );
nor ( n19395 , n19372 , n19394 );
nand ( n19396 , n13531 , n13536 );
and ( n19397 , n13545 , n16537 );
nor ( n19398 , n19397 , n16524 );
or ( n19399 , n19396 , n19398 );
not ( n19400 , n13536 );
nand ( n19401 , n239 , n19400 );
not ( n19402 , n19401 );
nand ( n19403 , n19402 , n15377 , n15378 );
not ( n19404 , n19396 );
nand ( n19405 , n16537 , n13538 , n19404 );
nand ( n19406 , n19399 , n19403 , n19405 );
not ( n19407 , n716 );
nor ( n19408 , n1611 , n1618 );
not ( n19409 , n19408 );
or ( n19410 , n19407 , n19409 );
or ( n19411 , n1618 , n16402 );
nand ( n19412 , n19410 , n19411 );
not ( n19413 , n751 );
or ( n19414 , n19413 , n1611 );
and ( n19415 , n1597 , n15718 );
nor ( n19416 , n19415 , n1584 );
or ( n19417 , n15719 , n1597 );
nand ( n19418 , n19417 , n15788 );
or ( n19419 , n19416 , n19418 );
or ( n19420 , n15727 , n1550 );
or ( n19421 , n15716 , n1585 );
nand ( n19422 , n597 , n691 );
nor ( n19423 , n1550 , n1585 );
not ( n19424 , n19423 );
nand ( n19425 , n19420 , n19421 , n19422 , n19424 );
nand ( n19426 , n19419 , n19425 );
not ( n19427 , n19426 );
or ( n19428 , n1585 , n19422 );
or ( n19429 , n15716 , n1550 );
nand ( n19430 , n19428 , n19429 );
not ( n19431 , n1584 );
nand ( n19432 , n19431 , n19418 , n19425 );
nand ( n19433 , n691 , n19423 );
not ( n19434 , n1597 );
nand ( n19435 , n19434 , n509 , n19425 );
nand ( n19436 , n19432 , n19433 , n19435 );
nor ( n19437 , n19430 , n19436 );
not ( n19438 , n19437 );
or ( n19439 , n19427 , n19438 );
or ( n19440 , n15721 , n1619 );
or ( n19441 , n15739 , n1583 );
nand ( n19442 , n19440 , n19441 );
nor ( n19443 , n1583 , n1619 );
not ( n19444 , n19443 );
nand ( n19445 , n19444 , n16400 );
nor ( n19446 , n19442 , n19445 );
or ( n19447 , n1642 , n15741 , n19446 );
and ( n19448 , n614 , n19443 );
not ( n19449 , n1642 );
nand ( n19450 , n696 , n19449 );
nand ( n19451 , n15792 , n19450 );
not ( n19452 , n19451 );
or ( n19453 , n1617 , n19452 , n19446 );
or ( n19454 , n1619 , n16400 );
nand ( n19455 , n19453 , n19454 );
nor ( n19456 , n15721 , n1583 );
nor ( n19457 , n19448 , n19455 , n19456 );
nand ( n19458 , n19447 , n19457 , n19437 );
nand ( n19459 , n19439 , n19458 );
or ( n19460 , n19413 , n1618 );
or ( n19461 , n15750 , n1611 );
nand ( n19462 , n19460 , n19461 );
not ( n19463 , n16402 );
or ( n19464 , n19462 , n19463 , n19408 );
not ( n19465 , n15754 );
not ( n19466 , n1766 );
and ( n19467 , n19465 , n19466 );
nor ( n19468 , n19467 , n635 );
and ( n19469 , n1807 , n19468 );
and ( n19470 , n1766 , n15754 );
nor ( n19471 , n19469 , n19470 );
nand ( n19472 , n19464 , n19471 );
nand ( n19473 , n19414 , n19459 , n19472 );
or ( n19474 , n19412 , n19473 );
and ( n19475 , n1642 , n15741 );
nor ( n19476 , n19475 , n1617 );
nor ( n19477 , n19476 , n19451 );
or ( n19478 , n19477 , n19446 , n19426 );
nand ( n19479 , n19478 , n19459 );
nand ( n19480 , n19474 , n19479 );
not ( n19481 , n782 );
nor ( n19482 , n1654 , n1665 );
not ( n19483 , n19482 );
or ( n19484 , n19481 , n19483 );
or ( n19485 , n1665 , n15192 );
nand ( n19486 , n19484 , n19485 );
or ( n19487 , n15119 , n1654 );
and ( n19488 , n1565 , n15103 );
nor ( n19489 , n19488 , n1615 );
or ( n19490 , n15107 , n1565 );
nand ( n19491 , n19490 , n15837 );
or ( n19492 , n19489 , n19491 );
or ( n19493 , n15811 , n1570 );
not ( n19494 , n1578 );
nand ( n19495 , n19494 , n774 );
nor ( n19496 , n1570 , n1578 );
not ( n19497 , n19496 );
nand ( n19498 , n19493 , n19495 , n18953 , n19497 );
nand ( n19499 , n19492 , n19498 );
not ( n19500 , n19499 );
or ( n19501 , n1570 , n18953 );
or ( n19502 , n15811 , n1578 );
nand ( n19503 , n19501 , n19502 );
not ( n19504 , n1615 );
nand ( n19505 , n19504 , n19491 , n19498 );
nand ( n19506 , n774 , n19496 );
not ( n19507 , n1565 );
nand ( n19508 , n19507 , n487 , n19498 );
nand ( n19509 , n19505 , n19506 , n19508 );
nor ( n19510 , n19503 , n19509 );
not ( n19511 , n19510 );
or ( n19512 , n19500 , n19511 );
or ( n19513 , n15168 , n1613 );
not ( n19514 , n1604 );
nand ( n19515 , n19514 , n695 );
nand ( n19516 , n19513 , n19515 );
nor ( n19517 , n1604 , n1613 );
not ( n19518 , n19517 );
nand ( n19519 , n19518 , n15189 );
nor ( n19520 , n19516 , n19519 );
or ( n19521 , n1644 , n15113 , n19520 );
and ( n19522 , n698 , n19517 );
not ( n19523 , n1644 );
nand ( n19524 , n779 , n19523 );
nand ( n19525 , n15839 , n19524 );
not ( n19526 , n19525 );
or ( n19527 , n1664 , n19526 , n19520 );
or ( n19528 , n1604 , n15189 );
nand ( n19529 , n19527 , n19528 );
nor ( n19530 , n15174 , n1613 );
nor ( n19531 , n19522 , n19529 , n19530 );
nand ( n19532 , n19521 , n19531 , n19510 );
nand ( n19533 , n19512 , n19532 );
or ( n19534 , n15119 , n1665 );
or ( n19535 , n15122 , n1654 );
nand ( n19536 , n19534 , n19535 );
not ( n19537 , n15192 );
or ( n19538 , n19536 , n19537 , n19482 );
not ( n19539 , n1696 );
and ( n19540 , n791 , n19539 );
nor ( n19541 , n19540 , n715 );
and ( n19542 , n1832 , n19541 );
and ( n19543 , n1696 , n15126 );
nor ( n19544 , n19542 , n19543 );
nand ( n19545 , n19538 , n19544 );
nand ( n19546 , n19487 , n19533 , n19545 );
or ( n19547 , n19486 , n19546 );
and ( n19548 , n1644 , n15113 );
nor ( n19549 , n19548 , n1664 );
nor ( n19550 , n19549 , n19525 );
or ( n19551 , n19550 , n19520 , n19499 );
nand ( n19552 , n19551 , n19533 );
nand ( n19553 , n19547 , n19552 );
not ( n19554 , n637 );
nor ( n19555 , n1626 , n1638 );
not ( n19556 , n19555 );
or ( n19557 , n19554 , n19556 );
or ( n19558 , n1638 , n15077 );
nand ( n19559 , n19557 , n19558 );
or ( n19560 , n15002 , n1626 );
and ( n19561 , n1564 , n14986 );
nor ( n19562 , n19561 , n1591 );
or ( n19563 , n14990 , n1564 );
nand ( n19564 , n19563 , n15882 );
or ( n19565 , n19562 , n19564 );
or ( n19566 , n15860 , n1563 );
or ( n19567 , n15857 , n1567 );
nand ( n19568 , n510 , n599 );
nor ( n19569 , n1563 , n1567 );
not ( n19570 , n19569 );
nand ( n19571 , n19566 , n19567 , n19568 , n19570 );
nand ( n19572 , n19565 , n19571 );
not ( n19573 , n19572 );
or ( n19574 , n1567 , n19568 );
or ( n19575 , n15857 , n1563 );
nand ( n19576 , n19574 , n19575 );
not ( n19577 , n1591 );
nand ( n19578 , n19577 , n19564 , n19571 );
nand ( n19579 , n599 , n19569 );
not ( n19580 , n1564 );
nand ( n19581 , n19580 , n508 , n19571 );
nand ( n19582 , n19578 , n19579 , n19581 );
nor ( n19583 , n19576 , n19582 );
not ( n19584 , n19583 );
or ( n19585 , n19573 , n19584 );
or ( n19586 , n15058 , n1603 );
or ( n19587 , n15052 , n1590 );
nand ( n19588 , n19586 , n19587 );
nor ( n19589 , n1590 , n1603 );
not ( n19590 , n19589 );
nand ( n19591 , n19590 , n15073 );
nor ( n19592 , n19588 , n19591 );
or ( n19593 , n1641 , n14996 , n19592 );
and ( n19594 , n516 , n19589 );
not ( n19595 , n1641 );
nand ( n19596 , n613 , n19595 );
nand ( n19597 , n15886 , n19596 );
not ( n19598 , n19597 );
or ( n19599 , n1636 , n19598 , n19592 );
or ( n19600 , n1603 , n15073 );
nand ( n19601 , n19599 , n19600 );
nor ( n19602 , n15058 , n1590 );
nor ( n19603 , n19594 , n19601 , n19602 );
nand ( n19604 , n19593 , n19603 , n19583 );
nand ( n19605 , n19585 , n19604 );
or ( n19606 , n15002 , n1638 );
or ( n19607 , n15005 , n1626 );
nand ( n19608 , n19606 , n19607 );
or ( n19609 , n19608 , n15078 , n19555 );
not ( n19610 , n1694 );
and ( n19611 , n636 , n19610 );
nor ( n19612 , n19611 , n537 );
and ( n19613 , n1831 , n19612 );
not ( n19614 , n636 );
and ( n19615 , n1694 , n19614 );
nor ( n19616 , n19613 , n19615 );
nand ( n19617 , n19609 , n19616 );
nand ( n19618 , n19560 , n19605 , n19617 );
or ( n19619 , n19559 , n19618 );
and ( n19620 , n1641 , n14996 );
nor ( n19621 , n19620 , n1636 );
nor ( n19622 , n19621 , n19597 );
or ( n19623 , n19622 , n19592 , n19572 );
nand ( n19624 , n19623 , n19605 );
nand ( n19625 , n19619 , n19624 );
not ( n19626 , n848 );
nor ( n19627 , n1653 , n1674 );
not ( n19628 , n19627 );
or ( n19629 , n19626 , n19628 );
not ( n19630 , n16361 );
not ( n19631 , n19630 );
or ( n19632 , n1674 , n19631 );
nand ( n19633 , n19629 , n19632 );
or ( n19634 , n16277 , n1653 );
and ( n19635 , n1596 , n16415 );
nor ( n19636 , n19635 , n1614 );
or ( n19637 , n16294 , n1596 );
nand ( n19638 , n19637 , n16437 );
or ( n19639 , n19636 , n19638 );
or ( n19640 , n16426 , n1577 );
not ( n19641 , n1598 );
nand ( n19642 , n19641 , n794 );
nor ( n19643 , n1577 , n1598 );
not ( n19644 , n19643 );
nand ( n19645 , n19640 , n19642 , n19034 , n19644 );
nand ( n19646 , n19639 , n19645 );
not ( n19647 , n19646 );
or ( n19648 , n1598 , n19034 );
or ( n19649 , n19027 , n1577 );
nand ( n19650 , n19648 , n19649 );
not ( n19651 , n1614 );
nand ( n19652 , n19651 , n19638 , n19645 );
nand ( n19653 , n793 , n19643 );
not ( n19654 , n1596 );
nand ( n19655 , n19654 , n488 , n19645 );
nand ( n19656 , n19652 , n19653 , n19655 );
nor ( n19657 , n19650 , n19656 );
not ( n19658 , n19657 );
or ( n19659 , n19647 , n19658 );
or ( n19660 , n16292 , n1643 );
or ( n19661 , n16332 , n1612 );
nand ( n19662 , n19660 , n19661 );
nor ( n19663 , n1612 , n1643 );
not ( n19664 , n19663 );
nand ( n19665 , n19664 , n16355 );
nor ( n19666 , n19662 , n19665 );
or ( n19667 , n1666 , n16297 , n19666 );
and ( n19668 , n807 , n19663 );
not ( n19669 , n1666 );
nand ( n19670 , n846 , n19669 );
nand ( n19671 , n16439 , n19670 );
not ( n19672 , n19671 );
or ( n19673 , n1662 , n19672 , n19666 );
or ( n19674 , n1643 , n16355 );
nand ( n19675 , n19673 , n19674 );
nor ( n19676 , n16292 , n1612 );
nor ( n19677 , n19668 , n19675 , n19676 );
nand ( n19678 , n19667 , n19677 , n19657 );
nand ( n19679 , n19659 , n19678 );
or ( n19680 , n16277 , n1674 );
or ( n19681 , n16281 , n1653 );
nand ( n19682 , n19680 , n19681 );
or ( n19683 , n19682 , n19630 , n19627 );
not ( n19684 , n16285 );
not ( n19685 , n1695 );
and ( n19686 , n19684 , n19685 );
nor ( n19687 , n19686 , n826 );
and ( n19688 , n1833 , n19687 );
and ( n19689 , n1695 , n16285 );
nor ( n19690 , n19688 , n19689 );
nand ( n19691 , n19683 , n19690 );
nand ( n19692 , n19634 , n19679 , n19691 );
or ( n19693 , n19633 , n19692 );
and ( n19694 , n1666 , n16297 );
nor ( n19695 , n19694 , n1662 );
nor ( n19696 , n19695 , n19671 );
or ( n19697 , n19696 , n19666 , n19646 );
nand ( n19698 , n19697 , n19679 );
nand ( n19699 , n19693 , n19698 );
and ( n19700 , n1679 , n19369 );
and ( n19701 , n912 , n19368 );
nor ( n19702 , n19700 , n19701 );
nor ( n19703 , n19702 , n19394 );
or ( n19704 , n614 , n15796 );
nand ( n19705 , n19704 , n1808 , n15797 );
nor ( n19706 , n15739 , n15712 );
nand ( n19707 , n15740 , n15770 );
nor ( n19708 , n17171 , n17185 );
and ( n19709 , n19707 , n19708 );
or ( n19710 , n19707 , n19708 );
nand ( n19711 , n19710 , n17197 );
nor ( n19712 , n19709 , n19711 );
or ( n19713 , n19706 , n19712 );
nand ( n19714 , n19713 , n15704 );
and ( n19715 , n19705 , n19714 );
nor ( n19716 , n19715 , n15703 );
nor ( n19717 , n15246 , n15247 );
or ( n19718 , n19717 , n15271 , n15236 );
nand ( n19719 , n15249 , n15271 );
or ( n19720 , n19719 , n15248 , n748 );
nand ( n19721 , n19718 , n19720 );
not ( n19722 , n779 );
not ( n19723 , n15098 );
or ( n19724 , n19722 , n19723 );
nor ( n19725 , n15152 , n16799 );
or ( n19726 , n19725 , n16796 );
and ( n19727 , n19725 , n16796 );
nor ( n19728 , n19727 , n15829 );
nand ( n19729 , n19726 , n19728 );
nand ( n19730 , n19724 , n19729 );
and ( n19731 , n15090 , n19730 );
not ( n19732 , n779 );
not ( n19733 , n15841 );
or ( n19734 , n19732 , n19733 );
or ( n19735 , n779 , n15841 );
nand ( n19736 , n19734 , n19735 );
and ( n19737 , n1826 , n19736 );
nor ( n19738 , n19731 , n19737 );
nor ( n19739 , n15089 , n19738 );
and ( n19740 , n508 , n16908 );
and ( n19741 , n595 , n16905 );
nor ( n19742 , n19740 , n19741 );
nor ( n19743 , n1211 , n1305 );
not ( n19744 , n19743 );
and ( n19745 , n19742 , n15884 , n19744 );
and ( n19746 , n599 , n19186 );
and ( n19747 , n510 , n16901 );
nor ( n19748 , n19746 , n19747 );
nand ( n19749 , n16901 , n19186 );
and ( n19750 , n19748 , n19568 , n19749 );
nor ( n19751 , n19745 , n19750 );
not ( n19752 , n516 );
not ( n19753 , n16910 );
or ( n19754 , n19752 , n19753 );
nand ( n19755 , n19754 , n15073 );
and ( n19756 , n16912 , n19755 );
and ( n19757 , n515 , n16910 );
nor ( n19758 , n19756 , n19757 );
and ( n19759 , n609 , n16928 );
nor ( n19760 , n1222 , n1303 );
nor ( n19761 , n19759 , n19760 );
and ( n19762 , n1218 , n15058 );
nor ( n19763 , n19762 , n1304 );
nor ( n19764 , n19763 , n19755 );
nor ( n19765 , n19761 , n19764 );
and ( n19766 , n613 , n19765 );
nor ( n19767 , n1222 , n14996 , n19764 );
nor ( n19768 , n19766 , n19767 );
nand ( n19769 , n19758 , n19768 );
nand ( n19770 , n19751 , n19769 );
not ( n19771 , n1385 );
nor ( n19772 , n19771 , n1386 );
or ( n19773 , n1302 , n15077 );
nor ( n19774 , n1216 , n1302 );
and ( n19775 , n637 , n19774 );
and ( n19776 , n638 , n16931 );
nor ( n19777 , n19775 , n19776 );
or ( n19778 , n16937 , n636 );
and ( n19779 , n638 , n16934 );
and ( n19780 , n637 , n16931 );
nor ( n19781 , n19779 , n19780 );
not ( n19782 , n19774 );
and ( n19783 , n19781 , n15077 , n19782 );
and ( n19784 , n636 , n16937 );
nor ( n19785 , n19784 , n16941 , n537 );
nor ( n19786 , n19783 , n19785 );
nand ( n19787 , n19778 , n19786 );
nand ( n19788 , n19773 , n19777 , n19787 );
not ( n19789 , n613 );
or ( n19790 , n19789 , n1222 );
nand ( n19791 , n19790 , n15886 , n19761 );
not ( n19792 , n19764 );
nand ( n19793 , n19788 , n19791 , n19792 , n19751 );
nand ( n19794 , n19770 , n19772 , n19793 );
and ( n19795 , n16908 , n15883 );
and ( n19796 , n595 , n19743 );
and ( n19797 , n508 , n16905 );
nor ( n19798 , n19795 , n19796 , n19797 );
or ( n19799 , n19750 , n19798 );
or ( n19800 , n1306 , n19568 );
not ( n19801 , n19749 );
and ( n19802 , n599 , n19801 );
and ( n19803 , n510 , n19186 );
nor ( n19804 , n19802 , n19803 );
nand ( n19805 , n19799 , n19800 , n19804 );
or ( n19806 , n19794 , n14973 , n19805 );
nand ( n19807 , n1386 , n19771 );
not ( n19808 , n17880 );
nand ( n19809 , n19808 , n17321 , n16899 , n17328 );
nor ( n19810 , n539 , n18059 , n19809 );
or ( n19811 , n14973 , n19807 , n19810 );
nand ( n19812 , n19806 , n19811 );
not ( n19813 , n19812 );
nor ( n19814 , n19813 , n1819 , n1863 , n1736 );
not ( n19815 , n2 );
or ( n19816 , n15246 , n19815 , n15263 );
or ( n19817 , n831 , n15244 );
nand ( n19818 , n19817 , n18683 , n15240 );
not ( n19819 , n2 );
not ( n19820 , n18686 );
or ( n19821 , n19818 , n19819 , n19820 );
nand ( n19822 , n19816 , n19821 );
and ( n19823 , n662 , n16976 );
and ( n19824 , n509 , n16979 );
nor ( n19825 , n19823 , n19824 );
nor ( n19826 , n1328 , n1378 );
not ( n19827 , n19826 );
and ( n19828 , n19825 , n15790 , n19827 );
and ( n19829 , n597 , n16972 );
and ( n19830 , n691 , n19230 );
nor ( n19831 , n19829 , n19830 );
nand ( n19832 , n19230 , n16972 );
and ( n19833 , n19831 , n19422 , n19832 );
nor ( n19834 , n19828 , n19833 );
not ( n19835 , n614 );
not ( n19836 , n16981 );
or ( n19837 , n19835 , n19836 );
nand ( n19838 , n19837 , n16400 );
and ( n19839 , n16983 , n19838 );
and ( n19840 , n612 , n16981 );
nor ( n19841 , n19839 , n19840 );
and ( n19842 , n678 , n16999 );
nor ( n19843 , n1325 , n1393 );
nor ( n19844 , n19842 , n19843 );
and ( n19845 , n1327 , n15721 );
nor ( n19846 , n19845 , n1326 );
nor ( n19847 , n19846 , n19838 );
nor ( n19848 , n19844 , n19847 );
and ( n19849 , n696 , n19848 );
nor ( n19850 , n1393 , n15741 , n19847 );
nor ( n19851 , n19849 , n19850 );
nand ( n19852 , n19841 , n19851 );
nand ( n19853 , n19834 , n19852 );
not ( n19854 , n1209 );
nor ( n19855 , n19854 , n1261 );
or ( n19856 , n1323 , n16402 );
nor ( n19857 , n1323 , n1324 );
and ( n19858 , n716 , n19857 );
and ( n19859 , n751 , n17002 );
nor ( n19860 , n19858 , n19859 );
or ( n19861 , n17008 , n747 );
and ( n19862 , n716 , n17002 );
and ( n19863 , n751 , n17005 );
nor ( n19864 , n19862 , n19863 );
not ( n19865 , n19857 );
and ( n19866 , n19864 , n16402 , n19865 );
and ( n19867 , n747 , n17008 );
nor ( n19868 , n19867 , n17011 , n635 );
nor ( n19869 , n19866 , n19868 );
nand ( n19870 , n19861 , n19869 );
nand ( n19871 , n19856 , n19860 , n19870 );
or ( n19872 , n15733 , n1393 );
nand ( n19873 , n19872 , n15792 , n19844 );
not ( n19874 , n19847 );
nand ( n19875 , n19871 , n19873 , n19874 , n19834 );
nand ( n19876 , n19853 , n19855 , n19875 );
and ( n19877 , n16979 , n15789 );
and ( n19878 , n662 , n19826 );
and ( n19879 , n509 , n16976 );
nor ( n19880 , n19877 , n19878 , n19879 );
or ( n19881 , n19833 , n19880 );
or ( n19882 , n1330 , n19422 );
not ( n19883 , n19832 );
and ( n19884 , n691 , n19883 );
and ( n19885 , n597 , n19230 );
nor ( n19886 , n19884 , n19885 );
nand ( n19887 , n19881 , n19882 , n19886 );
or ( n19888 , n19876 , n15703 , n19887 );
nand ( n19889 , n1261 , n19854 );
not ( n19890 , n17929 );
nand ( n19891 , n19890 , n17402 , n16970 , n17409 );
nor ( n19892 , n640 , n18112 , n19891 );
or ( n19893 , n15703 , n19889 , n19892 );
nand ( n19894 , n19888 , n19893 );
not ( n19895 , n19894 );
nor ( n19896 , n19895 , n1808 , n1859 , n1737 );
not ( n19897 , n846 );
not ( n19898 , n16347 );
or ( n19899 , n19897 , n19898 );
nor ( n19900 , n16274 , n16733 );
or ( n19901 , n19900 , n16730 );
and ( n19902 , n19900 , n16730 );
nor ( n19903 , n19902 , n16265 );
nand ( n19904 , n19901 , n19903 );
nand ( n19905 , n19899 , n19904 );
and ( n19906 , n16258 , n19905 );
not ( n19907 , n846 );
not ( n19908 , n16441 );
or ( n19909 , n19907 , n19908 );
or ( n19910 , n846 , n16441 );
nand ( n19911 , n19909 , n19910 );
and ( n19912 , n1828 , n19911 );
nor ( n19913 , n19906 , n19912 );
nor ( n19914 , n16257 , n19913 );
nand ( n19915 , n890 , n916 );
not ( n19916 , n19915 );
or ( n19917 , n917 , n19916 );
nand ( n19918 , n19917 , n912 , n19393 );
nor ( n19919 , n894 , n895 );
not ( n19920 , n19919 );
nor ( n19921 , n893 , n919 );
not ( n19922 , n19921 );
or ( n19923 , n19920 , n19922 );
nand ( n19924 , n19923 , n19393 );
nand ( n19925 , n19918 , n19924 );
not ( n19926 , n369 );
nand ( n19927 , n936 , n19926 );
and ( n19928 , n13660 , n19927 );
or ( n19929 , n14591 , n936 );
nand ( n19930 , n368 , n369 );
nand ( n19931 , n19929 , n19930 );
nor ( n19932 , n19928 , n19931 );
not ( n19933 , n370 );
nand ( n19934 , n937 , n19933 );
and ( n19935 , n18835 , n19934 );
or ( n19936 , n12640 , n937 );
nand ( n19937 , n350 , n370 );
nand ( n19938 , n19936 , n19937 );
nor ( n19939 , n19935 , n19938 );
not ( n19940 , n353 );
nand ( n19941 , n19940 , n939 );
and ( n19942 , n13633 , n19941 );
or ( n19943 , n14543 , n939 );
nand ( n19944 , n353 , n371 );
nand ( n19945 , n19943 , n19944 );
or ( n19946 , n19942 , n19945 );
not ( n19947 , n18815 );
not ( n19948 , n365 );
nand ( n19949 , n1006 , n19948 );
not ( n19950 , n19949 );
or ( n19951 , n19947 , n19950 );
nand ( n19952 , n372 , n19949 );
nand ( n19953 , n19951 , n19952 );
nand ( n19954 , n19946 , n19953 );
nor ( n19955 , n19932 , n19939 , n19954 );
not ( n19956 , n19954 );
not ( n19957 , n888 );
not ( n19958 , n19952 );
and ( n19959 , n19957 , n19958 );
nor ( n19960 , n14552 , n939 );
and ( n19961 , n19960 , n19953 );
nor ( n19962 , n19959 , n19961 );
nand ( n19963 , n365 , n12538 );
nand ( n19964 , n13633 , n19945 , n19953 );
and ( n19965 , n19962 , n19963 , n19964 );
not ( n19966 , n19965 );
or ( n19967 , n19956 , n19966 );
and ( n19968 , n13660 , n19931 );
and ( n19969 , n369 , n13675 );
nor ( n19970 , n19968 , n19969 );
or ( n19971 , n19970 , n19939 );
and ( n19972 , n18835 , n19938 );
nor ( n19973 , n19933 , n937 );
nor ( n19974 , n19972 , n19973 );
nand ( n19975 , n19971 , n19974 , n19965 );
nand ( n19976 , n19967 , n19975 );
not ( n19977 , n19976 );
or ( n19978 , n1002 , n19955 , n19977 );
nor ( n19979 , n879 , n933 );
nand ( n19980 , n366 , n19979 );
not ( n19981 , n386 );
nand ( n19982 , n988 , n19981 );
and ( n19983 , n366 , n13664 );
not ( n19984 , n879 );
and ( n19985 , n367 , n19984 );
nor ( n19986 , n19983 , n19985 );
and ( n19987 , n366 , n367 );
not ( n19988 , n19987 );
not ( n19989 , n19979 );
nand ( n19990 , n19986 , n19988 , n19989 );
and ( n19991 , n19982 , n19990 );
and ( n19992 , n19984 , n19987 );
nor ( n19993 , n19991 , n19992 );
nand ( n19994 , n19980 , n19993 , n19976 );
nor ( n19995 , n14593 , n933 );
or ( n19996 , n19994 , n1002 , n19995 );
nand ( n19997 , n19978 , n19996 );
and ( n19998 , n1802 , n19369 );
and ( n19999 , n890 , n19368 );
nor ( n20000 , n19998 , n19999 );
nor ( n20001 , n20000 , n19394 );
not ( n20002 , n892 );
nand ( n20003 , n920 , n921 );
not ( n20004 , n20003 );
and ( n20005 , n20002 , n20004 );
and ( n20006 , n892 , n20003 );
nor ( n20007 , n20005 , n20006 );
not ( n20008 , n1794 );
nand ( n20009 , n20008 , n1474 , n19393 );
nor ( n20010 , n20007 , n20009 );
and ( n20011 , n1661 , n19369 );
and ( n20012 , n893 , n19368 );
nor ( n20013 , n20011 , n20012 );
nor ( n20014 , n20013 , n19394 );
and ( n20015 , n1656 , n19369 );
and ( n20016 , n894 , n19368 );
nor ( n20017 , n20015 , n20016 );
nor ( n20018 , n20017 , n19394 );
and ( n20019 , n1651 , n19369 );
and ( n20020 , n895 , n19368 );
nor ( n20021 , n20019 , n20020 );
nor ( n20022 , n20021 , n19394 );
and ( n20023 , n1675 , n19369 );
and ( n20024 , n919 , n19368 );
nor ( n20025 , n20023 , n20024 );
nor ( n20026 , n20025 , n19394 );
nor ( n20027 , n920 , n20009 );
not ( n20028 , n921 );
xor ( n20029 , n920 , n20028 );
nor ( n20030 , n20029 , n20009 );
not ( n20031 , n922 );
not ( n20032 , n20003 );
nand ( n20033 , n20032 , n892 );
not ( n20034 , n20033 );
and ( n20035 , n20031 , n20034 );
and ( n20036 , n922 , n20033 );
nor ( n20037 , n20035 , n20036 );
nor ( n20038 , n20037 , n20009 );
not ( n20039 , n1092 );
or ( n20040 , n20039 , n1048 );
nand ( n20041 , n1048 , n20039 );
nand ( n20042 , n20040 , n20041 );
not ( n20043 , n1799 );
not ( n20044 , n902 );
nor ( n20045 , n20044 , n1066 );
not ( n20046 , n15589 );
not ( n20047 , n15587 );
nand ( n20048 , n20047 , n15584 );
nor ( n20049 , n20046 , n20048 );
nand ( n20050 , n20045 , n15603 , n20049 );
nand ( n20051 , n1066 , n20044 , n15603 , n20049 );
not ( n20052 , n20051 );
nand ( n20053 , n20043 , n19377 , n20050 , n20052 );
not ( n20054 , n1866 );
nor ( n20055 , n20054 , n1868 );
nand ( n20056 , n1803 , n20055 );
not ( n20057 , n20056 );
not ( n20058 , n20050 );
nand ( n20059 , n20043 , n20057 , n20051 , n20058 );
and ( n20060 , n20053 , n20059 );
not ( n20061 , n20060 );
and ( n20062 , n20042 , n20061 );
and ( n20063 , n1048 , n20060 );
nor ( n20064 , n20062 , n20063 );
nor ( n20065 , n1113 , n20064 );
not ( n20066 , n1050 );
nand ( n20067 , n1048 , n1092 );
not ( n20068 , n20067 );
or ( n20069 , n20066 , n20068 );
or ( n20070 , n1050 , n20067 );
nand ( n20071 , n20069 , n20070 );
and ( n20072 , n20071 , n20061 );
and ( n20073 , n1050 , n20060 );
nor ( n20074 , n20072 , n20073 );
nor ( n20075 , n1113 , n20074 );
and ( n20076 , n1092 , n20060 );
not ( n20077 , n1092 );
and ( n20078 , n20077 , n20061 );
nor ( n20079 , n20076 , n20078 );
nor ( n20080 , n1113 , n20079 );
not ( n20081 , n918 );
nor ( n20082 , n20081 , n18491 );
and ( n20083 , n1760 , n19369 );
and ( n20084 , n917 , n19368 );
nor ( n20085 , n20083 , n20084 );
nor ( n20086 , n20085 , n19394 );
not ( n20087 , n839 );
not ( n20088 , n16347 );
or ( n20089 , n20087 , n20088 );
nand ( n20090 , n17565 , n17537 );
not ( n20091 , n17705 );
or ( n20092 , n20090 , n20091 );
nand ( n20093 , n20090 , n20091 );
nand ( n20094 , n20092 , n20093 , n16268 );
nand ( n20095 , n20089 , n20094 );
and ( n20096 , n16258 , n20095 );
not ( n20097 , n16884 );
not ( n20098 , n17598 );
or ( n20099 , n20097 , n20098 );
or ( n20100 , n16884 , n17598 );
nand ( n20101 , n20099 , n20100 );
and ( n20102 , n1828 , n20101 );
nor ( n20103 , n20096 , n20102 );
nor ( n20104 , n16257 , n20103 );
not ( n20105 , n836 );
not ( n20106 , n16268 );
not ( n20107 , n20106 );
or ( n20108 , n20105 , n20107 );
not ( n20109 , n17568 );
nor ( n20110 , n20109 , n17541 );
nand ( n20111 , n18290 , n18295 );
or ( n20112 , n20110 , n20111 );
and ( n20113 , n20110 , n20111 );
nor ( n20114 , n20113 , n16267 );
nand ( n20115 , n20112 , n20114 );
nand ( n20116 , n20108 , n20115 );
and ( n20117 , n16258 , n20116 );
or ( n20118 , n17594 , n18310 );
nand ( n20119 , n20118 , n18311 );
and ( n20120 , n1828 , n20119 );
nor ( n20121 , n20117 , n20120 );
nor ( n20122 , n16257 , n20121 );
and ( n20123 , n14500 , n14486 );
not ( n20124 , n20123 );
not ( n20125 , n14495 );
not ( n20126 , n20125 );
or ( n20127 , n20124 , n20126 );
or ( n20128 , n20123 , n20125 );
nand ( n20129 , n20127 , n20128 );
nor ( n20130 , n13527 , n15399 , n13577 );
not ( n20131 , n784 );
not ( n20132 , n15098 );
or ( n20133 , n20131 , n20132 );
not ( n20134 , n17647 );
nor ( n20135 , n20134 , n17620 );
nand ( n20136 , n18176 , n18181 );
or ( n20137 , n20135 , n20136 );
and ( n20138 , n20135 , n20136 );
nor ( n20139 , n20138 , n15829 );
nand ( n20140 , n20137 , n20139 );
nand ( n20141 , n20133 , n20140 );
and ( n20142 , n15090 , n20141 );
or ( n20143 , n18193 , n18197 );
nand ( n20144 , n20143 , n18198 );
and ( n20145 , n1826 , n20144 );
nor ( n20146 , n20142 , n20145 );
nor ( n20147 , n15089 , n20146 );
nand ( n20148 , n13349 , n13352 );
not ( n20149 , n20148 );
not ( n20150 , n13371 );
or ( n20151 , n20149 , n20150 );
or ( n20152 , n20148 , n13371 );
nand ( n20153 , n20151 , n20152 );
not ( n20154 , n438 );
buf ( n20155 , n12868 );
not ( n20156 , n20155 );
buf ( n20157 , n12830 );
nand ( n20158 , n20156 , n20157 );
not ( n20159 , n20158 );
or ( n20160 , n20154 , n20159 );
nor ( n20161 , n267 , n1676 );
nand ( n20162 , n20160 , n20161 );
and ( n20163 , n1499 , n15209 , n15220 );
and ( n20164 , n20162 , n20163 );
and ( n20165 , n438 , n15203 );
nor ( n20166 , n20165 , n267 );
and ( n20167 , n15206 , n15211 );
nand ( n20168 , n1219 , n15205 , n20167 );
or ( n20169 , n20166 , n20168 );
not ( n20170 , n15205 );
not ( n20171 , n1538 );
and ( n20172 , n20170 , n20171 );
nor ( n20173 , n20172 , n267 );
not ( n20174 , n15210 );
nand ( n20175 , n789 , n15206 , n15215 , n20174 );
or ( n20176 , n20173 , n20175 );
nand ( n20177 , n20169 , n20176 );
not ( n20178 , n2 );
nor ( n20179 , n20164 , n20177 , n20178 );
nand ( n20180 , n15217 , n15207 , n538 , n15220 );
not ( n20181 , n20180 );
nand ( n20182 , n226 , n15377 );
not ( n20183 , n225 );
and ( n20184 , n15377 , n250 , n20183 );
not ( n20185 , n1219 );
nand ( n20186 , n20185 , n438 , n20167 );
nor ( n20187 , n20184 , n20186 );
nand ( n20188 , n438 , n20182 , n20187 );
not ( n20189 , n20188 );
or ( n20190 , n20181 , n20189 );
or ( n20191 , n438 , n1230 );
nand ( n20192 , n20190 , n20191 );
not ( n20193 , n20166 );
not ( n20194 , n15222 );
and ( n20195 , n20193 , n20194 );
not ( n20196 , n267 );
not ( n20197 , n438 );
not ( n20198 , n1379 );
and ( n20199 , n20197 , n20198 );
nor ( n20200 , n20199 , n387 );
not ( n20201 , n20200 );
and ( n20202 , n20196 , n20201 );
nand ( n20203 , n465 , n15215 , n15211 );
nor ( n20204 , n20202 , n20203 );
nor ( n20205 , n20195 , n20204 );
nand ( n20206 , n20179 , n20192 , n20205 );
not ( n20207 , n571 );
not ( n20208 , n14981 );
or ( n20209 , n20207 , n20208 );
nand ( n20210 , n17300 , n17272 );
not ( n20211 , n17861 );
or ( n20212 , n20210 , n20211 );
nand ( n20213 , n20210 , n20211 );
nand ( n20214 , n20212 , n20213 , n15874 );
nand ( n20215 , n20209 , n20214 );
and ( n20216 , n14974 , n20215 );
not ( n20217 , n16957 );
not ( n20218 , n17333 );
or ( n20219 , n20217 , n20218 );
or ( n20220 , n16957 , n17333 );
nand ( n20221 , n20219 , n20220 );
and ( n20222 , n1819 , n20221 );
nor ( n20223 , n20216 , n20222 );
nor ( n20224 , n14973 , n20223 );
nor ( n20225 , n594 , n1800 );
and ( n20226 , n607 , n608 );
not ( n20227 , n596 );
nand ( n20228 , n605 , n606 );
not ( n20229 , n562 );
nand ( n20230 , n598 , n603 );
nor ( n20231 , n20229 , n20230 );
nand ( n20232 , n604 , n20231 );
nor ( n20233 , n20228 , n20232 );
nand ( n20234 , n577 , n20233 );
nor ( n20235 , n20227 , n20234 );
nand ( n20236 , n602 , n20226 , n20235 );
and ( n20237 , n594 , n20236 );
or ( n20238 , n594 , n20236 );
nand ( n20239 , n20238 , n1800 );
nor ( n20240 , n20237 , n20239 );
nor ( n20241 , n834 , n20225 , n20240 );
not ( n20242 , n639 );
not ( n20243 , n14981 );
or ( n20244 , n20242 , n20243 );
not ( n20245 , n17303 );
nor ( n20246 , n20245 , n17277 );
nand ( n20247 , n18039 , n18044 );
or ( n20248 , n20246 , n20247 );
and ( n20249 , n20246 , n20247 );
not ( n20250 , n14980 );
nor ( n20251 , n20249 , n20250 );
nand ( n20252 , n20248 , n20251 );
nand ( n20253 , n20244 , n20252 );
and ( n20254 , n14974 , n20253 );
or ( n20255 , n18056 , n18060 );
nand ( n20256 , n20255 , n18061 );
and ( n20257 , n1819 , n20256 );
nor ( n20258 , n20254 , n20257 );
nor ( n20259 , n14973 , n20258 );
not ( n20260 , n670 );
not ( n20261 , n16393 );
or ( n20262 , n20260 , n20261 );
nand ( n20263 , n17381 , n17353 );
not ( n20264 , n17912 );
or ( n20265 , n20263 , n20264 );
nand ( n20266 , n20263 , n20264 );
nand ( n20267 , n20265 , n20266 , n17197 );
nand ( n20268 , n20262 , n20267 );
and ( n20269 , n15704 , n20268 );
not ( n20270 , n17028 );
not ( n20271 , n17414 );
or ( n20272 , n20270 , n20271 );
or ( n20273 , n17028 , n17414 );
nand ( n20274 , n20272 , n20273 );
and ( n20275 , n1808 , n20274 );
nor ( n20276 , n20269 , n20275 );
nor ( n20277 , n15703 , n20276 );
not ( n20278 , n696 );
not ( n20279 , n16393 );
or ( n20280 , n20278 , n20279 );
not ( n20281 , n15734 );
nor ( n20282 , n20281 , n15732 );
or ( n20283 , n20282 , n17222 );
and ( n20284 , n20282 , n17222 );
nor ( n20285 , n20284 , n17196 );
nand ( n20286 , n20283 , n20285 );
nand ( n20287 , n20280 , n20286 );
and ( n20288 , n15704 , n20287 );
not ( n20289 , n696 );
not ( n20290 , n15795 );
or ( n20291 , n20289 , n20290 );
or ( n20292 , n696 , n15795 );
nand ( n20293 , n20291 , n20292 );
and ( n20294 , n1808 , n20293 );
nor ( n20295 , n20288 , n20294 );
nor ( n20296 , n15703 , n20295 );
not ( n20297 , n717 );
not ( n20298 , n17198 );
or ( n20299 , n20297 , n20298 );
not ( n20300 , n17384 );
nor ( n20301 , n20300 , n17358 );
nand ( n20302 , n18092 , n18097 );
or ( n20303 , n20301 , n20302 );
and ( n20304 , n20301 , n20302 );
nor ( n20305 , n20304 , n18162 );
nand ( n20306 , n20303 , n20305 );
nand ( n20307 , n20299 , n20306 );
and ( n20308 , n15704 , n20307 );
or ( n20309 , n18109 , n18113 );
nand ( n20310 , n20309 , n18114 );
and ( n20311 , n1808 , n20310 );
nor ( n20312 , n20308 , n20311 );
nor ( n20313 , n15703 , n20312 );
not ( n20314 , n756 );
not ( n20315 , n18627 );
or ( n20316 , n20314 , n20315 );
nand ( n20317 , n17644 , n17616 );
not ( n20318 , n17767 );
or ( n20319 , n20317 , n20318 );
nand ( n20320 , n20317 , n20318 );
nand ( n20321 , n20319 , n20320 , n15097 );
nand ( n20322 , n20316 , n20321 );
and ( n20323 , n15090 , n20322 );
not ( n20324 , n17615 );
not ( n20325 , n17678 );
or ( n20326 , n20324 , n20325 );
or ( n20327 , n17615 , n17678 );
nand ( n20328 , n20326 , n20327 );
and ( n20329 , n1826 , n20328 );
nor ( n20330 , n20323 , n20329 );
nor ( n20331 , n15089 , n20330 );
and ( n20332 , n763 , n15263 );
not ( n20333 , n2 );
and ( n20334 , n15248 , n806 , n18895 );
nor ( n20335 , n20334 , n763 );
nor ( n20336 , n20332 , n20333 , n20335 );
and ( n20337 , n13633 , n19979 , n13620 );
nor ( n20338 , n1006 , n13683 , n13528 );
nand ( n20339 , n13660 , n13623 , n20337 , n20338 );
nor ( n20340 , n20339 , n988 , n13577 );
or ( n20341 , n1173 , n1275 );
nand ( n20342 , n1173 , n1275 );
nand ( n20343 , n20341 , n20342 );
or ( n20344 , n1277 , n1446 );
nand ( n20345 , n1277 , n1446 );
nand ( n20346 , n20344 , n20345 );
or ( n20347 , n1382 , n1442 );
nand ( n20348 , n1382 , n1442 );
nand ( n20349 , n20347 , n20348 );
not ( n20350 , n1276 );
and ( n20351 , n1447 , n20350 );
not ( n20352 , n1447 );
and ( n20353 , n20352 , n1276 );
nor ( n20354 , n20351 , n20353 );
nand ( n20355 , n20343 , n20346 , n20349 , n20354 );
not ( n20356 , n1173 );
not ( n20357 , n1244 );
or ( n20358 , n20356 , n20357 );
or ( n20359 , n1173 , n1244 );
nand ( n20360 , n20358 , n20359 );
not ( n20361 , n1245 );
not ( n20362 , n1442 );
or ( n20363 , n20361 , n20362 );
or ( n20364 , n1245 , n1442 );
nand ( n20365 , n20363 , n20364 );
not ( n20366 , n1246 );
not ( n20367 , n1446 );
or ( n20368 , n20366 , n20367 );
or ( n20369 , n1246 , n1446 );
nand ( n20370 , n20368 , n20369 );
not ( n20371 , n1199 );
not ( n20372 , n1447 );
or ( n20373 , n20371 , n20372 );
or ( n20374 , n1199 , n1447 );
nand ( n20375 , n20373 , n20374 );
nand ( n20376 , n20360 , n20365 , n20370 , n20375 );
xor ( n20377 , n1173 , n1183 );
xor ( n20378 , n1264 , n1446 );
nor ( n20379 , n20377 , n20378 );
not ( n20380 , n1263 );
not ( n20381 , n1442 );
and ( n20382 , n20380 , n20381 );
and ( n20383 , n1263 , n1442 );
nor ( n20384 , n20382 , n20383 );
not ( n20385 , n1265 );
not ( n20386 , n1447 );
and ( n20387 , n20385 , n20386 );
and ( n20388 , n1265 , n1447 );
nor ( n20389 , n20387 , n20388 );
nor ( n20390 , n20384 , n20389 );
nand ( n20391 , n20379 , n20390 );
nand ( n20392 , n1389 , n1442 );
not ( n20393 , n20392 );
nor ( n20394 , n1389 , n1442 );
nor ( n20395 , n20393 , n20394 );
nand ( n20396 , n1252 , n1446 );
not ( n20397 , n20396 );
nor ( n20398 , n1252 , n1446 );
nor ( n20399 , n20397 , n20398 );
nor ( n20400 , n20395 , n20399 );
xor ( n20401 , n1155 , n1173 );
and ( n20402 , n1391 , n1447 );
not ( n20403 , n1391 );
and ( n20404 , n20403 , n15467 );
nor ( n20405 , n20402 , n20404 );
nor ( n20406 , n20401 , n20405 );
nand ( n20407 , n20400 , n20406 );
and ( n20408 , n20391 , n20407 );
and ( n20409 , n20355 , n20376 , n20408 );
not ( n20410 , n20409 );
buf ( n20411 , n20410 );
not ( n20412 , n20411 );
and ( n20413 , n883 , n20412 );
not ( n20414 , n20355 );
nand ( n20415 , n20414 , n20408 );
not ( n20416 , n20415 );
not ( n20417 , n20416 );
not ( n20418 , n20417 );
and ( n20419 , n702 , n20418 );
nor ( n20420 , n20413 , n20419 );
not ( n20421 , n20376 );
and ( n20422 , n20355 , n20421 , n20408 );
not ( n20423 , n20422 );
buf ( n20424 , n20423 );
not ( n20425 , n20424 );
and ( n20426 , n800 , n20425 );
not ( n20427 , n20391 );
and ( n20428 , n20407 , n20427 );
not ( n20429 , n20428 );
not ( n20430 , n20429 );
and ( n20431 , n620 , n20430 );
not ( n20432 , n20407 );
not ( n20433 , n20432 );
not ( n20434 , n20433 );
and ( n20435 , n559 , n20434 );
nor ( n20436 , n20426 , n20431 , n20435 );
nand ( n20437 , n20420 , n20436 );
buf ( n20438 , n20409 );
and ( n20439 , n901 , n20438 );
not ( n20440 , n20416 );
not ( n20441 , n20440 );
and ( n20442 , n656 , n20441 );
nor ( n20443 , n20439 , n20442 );
not ( n20444 , n20424 );
and ( n20445 , n673 , n20444 );
not ( n20446 , n20428 );
not ( n20447 , n20446 );
and ( n20448 , n551 , n20447 );
not ( n20449 , n20432 );
not ( n20450 , n20449 );
and ( n20451 , n474 , n20450 );
nor ( n20452 , n20445 , n20448 , n20451 );
nand ( n20453 , n20443 , n20452 );
nor ( n20454 , n890 , n912 , n916 , n917 );
and ( n20455 , n19919 , n20454 );
nand ( n20456 , n893 , n919 );
nand ( n20457 , n20456 , n19919 );
not ( n20458 , n20457 );
not ( n20459 , n19393 );
nor ( n20460 , n20455 , n20458 , n20459 );
and ( n20461 , n926 , n20438 );
and ( n20462 , n1384 , n20441 );
nor ( n20463 , n20461 , n20462 );
and ( n20464 , n1180 , n20444 );
not ( n20465 , n20428 );
not ( n20466 , n20465 );
and ( n20467 , n1262 , n20466 );
not ( n20468 , n20449 );
and ( n20469 , n1154 , n20468 );
nor ( n20470 , n20464 , n20467 , n20469 );
nand ( n20471 , n20463 , n20470 );
not ( n20472 , n20411 );
and ( n20473 , n929 , n20472 );
and ( n20474 , n1390 , n20441 );
nor ( n20475 , n20473 , n20474 );
and ( n20476 , n1203 , n20444 );
and ( n20477 , n1159 , n20466 );
and ( n20478 , n1381 , n20468 );
nor ( n20479 , n20476 , n20477 , n20478 );
nand ( n20480 , n20475 , n20479 );
and ( n20481 , n934 , n20472 );
buf ( n20482 , n20415 );
not ( n20483 , n20482 );
and ( n20484 , n1097 , n20483 );
nor ( n20485 , n20481 , n20484 );
and ( n20486 , n1122 , n20444 );
not ( n20487 , n20465 );
and ( n20488 , n1070 , n20487 );
and ( n20489 , n991 , n20450 );
nor ( n20490 , n20486 , n20488 , n20489 );
nand ( n20491 , n20485 , n20490 );
not ( n20492 , n20411 );
and ( n20493 , n940 , n20492 );
not ( n20494 , n20417 );
and ( n20495 , n649 , n20494 );
nor ( n20496 , n20493 , n20495 );
not ( n20497 , n20424 );
and ( n20498 , n722 , n20497 );
not ( n20499 , n20428 );
not ( n20500 , n20499 );
and ( n20501 , n741 , n20500 );
and ( n20502 , n466 , n20434 );
nor ( n20503 , n20498 , n20501 , n20502 );
nand ( n20504 , n20496 , n20503 );
and ( n20505 , n959 , n20438 );
and ( n20506 , n761 , n20418 );
nor ( n20507 , n20505 , n20506 );
and ( n20508 , n686 , n20497 );
and ( n20509 , n688 , n20430 );
not ( n20510 , n20433 );
and ( n20511 , n587 , n20510 );
nor ( n20512 , n20508 , n20509 , n20511 );
nand ( n20513 , n20507 , n20512 );
and ( n20514 , n969 , n20438 );
and ( n20515 , n701 , n20483 );
nor ( n20516 , n20514 , n20515 );
and ( n20517 , n810 , n20444 );
and ( n20518 , n618 , n20487 );
not ( n20519 , n20432 );
not ( n20520 , n20519 );
and ( n20521 , n520 , n20520 );
nor ( n20522 , n20517 , n20518 , n20521 );
nand ( n20523 , n20516 , n20522 );
and ( n20524 , n982 , n20412 );
not ( n20525 , n20440 );
and ( n20526 , n634 , n20525 );
nor ( n20527 , n20524 , n20526 );
and ( n20528 , n781 , n20497 );
not ( n20529 , n20428 );
not ( n20530 , n20529 );
and ( n20531 , n536 , n20530 );
and ( n20532 , n464 , n20510 );
nor ( n20533 , n20528 , n20531 , n20532 );
nand ( n20534 , n20527 , n20533 );
and ( n20535 , n986 , n20412 );
and ( n20536 , n713 , n20525 );
nor ( n20537 , n20535 , n20536 );
and ( n20538 , n823 , n20497 );
and ( n20539 , n632 , n20530 );
and ( n20540 , n533 , n20520 );
nor ( n20541 , n20538 , n20539 , n20540 );
nand ( n20542 , n20537 , n20541 );
and ( n20543 , n988 , n20492 );
and ( n20544 , n1160 , n20525 );
nor ( n20545 , n20543 , n20544 );
and ( n20546 , n1366 , n20425 );
and ( n20547 , n1255 , n20500 );
and ( n20548 , n1364 , n20520 );
nor ( n20549 , n20546 , n20547 , n20548 );
nand ( n20550 , n20545 , n20549 );
and ( n20551 , n989 , n20438 );
and ( n20552 , n1402 , n20525 );
nor ( n20553 , n20551 , n20552 );
and ( n20554 , n1372 , n20425 );
and ( n20555 , n1257 , n20500 );
and ( n20556 , n1397 , n20510 );
nor ( n20557 , n20554 , n20555 , n20556 );
nand ( n20558 , n20553 , n20557 );
and ( n20559 , n1002 , n20438 );
and ( n20560 , n1274 , n20525 );
nor ( n20561 , n20559 , n20560 );
and ( n20562 , n1243 , n20425 );
not ( n20563 , n20429 );
and ( n20564 , n1207 , n20563 );
and ( n20565 , n1153 , n20434 );
nor ( n20566 , n20562 , n20564 , n20565 );
nand ( n20567 , n20561 , n20566 );
not ( n20568 , n2 );
or ( n20569 , n20568 , n1569 );
nand ( n20570 , n141 , n224 );
not ( n20571 , n13222 );
nor ( n20572 , n1640 , n20570 , n20571 );
and ( n20573 , n1559 , n20572 );
nor ( n20574 , n20573 , n1087 );
nor ( n20575 , n20569 , n20574 );
not ( n20576 , n2 );
or ( n20577 , n20576 , n1566 );
and ( n20578 , n1576 , n20572 );
nor ( n20579 , n20578 , n1088 );
nor ( n20580 , n20577 , n20579 );
not ( n20581 , n2 );
or ( n20582 , n20581 , n1602 );
and ( n20583 , n1609 , n20572 );
nor ( n20584 , n20583 , n1086 );
nor ( n20585 , n20582 , n20584 );
not ( n20586 , n2 );
or ( n20587 , n20586 , n1568 );
and ( n20588 , n1588 , n20572 );
nor ( n20589 , n20588 , n1099 );
nor ( n20590 , n20587 , n20589 );
not ( n20591 , n20423 );
and ( n20592 , n762 , n20591 );
not ( n20593 , n20440 );
and ( n20594 , n590 , n20593 );
nor ( n20595 , n20592 , n20594 );
not ( n20596 , n20410 );
and ( n20597 , n985 , n20596 );
not ( n20598 , n20446 );
and ( n20599 , n486 , n20598 );
not ( n20600 , n20433 );
and ( n20601 , n456 , n20600 );
nor ( n20602 , n20597 , n20599 , n20601 );
nand ( n20603 , n20595 , n20602 );
or ( n20604 , n16525 , n13538 , n19396 );
not ( n20605 , n754 );
nand ( n20606 , n135 , n137 , n1608 );
not ( n20607 , n20606 );
and ( n20608 , n20605 , n20607 );
not ( n20609 , n15378 );
nor ( n20610 , n20608 , n20609 );
or ( n20611 , n267 , n20610 , n19401 );
nand ( n20612 , n20604 , n20611 );
buf ( n20613 , n13222 );
and ( n20614 , n905 , n20613 );
nor ( n20615 , n20614 , n1599 );
not ( n20616 , n13573 );
buf ( n20617 , n18010 );
not ( n20618 , n20613 );
nand ( n20619 , n153 , n20617 , n20618 );
nand ( n20620 , n20615 , n20616 , n20619 );
and ( n20621 , n394 , n20494 );
and ( n20622 , n393 , n20520 );
nor ( n20623 , n20621 , n20622 );
buf ( n20624 , n20409 );
and ( n20625 , n254 , n20624 );
not ( n20626 , n20423 );
and ( n20627 , n395 , n20626 );
not ( n20628 , n20499 );
and ( n20629 , n378 , n20628 );
nor ( n20630 , n20625 , n20627 , n20629 );
nand ( n20631 , n20623 , n20630 );
buf ( n20632 , n1003 );
buf ( n20633 , n20632 );
not ( n20634 , n20633 );
not ( n20635 , n20634 );
not ( n20636 , n20635 );
nand ( n20637 , n365 , n20636 );
nor ( n20638 , n14593 , n14572 );
not ( n20639 , n20638 );
nor ( n20640 , n19930 , n20639 );
nand ( n20641 , n350 , n20640 );
not ( n20642 , n20641 );
nand ( n20643 , n20642 , n370 );
nor ( n20644 , n14549 , n19944 , n20643 );
or ( n20645 , n365 , n20644 );
and ( n20646 , n365 , n20644 );
not ( n20647 , n20635 );
nor ( n20648 , n20646 , n20647 );
nand ( n20649 , n20645 , n20648 );
and ( n20650 , n20637 , n20649 );
not ( n20651 , n2 );
or ( n20652 , n20651 , n226 );
nor ( n20653 , n20650 , n20652 );
and ( n20654 , n514 , n20472 );
and ( n20655 , n1026 , n20520 );
nor ( n20656 , n20654 , n20655 );
not ( n20657 , n20417 );
and ( n20658 , n1028 , n20657 );
and ( n20659 , n1027 , n20626 );
not ( n20660 , n20429 );
and ( n20661 , n1025 , n20660 );
nor ( n20662 , n20658 , n20659 , n20661 );
nand ( n20663 , n20656 , n20662 );
not ( n20664 , n17311 );
nor ( n20665 , n20664 , n17268 );
or ( n20666 , n20665 , n17308 );
and ( n20667 , n20665 , n17308 );
nor ( n20668 , n20667 , n14981 );
and ( n20669 , n20666 , n20668 );
and ( n20670 , n611 , n14981 );
nor ( n20671 , n20669 , n20670 );
or ( n20672 , n1819 , n20671 );
and ( n20673 , n611 , n17334 );
nor ( n20674 , n20673 , n17335 );
or ( n20675 , n14974 , n20674 );
nand ( n20676 , n20672 , n20675 );
and ( n20677 , n1251 , n20676 );
or ( n20678 , n15002 , n15874 );
and ( n20679 , n15003 , n15023 );
or ( n20680 , n20679 , n15865 );
and ( n20681 , n20679 , n15865 );
nor ( n20682 , n20681 , n14979 );
nand ( n20683 , n20680 , n20682 );
nand ( n20684 , n20678 , n20683 );
and ( n20685 , n14974 , n20684 );
and ( n20686 , n15887 , n638 );
not ( n20687 , n15887 );
and ( n20688 , n20687 , n15002 );
nor ( n20689 , n20686 , n20688 );
and ( n20690 , n1819 , n20689 );
nor ( n20691 , n20685 , n20690 );
nor ( n20692 , n14973 , n20691 );
and ( n20693 , n887 , n20438 );
and ( n20694 , n585 , n20494 );
nor ( n20695 , n20693 , n20694 );
not ( n20696 , n20423 );
and ( n20697 , n765 , n20696 );
and ( n20698 , n498 , n20563 );
and ( n20699 , n451 , n20510 );
nor ( n20700 , n20697 , n20698 , n20699 );
nand ( n20701 , n20695 , n20700 );
not ( n20702 , n17392 );
nor ( n20703 , n20702 , n17348 );
or ( n20704 , n20703 , n17389 );
and ( n20705 , n20703 , n17389 );
nor ( n20706 , n20705 , n15711 );
and ( n20707 , n20704 , n20706 );
and ( n20708 , n694 , n17198 );
nor ( n20709 , n20707 , n20708 );
or ( n20710 , n1808 , n20709 );
and ( n20711 , n694 , n17415 );
nor ( n20712 , n20711 , n17416 );
or ( n20713 , n15704 , n20712 );
nand ( n20714 , n20710 , n20713 );
and ( n20715 , n1260 , n20714 );
or ( n20716 , n19413 , n17197 );
and ( n20717 , n15746 , n15737 );
or ( n20718 , n20717 , n15767 );
and ( n20719 , n20717 , n15767 );
nor ( n20720 , n20719 , n17196 );
nand ( n20721 , n20718 , n20720 );
nand ( n20722 , n20716 , n20721 );
and ( n20723 , n15704 , n20722 );
and ( n20724 , n15794 , n751 );
not ( n20725 , n15794 );
and ( n20726 , n20725 , n19413 );
nor ( n20727 , n20724 , n20726 );
and ( n20728 , n1808 , n20727 );
nor ( n20729 , n20723 , n20728 );
nor ( n20730 , n15703 , n20729 );
not ( n20731 , n17655 );
nor ( n20732 , n20731 , n17610 );
or ( n20733 , n20732 , n17652 );
and ( n20734 , n20732 , n17652 );
nor ( n20735 , n20734 , n18627 );
and ( n20736 , n20733 , n20735 );
and ( n20737 , n760 , n15098 );
nor ( n20738 , n20736 , n20737 );
or ( n20739 , n1826 , n20738 );
and ( n20740 , n760 , n17679 );
nor ( n20741 , n20740 , n17680 );
or ( n20742 , n15090 , n20741 );
nand ( n20743 , n20739 , n20742 );
and ( n20744 , n1272 , n20743 );
not ( n20745 , n20416 );
not ( n20746 , n20745 );
and ( n20747 , n588 , n20746 );
not ( n20748 , n20428 );
not ( n20749 , n20748 );
and ( n20750 , n500 , n20749 );
not ( n20751 , n20432 );
not ( n20752 , n20751 );
and ( n20753 , n453 , n20752 );
nor ( n20754 , n20747 , n20750 , n20753 );
buf ( n20755 , n20423 );
not ( n20756 , n20755 );
and ( n20757 , n687 , n20756 );
and ( n20758 , n886 , n20438 );
nor ( n20759 , n20757 , n20758 );
nand ( n20760 , n20754 , n20759 );
or ( n20761 , n15119 , n15097 );
and ( n20762 , n15120 , n15139 );
or ( n20763 , n20762 , n15819 );
and ( n20764 , n20762 , n15819 );
nor ( n20765 , n20764 , n15096 );
nand ( n20766 , n20763 , n20765 );
nand ( n20767 , n20761 , n20766 );
and ( n20768 , n15090 , n20767 );
and ( n20769 , n15840 , n783 );
not ( n20770 , n15840 );
and ( n20771 , n20770 , n15119 );
nor ( n20772 , n20769 , n20771 );
and ( n20773 , n1826 , n20772 );
nor ( n20774 , n20768 , n20773 );
nor ( n20775 , n15089 , n20774 );
and ( n20776 , n975 , n13633 );
and ( n20777 , n976 , n13623 );
nor ( n20778 , n20776 , n20777 );
nand ( n20779 , n975 , n976 );
and ( n20780 , n20778 , n20779 , n13690 );
and ( n20781 , n880 , n18833 );
and ( n20782 , n974 , n18835 );
nor ( n20783 , n20781 , n20782 );
nand ( n20784 , n880 , n974 );
not ( n20785 , n20784 );
and ( n20786 , n13675 , n20785 );
and ( n20787 , n974 , n13675 );
and ( n20788 , n880 , n18835 );
nor ( n20789 , n20787 , n20788 );
and ( n20790 , n20789 , n20784 , n13683 );
not ( n20791 , n13668 );
and ( n20792 , n971 , n20791 );
and ( n20793 , n971 , n13660 );
and ( n20794 , n973 , n13664 );
nor ( n20795 , n20793 , n20794 );
nand ( n20796 , n971 , n973 );
and ( n20797 , n20795 , n20796 , n13668 );
not ( n20798 , n883 );
nand ( n20799 , n879 , n20798 );
and ( n20800 , n970 , n20799 );
and ( n20801 , n883 , n13643 );
nor ( n20802 , n20800 , n20801 , n13641 );
nor ( n20803 , n20797 , n20802 );
or ( n20804 , n933 , n20796 );
not ( n20805 , n973 );
or ( n20806 , n20805 , n935 );
nand ( n20807 , n20804 , n20806 );
nor ( n20808 , n20792 , n20803 , n20807 );
nor ( n20809 , n20790 , n20808 );
nor ( n20810 , n20786 , n20809 );
and ( n20811 , n20783 , n20810 );
nor ( n20812 , n20780 , n20811 );
not ( n20813 , n978 );
nand ( n20814 , n20813 , n1006 );
not ( n20815 , n13285 );
not ( n20816 , n939 );
and ( n20817 , n20815 , n20816 );
not ( n20818 , n877 );
nor ( n20819 , n20818 , n888 );
nor ( n20820 , n20817 , n20819 );
nand ( n20821 , n877 , n977 );
nand ( n20822 , n20820 , n20821 , n18807 );
and ( n20823 , n20812 , n20814 , n20822 );
nor ( n20824 , n979 , n981 );
or ( n20825 , n939 , n20821 );
or ( n20826 , n13285 , n888 );
or ( n20827 , n13307 , n13690 );
or ( n20828 , n937 , n20779 );
not ( n20829 , n976 );
or ( n20830 , n20829 , n938 );
nand ( n20831 , n20827 , n20828 , n20830 );
and ( n20832 , n20822 , n20831 );
and ( n20833 , n877 , n13620 );
nor ( n20834 , n20832 , n20833 );
nand ( n20835 , n20825 , n20826 , n20834 );
and ( n20836 , n20814 , n20835 );
and ( n20837 , n978 , n12538 );
nor ( n20838 , n20836 , n20837 , n878 );
nand ( n20839 , n20824 , n20838 );
nor ( n20840 , n20823 , n20839 );
not ( n20841 , n16267 );
or ( n20842 , n16277 , n20841 );
not ( n20843 , n16278 );
nor ( n20844 , n20843 , n16725 );
or ( n20845 , n20844 , n16421 );
and ( n20846 , n20844 , n16421 );
nor ( n20847 , n20846 , n16265 );
nand ( n20848 , n20845 , n20847 );
nand ( n20849 , n20842 , n20848 );
and ( n20850 , n16258 , n20849 );
and ( n20851 , n16440 , n837 );
not ( n20852 , n16440 );
and ( n20853 , n20852 , n16277 );
nor ( n20854 , n20851 , n20853 );
and ( n20855 , n1828 , n20854 );
nor ( n20856 , n20850 , n20855 );
nor ( n20857 , n16257 , n20856 );
not ( n20858 , n17576 );
nor ( n20859 , n20858 , n17533 );
or ( n20860 , n20859 , n17573 );
and ( n20861 , n20859 , n17573 );
nor ( n20862 , n20861 , n16347 );
and ( n20863 , n20860 , n20862 );
and ( n20864 , n849 , n20106 );
nor ( n20865 , n20863 , n20864 );
or ( n20866 , n1828 , n20865 );
and ( n20867 , n849 , n17599 );
nor ( n20868 , n20867 , n17600 );
or ( n20869 , n16258 , n20868 );
nand ( n20870 , n20866 , n20869 );
and ( n20871 , n1240 , n20870 );
and ( n20872 , n710 , n20746 );
not ( n20873 , n20529 );
and ( n20874 , n630 , n20873 );
not ( n20875 , n20449 );
and ( n20876 , n506 , n20875 );
nor ( n20877 , n20872 , n20874 , n20876 );
not ( n20878 , n20755 );
and ( n20879 , n833 , n20878 );
and ( n20880 , n878 , n20624 );
nor ( n20881 , n20879 , n20880 );
nand ( n20882 , n20877 , n20881 );
not ( n20883 , n177 );
not ( n20884 , n12852 );
not ( n20885 , n20884 );
or ( n20886 , n20883 , n20885 );
and ( n20887 , n876 , n12852 );
nor ( n20888 , n20887 , n13199 );
nand ( n20889 , n20886 , n20888 );
not ( n20890 , n20482 );
and ( n20891 , n709 , n20890 );
not ( n20892 , n20748 );
and ( n20893 , n626 , n20892 );
not ( n20894 , n20751 );
and ( n20895 , n527 , n20894 );
nor ( n20896 , n20891 , n20893 , n20895 );
and ( n20897 , n796 , n20756 );
and ( n20898 , n877 , n20438 );
nor ( n20899 , n20897 , n20898 );
nand ( n20900 , n20896 , n20899 );
and ( n20901 , n879 , n20438 );
and ( n20902 , n1400 , n20483 );
nor ( n20903 , n20901 , n20902 );
not ( n20904 , n20423 );
and ( n20905 , n1233 , n20904 );
and ( n20906 , n1221 , n20447 );
and ( n20907 , n1409 , n20468 );
nor ( n20908 , n20905 , n20906 , n20907 );
nand ( n20909 , n20903 , n20908 );
not ( n20910 , n20482 );
and ( n20911 , n707 , n20910 );
not ( n20912 , n20429 );
and ( n20913 , n623 , n20912 );
not ( n20914 , n20751 );
and ( n20915 , n507 , n20914 );
nor ( n20916 , n20911 , n20913 , n20915 );
and ( n20917 , n797 , n20878 );
and ( n20918 , n880 , n20438 );
nor ( n20919 , n20917 , n20918 );
nand ( n20920 , n20916 , n20919 );
not ( n20921 , n20755 );
and ( n20922 , n764 , n20921 );
and ( n20923 , n583 , n20483 );
nor ( n20924 , n20922 , n20923 );
not ( n20925 , n20409 );
not ( n20926 , n20925 );
and ( n20927 , n881 , n20926 );
not ( n20928 , n20465 );
and ( n20929 , n495 , n20928 );
not ( n20930 , n20432 );
not ( n20931 , n20930 );
and ( n20932 , n447 , n20931 );
nor ( n20933 , n20927 , n20929 , n20932 );
nand ( n20934 , n20924 , n20933 );
and ( n20935 , n884 , n20472 );
and ( n20936 , n1387 , n20441 );
nor ( n20937 , n20935 , n20936 );
and ( n20938 , n1236 , n20904 );
and ( n20939 , n1157 , n20466 );
not ( n20940 , n20930 );
and ( n20941 , n1401 , n20940 );
nor ( n20942 , n20938 , n20939 , n20941 );
nand ( n20943 , n20937 , n20942 );
and ( n20944 , n885 , n20412 );
and ( n20945 , n660 , n20657 );
nor ( n20946 , n20944 , n20945 );
and ( n20947 , n738 , n20696 );
and ( n20948 , n554 , n20563 );
and ( n20949 , n477 , n20434 );
nor ( n20950 , n20947 , n20948 , n20949 );
nand ( n20951 , n20946 , n20950 );
and ( n20952 , n888 , n20438 );
and ( n20953 , n1163 , n20483 );
nor ( n20954 , n20952 , n20953 );
and ( n20955 , n1239 , n20904 );
and ( n20956 , n1158 , n20466 );
and ( n20957 , n1396 , n20450 );
nor ( n20958 , n20955 , n20956 , n20957 );
nand ( n20959 , n20954 , n20958 );
and ( n20960 , n671 , n20921 );
and ( n20961 , n657 , n20483 );
nor ( n20962 , n20960 , n20961 );
not ( n20963 , n20925 );
and ( n20964 , n891 , n20963 );
and ( n20965 , n745 , n20928 );
and ( n20966 , n648 , n20940 );
nor ( n20967 , n20964 , n20965 , n20966 );
nand ( n20968 , n20962 , n20967 );
and ( n20969 , n1121 , n20921 );
and ( n20970 , n1096 , n20483 );
nor ( n20971 , n20969 , n20970 );
and ( n20972 , n896 , n20926 );
and ( n20973 , n1067 , n20928 );
and ( n20974 , n990 , n20940 );
nor ( n20975 , n20972 , n20973 , n20974 );
nand ( n20976 , n20971 , n20975 );
not ( n20977 , n179 );
not ( n20978 , n20884 );
or ( n20979 , n20977 , n20978 );
and ( n20980 , n906 , n12852 );
nor ( n20981 , n20980 , n13199 );
nand ( n20982 , n20979 , n20981 );
not ( n20983 , n189 );
not ( n20984 , n20884 );
or ( n20985 , n20983 , n20984 );
and ( n20986 , n907 , n12852 );
nor ( n20987 , n20986 , n13199 );
nand ( n20988 , n20985 , n20987 );
not ( n20989 , n181 );
not ( n20990 , n20884 );
or ( n20991 , n20989 , n20990 );
and ( n20992 , n908 , n12852 );
nor ( n20993 , n20992 , n13199 );
nand ( n20994 , n20991 , n20993 );
and ( n20995 , n909 , n20492 );
and ( n20996 , n1354 , n20525 );
nor ( n20997 , n20995 , n20996 );
and ( n20998 , n1293 , n20696 );
and ( n20999 , n1335 , n20430 );
and ( n21000 , n1313 , n20434 );
nor ( n21001 , n20998 , n20999 , n21000 );
nand ( n21002 , n20997 , n21001 );
and ( n21003 , n1272 , n20910 );
and ( n21004 , n1260 , n20749 );
not ( n21005 , n20449 );
and ( n21006 , n1251 , n21005 );
nor ( n21007 , n21003 , n21004 , n21006 );
and ( n21008 , n1240 , n20756 );
and ( n21009 , n925 , n20438 );
nor ( n21010 , n21008 , n21009 );
nand ( n21011 , n21007 , n21010 );
not ( n21012 , n20482 );
and ( n21013 , n1269 , n21012 );
not ( n21014 , n20499 );
and ( n21015 , n1213 , n21014 );
not ( n21016 , n20519 );
and ( n21017 , n1249 , n21016 );
nor ( n21018 , n21013 , n21015 , n21017 );
and ( n21019 , n1232 , n20921 );
not ( n21020 , n20925 );
and ( n21021 , n924 , n21020 );
nor ( n21022 , n21019 , n21021 );
nand ( n21023 , n21018 , n21022 );
and ( n21024 , n1467 , n20591 );
and ( n21025 , n1471 , n20593 );
nor ( n21026 , n21024 , n21025 );
and ( n21027 , n935 , n20596 );
and ( n21028 , n1439 , n20598 );
and ( n21029 , n1406 , n20600 );
nor ( n21030 , n21027 , n21028 , n21029 );
nand ( n21031 , n21026 , n21030 );
and ( n21032 , n936 , n20438 );
and ( n21033 , n1270 , n20483 );
nor ( n21034 , n21032 , n21033 );
and ( n21035 , n1235 , n20904 );
and ( n21036 , n1258 , n20487 );
and ( n21037 , n1152 , n20450 );
nor ( n21038 , n21035 , n21036 , n21037 );
nand ( n21039 , n21034 , n21038 );
and ( n21040 , n938 , n20492 );
and ( n21041 , n1271 , n20494 );
nor ( n21042 , n21040 , n21041 );
and ( n21043 , n1210 , n20696 );
and ( n21044 , n1259 , n20563 );
and ( n21045 , n1403 , n20434 );
nor ( n21046 , n21043 , n21044 , n21045 );
nand ( n21047 , n21042 , n21046 );
not ( n21048 , n20755 );
and ( n21049 , n1238 , n21048 );
and ( n21050 , n1394 , n20483 );
nor ( n21051 , n21049 , n21050 );
and ( n21052 , n939 , n20624 );
and ( n21053 , n1205 , n20447 );
and ( n21054 , n1399 , n20931 );
nor ( n21055 , n21052 , n21053 , n21054 );
nand ( n21056 , n21051 , n21055 );
not ( n21057 , n20745 );
and ( n21058 , n580 , n21057 );
not ( n21059 , n20429 );
and ( n21060 , n493 , n21059 );
and ( n21061 , n445 , n21005 );
nor ( n21062 , n21058 , n21060 , n21061 );
and ( n21063 , n680 , n20878 );
and ( n21064 , n941 , n20438 );
nor ( n21065 , n21063 , n21064 );
nand ( n21066 , n21062 , n21065 );
and ( n21067 , n943 , n20472 );
and ( n21068 , n568 , n20441 );
nor ( n21069 , n21067 , n21068 );
and ( n21070 , n730 , n20904 );
and ( n21071 , n742 , n20487 );
and ( n21072 , n645 , n20468 );
nor ( n21073 , n21070 , n21071 , n21072 );
nand ( n21074 , n21069 , n21073 );
and ( n21075 , n683 , n21048 );
and ( n21076 , n582 , n20483 );
nor ( n21077 , n21075 , n21076 );
and ( n21078 , n944 , n20963 );
and ( n21079 , n494 , n20447 );
and ( n21080 , n446 , n20931 );
nor ( n21081 , n21078 , n21079 , n21080 );
nand ( n21082 , n21077 , n21081 );
and ( n21083 , n685 , n21048 );
and ( n21084 , n584 , n20483 );
nor ( n21085 , n21083 , n21084 );
and ( n21086 , n945 , n20624 );
not ( n21087 , n20465 );
and ( n21088 , n497 , n21087 );
and ( n21089 , n449 , n20940 );
nor ( n21090 , n21086 , n21088 , n21089 );
nand ( n21091 , n21085 , n21090 );
and ( n21092 , n650 , n20746 );
not ( n21093 , n20529 );
and ( n21094 , n543 , n21093 );
and ( n21095 , n646 , n21005 );
nor ( n21096 , n21092 , n21094 , n21095 );
and ( n21097 , n724 , n20591 );
and ( n21098 , n946 , n20438 );
nor ( n21099 , n21097 , n21098 );
nand ( n21100 , n21096 , n21099 );
and ( n21101 , n947 , n20438 );
and ( n21102 , n651 , n20418 );
nor ( n21103 , n21101 , n21102 );
and ( n21104 , n725 , n20696 );
and ( n21105 , n743 , n20500 );
and ( n21106 , n647 , n20510 );
nor ( n21107 , n21104 , n21105 , n21106 );
nand ( n21108 , n21103 , n21107 );
not ( n21109 , n20745 );
and ( n21110 , n573 , n21109 );
and ( n21111 , n545 , n21014 );
and ( n21112 , n468 , n21016 );
nor ( n21113 , n21110 , n21111 , n21112 );
and ( n21114 , n727 , n21048 );
and ( n21115 , n948 , n21020 );
nor ( n21116 , n21114 , n21115 );
nand ( n21117 , n21113 , n21116 );
not ( n21118 , n20482 );
and ( n21119 , n658 , n21118 );
and ( n21120 , n546 , n21059 );
and ( n21121 , n469 , n20752 );
nor ( n21122 , n21119 , n21120 , n21121 );
and ( n21123 , n728 , n20878 );
and ( n21124 , n949 , n20438 );
nor ( n21125 , n21123 , n21124 );
nand ( n21126 , n21122 , n21125 );
and ( n21127 , n733 , n20591 );
and ( n21128 , n654 , n20657 );
nor ( n21129 , n21127 , n21128 );
and ( n21130 , n951 , n20596 );
and ( n21131 , n665 , n20598 );
not ( n21132 , n20930 );
and ( n21133 , n567 , n21132 );
nor ( n21134 , n21130 , n21131 , n21133 );
nand ( n21135 , n21129 , n21134 );
and ( n21136 , n786 , n20910 );
and ( n21137 , n549 , n20628 );
and ( n21138 , n472 , n20894 );
nor ( n21139 , n21136 , n21137 , n21138 );
and ( n21140 , n731 , n20878 );
and ( n21141 , n952 , n20624 );
nor ( n21142 , n21140 , n21141 );
nand ( n21143 , n21139 , n21142 );
and ( n21144 , n735 , n21048 );
and ( n21145 , n758 , n20483 );
nor ( n21146 , n21144 , n21145 );
and ( n21147 , n954 , n20963 );
and ( n21148 , n561 , n21087 );
and ( n21149 , n475 , n20940 );
nor ( n21150 , n21147 , n21148 , n21149 );
nand ( n21151 , n21146 , n21150 );
and ( n21152 , n955 , n20438 );
and ( n21153 , n787 , n20418 );
nor ( n21154 , n21152 , n21153 );
and ( n21155 , n734 , n20696 );
and ( n21156 , n552 , n20530 );
and ( n21157 , n443 , n20520 );
nor ( n21158 , n21155 , n21156 , n21157 );
nand ( n21159 , n21154 , n21158 );
and ( n21160 , n556 , n21109 );
and ( n21161 , n479 , n21014 );
not ( n21162 , n20519 );
and ( n21163 , n440 , n21162 );
nor ( n21164 , n21160 , n21161 , n21163 );
and ( n21165 , n644 , n20921 );
and ( n21166 , n956 , n21020 );
nor ( n21167 , n21165 , n21166 );
nand ( n21168 , n21164 , n21167 );
not ( n21169 , n20482 );
and ( n21170 , n755 , n21169 );
and ( n21171 , n663 , n20628 );
not ( n21172 , n20751 );
and ( n21173 , n564 , n21172 );
nor ( n21174 , n21170 , n21171 , n21173 );
and ( n21175 , n736 , n20756 );
and ( n21176 , n957 , n20624 );
nor ( n21177 , n21175 , n21176 );
nand ( n21178 , n21174 , n21177 );
not ( n21179 , n20482 );
and ( n21180 , n769 , n21179 );
and ( n21181 , n677 , n20873 );
and ( n21182 , n576 , n21172 );
nor ( n21183 , n21180 , n21181 , n21182 );
and ( n21184 , n676 , n20756 );
and ( n21185 , n960 , n20438 );
nor ( n21186 , n21184 , n21185 );
nand ( n21187 , n21183 , n21186 );
and ( n21188 , n578 , n21012 );
not ( n21189 , n20446 );
and ( n21190 , n491 , n21189 );
and ( n21191 , n450 , n21016 );
nor ( n21192 , n21188 , n21190 , n21191 );
and ( n21193 , n679 , n21048 );
and ( n21194 , n961 , n21020 );
nor ( n21195 , n21193 , n21194 );
nand ( n21196 , n21192 , n21195 );
and ( n21197 , n740 , n20921 );
and ( n21198 , n788 , n20441 );
nor ( n21199 , n21197 , n21198 );
and ( n21200 , n963 , n20926 );
and ( n21201 , n555 , n21087 );
and ( n21202 , n442 , n20931 );
nor ( n21203 , n21200 , n21201 , n21202 );
nand ( n21204 , n21199 , n21203 );
and ( n21205 , n699 , n21057 );
and ( n21206 , n616 , n20749 );
and ( n21207 , n518 , n20875 );
nor ( n21208 , n21205 , n21206 , n21207 );
and ( n21209 , n799 , n20756 );
and ( n21210 , n964 , n20624 );
nor ( n21211 , n21209 , n21210 );
nand ( n21212 , n21208 , n21211 );
not ( n21213 , n20482 );
and ( n21214 , n589 , n21213 );
and ( n21215 , n501 , n20530 );
and ( n21216 , n454 , n21162 );
nor ( n21217 , n21214 , n21215 , n21216 );
and ( n21218 , n767 , n20921 );
and ( n21219 , n965 , n21020 );
nor ( n21220 , n21218 , n21219 );
nand ( n21221 , n21217 , n21220 );
and ( n21222 , n672 , n21109 );
and ( n21223 , n619 , n21189 );
and ( n21224 , n521 , n21162 );
nor ( n21225 , n21222 , n21223 , n21224 );
and ( n21226 , n811 , n21048 );
and ( n21227 , n970 , n21020 );
nor ( n21228 , n21226 , n21227 );
nand ( n21229 , n21225 , n21228 );
and ( n21230 , n704 , n21109 );
and ( n21231 , n569 , n21189 );
and ( n21232 , n523 , n21162 );
nor ( n21233 , n21230 , n21231 , n21232 );
and ( n21234 , n813 , n20921 );
and ( n21235 , n972 , n21020 );
nor ( n21236 , n21234 , n21235 );
nand ( n21237 , n21233 , n21236 );
and ( n21238 , n705 , n21109 );
and ( n21239 , n624 , n21189 );
and ( n21240 , n525 , n21162 );
nor ( n21241 , n21238 , n21239 , n21240 );
and ( n21242 , n815 , n21048 );
and ( n21243 , n974 , n21020 );
nor ( n21244 , n21242 , n21243 );
nand ( n21245 , n21241 , n21244 );
and ( n21246 , n816 , n21048 );
and ( n21247 , n706 , n20494 );
nor ( n21248 , n21246 , n21247 );
and ( n21249 , n975 , n20624 );
and ( n21250 , n575 , n21087 );
and ( n21251 , n528 , n20940 );
nor ( n21252 , n21249 , n21250 , n21251 );
nand ( n21253 , n21248 , n21252 );
and ( n21254 , n708 , n21169 );
and ( n21255 , n627 , n21093 );
and ( n21256 , n530 , n21172 );
nor ( n21257 , n21254 , n21255 , n21256 );
and ( n21258 , n819 , n20878 );
and ( n21259 , n977 , n20438 );
nor ( n21260 , n21258 , n21259 );
nand ( n21261 , n21257 , n21260 );
and ( n21262 , n668 , n21012 );
and ( n21263 , n574 , n21014 );
and ( n21264 , n529 , n21016 );
nor ( n21265 , n21262 , n21263 , n21264 );
and ( n21266 , n818 , n20921 );
and ( n21267 , n978 , n21020 );
nor ( n21268 , n21266 , n21267 );
nand ( n21269 , n21265 , n21268 );
and ( n21270 , n669 , n21213 );
and ( n21271 , n625 , n21014 );
and ( n21272 , n526 , n21016 );
nor ( n21273 , n21270 , n21271 , n21272 );
and ( n21274 , n817 , n21048 );
and ( n21275 , n976 , n21020 );
nor ( n21276 , n21274 , n21275 );
nand ( n21277 , n21273 , n21276 );
and ( n21278 , n633 , n21213 );
and ( n21279 , n535 , n21014 );
and ( n21280 , n463 , n21016 );
nor ( n21281 , n21278 , n21279 , n21280 );
and ( n21282 , n780 , n20921 );
and ( n21283 , n979 , n21020 );
nor ( n21284 , n21282 , n21283 );
nand ( n21285 , n21281 , n21284 );
and ( n21286 , n770 , n21048 );
and ( n21287 , n591 , n20494 );
nor ( n21288 , n21286 , n21287 );
and ( n21289 , n983 , n20926 );
and ( n21290 , n503 , n20447 );
and ( n21291 , n457 , n20931 );
nor ( n21292 , n21289 , n21290 , n21291 );
nand ( n21293 , n21288 , n21292 );
and ( n21294 , n652 , n21057 );
and ( n21295 , n544 , n20628 );
and ( n21296 , n467 , n20914 );
nor ( n21297 , n21294 , n21295 , n21296 );
and ( n21298 , n726 , n20591 );
and ( n21299 , n1000 , n20438 );
nor ( n21300 , n21298 , n21299 );
nand ( n21301 , n21297 , n21300 );
not ( n21302 , n895 );
not ( n21303 , n919 );
and ( n21304 , n21303 , n20454 );
not ( n21305 , n894 );
nor ( n21306 , n21304 , n21305 , n19921 );
not ( n21307 , n21306 );
and ( n21308 , n21302 , n21307 );
nor ( n21309 , n21308 , n20459 );
not ( n21310 , n180 );
not ( n21311 , n20884 );
or ( n21312 , n21310 , n21311 );
and ( n21313 , n1007 , n12852 );
nor ( n21314 , n21313 , n13199 );
nand ( n21315 , n21312 , n21314 );
and ( n21316 , n593 , n20746 );
and ( n21317 , n504 , n21059 );
and ( n21318 , n459 , n20914 );
nor ( n21319 , n21316 , n21317 , n21318 );
and ( n21320 , n753 , n20878 );
and ( n21321 , n1008 , n20438 );
nor ( n21322 , n21320 , n21321 );
nand ( n21323 , n21319 , n21322 );
and ( n21324 , n832 , n21048 );
and ( n21325 , n666 , n20483 );
nor ( n21326 , n21324 , n21325 );
and ( n21327 , n1009 , n20963 );
and ( n21328 , n631 , n20447 );
and ( n21329 , n489 , n20520 );
nor ( n21330 , n21327 , n21328 , n21329 );
nand ( n21331 , n21326 , n21330 );
and ( n21332 , n714 , n21169 );
and ( n21333 , n572 , n20892 );
not ( n21334 , n20449 );
and ( n21335 , n534 , n21334 );
nor ( n21336 , n21332 , n21333 , n21335 );
and ( n21337 , n822 , n20921 );
and ( n21338 , n987 , n20438 );
nor ( n21339 , n21337 , n21338 );
nand ( n21340 , n21336 , n21339 );
not ( n21341 , n2 );
or ( n21342 , n21341 , n88 );
not ( n21343 , n1083 );
not ( n21344 , n19378 );
or ( n21345 , n21343 , n21344 );
nand ( n21346 , n21345 , n15668 );
and ( n21347 , n21346 , n15676 );
or ( n21348 , n19389 , n406 , n15678 );
nand ( n21349 , n1001 , n1812 );
and ( n21350 , n1083 , n21349 , n20056 );
nor ( n21351 , n21350 , n15651 );
or ( n21352 , n21351 , n15606 );
nand ( n21353 , n21348 , n21352 );
nand ( n21354 , n1083 , n15616 , n15617 );
and ( n21355 , n15622 , n21354 );
nor ( n21356 , n21355 , n19381 );
nor ( n21357 , n21347 , n21353 , n21356 );
nor ( n21358 , n21342 , n21357 );
nor ( n21359 , n20457 , n20459 );
not ( n21360 , n19200 );
nand ( n21361 , n19204 , n19211 );
nand ( n21362 , n19217 , n21361 );
not ( n21363 , n21362 );
or ( n21364 , n21360 , n21363 );
nand ( n21365 , n21364 , n19222 );
and ( n21366 , n19199 , n21365 );
nor ( n21367 , n21366 , n19194 );
or ( n21368 , n16923 , n21367 );
and ( n21369 , n16923 , n16906 );
not ( n21370 , n19207 );
and ( n21371 , n19204 , n21370 );
nand ( n21372 , n19199 , n19200 , n21371 );
or ( n21373 , n21369 , n21372 );
and ( n21374 , n21367 , n21369 , n21372 );
not ( n21375 , n21367 );
and ( n21376 , n16907 , n21375 );
nor ( n21377 , n21374 , n21376 );
nand ( n21378 , n21368 , n21373 , n21377 );
not ( n21379 , n19244 );
nand ( n21380 , n19248 , n19255 );
nand ( n21381 , n19261 , n21380 );
not ( n21382 , n21381 );
or ( n21383 , n21379 , n21382 );
nand ( n21384 , n21383 , n19266 );
and ( n21385 , n19243 , n21384 );
nor ( n21386 , n21385 , n19238 );
or ( n21387 , n16994 , n21386 );
and ( n21388 , n16994 , n16977 );
not ( n21389 , n19251 );
and ( n21390 , n19248 , n21389 );
nand ( n21391 , n21390 , n19243 , n19244 );
or ( n21392 , n21388 , n21391 );
and ( n21393 , n21386 , n21388 , n21391 );
not ( n21394 , n21386 );
and ( n21395 , n16978 , n21394 );
nor ( n21396 , n21393 , n21395 );
nand ( n21397 , n21387 , n21392 , n21396 );
not ( n21398 , n19332 );
nand ( n21399 , n19336 , n19343 );
nand ( n21400 , n19349 , n21399 );
not ( n21401 , n21400 );
or ( n21402 , n21398 , n21401 );
nand ( n21403 , n21402 , n19354 );
and ( n21404 , n19331 , n21403 );
nor ( n21405 , n21404 , n19326 );
or ( n21406 , n17064 , n21405 );
and ( n21407 , n17064 , n17061 );
not ( n21408 , n19339 );
and ( n21409 , n19336 , n21408 );
nand ( n21410 , n21409 , n19332 , n19331 );
or ( n21411 , n21407 , n21410 );
not ( n21412 , n17061 );
not ( n21413 , n21405 );
and ( n21414 , n21412 , n21413 );
and ( n21415 , n21405 , n21407 , n21410 );
nor ( n21416 , n21414 , n21415 );
nand ( n21417 , n21406 , n21411 , n21416 );
not ( n21418 , n13749 );
nand ( n21419 , n932 , n21418 );
nand ( n21420 , n989 , n1608 );
nor ( n21421 , n931 , n21420 );
nand ( n21422 , n900 , n928 );
nand ( n21423 , n924 , n1608 );
nor ( n21424 , n21421 , n21422 , n21423 );
nor ( n21425 , n13516 , n21424 );
not ( n21426 , n21420 );
not ( n21427 , n932 );
not ( n21428 , n21423 );
nand ( n21429 , n21426 , n21427 , n21428 );
nor ( n21430 , n21422 , n21429 );
not ( n21431 , n21430 );
not ( n21432 , n13516 );
not ( n21433 , n21422 );
nand ( n21434 , n989 , n1608 );
nor ( n21435 , n21427 , n21434 );
nand ( n21436 , n21428 , n21433 , n21435 );
nand ( n21437 , n21432 , n21436 );
nand ( n21438 , n21431 , n21437 );
nor ( n21439 , n21425 , n21438 );
and ( n21440 , n21419 , n21439 );
and ( n21441 , n17119 , n21430 );
nor ( n21442 , n21425 , n21437 );
and ( n21443 , n21441 , n21442 );
nor ( n21444 , n21440 , n21443 );
nand ( n21445 , n1623 , n21439 );
not ( n21446 , n21429 );
not ( n21447 , n21442 );
not ( n21448 , n21430 );
not ( n21449 , n21437 );
not ( n21450 , n21449 );
or ( n21451 , n21448 , n21450 );
nand ( n21452 , n21451 , n21438 );
not ( n21453 , n21452 );
and ( n21454 , n16462 , n21446 , n21447 , n21453 );
not ( n21455 , n900 );
nand ( n21456 , n21454 , n931 , n21455 );
nand ( n21457 , n21444 , n21445 , n21456 );
nor ( n21458 , n16840 , n16891 );
not ( n21459 , n21458 );
not ( n21460 , n16889 );
or ( n21461 , n21459 , n21460 );
or ( n21462 , n21458 , n16889 );
nand ( n21463 , n21461 , n21462 );
not ( n21464 , n16924 );
nor ( n21465 , n21464 , n16913 );
not ( n21466 , n21465 );
not ( n21467 , n16962 );
or ( n21468 , n21466 , n21467 );
or ( n21469 , n21465 , n16962 );
nand ( n21470 , n21468 , n21469 );
not ( n21471 , n16995 );
nor ( n21472 , n21471 , n16984 );
not ( n21473 , n21472 );
not ( n21474 , n17033 );
or ( n21475 , n21473 , n21474 );
or ( n21476 , n21472 , n17033 );
nand ( n21477 , n21475 , n21476 );
not ( n21478 , n17065 );
nor ( n21479 , n21478 , n17054 );
not ( n21480 , n21479 );
not ( n21481 , n17103 );
or ( n21482 , n21480 , n21481 );
or ( n21483 , n21479 , n17103 );
nand ( n21484 , n21482 , n21483 );
and ( n21485 , n1371 , n21012 );
and ( n21486 , n1266 , n21189 );
and ( n21487 , n1253 , n21132 );
nor ( n21488 , n21485 , n21486 , n21487 );
and ( n21489 , n1247 , n20921 );
and ( n21490 , n928 , n21020 );
nor ( n21491 , n21489 , n21490 );
nand ( n21492 , n21488 , n21491 );
and ( n21493 , n712 , n20890 );
and ( n21494 , n629 , n21093 );
and ( n21495 , n532 , n20752 );
nor ( n21496 , n21493 , n21494 , n21495 );
and ( n21497 , n820 , n20878 );
and ( n21498 , n981 , n20438 );
nor ( n21499 , n21497 , n21498 );
nand ( n21500 , n21496 , n21499 );
and ( n21501 , n700 , n21057 );
and ( n21502 , n617 , n20873 );
and ( n21503 , n519 , n21334 );
nor ( n21504 , n21501 , n21502 , n21503 );
and ( n21505 , n809 , n20591 );
and ( n21506 , n966 , n20438 );
nor ( n21507 , n21505 , n21506 );
nand ( n21508 , n21504 , n21507 );
and ( n21509 , n962 , n20438 );
and ( n21510 , n565 , n20418 );
nor ( n21511 , n21509 , n21510 );
and ( n21512 , n739 , n20696 );
and ( n21513 , n485 , n20430 );
and ( n21514 , n478 , n20510 );
nor ( n21515 , n21512 , n21513 , n21514 );
nand ( n21516 , n21511 , n21515 );
not ( n21517 , n1045 );
nor ( n21518 , n21517 , n15618 , n19381 );
and ( n21519 , n21518 , n15616 , n15622 );
not ( n21520 , n889 );
nand ( n21521 , n1150 , n21520 );
not ( n21522 , n21521 );
and ( n21523 , n15588 , n15603 );
not ( n21524 , n20048 );
nand ( n21525 , n21522 , n21523 , n21524 );
or ( n21526 , n312 , n1045 );
nand ( n21527 , n21526 , n19391 );
or ( n21528 , n405 , n1045 );
and ( n21529 , n1124 , n15631 , n15582 , n15634 );
nand ( n21530 , n21528 , n21529 );
or ( n21531 , n1045 , n15649 );
not ( n21532 , n1150 );
nand ( n21533 , n889 , n21532 );
not ( n21534 , n21533 );
nand ( n21535 , n21534 , n21523 , n21524 );
not ( n21536 , n21535 );
nand ( n21537 , n21531 , n21536 );
nand ( n21538 , n21525 , n21527 , n21530 , n21537 );
nor ( n21539 , n21519 , n21538 );
nor ( n21540 , n21342 , n21539 );
and ( n21541 , n566 , n21048 );
and ( n21542 , n557 , n20494 );
nor ( n21543 , n21541 , n21542 );
and ( n21544 , n958 , n20624 );
and ( n21545 , n480 , n20928 );
and ( n21546 , n441 , n20931 );
nor ( n21547 , n21544 , n21545 , n21546 );
nand ( n21548 , n21543 , n21547 );
and ( n21549 , n579 , n21213 );
and ( n21550 , n496 , n20530 );
and ( n21551 , n448 , n21132 );
nor ( n21552 , n21549 , n21550 , n21551 );
and ( n21553 , n684 , n20921 );
and ( n21554 , n942 , n21020 );
nor ( n21555 , n21553 , n21554 );
nand ( n21556 , n21552 , n21555 );
and ( n21557 , n729 , n20591 );
and ( n21558 , n653 , n20657 );
nor ( n21559 , n21557 , n21558 );
and ( n21560 , n950 , n20596 );
and ( n21561 , n547 , n20500 );
and ( n21562 , n470 , n20600 );
nor ( n21563 , n21560 , n21561 , n21562 );
nand ( n21564 , n21559 , n21563 );
and ( n21565 , n1588 , n1655 );
buf ( n21566 , n21565 );
and ( n21567 , n1342 , n21566 );
not ( n21568 , n461 );
not ( n21569 , n15094 );
not ( n21570 , n21569 );
not ( n21571 , n21570 );
and ( n21572 , n21568 , n21571 );
buf ( n21573 , n21569 );
nor ( n21574 , n573 , n21573 );
nor ( n21575 , n21572 , n21574 , n21565 );
nor ( n21576 , n21567 , n21575 );
not ( n21577 , n18 );
nand ( n21578 , n21577 , n17 );
not ( n21579 , n21578 );
not ( n21580 , n21579 );
buf ( n21581 , n21580 );
buf ( n21582 , n21581 );
not ( n21583 , n21582 );
nand ( n21584 , n14 , n15 );
not ( n21585 , n16 );
nor ( n21586 , n12 , n13 );
nand ( n21587 , n21585 , n21586 );
nor ( n21588 , n21584 , n21587 );
nand ( n21589 , n18682 , n15273 );
not ( n21590 , n21589 );
nand ( n21591 , n21588 , n21590 );
not ( n21592 , n21591 );
and ( n21593 , n21583 , n21592 );
buf ( n21594 , n21593 );
not ( n21595 , n21594 );
not ( n21596 , n21595 );
or ( n21597 , n21576 , n21596 );
buf ( n21598 , n21593 );
nand ( n21599 , n33 , n21598 );
nand ( n21600 , n21597 , n2 , n21599 );
not ( n21601 , n19288 );
nand ( n21602 , n19292 , n19299 );
nand ( n21603 , n19306 , n21602 );
not ( n21604 , n21603 );
or ( n21605 , n21601 , n21604 );
nand ( n21606 , n21605 , n19311 );
and ( n21607 , n19287 , n21606 );
nor ( n21608 , n21607 , n19281 );
or ( n21609 , n16852 , n21608 );
not ( n21610 , n16849 );
not ( n21611 , n21608 );
and ( n21612 , n21610 , n21611 );
nand ( n21613 , n16852 , n16849 );
not ( n21614 , n19295 );
and ( n21615 , n19292 , n21614 );
and ( n21616 , n19287 , n19288 , n21615 );
and ( n21617 , n21613 , n21616 );
nor ( n21618 , n21612 , n21617 );
nor ( n21619 , n21613 , n21616 );
nand ( n21620 , n21619 , n21608 );
nand ( n21621 , n21609 , n21618 , n21620 );
and ( n21622 , n391 , n1148 );
nor ( n21623 , n1095 , n1100 );
and ( n21624 , n15629 , n21623 );
nand ( n21625 , n15610 , n21624 );
and ( n21626 , n21517 , n15585 );
nor ( n21627 , n1124 , n1174 );
and ( n21628 , n15594 , n21627 );
nand ( n21629 , n19389 , n21626 , n21628 );
nor ( n21630 , n1095 , n21625 , n21629 );
not ( n21631 , n1066 );
nor ( n21632 , n902 , n1113 );
and ( n21633 , n21631 , n21532 , n21632 );
and ( n21634 , n21630 , n889 , n21633 );
not ( n21635 , n1095 );
nand ( n21636 , n1608 , n15647 );
nor ( n21637 , n21635 , n21636 );
nor ( n21638 , n21634 , n21637 );
and ( n21639 , n21517 , n21622 , n21638 );
and ( n21640 , n1029 , n21638 );
nor ( n21641 , n21639 , n21640 );
nand ( n21642 , n15619 , n15622 );
nor ( n21643 , n21517 , n21642 );
and ( n21644 , n15629 , n21643 , n21638 );
nand ( n21645 , n21520 , n21633 );
not ( n21646 , n21645 );
and ( n21647 , n15631 , n15586 );
or ( n21648 , n1045 , n1148 );
or ( n21649 , n21517 , n15629 );
nand ( n21650 , n21648 , n21649 );
and ( n21651 , n15601 , n21647 , n15599 , n21650 );
not ( n21652 , n1174 );
nand ( n21653 , n21646 , n21651 , n1806 , n21652 );
and ( n21654 , n15586 , n21624 );
or ( n21655 , n1806 , n19389 , n21645 );
nand ( n21656 , n1150 , n15585 );
nor ( n21657 , n889 , n1066 );
nand ( n21658 , n21657 , n21632 );
or ( n21659 , n21656 , n1083 , n21658 );
nand ( n21660 , n21655 , n21659 );
nand ( n21661 , n21628 , n21654 , n21650 , n21660 );
nand ( n21662 , n21653 , n21661 );
and ( n21663 , n21638 , n21662 );
nor ( n21664 , n21644 , n21663 );
nand ( n21665 , n21641 , n21664 );
not ( n21666 , n21430 );
nand ( n21667 , n21666 , n17119 );
or ( n21668 , n21667 , n21447 );
nand ( n21669 , n931 , n13749 );
and ( n21670 , n21669 , n21439 );
and ( n21671 , n21437 , n21667 );
or ( n21672 , n21437 , n21441 );
nand ( n21673 , n21672 , n21425 );
nor ( n21674 , n21671 , n21673 );
not ( n21675 , n931 );
not ( n21676 , n928 );
not ( n21677 , n930 );
and ( n21678 , n21675 , n21676 , n21677 );
nor ( n21679 , n929 , n931 );
not ( n21680 , n21435 );
nand ( n21681 , n21679 , n21680 );
or ( n21682 , n21681 , n900 , n21423 );
or ( n21683 , n931 , n900 , n928 );
nand ( n21684 , n21682 , n21683 );
nor ( n21685 , n21678 , n21684 );
nor ( n21686 , n21685 , n21442 , n21452 );
nor ( n21687 , n21670 , n21674 , n21686 );
nand ( n21688 , n21668 , n21687 , n21445 );
and ( n21689 , n682 , n20904 );
and ( n21690 , n581 , n20593 );
nor ( n21691 , n21689 , n21690 );
and ( n21692 , n999 , n20624 );
and ( n21693 , n492 , n21189 );
and ( n21694 , n444 , n20600 );
nor ( n21695 , n21692 , n21693 , n21694 );
nand ( n21696 , n21691 , n21695 );
and ( n21697 , n711 , n20910 );
and ( n21698 , n628 , n21059 );
and ( n21699 , n531 , n20894 );
nor ( n21700 , n21697 , n21698 , n21699 );
and ( n21701 , n821 , n20591 );
and ( n21702 , n980 , n20438 );
nor ( n21703 , n21701 , n21702 );
nand ( n21704 , n21700 , n21703 );
and ( n21705 , n703 , n21118 );
and ( n21706 , n621 , n20873 );
and ( n21707 , n522 , n20752 );
nor ( n21708 , n21705 , n21706 , n21707 );
and ( n21709 , n812 , n20591 );
and ( n21710 , n971 , n20438 );
nor ( n21711 , n21709 , n21710 );
nand ( n21712 , n21708 , n21711 );
and ( n21713 , n661 , n21179 );
and ( n21714 , n502 , n20912 );
and ( n21715 , n455 , n21005 );
nor ( n21716 , n21713 , n21714 , n21715 );
and ( n21717 , n768 , n20591 );
and ( n21718 , n968 , n20438 );
nor ( n21719 , n21717 , n21718 );
nand ( n21720 , n21716 , n21719 );
and ( n21721 , n1241 , n20591 );
and ( n21722 , n1273 , n20593 );
nor ( n21723 , n21721 , n21722 );
and ( n21724 , n930 , n20624 );
and ( n21725 , n1209 , n20500 );
and ( n21726 , n1385 , n21132 );
nor ( n21727 , n21724 , n21725 , n21726 );
nand ( n21728 , n21723 , n21727 );
and ( n21729 , n1098 , n21179 );
and ( n21730 , n1068 , n20749 );
and ( n21731 , n992 , n20894 );
nor ( n21732 , n21729 , n21730 , n21731 );
and ( n21733 , n1123 , n20591 );
and ( n21734 , n931 , n20438 );
nor ( n21735 , n21733 , n21734 );
nand ( n21736 , n21732 , n21735 );
not ( n21737 , n2 );
nand ( n21738 , n18 , n15957 );
not ( n21739 , n21738 );
not ( n21740 , n21739 );
buf ( n21741 , n21740 );
not ( n21742 , n21741 );
buf ( n21743 , n21742 );
nand ( n21744 , n16 , n21586 );
not ( n21745 , n21744 );
and ( n21746 , n14 , n15947 );
nand ( n21747 , n21745 , n21746 );
not ( n21748 , n21747 );
nand ( n21749 , n21748 , n21590 );
not ( n21750 , n21749 );
nand ( n21751 , n21743 , n21750 );
buf ( n21752 , n21751 );
not ( n21753 , n21752 );
and ( n21754 , n23 , n21753 );
and ( n21755 , n1481 , n21752 );
nor ( n21756 , n21754 , n21755 );
nor ( n21757 , n21737 , n21756 );
not ( n21758 , n2 );
nor ( n21759 , n21584 , n21744 );
nand ( n21760 , n21759 , n21590 );
not ( n21761 , n21760 );
nand ( n21762 , n21743 , n21761 );
buf ( n21763 , n21762 );
not ( n21764 , n21763 );
and ( n21765 , n23 , n21764 );
and ( n21766 , n1485 , n21763 );
nor ( n21767 , n21765 , n21766 );
nor ( n21768 , n21758 , n21767 );
and ( n21769 , n1234 , n20591 );
and ( n21770 , n1161 , n20593 );
nor ( n21771 , n21769 , n21770 );
and ( n21772 , n933 , n20624 );
and ( n21773 , n1156 , n20598 );
and ( n21774 , n1151 , n21132 );
nor ( n21775 , n21772 , n21773 , n21774 );
nand ( n21776 , n21771 , n21775 );
not ( n21777 , n153 );
not ( n21778 , n20618 );
not ( n21779 , n21778 );
or ( n21780 , n21777 , n21779 );
not ( n21781 , n20613 );
and ( n21782 , n801 , n21781 );
nor ( n21783 , n21782 , n1600 );
nand ( n21784 , n21780 , n21783 );
and ( n21785 , n940 , n1228 );
and ( n21786 , n141 , n896 );
nor ( n21787 , n141 , n896 );
nor ( n21788 , n21786 , n21787 , n18011 );
nor ( n21789 , n21785 , n21788 );
or ( n21790 , n16506 , n21789 );
or ( n21791 , n1024 , n12691 );
nand ( n21792 , n21791 , n16506 , n12692 );
nand ( n21793 , n21790 , n21792 );
not ( n21794 , n2 );
not ( n21795 , n21587 );
nand ( n21796 , n21746 , n21795 );
not ( n21797 , n21796 );
nand ( n21798 , n21797 , n21590 );
not ( n21799 , n21798 );
nand ( n21800 , n21743 , n21799 );
buf ( n21801 , n21800 );
not ( n21802 , n21801 );
and ( n21803 , n28 , n21802 );
and ( n21804 , n1533 , n21801 );
nor ( n21805 , n21803 , n21804 );
nor ( n21806 , n21794 , n21805 );
not ( n21807 , n2 );
and ( n21808 , n34 , n21753 );
and ( n21809 , n1537 , n21752 );
nor ( n21810 , n21808 , n21809 );
nor ( n21811 , n21807 , n21810 );
buf ( n21812 , n14978 );
not ( n21813 , n21812 );
buf ( n21814 , n21813 );
and ( n21815 , n1211 , n21814 );
not ( n21816 , n1801 );
buf ( n21817 , n14977 );
not ( n21818 , n21817 );
and ( n21819 , n21816 , n21818 );
not ( n21820 , n21817 );
nor ( n21821 , n440 , n21820 );
not ( n21822 , n21812 );
nor ( n21823 , n21819 , n21821 , n21822 );
nor ( n21824 , n21815 , n21823 );
and ( n21825 , n21583 , n21799 );
not ( n21826 , n21825 );
buf ( n21827 , n21826 );
not ( n21828 , n21827 );
or ( n21829 , n21824 , n21828 );
buf ( n21830 , n21825 );
nand ( n21831 , n24 , n21830 );
nand ( n21832 , n21829 , n2 , n21831 );
and ( n21833 , n1204 , n21814 );
not ( n21834 , n1795 );
not ( n21835 , n21817 );
and ( n21836 , n21834 , n21835 );
not ( n21837 , n21817 );
nor ( n21838 , n441 , n21837 );
not ( n21839 , n21812 );
nor ( n21840 , n21836 , n21838 , n21839 );
nor ( n21841 , n21833 , n21840 );
not ( n21842 , n21827 );
or ( n21843 , n21841 , n21842 );
buf ( n21844 , n21825 );
nand ( n21845 , n21 , n21844 );
nand ( n21846 , n21843 , n2 , n21845 );
and ( n21847 , n1311 , n21814 );
not ( n21848 , n151 );
not ( n21849 , n21817 );
and ( n21850 , n21848 , n21849 );
not ( n21851 , n21817 );
nor ( n21852 , n442 , n21851 );
nor ( n21853 , n21850 , n21852 , n21839 );
nor ( n21854 , n21847 , n21853 );
or ( n21855 , n21854 , n21842 );
nand ( n21856 , n43 , n21844 );
nand ( n21857 , n21855 , n2 , n21856 );
not ( n21858 , n21812 );
not ( n21859 , n21858 );
not ( n21860 , n21817 );
and ( n21861 , n253 , n21860 );
and ( n21862 , n443 , n21817 );
nor ( n21863 , n21861 , n21862 );
not ( n21864 , n21863 );
and ( n21865 , n21859 , n21864 );
buf ( n21866 , n21858 );
and ( n21867 , n1305 , n21866 );
nor ( n21868 , n21865 , n21867 );
or ( n21869 , n21868 , n21830 );
not ( n21870 , n21826 );
nand ( n21871 , n25 , n21870 );
nand ( n21872 , n21869 , n2 , n21871 );
and ( n21873 , n1298 , n21866 );
not ( n21874 , n140 );
not ( n21875 , n21817 );
and ( n21876 , n21874 , n21875 );
not ( n21877 , n21817 );
nor ( n21878 , n444 , n21877 );
nor ( n21879 , n21876 , n21878 , n21813 );
nor ( n21880 , n21873 , n21879 );
not ( n21881 , n21827 );
or ( n21882 , n21880 , n21881 );
nand ( n21883 , n38 , n21870 );
nand ( n21884 , n21882 , n2 , n21883 );
and ( n21885 , n1295 , n21866 );
not ( n21886 , n145 );
not ( n21887 , n21817 );
and ( n21888 , n21886 , n21887 );
not ( n21889 , n21817 );
nor ( n21890 , n445 , n21889 );
not ( n21891 , n21812 );
nor ( n21892 , n21888 , n21890 , n21891 );
nor ( n21893 , n21885 , n21892 );
not ( n21894 , n21827 );
or ( n21895 , n21893 , n21894 );
nand ( n21896 , n42 , n21830 );
nand ( n21897 , n21895 , n2 , n21896 );
and ( n21898 , n1368 , n21814 );
not ( n21899 , n136 );
and ( n21900 , n21899 , n21835 );
nor ( n21901 , n446 , n21837 );
nor ( n21902 , n21900 , n21901 , n21822 );
nor ( n21903 , n21898 , n21902 );
or ( n21904 , n21903 , n21881 );
nand ( n21905 , n39 , n21844 );
nand ( n21906 , n21904 , n2 , n21905 );
and ( n21907 , n1296 , n21866 );
not ( n21908 , n148 );
and ( n21909 , n21908 , n21818 );
nor ( n21910 , n448 , n21851 );
nor ( n21911 , n21909 , n21910 , n21839 );
nor ( n21912 , n21907 , n21911 );
or ( n21913 , n21912 , n21842 );
nand ( n21914 , n41 , n21830 );
nand ( n21915 , n21913 , n2 , n21914 );
and ( n21916 , n1375 , n21866 );
not ( n21917 , n147 );
not ( n21918 , n21817 );
and ( n21919 , n21917 , n21918 );
not ( n21920 , n21817 );
nor ( n21921 , n449 , n21920 );
not ( n21922 , n21812 );
nor ( n21923 , n21919 , n21921 , n21922 );
nor ( n21924 , n21916 , n21923 );
or ( n21925 , n21924 , n21842 );
nand ( n21926 , n37 , n21844 );
nand ( n21927 , n21925 , n2 , n21926 );
and ( n21928 , n1202 , n21814 );
not ( n21929 , n152 );
and ( n21930 , n21929 , n21849 );
nor ( n21931 , n450 , n21837 );
nor ( n21932 , n21930 , n21931 , n21891 );
nor ( n21933 , n21928 , n21932 );
not ( n21934 , n21827 );
or ( n21935 , n21933 , n21934 );
nand ( n21936 , n46 , n21844 );
nand ( n21937 , n21935 , n2 , n21936 );
and ( n21938 , n1182 , n21814 );
not ( n21939 , n159 );
and ( n21940 , n21939 , n21918 );
not ( n21941 , n21817 );
nor ( n21942 , n453 , n21941 );
nor ( n21943 , n21940 , n21942 , n21822 );
nor ( n21944 , n21938 , n21943 );
or ( n21945 , n21944 , n21881 );
nand ( n21946 , n45 , n21844 );
nand ( n21947 , n21945 , n2 , n21946 );
and ( n21948 , n1383 , n21814 );
not ( n21949 , n193 );
and ( n21950 , n21949 , n21818 );
nor ( n21951 , n466 , n21941 );
not ( n21952 , n21812 );
nor ( n21953 , n21950 , n21951 , n21952 );
nor ( n21954 , n21948 , n21953 );
not ( n21955 , n21827 );
or ( n21956 , n21954 , n21955 );
nand ( n21957 , n52 , n21844 );
nand ( n21958 , n21956 , n2 , n21957 );
and ( n21959 , n1300 , n21866 );
not ( n21960 , n439 );
and ( n21961 , n21960 , n21918 );
nor ( n21962 , n467 , n21920 );
nor ( n21963 , n21961 , n21962 , n21822 );
nor ( n21964 , n21959 , n21963 );
or ( n21965 , n21964 , n21881 );
nand ( n21966 , n34 , n21844 );
nand ( n21967 , n21965 , n2 , n21966 );
and ( n21968 , n1370 , n21866 );
and ( n21969 , n21568 , n21875 );
nor ( n21970 , n468 , n21889 );
nor ( n21971 , n21969 , n21970 , n21839 );
nor ( n21972 , n21968 , n21971 );
or ( n21973 , n21972 , n21828 );
nand ( n21974 , n33 , n21830 );
nand ( n21975 , n21973 , n2 , n21974 );
and ( n21976 , n1301 , n21814 );
not ( n21977 , n186 );
and ( n21978 , n21977 , n21887 );
nor ( n21979 , n469 , n21920 );
not ( n21980 , n21812 );
nor ( n21981 , n21978 , n21979 , n21980 );
nor ( n21982 , n21976 , n21981 );
or ( n21983 , n21982 , n21828 );
nand ( n21984 , n51 , n21844 );
nand ( n21985 , n21983 , n2 , n21984 );
and ( n21986 , n1206 , n21814 );
not ( n21987 , n428 );
and ( n21988 , n21987 , n21875 );
nor ( n21989 , n470 , n21877 );
nor ( n21990 , n21988 , n21989 , n21922 );
nor ( n21991 , n21986 , n21990 );
or ( n21992 , n21991 , n21894 );
nand ( n21993 , n32 , n21830 );
nand ( n21994 , n21992 , n2 , n21993 );
and ( n21995 , n1302 , n21814 );
not ( n21996 , n415 );
and ( n21997 , n21996 , n21918 );
nor ( n21998 , n471 , n21851 );
nor ( n21999 , n21997 , n21998 , n21891 );
nor ( n22000 , n21995 , n21999 );
or ( n22001 , n22000 , n21894 );
nand ( n22002 , n31 , n21830 );
nand ( n22003 , n22001 , n2 , n22002 );
and ( n22004 , n1303 , n21866 );
not ( n22005 , n383 );
and ( n22006 , n22005 , n21875 );
nor ( n22007 , n472 , n21820 );
nor ( n22008 , n22006 , n22007 , n21980 );
nor ( n22009 , n22004 , n22008 );
or ( n22010 , n22009 , n21894 );
nand ( n22011 , n29 , n21870 );
nand ( n22012 , n22010 , n2 , n22011 );
and ( n22013 , n1222 , n21866 );
not ( n22014 , n352 );
and ( n22015 , n22014 , n21849 );
nor ( n22016 , n473 , n21877 );
nor ( n22017 , n22015 , n22016 , n21922 );
nor ( n22018 , n22013 , n22017 );
not ( n22019 , n21827 );
or ( n22020 , n22018 , n22019 );
nand ( n22021 , n28 , n21830 );
nand ( n22022 , n22020 , n2 , n22021 );
and ( n22023 , n1218 , n21814 );
not ( n22024 , n284 );
and ( n22025 , n22024 , n21835 );
nor ( n22026 , n475 , n21820 );
nor ( n22027 , n22025 , n22026 , n21980 );
nor ( n22028 , n22023 , n22027 );
or ( n22029 , n22028 , n21830 );
nand ( n22030 , n26 , n21870 );
nand ( n22031 , n22029 , n2 , n22030 );
and ( n22032 , n1308 , n21814 );
not ( n22033 , n192 );
and ( n22034 , n22033 , n21835 );
nor ( n22035 , n476 , n21820 );
nor ( n22036 , n22034 , n22035 , n21891 );
nor ( n22037 , n22032 , n22036 );
or ( n22038 , n22037 , n22019 );
nand ( n22039 , n22 , n21830 );
nand ( n22040 , n22038 , n2 , n22039 );
and ( n22041 , n1309 , n21866 );
not ( n22042 , n178 );
and ( n22043 , n22042 , n21887 );
nor ( n22044 , n477 , n21837 );
nor ( n22045 , n22043 , n22044 , n21952 );
nor ( n22046 , n22041 , n22045 );
or ( n22047 , n22046 , n21828 );
nand ( n22048 , n49 , n21844 );
nand ( n22049 , n22047 , n2 , n22048 );
and ( n22050 , n1184 , n21866 );
not ( n22051 , n156 );
and ( n22052 , n22051 , n21860 );
nor ( n22053 , n478 , n21941 );
nor ( n22054 , n22052 , n22053 , n21922 );
nor ( n22055 , n22050 , n22054 );
or ( n22056 , n22055 , n22019 );
nand ( n22057 , n44 , n21830 );
nand ( n22058 , n22056 , n2 , n22057 );
not ( n22059 , n15708 );
and ( n22060 , n1378 , n22059 );
not ( n22061 , n15707 );
and ( n22062 , n21816 , n22061 );
nor ( n22063 , n479 , n22061 );
nor ( n22064 , n22062 , n22063 , n22059 );
nor ( n22065 , n22060 , n22064 );
and ( n22066 , n21583 , n21750 );
not ( n22067 , n22066 );
buf ( n22068 , n22067 );
not ( n22069 , n22068 );
or ( n22070 , n22065 , n22069 );
buf ( n22071 , n22066 );
nand ( n22072 , n24 , n22071 );
nand ( n22073 , n22070 , n2 , n22072 );
and ( n22074 , n1367 , n22059 );
and ( n22075 , n21834 , n22061 );
nor ( n22076 , n480 , n22061 );
nor ( n22077 , n22075 , n22076 , n22059 );
nor ( n22078 , n22074 , n22077 );
not ( n22079 , n22068 );
or ( n22080 , n22078 , n22079 );
nand ( n22081 , n21 , n22071 );
nand ( n22082 , n22080 , n2 , n22081 );
and ( n22083 , n1374 , n22059 );
and ( n22084 , n22051 , n22061 );
nor ( n22085 , n485 , n22061 );
nor ( n22086 , n22084 , n22085 , n22059 );
nor ( n22087 , n22083 , n22086 );
not ( n22088 , n22068 );
or ( n22089 , n22087 , n22088 );
nand ( n22090 , n44 , n22071 );
nand ( n22091 , n22089 , n2 , n22090 );
not ( n22092 , n13367 );
not ( n22093 , n22092 );
and ( n22094 , n13370 , n13360 );
not ( n22095 , n22094 );
or ( n22096 , n22093 , n22095 );
or ( n22097 , n22092 , n22094 );
nand ( n22098 , n22096 , n22097 );
and ( n22099 , n1373 , n22059 );
and ( n22100 , n21929 , n22061 );
nor ( n22101 , n491 , n22061 );
nor ( n22102 , n22100 , n22101 , n22059 );
nor ( n22103 , n22099 , n22102 );
or ( n22104 , n22103 , n22069 );
buf ( n22105 , n22066 );
nand ( n22106 , n46 , n22105 );
nand ( n22107 , n22104 , n2 , n22106 );
and ( n22108 , n1317 , n22059 );
and ( n22109 , n21874 , n22061 );
nor ( n22110 , n492 , n22061 );
nor ( n22111 , n22109 , n22110 , n22059 );
nor ( n22112 , n22108 , n22111 );
or ( n22113 , n22112 , n22088 );
nand ( n22114 , n38 , n22071 );
nand ( n22115 , n22113 , n2 , n22114 );
and ( n22116 , n1314 , n22059 );
and ( n22117 , n21886 , n22061 );
nor ( n22118 , n493 , n22061 );
nor ( n22119 , n22117 , n22118 , n22059 );
nor ( n22120 , n22116 , n22119 );
or ( n22121 , n22120 , n22079 );
not ( n22122 , n22067 );
nand ( n22123 , n42 , n22122 );
nand ( n22124 , n22121 , n2 , n22123 );
and ( n22125 , n1192 , n22059 );
and ( n22126 , n21899 , n22061 );
nor ( n22127 , n494 , n22061 );
nor ( n22128 , n22126 , n22127 , n22059 );
nor ( n22129 , n22125 , n22128 );
or ( n22130 , n22129 , n22079 );
nand ( n22131 , n39 , n22105 );
nand ( n22132 , n22130 , n2 , n22131 );
and ( n22133 , n1315 , n22059 );
and ( n22134 , n21908 , n22061 );
nor ( n22135 , n496 , n22061 );
nor ( n22136 , n22134 , n22135 , n22059 );
nor ( n22137 , n22133 , n22136 );
not ( n22138 , n22068 );
or ( n22139 , n22137 , n22138 );
nand ( n22140 , n41 , n22071 );
nand ( n22141 , n22139 , n2 , n22140 );
and ( n22142 , n1318 , n22059 );
and ( n22143 , n21917 , n22061 );
nor ( n22144 , n497 , n22061 );
nor ( n22145 , n22143 , n22144 , n22059 );
nor ( n22146 , n22142 , n22145 );
or ( n22147 , n22146 , n22088 );
nand ( n22148 , n37 , n22105 );
nand ( n22149 , n22147 , n2 , n22148 );
nand ( n22150 , n17 , n18 );
not ( n22151 , n22150 );
buf ( n22152 , n22151 );
not ( n22153 , n22152 );
not ( n22154 , n22153 );
buf ( n22155 , n22154 );
and ( n22156 , n22155 , n21750 );
buf ( n22157 , n22156 );
not ( n22158 , n22157 );
or ( n22159 , n16033 , n22158 );
not ( n22160 , n1125 );
not ( n22161 , n1576 );
or ( n22162 , n22160 , n22161 );
nand ( n22163 , n1576 , n1858 );
nand ( n22164 , n22162 , n22163 );
not ( n22165 , n22164 );
or ( n22166 , n136 , n22165 );
or ( n22167 , n499 , n22164 );
not ( n22168 , n22157 );
nand ( n22169 , n22166 , n22167 , n22168 );
nand ( n22170 , n22159 , n2 , n22169 );
and ( n22171 , n1334 , n22059 );
and ( n22172 , n21939 , n22061 );
nor ( n22173 , n500 , n22061 );
nor ( n22174 , n22172 , n22173 , n22059 );
nor ( n22175 , n22171 , n22174 );
or ( n22176 , n22175 , n22088 );
nand ( n22177 , n45 , n22105 );
nand ( n22178 , n22176 , n2 , n22177 );
and ( n22179 , n501 , n22165 );
and ( n22180 , n148 , n22164 );
nor ( n22181 , n22179 , n22180 );
not ( n22182 , n22157 );
not ( n22183 , n22182 );
or ( n22184 , n22181 , n22183 );
not ( n22185 , n22157 );
or ( n22186 , n16041 , n22185 );
nand ( n22187 , n22184 , n22186 , n2 );
and ( n22188 , n502 , n22165 );
and ( n22189 , n147 , n22164 );
nor ( n22190 , n22188 , n22189 );
or ( n22191 , n22190 , n22183 );
not ( n22192 , n22157 );
or ( n22193 , n16025 , n22192 );
nand ( n22194 , n22191 , n22193 , n2 );
not ( n22195 , n22157 );
or ( n22196 , n16057 , n22195 );
or ( n22197 , n159 , n22165 );
or ( n22198 , n504 , n22164 );
not ( n22199 , n22157 );
nand ( n22200 , n22197 , n22198 , n22199 );
nand ( n22201 , n22196 , n2 , n22200 );
and ( n22202 , n535 , n22165 );
and ( n22203 , n1801 , n22164 );
nor ( n22204 , n22202 , n22203 );
or ( n22205 , n22204 , n22183 );
or ( n22206 , n16065 , n22182 );
nand ( n22207 , n22205 , n22206 , n2 );
and ( n22208 , n542 , n18078 );
not ( n22209 , n17274 );
nand ( n22210 , n22209 , n17295 );
not ( n22211 , n17292 );
and ( n22212 , n22210 , n22211 );
or ( n22213 , n22210 , n22211 );
not ( n22214 , n14979 );
nand ( n22215 , n22213 , n22214 );
nor ( n22216 , n22212 , n22215 );
nor ( n22217 , n22208 , n22216 );
or ( n22218 , n1819 , n22217 );
and ( n22219 , n542 , n17332 );
nor ( n22220 , n22219 , n17333 );
or ( n22221 , n14974 , n22220 );
nand ( n22222 , n22218 , n22221 );
and ( n22223 , n1251 , n22222 );
and ( n22224 , n1319 , n22059 );
not ( n22225 , n144 );
and ( n22226 , n22225 , n22061 );
nor ( n22227 , n543 , n22061 );
nor ( n22228 , n22226 , n22227 , n22059 );
nor ( n22229 , n22224 , n22228 );
not ( n22230 , n22068 );
or ( n22231 , n22229 , n22230 );
nand ( n22232 , n36 , n22105 );
nand ( n22233 , n22231 , n2 , n22232 );
and ( n22234 , n1320 , n22059 );
and ( n22235 , n21960 , n22061 );
nor ( n22236 , n544 , n22061 );
nor ( n22237 , n22235 , n22236 , n22059 );
nor ( n22238 , n22234 , n22237 );
buf ( n22239 , n22067 );
not ( n22240 , n22239 );
or ( n22241 , n22238 , n22240 );
nand ( n22242 , n34 , n22105 );
nand ( n22243 , n22241 , n2 , n22242 );
and ( n22244 , n1321 , n22059 );
and ( n22245 , n21568 , n22061 );
nor ( n22246 , n545 , n22061 );
nor ( n22247 , n22245 , n22246 , n22059 );
nor ( n22248 , n22244 , n22247 );
or ( n22249 , n22248 , n22069 );
nand ( n22250 , n33 , n22071 );
nand ( n22251 , n22249 , n2 , n22250 );
and ( n22252 , n1405 , n22059 );
and ( n22253 , n21987 , n22061 );
nor ( n22254 , n547 , n22061 );
nor ( n22255 , n22253 , n22254 , n22059 );
nor ( n22256 , n22252 , n22255 );
or ( n22257 , n22256 , n22230 );
nand ( n22258 , n32 , n22071 );
nand ( n22259 , n22257 , n2 , n22258 );
and ( n22260 , n1323 , n22059 );
and ( n22261 , n21996 , n22061 );
nor ( n22262 , n548 , n22061 );
nor ( n22263 , n22261 , n22262 , n22059 );
nor ( n22264 , n22260 , n22263 );
or ( n22265 , n22264 , n22230 );
nand ( n22266 , n31 , n22122 );
nand ( n22267 , n22265 , n2 , n22266 );
and ( n22268 , n1325 , n22059 );
and ( n22269 , n22005 , n22061 );
nor ( n22270 , n549 , n22061 );
nor ( n22271 , n22269 , n22270 , n22059 );
nor ( n22272 , n22268 , n22271 );
not ( n22273 , n22068 );
or ( n22274 , n22272 , n22273 );
nand ( n22275 , n29 , n22122 );
nand ( n22276 , n22274 , n2 , n22275 );
and ( n22277 , n1393 , n22059 );
and ( n22278 , n22014 , n22061 );
nor ( n22279 , n550 , n22061 );
nor ( n22280 , n22278 , n22279 , n22059 );
nor ( n22281 , n22277 , n22280 );
or ( n22282 , n22281 , n22273 );
nand ( n22283 , n28 , n22071 );
nand ( n22284 , n22282 , n2 , n22283 );
and ( n22285 , n1326 , n22059 );
not ( n22286 , n283 );
and ( n22287 , n22286 , n22061 );
nor ( n22288 , n551 , n22061 );
nor ( n22289 , n22287 , n22288 , n22059 );
nor ( n22290 , n22285 , n22289 );
or ( n22291 , n22290 , n22071 );
nand ( n22292 , n27 , n22122 );
nand ( n22293 , n22291 , n2 , n22292 );
and ( n22294 , n1165 , n22059 );
and ( n22295 , n22033 , n22061 );
nor ( n22296 , n553 , n22061 );
nor ( n22297 , n22295 , n22296 , n22059 );
nor ( n22298 , n22294 , n22297 );
not ( n22299 , n22068 );
or ( n22300 , n22298 , n22299 );
nand ( n22301 , n22 , n22071 );
nand ( n22302 , n22300 , n2 , n22301 );
and ( n22303 , n1331 , n22059 );
and ( n22304 , n22042 , n22061 );
nor ( n22305 , n554 , n22061 );
nor ( n22306 , n22304 , n22305 , n22059 );
nor ( n22307 , n22303 , n22306 );
not ( n22308 , n22068 );
or ( n22309 , n22307 , n22308 );
nand ( n22310 , n49 , n22105 );
nand ( n22311 , n22309 , n2 , n22310 );
buf ( n22312 , n21565 );
and ( n22313 , n1186 , n22312 );
not ( n22314 , n21569 );
not ( n22315 , n22314 );
and ( n22316 , n21816 , n22315 );
nor ( n22317 , n556 , n21573 );
nor ( n22318 , n22316 , n22317 , n21565 );
nor ( n22319 , n22313 , n22318 );
not ( n22320 , n21595 );
or ( n22321 , n22319 , n22320 );
nand ( n22322 , n24 , n21598 );
nand ( n22323 , n22321 , n2 , n22322 );
and ( n22324 , n1350 , n21566 );
not ( n22325 , n21570 );
and ( n22326 , n21834 , n22325 );
buf ( n22327 , n21569 );
nor ( n22328 , n557 , n22327 );
nor ( n22329 , n22326 , n22328 , n21565 );
nor ( n22330 , n22324 , n22329 );
not ( n22331 , n21594 );
not ( n22332 , n22331 );
or ( n22333 , n22330 , n22332 );
nand ( n22334 , n21 , n21598 );
nand ( n22335 , n22333 , n2 , n22334 );
and ( n22336 , n1143 , n20591 );
and ( n22337 , n1102 , n20657 );
nor ( n22338 , n22336 , n22337 );
and ( n22339 , n932 , n20624 );
and ( n22340 , n1071 , n20500 );
and ( n22341 , n1005 , n21162 );
nor ( n22342 , n22339 , n22340 , n22341 );
nand ( n22343 , n22338 , n22342 );
and ( n22344 , n1307 , n21866 );
not ( n22345 , n185 );
and ( n22346 , n22345 , n21818 );
nor ( n22347 , n564 , n21889 );
not ( n22348 , n21812 );
nor ( n22349 , n22346 , n22347 , n22348 );
nor ( n22350 , n22344 , n22349 );
or ( n22351 , n22350 , n21934 );
nand ( n22352 , n50 , n21844 );
nand ( n22353 , n22351 , n2 , n22352 );
and ( n22354 , n1408 , n21566 );
and ( n22355 , n22051 , n21573 );
nor ( n22356 , n565 , n21573 );
nor ( n22357 , n22355 , n22356 , n21565 );
nor ( n22358 , n22354 , n22357 );
not ( n22359 , n21595 );
or ( n22360 , n22358 , n22359 );
nand ( n22361 , n44 , n21598 );
nand ( n22362 , n22360 , n2 , n22361 );
and ( n22363 , n1216 , n21814 );
not ( n22364 , n1610 );
and ( n22365 , n22364 , n21849 );
nor ( n22366 , n567 , n21941 );
nor ( n22367 , n22365 , n22366 , n22348 );
nor ( n22368 , n22363 , n22367 );
or ( n22369 , n22368 , n21955 );
nand ( n22370 , n30 , n21870 );
nand ( n22371 , n22369 , n2 , n22370 );
and ( n22372 , n1215 , n21566 );
not ( n22373 , n143 );
and ( n22374 , n22373 , n21573 );
nor ( n22375 , n568 , n21573 );
nor ( n22376 , n22374 , n22375 , n21565 );
nor ( n22377 , n22372 , n22376 );
or ( n22378 , n22377 , n22359 );
nand ( n22379 , n40 , n21598 );
nand ( n22380 , n22378 , n2 , n22379 );
and ( n22381 , n569 , n22165 );
and ( n22382 , n186 , n22164 );
nor ( n22383 , n22381 , n22382 );
not ( n22384 , n22182 );
or ( n22385 , n22383 , n22384 );
or ( n22386 , n16077 , n22192 );
nand ( n22387 , n22385 , n22386 , n2 );
and ( n22388 , n1490 , n20591 );
and ( n22389 , n1542 , n20593 );
nor ( n22390 , n22388 , n22389 );
and ( n22391 , n927 , n20624 );
and ( n22392 , n1498 , n20598 );
and ( n22393 , n1489 , n20600 );
nor ( n22394 , n22391 , n22392 , n22393 );
nand ( n22395 , n22390 , n22394 );
not ( n22396 , n22157 );
or ( n22397 , n15977 , n22396 );
or ( n22398 , n253 , n22165 );
or ( n22399 , n574 , n22164 );
nand ( n22400 , n22398 , n22399 , n22168 );
nand ( n22401 , n22397 , n2 , n22400 );
or ( n22402 , n15993 , n22195 );
or ( n22403 , n383 , n22165 );
or ( n22404 , n575 , n22164 );
nand ( n22405 , n22403 , n22404 , n22199 );
nand ( n22406 , n22402 , n2 , n22405 );
and ( n22407 , n1310 , n21814 );
not ( n22408 , n157 );
not ( n22409 , n21817 );
and ( n22410 , n22408 , n22409 );
nor ( n22411 , n576 , n21889 );
nor ( n22412 , n22410 , n22411 , n21952 );
nor ( n22413 , n22407 , n22412 );
buf ( n22414 , n21826 );
not ( n22415 , n22414 );
or ( n22416 , n22413 , n22415 );
nand ( n22417 , n47 , n21844 );
nand ( n22418 , n22416 , n2 , n22417 );
not ( n22419 , n21565 );
and ( n22420 , n152 , n22327 );
and ( n22421 , n578 , n22314 );
nor ( n22422 , n22420 , n22421 );
not ( n22423 , n22422 );
and ( n22424 , n22419 , n22423 );
and ( n22425 , n1407 , n22312 );
nor ( n22426 , n22424 , n22425 );
not ( n22427 , n22331 );
or ( n22428 , n22426 , n22427 );
nand ( n22429 , n46 , n21598 );
nand ( n22430 , n22428 , n2 , n22429 );
and ( n22431 , n1337 , n21566 );
and ( n22432 , n21908 , n22325 );
nor ( n22433 , n579 , n21573 );
nor ( n22434 , n22432 , n22433 , n21565 );
nor ( n22435 , n22431 , n22434 );
not ( n22436 , n21595 );
or ( n22437 , n22435 , n22436 );
nand ( n22438 , n41 , n21598 );
nand ( n22439 , n22437 , n2 , n22438 );
and ( n22440 , n1214 , n22312 );
and ( n22441 , n21886 , n21573 );
nor ( n22442 , n580 , n21573 );
nor ( n22443 , n22441 , n22442 , n21565 );
nor ( n22444 , n22440 , n22443 );
or ( n22445 , n22444 , n22332 );
buf ( n22446 , n21593 );
nand ( n22447 , n42 , n22446 );
nand ( n22448 , n22445 , n2 , n22447 );
and ( n22449 , n1191 , n22312 );
and ( n22450 , n21874 , n21571 );
nor ( n22451 , n581 , n22327 );
nor ( n22452 , n22450 , n22451 , n21565 );
nor ( n22453 , n22449 , n22452 );
or ( n22454 , n22453 , n22332 );
nand ( n22455 , n38 , n21598 );
nand ( n22456 , n22454 , n2 , n22455 );
and ( n22457 , n1338 , n21566 );
and ( n22458 , n21899 , n22327 );
nor ( n22459 , n582 , n22327 );
nor ( n22460 , n22458 , n22459 , n21565 );
nor ( n22461 , n22457 , n22460 );
or ( n22462 , n22461 , n21596 );
nand ( n22463 , n39 , n21598 );
nand ( n22464 , n22462 , n2 , n22463 );
not ( n22465 , n21858 );
and ( n22466 , n175 , n21860 );
and ( n22467 , n587 , n21817 );
nor ( n22468 , n22466 , n22467 );
not ( n22469 , n22468 );
and ( n22470 , n22465 , n22469 );
and ( n22471 , n1196 , n21866 );
nor ( n22472 , n22470 , n22471 );
not ( n22473 , n21827 );
or ( n22474 , n22472 , n22473 );
nand ( n22475 , n48 , n21830 );
nand ( n22476 , n22474 , n2 , n22475 );
not ( n22477 , n1800 );
nand ( n22478 , n602 , n22477 );
nand ( n22479 , n577 , n596 );
not ( n22480 , n20233 );
nor ( n22481 , n22479 , n22480 );
and ( n22482 , n20226 , n22481 );
or ( n22483 , n602 , n22482 );
and ( n22484 , n602 , n22482 );
nor ( n22485 , n22484 , n22477 );
nand ( n22486 , n22483 , n22485 );
and ( n22487 , n22478 , n22486 );
nor ( n22488 , n22487 , n834 );
and ( n22489 , n659 , n21118 );
and ( n22490 , n553 , n20628 );
and ( n22491 , n476 , n21334 );
nor ( n22492 , n22489 , n22490 , n22491 );
and ( n22493 , n737 , n20591 );
and ( n22494 , n897 , n20438 );
nor ( n22495 , n22493 , n22494 );
nand ( n22496 , n22492 , n22495 );
not ( n22497 , n22477 );
not ( n22498 , n608 );
not ( n22499 , n605 );
nor ( n22500 , n22499 , n20232 );
nand ( n22501 , n606 , n22500 );
nor ( n22502 , n22498 , n22479 , n22501 );
nand ( n22503 , n22497 , n22502 );
xor ( n22504 , n22503 , n607 );
nor ( n22505 , n834 , n22504 );
and ( n22506 , n616 , n22165 );
and ( n22507 , n193 , n22164 );
nor ( n22508 , n22506 , n22507 );
or ( n22509 , n22508 , n22183 );
not ( n22510 , n22157 );
or ( n22511 , n16089 , n22510 );
nand ( n22512 , n22509 , n22511 , n2 );
or ( n22513 , n16021 , n22195 );
or ( n22514 , n144 , n22165 );
or ( n22515 , n618 , n22164 );
nand ( n22516 , n22514 , n22515 , n22168 );
nand ( n22517 , n22513 , n2 , n22516 );
or ( n22518 , n16017 , n22396 );
or ( n22519 , n1082 , n22165 );
or ( n22520 , n619 , n22164 );
not ( n22521 , n22157 );
nand ( n22522 , n22519 , n22520 , n22521 );
nand ( n22523 , n22518 , n2 , n22522 );
or ( n22524 , n16013 , n22195 );
or ( n22525 , n439 , n22165 );
or ( n22526 , n620 , n22164 );
nand ( n22527 , n22525 , n22526 , n22521 );
nand ( n22528 , n22524 , n2 , n22527 );
and ( n22529 , n621 , n22165 );
and ( n22530 , n461 , n22164 );
nor ( n22531 , n22529 , n22530 );
or ( n22532 , n22531 , n22384 );
not ( n22533 , n22157 );
or ( n22534 , n16009 , n22533 );
nand ( n22535 , n22532 , n22534 , n2 );
and ( n22536 , n622 , n22165 );
and ( n22537 , n428 , n22164 );
nor ( n22538 , n22536 , n22537 );
or ( n22539 , n22538 , n22384 );
not ( n22540 , n22157 );
or ( n22541 , n16005 , n22540 );
nand ( n22542 , n22539 , n22541 , n2 );
and ( n22543 , n625 , n22165 );
and ( n22544 , n352 , n22164 );
nor ( n22545 , n22543 , n22544 );
or ( n22546 , n22545 , n22384 );
or ( n22547 , n15989 , n22510 );
nand ( n22548 , n22546 , n22547 , n2 );
not ( n22549 , n20904 );
or ( n22550 , n19062 , n22549 );
not ( n22551 , n900 );
not ( n22552 , n20624 );
or ( n22553 , n22551 , n22552 );
and ( n22554 , n1388 , n20416 );
and ( n22555 , n1261 , n20428 );
and ( n22556 , n1386 , n20432 );
nor ( n22557 , n22554 , n22555 , n22556 );
nand ( n22558 , n22550 , n22553 , n22557 );
or ( n22559 , n15985 , n22396 );
or ( n22560 , n283 , n22165 );
or ( n22561 , n626 , n22164 );
nand ( n22562 , n22560 , n22561 , n22521 );
nand ( n22563 , n22559 , n2 , n22562 );
or ( n22564 , n15981 , n22158 );
or ( n22565 , n284 , n22165 );
or ( n22566 , n627 , n22164 );
nand ( n22567 , n22565 , n22566 , n22199 );
nand ( n22568 , n22564 , n2 , n22567 );
or ( n22569 , n15969 , n22396 );
or ( n22570 , n192 , n22165 );
or ( n22571 , n629 , n22164 );
nand ( n22572 , n22570 , n22571 , n22168 );
nand ( n22573 , n22569 , n2 , n22572 );
or ( n22574 , n16053 , n22158 );
or ( n22575 , n156 , n22165 );
or ( n22576 , n632 , n22164 );
nand ( n22577 , n22575 , n22576 , n22521 );
nand ( n22578 , n22574 , n2 , n22577 );
or ( n22579 , n15005 , n14980 );
and ( n22580 , n15006 , n15032 );
or ( n22581 , n22580 , n16674 );
and ( n22582 , n22580 , n16674 );
nor ( n22583 , n22582 , n14979 );
nand ( n22584 , n22581 , n22583 );
nand ( n22585 , n22579 , n22584 );
and ( n22586 , n14974 , n22585 );
and ( n22587 , n15075 , n15005 );
not ( n22588 , n15075 );
and ( n22589 , n22588 , n637 );
nor ( n22590 , n22587 , n22589 );
and ( n22591 , n1819 , n22590 );
nor ( n22592 , n22586 , n22591 );
nor ( n22593 , n14973 , n22592 );
and ( n22594 , n643 , n18162 );
not ( n22595 , n17355 );
nand ( n22596 , n22595 , n17376 );
not ( n22597 , n17373 );
and ( n22598 , n22596 , n22597 );
or ( n22599 , n22596 , n22597 );
nand ( n22600 , n22599 , n15709 );
nor ( n22601 , n22598 , n22600 );
nor ( n22602 , n22594 , n22601 );
or ( n22603 , n1808 , n22602 );
and ( n22604 , n643 , n17413 );
nor ( n22605 , n22604 , n17414 );
or ( n22606 , n15704 , n22605 );
nand ( n22607 , n22603 , n22606 );
and ( n22608 , n1260 , n22607 );
buf ( n22609 , n16264 );
not ( n22610 , n22609 );
buf ( n22611 , n22610 );
and ( n22612 , n1288 , n22611 );
buf ( n22613 , n16262 );
not ( n22614 , n22613 );
not ( n22615 , n22614 );
and ( n22616 , n21816 , n22615 );
buf ( n22617 , n22613 );
nor ( n22618 , n644 , n22617 );
not ( n22619 , n22609 );
nor ( n22620 , n22616 , n22618 , n22619 );
nor ( n22621 , n22612 , n22620 );
and ( n22622 , n21583 , n21761 );
buf ( n22623 , n22622 );
not ( n22624 , n22623 );
not ( n22625 , n22624 );
or ( n22626 , n22621 , n22625 );
buf ( n22627 , n22622 );
nand ( n22628 , n24 , n22627 );
nand ( n22629 , n22626 , n2 , n22628 );
and ( n22630 , n1376 , n21866 );
not ( n22631 , n1082 );
and ( n22632 , n22631 , n22409 );
nor ( n22633 , n647 , n21851 );
nor ( n22634 , n22632 , n22633 , n21952 );
nor ( n22635 , n22630 , n22634 );
or ( n22636 , n22635 , n22473 );
nand ( n22637 , n35 , n21830 );
nand ( n22638 , n22636 , n2 , n22637 );
not ( n22639 , n21565 );
and ( n22640 , n144 , n22327 );
and ( n22641 , n650 , n22314 );
nor ( n22642 , n22640 , n22641 );
not ( n22643 , n22642 );
and ( n22644 , n22639 , n22643 );
and ( n22645 , n1200 , n22312 );
nor ( n22646 , n22644 , n22645 );
not ( n22647 , n22331 );
or ( n22648 , n22646 , n22647 );
nand ( n22649 , n36 , n21598 );
nand ( n22650 , n22648 , n2 , n22649 );
and ( n22651 , n1340 , n22312 );
and ( n22652 , n22631 , n22315 );
nor ( n22653 , n651 , n21573 );
nor ( n22654 , n22652 , n22653 , n21565 );
nor ( n22655 , n22651 , n22654 );
or ( n22656 , n22655 , n22359 );
nand ( n22657 , n35 , n21598 );
nand ( n22658 , n22656 , n2 , n22657 );
and ( n22659 , n1341 , n22312 );
not ( n22660 , n21570 );
and ( n22661 , n21960 , n22660 );
nor ( n22662 , n652 , n21573 );
nor ( n22663 , n22661 , n22662 , n21565 );
nor ( n22664 , n22659 , n22663 );
or ( n22665 , n22664 , n22647 );
nand ( n22666 , n34 , n21598 );
nand ( n22667 , n22665 , n2 , n22666 );
and ( n22668 , n1343 , n22312 );
and ( n22669 , n21987 , n22660 );
nor ( n22670 , n653 , n21573 );
nor ( n22671 , n22669 , n22670 , n21565 );
nor ( n22672 , n22668 , n22671 );
or ( n22673 , n22672 , n21596 );
nand ( n22674 , n32 , n22446 );
nand ( n22675 , n22673 , n2 , n22674 );
and ( n22676 , n1345 , n22312 );
and ( n22677 , n22364 , n22325 );
nor ( n22678 , n654 , n21573 );
nor ( n22679 , n22677 , n22678 , n21565 );
nor ( n22680 , n22676 , n22679 );
not ( n22681 , n22331 );
or ( n22682 , n22680 , n22681 );
nand ( n22683 , n30 , n22446 );
nand ( n22684 , n22682 , n2 , n22683 );
not ( n22685 , n21565 );
and ( n22686 , n352 , n22327 );
and ( n22687 , n655 , n22314 );
nor ( n22688 , n22686 , n22687 );
not ( n22689 , n22688 );
and ( n22690 , n22685 , n22689 );
and ( n22691 , n1346 , n22312 );
nor ( n22692 , n22690 , n22691 );
or ( n22693 , n22692 , n22427 );
nand ( n22694 , n28 , n22446 );
nand ( n22695 , n22693 , n2 , n22694 );
and ( n22696 , n1347 , n22312 );
and ( n22697 , n22286 , n22325 );
nor ( n22698 , n656 , n21573 );
nor ( n22699 , n22697 , n22698 , n21565 );
nor ( n22700 , n22696 , n22699 );
or ( n22701 , n22700 , n22647 );
nand ( n22702 , n27 , n21598 );
nand ( n22703 , n22701 , n2 , n22702 );
and ( n22704 , n1361 , n21566 );
not ( n22705 , n323 );
not ( n22706 , n22314 );
and ( n22707 , n22705 , n22706 );
nor ( n22708 , n657 , n21573 );
nor ( n22709 , n22707 , n22708 , n21565 );
nor ( n22710 , n22704 , n22709 );
or ( n22711 , n22710 , n22436 );
nand ( n22712 , n23 , n21598 );
nand ( n22713 , n22711 , n2 , n22712 );
and ( n22714 , n1395 , n21566 );
and ( n22715 , n22033 , n22706 );
nor ( n22716 , n659 , n22327 );
nor ( n22717 , n22715 , n22716 , n21565 );
nor ( n22718 , n22714 , n22717 );
or ( n22719 , n22718 , n22681 );
nand ( n22720 , n22 , n21598 );
nand ( n22721 , n22719 , n2 , n22720 );
and ( n22722 , n1329 , n22059 );
and ( n22723 , n22345 , n22061 );
nor ( n22724 , n663 , n22061 );
nor ( n22725 , n22723 , n22724 , n22059 );
nor ( n22726 , n22722 , n22725 );
or ( n22727 , n22726 , n22308 );
nand ( n22728 , n50 , n22071 );
nand ( n22729 , n22727 , n2 , n22728 );
and ( n22730 , n1324 , n22059 );
and ( n22731 , n22364 , n22061 );
nor ( n22732 , n665 , n22061 );
nor ( n22733 , n22731 , n22732 , n22059 );
nor ( n22734 , n22730 , n22733 );
or ( n22735 , n22734 , n22299 );
nand ( n22736 , n30 , n22122 );
nand ( n22737 , n22735 , n2 , n22736 );
and ( n22738 , n1398 , n22611 );
not ( n22739 , n22613 );
not ( n22740 , n22739 );
and ( n22741 , n22705 , n22740 );
buf ( n22742 , n22613 );
nor ( n22743 , n671 , n22742 );
not ( n22744 , n22609 );
nor ( n22745 , n22741 , n22743 , n22744 );
nor ( n22746 , n22738 , n22745 );
not ( n22747 , n22624 );
or ( n22748 , n22746 , n22747 );
nand ( n22749 , n23 , n22627 );
nand ( n22750 , n22748 , n2 , n22749 );
not ( n22751 , n22609 );
buf ( n22752 , n22751 );
and ( n22753 , n1404 , n22752 );
and ( n22754 , n22286 , n22740 );
nor ( n22755 , n673 , n22742 );
not ( n22756 , n22609 );
nor ( n22757 , n22754 , n22755 , n22756 );
nor ( n22758 , n22753 , n22757 );
or ( n22759 , n22758 , n22747 );
nand ( n22760 , n27 , n22627 );
nand ( n22761 , n22759 , n2 , n22760 );
and ( n22762 , n1333 , n22059 );
and ( n22763 , n22408 , n22061 );
nor ( n22764 , n677 , n22061 );
nor ( n22765 , n22763 , n22764 , n22059 );
nor ( n22766 , n22762 , n22765 );
or ( n22767 , n22766 , n22069 );
nand ( n22768 , n47 , n22105 );
nand ( n22769 , n22767 , n2 , n22768 );
and ( n22770 , n1472 , n22611 );
and ( n22771 , n21929 , n22742 );
nor ( n22772 , n679 , n22742 );
not ( n22773 , n22609 );
nor ( n22774 , n22771 , n22772 , n22773 );
nor ( n22775 , n22770 , n22774 );
not ( n22776 , n22623 );
not ( n22777 , n22776 );
or ( n22778 , n22775 , n22777 );
nand ( n22779 , n46 , n22627 );
nand ( n22780 , n22778 , n2 , n22779 );
and ( n22781 , n1291 , n22752 );
and ( n22782 , n22408 , n22740 );
nor ( n22783 , n676 , n22617 );
not ( n22784 , n22609 );
nor ( n22785 , n22782 , n22783 , n22784 );
nor ( n22786 , n22781 , n22785 );
or ( n22787 , n22786 , n22747 );
nand ( n22788 , n47 , n22627 );
nand ( n22789 , n22787 , n2 , n22788 );
and ( n22790 , n1445 , n22611 );
and ( n22791 , n21886 , n22615 );
nor ( n22792 , n680 , n22617 );
nor ( n22793 , n22791 , n22792 , n22744 );
nor ( n22794 , n22790 , n22793 );
or ( n22795 , n22794 , n22777 );
nand ( n22796 , n42 , n22627 );
nand ( n22797 , n22795 , n2 , n22796 );
and ( n22798 , n1280 , n22752 );
not ( n22799 , n22739 );
and ( n22800 , n21874 , n22799 );
nor ( n22801 , n682 , n22617 );
not ( n22802 , n22609 );
nor ( n22803 , n22800 , n22801 , n22802 );
nor ( n22804 , n22798 , n22803 );
not ( n22805 , n22624 );
or ( n22806 , n22804 , n22805 );
nand ( n22807 , n38 , n22627 );
nand ( n22808 , n22806 , n2 , n22807 );
and ( n22809 , n1441 , n22611 );
not ( n22810 , n22614 );
and ( n22811 , n21899 , n22810 );
nor ( n22812 , n683 , n22617 );
not ( n22813 , n22609 );
nor ( n22814 , n22811 , n22812 , n22813 );
nor ( n22815 , n22809 , n22814 );
not ( n22816 , n22776 );
or ( n22817 , n22815 , n22816 );
nand ( n22818 , n39 , n22627 );
nand ( n22819 , n22817 , n2 , n22818 );
and ( n22820 , n1440 , n22752 );
not ( n22821 , n22614 );
and ( n22822 , n21908 , n22821 );
nor ( n22823 , n684 , n22617 );
nor ( n22824 , n22822 , n22823 , n22813 );
nor ( n22825 , n22820 , n22824 );
or ( n22826 , n22825 , n22805 );
nand ( n22827 , n41 , n22627 );
nand ( n22828 , n22826 , n2 , n22827 );
and ( n22829 , n1281 , n22752 );
and ( n22830 , n21917 , n22742 );
nor ( n22831 , n685 , n22617 );
nor ( n22832 , n22830 , n22831 , n22610 );
nor ( n22833 , n22829 , n22832 );
or ( n22834 , n22833 , n22777 );
buf ( n22835 , n22622 );
nand ( n22836 , n37 , n22835 );
nand ( n22837 , n22834 , n2 , n22836 );
and ( n22838 , n1461 , n22752 );
not ( n22839 , n175 );
and ( n22840 , n22839 , n22810 );
nor ( n22841 , n686 , n22617 );
nor ( n22842 , n22840 , n22841 , n22619 );
nor ( n22843 , n22838 , n22842 );
or ( n22844 , n22843 , n22777 );
nand ( n22845 , n48 , n22627 );
nand ( n22846 , n22844 , n2 , n22845 );
and ( n22847 , n1462 , n22611 );
and ( n22848 , n21939 , n22821 );
not ( n22849 , n22739 );
nor ( n22850 , n687 , n22849 );
nor ( n22851 , n22848 , n22850 , n22744 );
nor ( n22852 , n22847 , n22851 );
not ( n22853 , n22776 );
or ( n22854 , n22852 , n22853 );
nand ( n22855 , n45 , n22627 );
nand ( n22856 , n22854 , n2 , n22855 );
and ( n22857 , n1332 , n22059 );
and ( n22858 , n22839 , n22061 );
nor ( n22859 , n688 , n22061 );
nor ( n22860 , n22858 , n22859 , n22059 );
nor ( n22861 , n22857 , n22860 );
or ( n22862 , n22861 , n22299 );
nand ( n22863 , n48 , n22105 );
nand ( n22864 , n22862 , n2 , n22863 );
and ( n22865 , n720 , n18627 );
not ( n22866 , n17618 );
nand ( n22867 , n22866 , n17639 );
not ( n22868 , n17636 );
and ( n22869 , n22867 , n22868 );
or ( n22870 , n22867 , n22868 );
nand ( n22871 , n22870 , n15095 );
nor ( n22872 , n22869 , n22871 );
nor ( n22873 , n22865 , n22872 );
or ( n22874 , n1826 , n22873 );
and ( n22875 , n720 , n17677 );
nor ( n22876 , n22875 , n17678 );
or ( n22877 , n15090 , n22876 );
nand ( n22878 , n22874 , n22877 );
and ( n22879 , n1272 , n22878 );
and ( n22880 , n1278 , n22752 );
and ( n22881 , n21949 , n22799 );
nor ( n22882 , n722 , n22849 );
nor ( n22883 , n22881 , n22882 , n22744 );
nor ( n22884 , n22880 , n22883 );
or ( n22885 , n22884 , n22853 );
nand ( n22886 , n52 , n22627 );
nand ( n22887 , n22885 , n2 , n22886 );
and ( n22888 , n1282 , n22611 );
and ( n22889 , n22225 , n22810 );
nor ( n22890 , n724 , n22617 );
nor ( n22891 , n22889 , n22890 , n22802 );
nor ( n22892 , n22888 , n22891 );
or ( n22893 , n22892 , n22805 );
nand ( n22894 , n36 , n22627 );
nand ( n22895 , n22893 , n2 , n22894 );
not ( n22896 , n22751 );
and ( n22897 , n1082 , n22742 );
and ( n22898 , n725 , n22739 );
nor ( n22899 , n22897 , n22898 );
not ( n22900 , n22899 );
and ( n22901 , n22896 , n22900 );
and ( n22902 , n1434 , n22752 );
nor ( n22903 , n22901 , n22902 );
not ( n22904 , n22624 );
or ( n22905 , n22903 , n22904 );
nand ( n22906 , n35 , n22627 );
nand ( n22907 , n22905 , n2 , n22906 );
and ( n22908 , n1413 , n22752 );
and ( n22909 , n21960 , n22799 );
nor ( n22910 , n726 , n22617 );
nor ( n22911 , n22909 , n22910 , n22813 );
nor ( n22912 , n22908 , n22911 );
or ( n22913 , n22912 , n22805 );
nand ( n22914 , n34 , n22627 );
nand ( n22915 , n22913 , n2 , n22914 );
and ( n22916 , n1460 , n22752 );
not ( n22917 , n22614 );
and ( n22918 , n21568 , n22917 );
nor ( n22919 , n727 , n22742 );
nor ( n22920 , n22918 , n22919 , n22773 );
nor ( n22921 , n22916 , n22920 );
or ( n22922 , n22921 , n22747 );
nand ( n22923 , n33 , n22835 );
nand ( n22924 , n22922 , n2 , n22923 );
and ( n22925 , n1412 , n22611 );
and ( n22926 , n21987 , n22821 );
nor ( n22927 , n729 , n22849 );
nor ( n22928 , n22926 , n22927 , n22619 );
nor ( n22929 , n22925 , n22928 );
or ( n22930 , n22929 , n22816 );
nand ( n22931 , n32 , n22627 );
nand ( n22932 , n22930 , n2 , n22931 );
not ( n22933 , n22751 );
and ( n22934 , n143 , n22742 );
and ( n22935 , n730 , n22739 );
nor ( n22936 , n22934 , n22935 );
not ( n22937 , n22936 );
and ( n22938 , n22933 , n22937 );
and ( n22939 , n1279 , n22752 );
nor ( n22940 , n22938 , n22939 );
or ( n22941 , n22940 , n22904 );
nand ( n22942 , n40 , n22627 );
nand ( n22943 , n22941 , n2 , n22942 );
and ( n22944 , n1285 , n22752 );
and ( n22945 , n22005 , n22917 );
nor ( n22946 , n731 , n22742 );
nor ( n22947 , n22945 , n22946 , n22802 );
nor ( n22948 , n22944 , n22947 );
or ( n22949 , n22948 , n22816 );
nand ( n22950 , n29 , n22835 );
nand ( n22951 , n22949 , n2 , n22950 );
and ( n22952 , n1286 , n22752 );
and ( n22953 , n22014 , n22917 );
nor ( n22954 , n732 , n22617 );
nor ( n22955 , n22953 , n22954 , n22802 );
nor ( n22956 , n22952 , n22955 );
or ( n22957 , n22956 , n22816 );
nand ( n22958 , n28 , n22627 );
nand ( n22959 , n22957 , n2 , n22958 );
and ( n22960 , n1284 , n22611 );
and ( n22961 , n22364 , n22742 );
nor ( n22962 , n733 , n22617 );
nor ( n22963 , n22961 , n22962 , n22813 );
nor ( n22964 , n22960 , n22963 );
not ( n22965 , n22776 );
or ( n22966 , n22964 , n22965 );
nand ( n22967 , n30 , n22627 );
nand ( n22968 , n22966 , n2 , n22967 );
and ( n22969 , n785 , n21169 );
and ( n22970 , n548 , n21093 );
and ( n22971 , n471 , n20914 );
nor ( n22972 , n22969 , n22970 , n22971 );
and ( n22973 , n675 , n20591 );
and ( n22974 , n899 , n20438 );
nor ( n22975 , n22973 , n22974 );
nand ( n22976 , n22972 , n22975 );
and ( n22977 , n1475 , n22611 );
not ( n22978 , n253 );
and ( n22979 , n22978 , n22742 );
nor ( n22980 , n734 , n22849 );
nor ( n22981 , n22979 , n22980 , n22773 );
nor ( n22982 , n22977 , n22981 );
or ( n22983 , n22982 , n22965 );
nand ( n22984 , n25 , n22627 );
nand ( n22985 , n22983 , n2 , n22984 );
and ( n22986 , n1289 , n22611 );
and ( n22987 , n22033 , n22742 );
nor ( n22988 , n737 , n22849 );
nor ( n22989 , n22987 , n22988 , n22756 );
nor ( n22990 , n22986 , n22989 );
or ( n22991 , n22990 , n22625 );
nand ( n22992 , n22 , n22835 );
nand ( n22993 , n22991 , n2 , n22992 );
and ( n22994 , n1292 , n22611 );
and ( n22995 , n22051 , n22821 );
nor ( n22996 , n739 , n22617 );
nor ( n22997 , n22995 , n22996 , n22773 );
nor ( n22998 , n22994 , n22997 );
or ( n22999 , n22998 , n22965 );
nand ( n23000 , n44 , n22627 );
nand ( n23001 , n22999 , n2 , n23000 );
and ( n23002 , n1316 , n22059 );
and ( n23003 , n22373 , n22061 );
nor ( n23004 , n742 , n22061 );
nor ( n23005 , n23003 , n23004 , n22059 );
nor ( n23006 , n23002 , n23005 );
or ( n23007 , n23006 , n22299 );
nand ( n23008 , n40 , n22071 );
nand ( n23009 , n23007 , n2 , n23008 );
and ( n23010 , n1377 , n22059 );
and ( n23011 , n22631 , n22061 );
nor ( n23012 , n743 , n22061 );
nor ( n23013 , n23011 , n23012 , n22059 );
nor ( n23014 , n23010 , n23013 );
or ( n23015 , n23014 , n22079 );
nand ( n23016 , n35 , n22071 );
nand ( n23017 , n23015 , n2 , n23016 );
and ( n23018 , n1330 , n22059 );
and ( n23019 , n22705 , n22061 );
nor ( n23020 , n745 , n22061 );
nor ( n23021 , n23019 , n23020 , n22059 );
nor ( n23022 , n23018 , n23021 );
or ( n23023 , n23022 , n22138 );
nand ( n23024 , n23 , n22071 );
nand ( n23025 , n23023 , n2 , n23024 );
and ( n23026 , n1410 , n21566 );
and ( n23027 , n22408 , n22315 );
nor ( n23028 , n769 , n21573 );
nor ( n23029 , n23027 , n23028 , n21565 );
nor ( n23030 , n23026 , n23029 );
or ( n23031 , n23030 , n22332 );
nand ( n23032 , n47 , n21598 );
nand ( n23033 , n23031 , n2 , n23032 );
and ( n23034 , n1344 , n21566 );
and ( n23035 , n21996 , n22706 );
nor ( n23036 , n785 , n22327 );
nor ( n23037 , n23035 , n23036 , n21565 );
nor ( n23038 , n23034 , n23037 );
or ( n23039 , n23038 , n22647 );
nand ( n23040 , n31 , n22446 );
nand ( n23041 , n23039 , n2 , n23040 );
and ( n23042 , n1195 , n21566 );
and ( n23043 , n22005 , n22660 );
nor ( n23044 , n786 , n22327 );
nor ( n23045 , n23043 , n23044 , n21565 );
nor ( n23046 , n23042 , n23045 );
or ( n23047 , n23046 , n22320 );
nand ( n23048 , n29 , n21598 );
nand ( n23049 , n23047 , n2 , n23048 );
and ( n23050 , n1185 , n21566 );
and ( n23051 , n22978 , n21571 );
nor ( n23052 , n787 , n21573 );
nor ( n23053 , n23051 , n23052 , n21565 );
nor ( n23054 , n23050 , n23053 );
or ( n23055 , n23054 , n22320 );
nand ( n23056 , n25 , n21598 );
nand ( n23057 , n23055 , n2 , n23056 );
and ( n23058 , n1353 , n21566 );
and ( n23059 , n21848 , n21571 );
nor ( n23060 , n788 , n21573 );
nor ( n23061 , n23059 , n23060 , n21565 );
nor ( n23062 , n23058 , n23061 );
or ( n23063 , n23062 , n22320 );
nand ( n23064 , n43 , n21598 );
nand ( n23065 , n23063 , n2 , n23064 );
and ( n23066 , n798 , n16747 );
not ( n23067 , n17539 );
nand ( n23068 , n23067 , n17560 );
not ( n23069 , n17557 );
and ( n23070 , n23068 , n23069 );
or ( n23071 , n23068 , n23069 );
nand ( n23072 , n23071 , n16266 );
nor ( n23073 , n23070 , n23072 );
nor ( n23074 , n23066 , n23073 );
or ( n23075 , n1828 , n23074 );
and ( n23076 , n798 , n17597 );
nor ( n23077 , n23076 , n17598 );
or ( n23078 , n16258 , n23077 );
nand ( n23079 , n23075 , n23078 );
and ( n23080 , n1240 , n23079 );
not ( n23081 , n1231 );
or ( n23082 , n23081 , n22549 );
or ( n23083 , n12538 , n22552 );
and ( n23084 , n1268 , n20416 );
and ( n23085 , n1256 , n20428 );
and ( n23086 , n1248 , n20432 );
nor ( n23087 , n23084 , n23085 , n23086 );
nand ( n23088 , n23082 , n23083 , n23087 );
or ( n23089 , n19230 , n22308 );
nand ( n23090 , n23089 , n2 , n22301 );
or ( n23091 , n17047 , n22427 );
nand ( n23092 , n23091 , n2 , n23056 );
or ( n23093 , n17060 , n22681 );
nand ( n23094 , n23093 , n2 , n22322 );
or ( n23095 , n17098 , n22681 );
nand ( n23096 , n23095 , n2 , n23048 );
or ( n23097 , n16937 , n22473 );
nand ( n23098 , n23097 , n2 , n21993 );
or ( n23099 , n16905 , n21955 );
nand ( n23100 , n23099 , n2 , n21831 );
or ( n23101 , n16931 , n21955 );
nand ( n23102 , n23101 , n2 , n22370 );
or ( n23103 , n16910 , n22473 );
nand ( n23104 , n23103 , n2 , n22030 );
or ( n23105 , n16861 , n22904 );
nand ( n23106 , n31 , n22835 );
nand ( n23107 , n23105 , n2 , n23106 );
or ( n23108 , n16858 , n22625 );
nand ( n23109 , n23108 , n2 , n22967 );
or ( n23110 , n16855 , n22625 );
nand ( n23111 , n23110 , n2 , n22950 );
or ( n23112 , n16836 , n22904 );
nand ( n23113 , n26 , n22627 );
nand ( n23114 , n23112 , n2 , n23113 );
not ( n23115 , n2 );
not ( n23116 , n21801 );
and ( n23117 , n36 , n23116 );
and ( n23118 , n1526 , n21801 );
nor ( n23119 , n23117 , n23118 );
nor ( n23120 , n23115 , n23119 );
nand ( n23121 , n2 , n29 );
nor ( n23122 , n17 , n18 );
not ( n23123 , n23122 );
buf ( n23124 , n23123 );
not ( n23125 , n23124 );
not ( n23126 , n23125 );
or ( n23127 , n23126 , n21760 );
buf ( n23128 , n23127 );
not ( n23129 , n23128 );
not ( n23130 , n23129 );
or ( n23131 , n23121 , n23130 );
nand ( n23132 , n1181 , n1858 );
not ( n23133 , n2 );
not ( n23134 , n23127 );
nor ( n23135 , n23133 , n23134 );
nand ( n23136 , n1293 , n23132 , n23135 );
nand ( n23137 , n23131 , n23136 );
not ( n23138 , n21844 );
nand ( n23139 , n1298 , n23138 );
nand ( n23140 , n23139 , n2 , n21883 );
or ( n23141 , n16928 , n22415 );
nand ( n23142 , n23141 , n2 , n22011 );
or ( n23143 , n16912 , n21934 );
nand ( n23144 , n27 , n21830 );
nand ( n23145 , n23143 , n2 , n23144 );
or ( n23146 , n16908 , n22415 );
nand ( n23147 , n23146 , n2 , n21871 );
or ( n23148 , n16901 , n22019 );
nand ( n23149 , n23 , n21830 );
nand ( n23150 , n23148 , n2 , n23149 );
or ( n23151 , n19186 , n22415 );
nand ( n23152 , n23151 , n2 , n22039 );
buf ( n23153 , n23124 );
buf ( n23154 , n23153 );
or ( n23155 , n23154 , n21798 );
buf ( n23156 , n23155 );
not ( n23157 , n23156 );
not ( n23158 , n23157 );
or ( n23159 , n23121 , n23158 );
nand ( n23160 , n1254 , n1858 );
not ( n23161 , n2 );
not ( n23162 , n23155 );
nor ( n23163 , n23161 , n23162 );
nand ( n23164 , n1313 , n23160 , n23163 );
nand ( n23165 , n23159 , n23164 );
not ( n23166 , n22105 );
nand ( n23167 , n1314 , n23166 );
nand ( n23168 , n23167 , n2 , n22123 );
or ( n23169 , n17011 , n22273 );
nand ( n23170 , n23169 , n2 , n22250 );
or ( n23171 , n17005 , n22273 );
nand ( n23172 , n23171 , n2 , n22266 );
or ( n23173 , n17002 , n22071 );
nand ( n23174 , n23173 , n2 , n22736 );
or ( n23175 , n16999 , n22071 );
nand ( n23176 , n23175 , n2 , n22275 );
or ( n23177 , n16983 , n22138 );
nand ( n23178 , n23177 , n2 , n22292 );
or ( n23179 , n16981 , n22308 );
nand ( n23180 , n26 , n22071 );
nand ( n23181 , n23179 , n2 , n23180 );
or ( n23182 , n16979 , n22240 );
nand ( n23183 , n25 , n22071 );
nand ( n23184 , n23182 , n2 , n23183 );
or ( n23185 , n16972 , n22230 );
nand ( n23186 , n23185 , n2 , n23024 );
or ( n23187 , n23154 , n21749 );
buf ( n23188 , n23187 );
not ( n23189 , n23188 );
not ( n23190 , n23189 );
or ( n23191 , n23121 , n23190 );
nand ( n23192 , n1267 , n1858 );
not ( n23193 , n2 );
not ( n23194 , n23187 );
nor ( n23195 , n23193 , n23194 );
nand ( n23196 , n1335 , n23192 , n23195 );
nand ( n23197 , n23191 , n23196 );
or ( n23198 , n17067 , n22436 );
nand ( n23199 , n23198 , n2 , n22694 );
or ( n23200 , n17051 , n22427 );
nand ( n23201 , n26 , n21598 );
nand ( n23202 , n23200 , n2 , n23201 );
or ( n23203 , n23154 , n21591 );
buf ( n23204 , n23203 );
not ( n23205 , n23204 );
not ( n23206 , n23205 );
or ( n23207 , n23121 , n23206 );
nand ( n23208 , n1229 , n1858 );
not ( n23209 , n2 );
not ( n23210 , n23203 );
nor ( n23211 , n23209 , n23210 );
nand ( n23212 , n1354 , n23208 , n23211 );
nand ( n23213 , n23207 , n23212 );
or ( n23214 , n17043 , n21596 );
nand ( n23215 , n23214 , n2 , n22712 );
or ( n23216 , n16941 , n21934 );
nand ( n23217 , n23216 , n2 , n21974 );
or ( n23218 , n16976 , n22240 );
nand ( n23219 , n23218 , n2 , n22072 );
or ( n23220 , n16997 , n22240 );
nand ( n23221 , n23220 , n2 , n22283 );
or ( n23222 , n18949 , n22436 );
nand ( n23223 , n23222 , n2 , n22720 );
or ( n23224 , n16839 , n22965 );
nand ( n23225 , n23224 , n2 , n22760 );
or ( n23226 , n17008 , n22138 );
nand ( n23227 , n23226 , n2 , n22258 );
or ( n23228 , n16868 , n22853 );
nand ( n23229 , n23228 , n2 , n22923 );
or ( n23230 , n16832 , n22853 );
nand ( n23231 , n23230 , n2 , n22984 );
not ( n23232 , n2 );
and ( n23233 , n31 , n21764 );
and ( n23234 , n1476 , n21763 );
nor ( n23235 , n23233 , n23234 );
nor ( n23236 , n23232 , n23235 );
not ( n23237 , n2 );
not ( n23238 , n21763 );
and ( n23239 , n25 , n23238 );
and ( n23240 , n1477 , n21763 );
nor ( n23241 , n23239 , n23240 );
nor ( n23242 , n23237 , n23241 );
not ( n23243 , n2 );
not ( n23244 , n21752 );
and ( n23245 , n24 , n23244 );
and ( n23246 , n1478 , n21752 );
nor ( n23247 , n23245 , n23246 );
nor ( n23248 , n23243 , n23247 );
not ( n23249 , n2 );
and ( n23250 , n34 , n23238 );
and ( n23251 , n1479 , n21763 );
nor ( n23252 , n23250 , n23251 );
nor ( n23253 , n23249 , n23252 );
not ( n23254 , n2 );
and ( n23255 , n32 , n23238 );
and ( n23256 , n1480 , n21763 );
nor ( n23257 , n23255 , n23256 );
nor ( n23258 , n23254 , n23257 );
not ( n23259 , n2 );
not ( n23260 , n21763 );
and ( n23261 , n24 , n23260 );
and ( n23262 , n1482 , n21763 );
nor ( n23263 , n23261 , n23262 );
nor ( n23264 , n23259 , n23263 );
not ( n23265 , n2 );
and ( n23266 , n33 , n23260 );
and ( n23267 , n1483 , n21763 );
nor ( n23268 , n23266 , n23267 );
nor ( n23269 , n23265 , n23268 );
not ( n23270 , n2 );
and ( n23271 , n35 , n23260 );
and ( n23272 , n1484 , n21763 );
nor ( n23273 , n23271 , n23272 );
nor ( n23274 , n23270 , n23273 );
not ( n23275 , n2 );
and ( n23276 , n36 , n23260 );
and ( n23277 , n1486 , n21763 );
nor ( n23278 , n23276 , n23277 );
nor ( n23279 , n23275 , n23278 );
not ( n23280 , n2 );
not ( n23281 , n21752 );
and ( n23282 , n28 , n23281 );
and ( n23283 , n1488 , n21752 );
nor ( n23284 , n23282 , n23283 );
nor ( n23285 , n23280 , n23284 );
not ( n23286 , n2 );
and ( n23287 , n27 , n23281 );
and ( n23288 , n1491 , n21752 );
nor ( n23289 , n23287 , n23288 );
nor ( n23290 , n23286 , n23289 );
not ( n23291 , n2 );
and ( n23292 , n27 , n21764 );
and ( n23293 , n1492 , n21763 );
nor ( n23294 , n23292 , n23293 );
nor ( n23295 , n23291 , n23294 );
not ( n23296 , n2 );
and ( n23297 , n25 , n23281 );
and ( n23298 , n1493 , n21752 );
nor ( n23299 , n23297 , n23298 );
nor ( n23300 , n23296 , n23299 );
not ( n23301 , n2 );
nand ( n23302 , n21743 , n21592 );
buf ( n23303 , n23302 );
not ( n23304 , n23303 );
and ( n23305 , n27 , n23304 );
and ( n23306 , n1503 , n23303 );
nor ( n23307 , n23305 , n23306 );
nor ( n23308 , n23301 , n23307 );
not ( n23309 , n2 );
and ( n23310 , n25 , n23304 );
and ( n23311 , n1504 , n23303 );
nor ( n23312 , n23310 , n23311 );
nor ( n23313 , n23309 , n23312 );
not ( n23314 , n2 );
and ( n23315 , n23 , n23304 );
and ( n23316 , n1505 , n23303 );
nor ( n23317 , n23315 , n23316 );
nor ( n23318 , n23314 , n23317 );
not ( n23319 , n2 );
not ( n23320 , n23303 );
and ( n23321 , n36 , n23320 );
and ( n23322 , n1506 , n23303 );
nor ( n23323 , n23321 , n23322 );
nor ( n23324 , n23319 , n23323 );
not ( n23325 , n2 );
and ( n23326 , n35 , n23320 );
and ( n23327 , n1507 , n23303 );
nor ( n23328 , n23326 , n23327 );
nor ( n23329 , n23325 , n23328 );
not ( n23330 , n2 );
and ( n23331 , n32 , n23320 );
and ( n23332 , n1508 , n23303 );
nor ( n23333 , n23331 , n23332 );
nor ( n23334 , n23330 , n23333 );
not ( n23335 , n2 );
and ( n23336 , n28 , n23238 );
and ( n23337 , n1510 , n21763 );
nor ( n23338 , n23336 , n23337 );
nor ( n23339 , n23335 , n23338 );
not ( n23340 , n2 );
and ( n23341 , n26 , n21764 );
and ( n23342 , n1511 , n21763 );
nor ( n23343 , n23341 , n23342 );
nor ( n23344 , n23340 , n23343 );
not ( n23345 , n2 );
and ( n23346 , n27 , n23116 );
and ( n23347 , n1512 , n21801 );
nor ( n23348 , n23346 , n23347 );
nor ( n23349 , n23345 , n23348 );
not ( n23350 , n2 );
and ( n23351 , n25 , n21802 );
and ( n23352 , n1514 , n21801 );
nor ( n23353 , n23351 , n23352 );
nor ( n23354 , n23350 , n23353 );
not ( n23355 , n2 );
and ( n23356 , n23 , n23116 );
and ( n23357 , n1515 , n21801 );
nor ( n23358 , n23356 , n23357 );
nor ( n23359 , n23355 , n23358 );
not ( n23360 , n2 );
not ( n23361 , n21801 );
and ( n23362 , n35 , n23361 );
and ( n23363 , n1516 , n21801 );
nor ( n23364 , n23362 , n23363 );
nor ( n23365 , n23360 , n23364 );
not ( n23366 , n2 );
and ( n23367 , n33 , n23361 );
and ( n23368 , n1518 , n21801 );
nor ( n23369 , n23367 , n23368 );
nor ( n23370 , n23366 , n23369 );
not ( n23371 , n2 );
and ( n23372 , n26 , n23244 );
and ( n23373 , n1519 , n21752 );
nor ( n23374 , n23372 , n23373 );
nor ( n23375 , n23371 , n23374 );
not ( n23376 , n2 );
and ( n23377 , n32 , n23244 );
and ( n23378 , n1520 , n21752 );
nor ( n23379 , n23377 , n23378 );
nor ( n23380 , n23376 , n23379 );
not ( n23381 , n2 );
and ( n23382 , n31 , n23361 );
and ( n23383 , n1522 , n21801 );
nor ( n23384 , n23382 , n23383 );
nor ( n23385 , n23381 , n23384 );
not ( n23386 , n2 );
and ( n23387 , n36 , n23244 );
and ( n23388 , n1523 , n21752 );
nor ( n23389 , n23387 , n23388 );
nor ( n23390 , n23386 , n23389 );
not ( n23391 , n2 );
and ( n23392 , n34 , n21802 );
and ( n23393 , n1524 , n21801 );
nor ( n23394 , n23392 , n23393 );
nor ( n23395 , n23391 , n23394 );
not ( n23396 , n2 );
and ( n23397 , n24 , n21802 );
and ( n23398 , n1525 , n21801 );
nor ( n23399 , n23397 , n23398 );
nor ( n23400 , n23396 , n23399 );
not ( n23401 , n2 );
not ( n23402 , n23303 );
and ( n23403 , n28 , n23402 );
and ( n23404 , n1529 , n23303 );
nor ( n23405 , n23403 , n23404 );
nor ( n23406 , n23401 , n23405 );
not ( n23407 , n2 );
and ( n23408 , n35 , n21753 );
and ( n23409 , n1531 , n21752 );
nor ( n23410 , n23408 , n23409 );
nor ( n23411 , n23407 , n23410 );
not ( n23412 , n2 );
and ( n23413 , n31 , n23402 );
and ( n23414 , n1532 , n23303 );
nor ( n23415 , n23413 , n23414 );
nor ( n23416 , n23412 , n23415 );
not ( n23417 , n2 );
and ( n23418 , n34 , n23304 );
and ( n23419 , n1534 , n23303 );
nor ( n23420 , n23418 , n23419 );
nor ( n23421 , n23417 , n23420 );
not ( n23422 , n2 );
and ( n23423 , n26 , n23402 );
and ( n23424 , n1535 , n23303 );
nor ( n23425 , n23423 , n23424 );
nor ( n23426 , n23422 , n23425 );
not ( n23427 , n2 );
and ( n23428 , n24 , n23320 );
and ( n23429 , n1536 , n23303 );
nor ( n23430 , n23428 , n23429 );
nor ( n23431 , n23427 , n23430 );
not ( n23432 , n2 );
and ( n23433 , n33 , n23281 );
and ( n23434 , n1540 , n21752 );
nor ( n23435 , n23433 , n23434 );
nor ( n23436 , n23432 , n23435 );
not ( n23437 , n2 );
and ( n23438 , n31 , n21753 );
and ( n23439 , n1541 , n21752 );
nor ( n23440 , n23438 , n23439 );
nor ( n23441 , n23437 , n23440 );
and ( n23442 , n757 , n20591 );
and ( n23443 , n592 , n20418 );
nor ( n23444 , n23442 , n23443 );
and ( n23445 , n984 , n20624 );
and ( n23446 , n505 , n20598 );
and ( n23447 , n458 , n20600 );
nor ( n23448 , n23445 , n23446 , n23447 );
nand ( n23449 , n23444 , n23448 );
and ( n23450 , n586 , n21118 );
and ( n23451 , n499 , n20892 );
and ( n23452 , n452 , n20875 );
nor ( n23453 , n23450 , n23451 , n23452 );
and ( n23454 , n766 , n20591 );
and ( n23455 , n967 , n20438 );
nor ( n23456 , n23454 , n23455 );
nand ( n23457 , n23453 , n23456 );
not ( n23458 , n2 );
and ( n23459 , n32 , n23361 );
and ( n23460 , n1517 , n21801 );
nor ( n23461 , n23459 , n23460 );
nor ( n23462 , n23458 , n23461 );
not ( n23463 , n14490 );
nand ( n23464 , n14494 , n14488 );
not ( n23465 , n23464 );
or ( n23466 , n23463 , n23465 );
or ( n23467 , n14490 , n23464 );
nand ( n23468 , n23466 , n23467 );
and ( n23469 , n1351 , n22312 );
and ( n23470 , n22839 , n21573 );
nor ( n23471 , n761 , n21573 );
nor ( n23472 , n23470 , n23471 , n21565 );
nor ( n23473 , n23469 , n23472 );
or ( n23474 , n23473 , n22359 );
nand ( n23475 , n48 , n21598 );
nand ( n23476 , n23474 , n2 , n23475 );
and ( n23477 , n667 , n20890 );
and ( n23478 , n622 , n20912 );
and ( n23479 , n524 , n20875 );
nor ( n23480 , n23477 , n23478 , n23479 );
and ( n23481 , n814 , n20591 );
and ( n23482 , n973 , n20438 );
nor ( n23483 , n23481 , n23482 );
nand ( n23484 , n23480 , n23483 );
not ( n23485 , n2 );
and ( n23486 , n33 , n23402 );
and ( n23487 , n1509 , n23303 );
nor ( n23488 , n23486 , n23487 );
nor ( n23489 , n23485 , n23488 );
not ( n23490 , n2 );
and ( n23491 , n26 , n23116 );
and ( n23492 , n1513 , n21801 );
nor ( n23493 , n23491 , n23492 );
nor ( n23494 , n23490 , n23493 );
or ( n23495 , n16273 , n22549 );
or ( n23496 , n13623 , n22552 );
and ( n23497 , n1162 , n20416 );
and ( n23498 , n1212 , n20428 );
and ( n23499 , n1250 , n20432 );
nor ( n23500 , n23497 , n23498 , n23499 );
nand ( n23501 , n23495 , n23496 , n23500 );
and ( n23502 , n655 , n20890 );
and ( n23503 , n550 , n20912 );
and ( n23504 , n473 , n21172 );
nor ( n23505 , n23502 , n23503 , n23504 );
and ( n23506 , n732 , n20591 );
and ( n23507 , n953 , n20438 );
nor ( n23508 , n23506 , n23507 );
nand ( n23509 , n23505 , n23508 );
not ( n23510 , n2 );
not ( n23511 , n23204 );
and ( n23512 , n26 , n23511 );
and ( n23513 , n1273 , n23204 );
nor ( n23514 , n23512 , n23513 );
nor ( n23515 , n23510 , n23514 );
not ( n23516 , n2 );
not ( n23517 , n23204 );
and ( n23518 , n45 , n23517 );
and ( n23519 , n1271 , n23204 );
nor ( n23520 , n23518 , n23519 );
nor ( n23521 , n23516 , n23520 );
not ( n23522 , n2 );
not ( n23523 , n16 );
and ( n23524 , n23523 , n21739 );
nand ( n23525 , n15943 , n15947 , n21586 );
not ( n23526 , n23525 );
nand ( n23527 , n23526 , n21590 );
not ( n23528 , n23527 );
and ( n23529 , n23524 , n23528 );
and ( n23530 , n49 , n23529 );
not ( n23531 , n23529 );
and ( n23532 , n1198 , n23531 );
nor ( n23533 , n23530 , n23532 );
nor ( n23534 , n23522 , n23533 );
not ( n23535 , n2 );
not ( n23536 , n23204 );
and ( n23537 , n48 , n23536 );
and ( n23538 , n1270 , n23204 );
nor ( n23539 , n23537 , n23538 );
nor ( n23540 , n23535 , n23539 );
not ( n23541 , n2 );
and ( n23542 , n40 , n23517 );
and ( n23543 , n1269 , n23204 );
nor ( n23544 , n23542 , n23543 );
nor ( n23545 , n23541 , n23544 );
not ( n23546 , n2 );
not ( n23547 , n23188 );
and ( n23548 , n39 , n23547 );
and ( n23549 , n1267 , n23188 );
nor ( n23550 , n23548 , n23549 );
nor ( n23551 , n23546 , n23550 );
not ( n23552 , n2 );
not ( n23553 , n23188 );
and ( n23554 , n28 , n23553 );
and ( n23555 , n1266 , n23188 );
nor ( n23556 , n23554 , n23555 );
nor ( n23557 , n23552 , n23556 );
not ( n23558 , n2 );
not ( n23559 , n23188 );
and ( n23560 , n31 , n23559 );
and ( n23561 , n1265 , n23188 );
nor ( n23562 , n23560 , n23561 );
nor ( n23563 , n23558 , n23562 );
not ( n23564 , n2 );
not ( n23565 , n23188 );
and ( n23566 , n33 , n23565 );
and ( n23567 , n1263 , n23188 );
nor ( n23568 , n23566 , n23567 );
nor ( n23569 , n23564 , n23568 );
not ( n23570 , n2 );
not ( n23571 , n23188 );
and ( n23572 , n35 , n23571 );
and ( n23573 , n1262 , n23188 );
nor ( n23574 , n23572 , n23573 );
nor ( n23575 , n23570 , n23574 );
not ( n23576 , n21830 );
nand ( n23577 , n1182 , n23576 );
nand ( n23578 , n23577 , n2 , n21946 );
not ( n23579 , n22835 );
nand ( n23580 , n1392 , n23579 );
nand ( n23581 , n49 , n22627 );
nand ( n23582 , n23580 , n2 , n23581 );
not ( n23583 , n2 );
not ( n23584 , n23204 );
and ( n23585 , n43 , n23584 );
and ( n23586 , n1163 , n23204 );
nor ( n23587 , n23585 , n23586 );
nor ( n23588 , n23583 , n23587 );
not ( n23589 , n2 );
not ( n23590 , n23204 );
and ( n23591 , n25 , n23590 );
and ( n23592 , n1388 , n23204 );
nor ( n23593 , n23591 , n23592 );
nor ( n23594 , n23589 , n23593 );
not ( n23595 , n1125 );
not ( n23596 , n1559 );
or ( n23597 , n23595 , n23596 );
nand ( n23598 , n1559 , n1858 );
nand ( n23599 , n23597 , n23598 );
not ( n23600 , n23599 );
and ( n23601 , n455 , n23600 );
and ( n23602 , n147 , n23599 );
nor ( n23603 , n23601 , n23602 );
not ( n23604 , n22151 );
buf ( n23605 , n23604 );
not ( n23606 , n23605 );
not ( n23607 , n23606 );
or ( n23608 , n23607 , n21798 );
not ( n23609 , n23608 );
not ( n23610 , n23609 );
not ( n23611 , n23610 );
or ( n23612 , n23603 , n23611 );
or ( n23613 , n16025 , n23610 );
nand ( n23614 , n23612 , n23613 , n2 );
buf ( n23615 , n23609 );
not ( n23616 , n23615 );
or ( n23617 , n15901 , n23616 );
or ( n23618 , n152 , n23600 );
or ( n23619 , n456 , n23599 );
not ( n23620 , n23609 );
nand ( n23621 , n23618 , n23619 , n23620 );
nand ( n23622 , n23617 , n2 , n23621 );
not ( n23623 , n23615 );
or ( n23624 , n16085 , n23623 );
or ( n23625 , n175 , n23600 );
or ( n23626 , n457 , n23599 );
buf ( n23627 , n23608 );
nand ( n23628 , n23625 , n23626 , n23627 );
nand ( n23629 , n23624 , n2 , n23628 );
or ( n23630 , n16057 , n23623 );
or ( n23631 , n159 , n23600 );
or ( n23632 , n459 , n23599 );
nand ( n23633 , n23631 , n23632 , n23620 );
nand ( n23634 , n23630 , n2 , n23633 );
or ( n23635 , n16065 , n23623 );
or ( n23636 , n1801 , n23600 );
or ( n23637 , n463 , n23599 );
not ( n23638 , n23609 );
nand ( n23639 , n23636 , n23637 , n23638 );
nand ( n23640 , n23635 , n2 , n23639 );
nor ( n23641 , n267 , n1230 );
nand ( n23642 , n23641 , n20194 );
not ( n23643 , n23642 );
nand ( n23644 , n23643 , n465 );
not ( n23645 , n20175 );
nand ( n23646 , n23645 , n1538 , n15377 );
not ( n23647 , n387 );
nor ( n23648 , n1379 , n267 , n20203 );
nand ( n23649 , n23647 , n23648 , n465 );
and ( n23650 , n23644 , n23646 , n23649 );
not ( n23651 , n2 );
nor ( n23652 , n23650 , n23651 );
and ( n23653 , n1304 , n21814 );
and ( n23654 , n22286 , n21887 );
nor ( n23655 , n474 , n21837 );
nor ( n23656 , n23654 , n23655 , n22348 );
nor ( n23657 , n23653 , n23656 );
or ( n23658 , n23657 , n21830 );
nand ( n23659 , n23658 , n2 , n23144 );
and ( n23660 , n486 , n22165 );
and ( n23661 , n152 , n22164 );
nor ( n23662 , n23660 , n23661 );
buf ( n23663 , n22157 );
or ( n23664 , n23662 , n23663 );
or ( n23665 , n15901 , n22510 );
nand ( n23666 , n23664 , n23665 , n2 );
or ( n23667 , n16069 , n23627 );
or ( n23668 , n178 , n23600 );
or ( n23669 , n489 , n23599 );
nand ( n23670 , n23668 , n23669 , n23620 );
nand ( n23671 , n23667 , n2 , n23670 );
and ( n23672 , n495 , n22165 );
and ( n23673 , n140 , n22164 );
nor ( n23674 , n23672 , n23673 );
or ( n23675 , n23674 , n22157 );
or ( n23676 , n16029 , n22533 );
nand ( n23677 , n23675 , n23676 , n2 );
and ( n23678 , n498 , n22165 );
and ( n23679 , n145 , n22164 );
nor ( n23680 , n23678 , n23679 );
or ( n23681 , n23680 , n23663 );
or ( n23682 , n16045 , n22533 );
nand ( n23683 , n23681 , n23682 , n2 );
and ( n23684 , n503 , n22165 );
and ( n23685 , n175 , n22164 );
nor ( n23686 , n23684 , n23685 );
or ( n23687 , n23686 , n23663 );
or ( n23688 , n16085 , n22510 );
nand ( n23689 , n23687 , n23688 , n2 );
and ( n23690 , n505 , n22165 );
and ( n23691 , n157 , n22164 );
nor ( n23692 , n23690 , n23691 );
or ( n23693 , n23692 , n23663 );
or ( n23694 , n16061 , n22185 );
nand ( n23695 , n23693 , n23694 , n2 );
and ( n23696 , n506 , n23600 );
and ( n23697 , n323 , n23599 );
nor ( n23698 , n23696 , n23697 );
or ( n23699 , n23698 , n23611 );
or ( n23700 , n15973 , n23627 );
nand ( n23701 , n23699 , n23700 , n2 );
or ( n23702 , n16001 , n23623 );
or ( n23703 , n415 , n23600 );
or ( n23704 , n507 , n23599 );
nand ( n23705 , n23703 , n23704 , n23627 );
nand ( n23706 , n23702 , n2 , n23705 );
and ( n23707 , n518 , n23600 );
and ( n23708 , n193 , n23599 );
nor ( n23709 , n23707 , n23708 );
or ( n23710 , n23709 , n23611 );
or ( n23711 , n16089 , n23627 );
nand ( n23712 , n23710 , n23711 , n2 );
not ( n23713 , n23615 );
or ( n23714 , n16021 , n23713 );
or ( n23715 , n144 , n23600 );
or ( n23716 , n520 , n23599 );
nand ( n23717 , n23715 , n23716 , n23627 );
nand ( n23718 , n23714 , n2 , n23717 );
or ( n23719 , n16017 , n23713 );
or ( n23720 , n1082 , n23600 );
or ( n23721 , n521 , n23599 );
nand ( n23722 , n23720 , n23721 , n23620 );
nand ( n23723 , n23719 , n2 , n23722 );
or ( n23724 , n16077 , n23627 );
or ( n23725 , n186 , n23600 );
or ( n23726 , n523 , n23599 );
nand ( n23727 , n23725 , n23726 , n23620 );
nand ( n23728 , n23724 , n2 , n23727 );
or ( n23729 , n15997 , n23616 );
or ( n23730 , n1610 , n23600 );
or ( n23731 , n525 , n23599 );
nand ( n23732 , n23730 , n23731 , n23627 );
nand ( n23733 , n23729 , n2 , n23732 );
or ( n23734 , n15989 , n23616 );
or ( n23735 , n352 , n23600 );
or ( n23736 , n526 , n23599 );
nand ( n23737 , n23735 , n23736 , n23627 );
nand ( n23738 , n23734 , n2 , n23737 );
not ( n23739 , n23615 );
or ( n23740 , n15985 , n23739 );
or ( n23741 , n283 , n23600 );
or ( n23742 , n527 , n23599 );
nand ( n23743 , n23741 , n23742 , n23627 );
nand ( n23744 , n23740 , n2 , n23743 );
or ( n23745 , n15993 , n23739 );
or ( n23746 , n383 , n23600 );
or ( n23747 , n528 , n23599 );
nand ( n23748 , n23746 , n23747 , n23627 );
nand ( n23749 , n23745 , n2 , n23748 );
and ( n23750 , n529 , n23600 );
and ( n23751 , n253 , n23599 );
nor ( n23752 , n23750 , n23751 );
or ( n23753 , n23752 , n23611 );
or ( n23754 , n15977 , n23610 );
nand ( n23755 , n23753 , n23754 , n2 );
or ( n23756 , n15981 , n23739 );
or ( n23757 , n284 , n23600 );
or ( n23758 , n530 , n23599 );
nand ( n23759 , n23757 , n23758 , n23638 );
nand ( n23760 , n23756 , n2 , n23759 );
or ( n23761 , n16073 , n23627 );
or ( n23762 , n185 , n23600 );
or ( n23763 , n531 , n23599 );
nand ( n23764 , n23762 , n23763 , n23620 );
nand ( n23765 , n23761 , n2 , n23764 );
or ( n23766 , n15969 , n23616 );
or ( n23767 , n192 , n23600 );
or ( n23768 , n532 , n23599 );
nand ( n23769 , n23767 , n23768 , n23638 );
nand ( n23770 , n23766 , n2 , n23769 );
or ( n23771 , n16049 , n23713 );
or ( n23772 , n151 , n23600 );
or ( n23773 , n534 , n23599 );
nand ( n23774 , n23772 , n23773 , n23638 );
nand ( n23775 , n23771 , n2 , n23774 );
or ( n23776 , n16053 , n23739 );
or ( n23777 , n156 , n23600 );
or ( n23778 , n533 , n23599 );
nand ( n23779 , n23777 , n23778 , n23620 );
nand ( n23780 , n23776 , n2 , n23779 );
and ( n23781 , n536 , n22165 );
and ( n23782 , n1795 , n22164 );
nor ( n23783 , n23781 , n23782 );
or ( n23784 , n23783 , n22157 );
or ( n23785 , n15965 , n22540 );
nand ( n23786 , n23784 , n23785 , n2 );
not ( n23787 , n2 );
or ( n23788 , n1230 , n20180 );
nand ( n23789 , n23788 , n23642 );
and ( n23790 , n538 , n23789 );
not ( n23791 , n15219 );
not ( n23792 , n1379 );
and ( n23793 , n23791 , n23792 );
nor ( n23794 , n23793 , n387 );
nor ( n23795 , n267 , n23794 , n20203 );
nor ( n23796 , n23790 , n23795 );
nor ( n23797 , n23787 , n23796 );
and ( n23798 , n1322 , n22059 );
and ( n23799 , n21977 , n22061 );
nor ( n23800 , n546 , n22061 );
nor ( n23801 , n23799 , n23800 , n22059 );
nor ( n23802 , n23798 , n23801 );
or ( n23803 , n23802 , n22071 );
nand ( n23804 , n51 , n22105 );
nand ( n23805 , n23803 , n2 , n23804 );
and ( n23806 , n1328 , n22059 );
and ( n23807 , n22978 , n22061 );
nor ( n23808 , n552 , n22061 );
nor ( n23809 , n23807 , n23808 , n22059 );
nor ( n23810 , n23806 , n23809 );
or ( n23811 , n23810 , n22071 );
nand ( n23812 , n23811 , n2 , n23183 );
and ( n23813 , n1369 , n22059 );
and ( n23814 , n21848 , n22061 );
nor ( n23815 , n555 , n22061 );
nor ( n23816 , n23814 , n23815 , n22059 );
nor ( n23817 , n23813 , n23816 );
or ( n23818 , n23817 , n22071 );
nand ( n23819 , n43 , n22105 );
nand ( n23820 , n23818 , n2 , n23819 );
or ( n23821 , n16013 , n23713 );
or ( n23822 , n439 , n23600 );
or ( n23823 , n559 , n23599 );
nand ( n23824 , n23822 , n23823 , n23627 );
nand ( n23825 , n23821 , n2 , n23824 );
not ( n23826 , n2 );
not ( n23827 , n23128 );
and ( n23828 , n41 , n23827 );
and ( n23829 , n1372 , n23128 );
nor ( n23830 , n23828 , n23829 );
nor ( n23831 , n23826 , n23830 );
and ( n23832 , n1327 , n22059 );
and ( n23833 , n22024 , n22061 );
nor ( n23834 , n561 , n22061 );
nor ( n23835 , n23833 , n23834 , n22059 );
nor ( n23836 , n23832 , n23835 );
or ( n23837 , n23836 , n22071 );
nand ( n23838 , n23837 , n2 , n23180 );
and ( n23839 , n1290 , n22752 );
and ( n23840 , n21834 , n22740 );
nor ( n23841 , n566 , n22617 );
nor ( n23842 , n23840 , n23841 , n22784 );
nor ( n23843 , n23839 , n23842 );
or ( n23844 , n23843 , n22835 );
nand ( n23845 , n21 , n22627 );
nand ( n23846 , n23844 , n2 , n23845 );
and ( n23847 , n572 , n22165 );
and ( n23848 , n151 , n22164 );
nor ( n23849 , n23847 , n23848 );
or ( n23850 , n23849 , n22157 );
or ( n23851 , n16049 , n22540 );
nand ( n23852 , n23850 , n23851 , n2 );
nand ( n23853 , n22155 , n21592 );
not ( n23854 , n23853 );
not ( n23855 , n23854 );
or ( n23856 , n16029 , n23855 );
not ( n23857 , n1125 );
not ( n23858 , n1588 );
or ( n23859 , n23857 , n23858 );
nand ( n23860 , n1588 , n1858 );
nand ( n23861 , n23859 , n23860 );
not ( n23862 , n23861 );
or ( n23863 , n140 , n23862 );
or ( n23864 , n583 , n23861 );
buf ( n23865 , n23853 );
nand ( n23866 , n23863 , n23864 , n23865 );
nand ( n23867 , n23856 , n2 , n23866 );
and ( n23868 , n1339 , n21566 );
and ( n23869 , n21917 , n22706 );
nor ( n23870 , n584 , n22327 );
nor ( n23871 , n23869 , n23870 , n21565 );
nor ( n23872 , n23868 , n23871 );
or ( n23873 , n23872 , n22446 );
nand ( n23874 , n37 , n21598 );
nand ( n23875 , n23873 , n2 , n23874 );
not ( n23876 , n23854 );
or ( n23877 , n16045 , n23876 );
or ( n23878 , n145 , n23862 );
or ( n23879 , n585 , n23861 );
nand ( n23880 , n23878 , n23879 , n23865 );
nand ( n23881 , n23877 , n2 , n23880 );
and ( n23882 , n586 , n23862 );
and ( n23883 , n136 , n23861 );
nor ( n23884 , n23882 , n23883 );
not ( n23885 , n23865 );
or ( n23886 , n23884 , n23885 );
not ( n23887 , n23853 );
not ( n23888 , n23887 );
or ( n23889 , n16033 , n23888 );
nand ( n23890 , n23886 , n23889 , n2 );
and ( n23891 , n1352 , n22312 );
and ( n23892 , n21939 , n22315 );
nor ( n23893 , n588 , n22327 );
nor ( n23894 , n23892 , n23893 , n21565 );
nor ( n23895 , n23891 , n23894 );
or ( n23896 , n23895 , n22446 );
nand ( n23897 , n45 , n21598 );
nand ( n23898 , n23896 , n2 , n23897 );
or ( n23899 , n16041 , n23876 );
or ( n23900 , n148 , n23862 );
or ( n23901 , n589 , n23861 );
buf ( n23902 , n23853 );
nand ( n23903 , n23900 , n23901 , n23902 );
nand ( n23904 , n23899 , n2 , n23903 );
and ( n23905 , n590 , n23862 );
and ( n23906 , n152 , n23861 );
nor ( n23907 , n23905 , n23906 );
or ( n23908 , n23907 , n23885 );
not ( n23909 , n23887 );
or ( n23910 , n15901 , n23909 );
nand ( n23911 , n23908 , n23910 , n2 );
and ( n23912 , n591 , n23862 );
and ( n23913 , n175 , n23861 );
nor ( n23914 , n23912 , n23913 );
or ( n23915 , n23914 , n23885 );
or ( n23916 , n16085 , n23909 );
nand ( n23917 , n23915 , n23916 , n2 );
and ( n23918 , n592 , n23862 );
and ( n23919 , n157 , n23861 );
nor ( n23920 , n23918 , n23919 );
or ( n23921 , n23920 , n23885 );
not ( n23922 , n23887 );
or ( n23923 , n16061 , n23922 );
nand ( n23924 , n23921 , n23923 , n2 );
and ( n23925 , n593 , n23862 );
and ( n23926 , n159 , n23861 );
nor ( n23927 , n23925 , n23926 );
or ( n23928 , n23927 , n23885 );
not ( n23929 , n23887 );
or ( n23930 , n16057 , n23929 );
nand ( n23931 , n23928 , n23930 , n2 );
and ( n23932 , n617 , n22165 );
and ( n23933 , n143 , n22164 );
nor ( n23934 , n23932 , n23933 );
or ( n23935 , n23934 , n22157 );
or ( n23936 , n16081 , n22540 );
nand ( n23937 , n23935 , n23936 , n2 );
and ( n23938 , n623 , n22165 );
and ( n23939 , n415 , n22164 );
nor ( n23940 , n23938 , n23939 );
or ( n23941 , n23940 , n22157 );
or ( n23942 , n16001 , n22533 );
nand ( n23943 , n23941 , n23942 , n2 );
and ( n23944 , n624 , n22165 );
and ( n23945 , n1610 , n22164 );
nor ( n23946 , n23944 , n23945 );
or ( n23947 , n23946 , n22157 );
or ( n23948 , n15997 , n22192 );
nand ( n23949 , n23947 , n23948 , n2 );
and ( n23950 , n628 , n22165 );
and ( n23951 , n185 , n22164 );
nor ( n23952 , n23950 , n23951 );
or ( n23953 , n23952 , n23663 );
or ( n23954 , n16073 , n22192 );
nand ( n23955 , n23953 , n23954 , n2 );
and ( n23956 , n630 , n22165 );
and ( n23957 , n323 , n22164 );
nor ( n23958 , n23956 , n23957 );
or ( n23959 , n23958 , n22157 );
or ( n23960 , n15973 , n22185 );
nand ( n23961 , n23959 , n23960 , n2 );
and ( n23962 , n631 , n22165 );
and ( n23963 , n178 , n22164 );
nor ( n23964 , n23962 , n23963 );
or ( n23965 , n23964 , n23663 );
or ( n23966 , n16069 , n22185 );
nand ( n23967 , n23965 , n23966 , n2 );
not ( n23968 , n23854 );
or ( n23969 , n16065 , n23968 );
or ( n23970 , n1801 , n23862 );
or ( n23971 , n633 , n23861 );
nand ( n23972 , n23970 , n23971 , n23865 );
nand ( n23973 , n23969 , n2 , n23972 );
or ( n23974 , n15965 , n23855 );
or ( n23975 , n1795 , n23862 );
or ( n23976 , n634 , n23861 );
nand ( n23977 , n23975 , n23976 , n23865 );
nand ( n23978 , n23974 , n2 , n23977 );
not ( n23979 , n21858 );
and ( n23980 , n143 , n21860 );
and ( n23981 , n645 , n21817 );
nor ( n23982 , n23980 , n23981 );
not ( n23983 , n23982 );
and ( n23984 , n23979 , n23983 );
and ( n23985 , n1297 , n21866 );
nor ( n23986 , n23984 , n23985 );
or ( n23987 , n23986 , n21830 );
nand ( n23988 , n40 , n21830 );
nand ( n23989 , n23987 , n2 , n23988 );
and ( n23990 , n1299 , n21814 );
and ( n23991 , n22225 , n22409 );
nor ( n23992 , n646 , n21877 );
nor ( n23993 , n23991 , n23992 , n21980 );
nor ( n23994 , n23990 , n23993 );
or ( n23995 , n23994 , n21830 );
nand ( n23996 , n36 , n21830 );
nand ( n23997 , n23995 , n2 , n23996 );
and ( n23998 , n1336 , n21566 );
not ( n23999 , n21570 );
and ( n24000 , n21949 , n23999 );
nor ( n24001 , n649 , n21573 );
nor ( n24002 , n24000 , n24001 , n21565 );
nor ( n24003 , n23998 , n24002 );
or ( n24004 , n24003 , n22446 );
nand ( n24005 , n52 , n21598 );
nand ( n24006 , n24004 , n2 , n24005 );
and ( n24007 , n1306 , n21866 );
and ( n24008 , n22705 , n22409 );
nor ( n24009 , n648 , n21920 );
nor ( n24010 , n24008 , n24009 , n22348 );
nor ( n24011 , n24007 , n24010 );
or ( n24012 , n24011 , n21830 );
nand ( n24013 , n24012 , n2 , n23149 );
and ( n24014 , n1193 , n22312 );
and ( n24015 , n21977 , n23999 );
nor ( n24016 , n658 , n21573 );
nor ( n24017 , n24015 , n24016 , n21565 );
nor ( n24018 , n24014 , n24017 );
or ( n24019 , n24018 , n22446 );
nand ( n24020 , n51 , n21598 );
nand ( n24021 , n24019 , n2 , n24020 );
and ( n24022 , n1411 , n22312 );
and ( n24023 , n22042 , n23999 );
nor ( n24024 , n660 , n21573 );
nor ( n24025 , n24023 , n24024 , n21565 );
nor ( n24026 , n24022 , n24025 );
or ( n24027 , n24026 , n22446 );
nand ( n24028 , n49 , n21598 );
nand ( n24029 , n24027 , n2 , n24028 );
or ( n24030 , n16025 , n23968 );
or ( n24031 , n147 , n23862 );
or ( n24032 , n661 , n23861 );
nand ( n24033 , n24031 , n24032 , n23902 );
nand ( n24034 , n24030 , n2 , n24033 );
and ( n24035 , n666 , n23862 );
and ( n24036 , n178 , n23861 );
nor ( n24037 , n24035 , n24036 );
or ( n24038 , n24037 , n23885 );
or ( n24039 , n16069 , n23909 );
nand ( n24040 , n24038 , n24039 , n2 );
and ( n24041 , n667 , n23862 );
and ( n24042 , n428 , n23861 );
nor ( n24043 , n24041 , n24042 );
or ( n24044 , n24043 , n23885 );
or ( n24045 , n16005 , n23929 );
nand ( n24046 , n24044 , n24045 , n2 );
or ( n24047 , n15977 , n23855 );
or ( n24048 , n253 , n23862 );
or ( n24049 , n668 , n23861 );
nand ( n24050 , n24048 , n24049 , n23902 );
nand ( n24051 , n24047 , n2 , n24050 );
and ( n24052 , n669 , n23862 );
and ( n24053 , n352 , n23861 );
nor ( n24054 , n24052 , n24053 );
or ( n24055 , n24054 , n23885 );
or ( n24056 , n15989 , n23929 );
nand ( n24057 , n24055 , n24056 , n2 );
and ( n24058 , n672 , n23862 );
and ( n24059 , n1082 , n23861 );
nor ( n24060 , n24058 , n24059 );
or ( n24061 , n24060 , n23885 );
or ( n24062 , n16017 , n23929 );
nand ( n24063 , n24061 , n24062 , n2 );
not ( n24064 , n22751 );
and ( n24065 , n415 , n22742 );
and ( n24066 , n675 , n22739 );
nor ( n24067 , n24065 , n24066 );
not ( n24068 , n24067 );
and ( n24069 , n24064 , n24068 );
and ( n24070 , n1283 , n22752 );
nor ( n24071 , n24069 , n24070 );
or ( n24072 , n24071 , n22835 );
nand ( n24073 , n24072 , n2 , n23106 );
and ( n24074 , n699 , n23862 );
and ( n24075 , n193 , n23861 );
nor ( n24076 , n24074 , n24075 );
or ( n24077 , n24076 , n23885 );
or ( n24078 , n16089 , n23888 );
nand ( n24079 , n24077 , n24078 , n2 );
not ( n24080 , n23854 );
or ( n24081 , n16081 , n24080 );
or ( n24082 , n143 , n23862 );
or ( n24083 , n700 , n23861 );
nand ( n24084 , n24082 , n24083 , n23865 );
nand ( n24085 , n24081 , n2 , n24084 );
and ( n24086 , n701 , n23862 );
and ( n24087 , n144 , n23861 );
nor ( n24088 , n24086 , n24087 );
or ( n24089 , n24088 , n23885 );
or ( n24090 , n16021 , n23888 );
nand ( n24091 , n24089 , n24090 , n2 );
or ( n24092 , n16013 , n24080 );
or ( n24093 , n439 , n23862 );
or ( n24094 , n702 , n23861 );
nand ( n24095 , n24093 , n24094 , n23865 );
nand ( n24096 , n24092 , n2 , n24095 );
and ( n24097 , n703 , n23862 );
and ( n24098 , n461 , n23861 );
nor ( n24099 , n24097 , n24098 );
or ( n24100 , n24099 , n23885 );
not ( n24101 , n23854 );
or ( n24102 , n16009 , n24101 );
nand ( n24103 , n24100 , n24102 , n2 );
or ( n24104 , n16077 , n23855 );
or ( n24105 , n186 , n23862 );
or ( n24106 , n704 , n23861 );
nand ( n24107 , n24105 , n24106 , n23902 );
nand ( n24108 , n24104 , n2 , n24107 );
or ( n24109 , n15997 , n24080 );
or ( n24110 , n1610 , n23862 );
or ( n24111 , n705 , n23861 );
nand ( n24112 , n24110 , n24111 , n23865 );
nand ( n24113 , n24109 , n2 , n24112 );
and ( n24114 , n706 , n23862 );
and ( n24115 , n383 , n23861 );
nor ( n24116 , n24114 , n24115 );
or ( n24117 , n24116 , n23885 );
or ( n24118 , n15993 , n23888 );
nand ( n24119 , n24117 , n24118 , n2 );
or ( n24120 , n16001 , n24080 );
or ( n24121 , n415 , n23862 );
or ( n24122 , n707 , n23861 );
nand ( n24123 , n24121 , n24122 , n23865 );
nand ( n24124 , n24120 , n2 , n24123 );
or ( n24125 , n15981 , n23968 );
or ( n24126 , n284 , n23862 );
or ( n24127 , n708 , n23861 );
nand ( n24128 , n24126 , n24127 , n23865 );
nand ( n24129 , n24125 , n2 , n24128 );
or ( n24130 , n15985 , n23968 );
or ( n24131 , n283 , n23862 );
or ( n24132 , n709 , n23861 );
nand ( n24133 , n24131 , n24132 , n23902 );
nand ( n24134 , n24130 , n2 , n24133 );
and ( n24135 , n710 , n23862 );
and ( n24136 , n323 , n23861 );
nor ( n24137 , n24135 , n24136 );
or ( n24138 , n24137 , n23885 );
or ( n24139 , n15973 , n23909 );
nand ( n24140 , n24138 , n24139 , n2 );
or ( n24141 , n16073 , n23855 );
or ( n24142 , n185 , n23862 );
or ( n24143 , n711 , n23861 );
nand ( n24144 , n24142 , n24143 , n23865 );
nand ( n24145 , n24141 , n2 , n24144 );
or ( n24146 , n15969 , n23876 );
or ( n24147 , n192 , n23862 );
or ( n24148 , n712 , n23861 );
nand ( n24149 , n24147 , n24148 , n23865 );
nand ( n24150 , n24146 , n2 , n24149 );
and ( n24151 , n713 , n23862 );
and ( n24152 , n156 , n23861 );
nor ( n24153 , n24151 , n24152 );
or ( n24154 , n24153 , n23885 );
or ( n24155 , n16053 , n23922 );
nand ( n24156 , n24154 , n24155 , n2 );
or ( n24157 , n16049 , n23876 );
or ( n24158 , n151 , n23862 );
or ( n24159 , n714 , n23861 );
nand ( n24160 , n24158 , n24159 , n23902 );
nand ( n24161 , n24157 , n2 , n24160 );
and ( n24162 , n1421 , n22611 );
and ( n24163 , n21977 , n22799 );
nor ( n24164 , n728 , n22617 );
nor ( n24165 , n24163 , n24164 , n22784 );
nor ( n24166 , n24162 , n24165 );
or ( n24167 , n24166 , n22835 );
nand ( n24168 , n51 , n22627 );
nand ( n24169 , n24167 , n2 , n24168 );
and ( n24170 , n1287 , n22611 );
and ( n24171 , n22024 , n22917 );
nor ( n24172 , n735 , n22742 );
nor ( n24173 , n24171 , n24172 , n22619 );
nor ( n24174 , n24170 , n24173 );
or ( n24175 , n24174 , n22835 );
nand ( n24176 , n24175 , n2 , n23113 );
and ( n24177 , n1473 , n22611 );
and ( n24178 , n22345 , n22615 );
nor ( n24179 , n736 , n22617 );
nor ( n24180 , n24178 , n24179 , n22756 );
nor ( n24181 , n24177 , n24180 );
or ( n24182 , n24181 , n22835 );
nand ( n24183 , n50 , n22627 );
nand ( n24184 , n24182 , n2 , n24183 );
not ( n24185 , n2 );
not ( n24186 , n23188 );
and ( n24187 , n25 , n24186 );
and ( n24188 , n1261 , n23188 );
nor ( n24189 , n24187 , n24188 );
nor ( n24190 , n24185 , n24189 );
and ( n24191 , n1392 , n22611 );
and ( n24192 , n22042 , n22615 );
nor ( n24193 , n738 , n22742 );
nor ( n24194 , n24192 , n24193 , n22784 );
nor ( n24195 , n24191 , n24194 );
or ( n24196 , n24195 , n22835 );
nand ( n24197 , n24196 , n2 , n23581 );
and ( n24198 , n1312 , n22752 );
and ( n24199 , n21848 , n22810 );
nor ( n24200 , n740 , n22742 );
nor ( n24201 , n24199 , n24200 , n22756 );
nor ( n24202 , n24198 , n24201 );
or ( n24203 , n24202 , n22835 );
nand ( n24204 , n43 , n22627 );
nand ( n24205 , n24203 , n2 , n24204 );
and ( n24206 , n1194 , n22059 );
and ( n24207 , n21949 , n22061 );
nor ( n24208 , n741 , n22061 );
nor ( n24209 , n24207 , n24208 , n22059 );
nor ( n24210 , n24206 , n24209 );
or ( n24211 , n24210 , n22071 );
nand ( n24212 , n52 , n22105 );
nand ( n24213 , n24211 , n2 , n24212 );
not ( n24214 , n2 );
and ( n24215 , n45 , n23565 );
and ( n24216 , n1259 , n23188 );
nor ( n24217 , n24215 , n24216 );
nor ( n24218 , n24214 , n24217 );
and ( n24219 , n1349 , n21566 );
and ( n24220 , n22345 , n23999 );
nor ( n24221 , n755 , n21573 );
nor ( n24222 , n24220 , n24221 , n21565 );
nor ( n24223 , n24219 , n24222 );
or ( n24224 , n24223 , n22446 );
nand ( n24225 , n50 , n21598 );
nand ( n24226 , n24224 , n2 , n24225 );
not ( n24227 , n21565 );
and ( n24228 , n284 , n22327 );
and ( n24229 , n758 , n22314 );
nor ( n24230 , n24228 , n24229 );
not ( n24231 , n24230 );
and ( n24232 , n24227 , n24231 );
and ( n24233 , n1348 , n22312 );
nor ( n24234 , n24232 , n24233 );
or ( n24235 , n24234 , n22446 );
nand ( n24236 , n24235 , n2 , n23201 );
not ( n24237 , n2 );
nand ( n24238 , n789 , n15377 );
nand ( n24239 , n1230 , n15377 );
and ( n24240 , n24238 , n24239 );
nor ( n24241 , n24240 , n20168 );
or ( n24242 , n1538 , n24238 , n20175 );
not ( n24243 , n789 );
or ( n24244 , n24243 , n23642 );
nand ( n24245 , n24242 , n24244 );
nor ( n24246 , n24241 , n24245 );
nor ( n24247 , n24237 , n24246 );
not ( n24248 , n2 );
and ( n24249 , n48 , n24186 );
and ( n24250 , n1258 , n23188 );
nor ( n24251 , n24249 , n24250 );
nor ( n24252 , n24248 , n24251 );
not ( n24253 , n2 );
and ( n24254 , n41 , n23547 );
and ( n24255 , n1257 , n23188 );
nor ( n24256 , n24254 , n24255 );
nor ( n24257 , n24253 , n24256 );
not ( n24258 , n15649 );
nand ( n24259 , n889 , n24258 );
nor ( n24260 , n19377 , n24259 );
or ( n24261 , n1799 , n24260 );
nand ( n24262 , n24261 , n20052 );
and ( n24263 , n20057 , n21535 );
nor ( n24264 , n24263 , n24259 );
or ( n24265 , n1799 , n24264 );
or ( n24266 , n24259 , n21535 );
nand ( n24267 , n24266 , n20050 );
nand ( n24268 , n24265 , n24267 );
and ( n24269 , n24262 , n24268 );
nor ( n24270 , n24269 , n21342 );
not ( n24271 , n15649 );
and ( n24272 , n902 , n24271 );
nand ( n24273 , n20043 , n20056 , n24272 , n20058 );
or ( n24274 , n407 , n902 );
not ( n24275 , n15607 );
nand ( n24276 , n1113 , n15601 );
nor ( n24277 , n24275 , n24276 , n1174 , n15587 );
nand ( n24278 , n24274 , n24277 );
not ( n24279 , n24271 );
or ( n24280 , n19376 , n24279 );
not ( n24281 , n24272 );
nand ( n24282 , n24280 , n24281 );
nand ( n24283 , n24282 , n20043 , n20052 );
and ( n24284 , n24273 , n24278 , n24283 );
nor ( n24285 , n24284 , n21342 );
not ( n24286 , n13641 );
nand ( n24287 , n947 , n19984 );
or ( n24288 , n947 , n13643 );
nand ( n24289 , n24288 , n1000 );
nand ( n24290 , n24286 , n24287 , n24289 );
and ( n24291 , n948 , n13660 );
and ( n24292 , n950 , n13664 );
nor ( n24293 , n24291 , n24292 );
nand ( n24294 , n948 , n950 );
nand ( n24295 , n24293 , n24294 , n13668 );
and ( n24296 , n951 , n13675 );
and ( n24297 , n899 , n18835 );
nor ( n24298 , n24296 , n24297 );
nand ( n24299 , n899 , n951 );
nand ( n24300 , n24298 , n24299 , n13683 );
nand ( n24301 , n24290 , n24295 , n24300 );
and ( n24302 , n899 , n18833 );
and ( n24303 , n951 , n18835 );
nor ( n24304 , n24302 , n24303 );
or ( n24305 , n933 , n24294 );
and ( n24306 , n948 , n20791 );
and ( n24307 , n950 , n13660 );
nor ( n24308 , n24306 , n24307 );
nand ( n24309 , n24305 , n24308 );
and ( n24310 , n24300 , n24309 );
not ( n24311 , n24299 );
and ( n24312 , n13675 , n24311 );
nor ( n24313 , n24310 , n24312 );
and ( n24314 , n24301 , n24304 , n24313 );
and ( n24315 , n952 , n13633 );
and ( n24316 , n953 , n13623 );
nor ( n24317 , n24315 , n24316 );
nand ( n24318 , n952 , n953 );
and ( n24319 , n24317 , n24318 , n13690 );
nor ( n24320 , n24314 , n24319 );
not ( n24321 , n955 );
nand ( n24322 , n24321 , n1006 );
not ( n24323 , n13265 );
not ( n24324 , n888 );
and ( n24325 , n24323 , n24324 );
not ( n24326 , n954 );
nor ( n24327 , n24326 , n939 );
nor ( n24328 , n24325 , n24327 );
nand ( n24329 , n901 , n954 );
nand ( n24330 , n24328 , n24329 , n18807 );
and ( n24331 , n24320 , n24322 , n24330 );
nor ( n24332 , n897 , n956 );
or ( n24333 , n939 , n24329 );
and ( n24334 , n901 , n13620 );
and ( n24335 , n954 , n18815 );
nor ( n24336 , n24334 , n24335 );
not ( n24337 , n952 );
or ( n24338 , n24337 , n13690 );
or ( n24339 , n937 , n24318 );
or ( n24340 , n13296 , n938 );
nand ( n24341 , n24338 , n24339 , n24340 );
nand ( n24342 , n24330 , n24341 );
nand ( n24343 , n24333 , n24336 , n24342 );
and ( n24344 , n24322 , n24343 );
and ( n24345 , n955 , n12538 );
nor ( n24346 , n24344 , n24345 , n891 );
nand ( n24347 , n24332 , n24346 );
nor ( n24348 , n24331 , n24347 );
not ( n24349 , n2 );
not ( n24350 , n23156 );
and ( n24351 , n34 , n24350 );
and ( n24352 , n1155 , n23156 );
nor ( n24353 , n24351 , n24352 );
nor ( n24354 , n24349 , n24353 );
not ( n24355 , n2 );
and ( n24356 , n52 , n24186 );
and ( n24357 , n1255 , n23188 );
nor ( n24358 , n24356 , n24357 );
nor ( n24359 , n24355 , n24358 );
not ( n24360 , n2 );
and ( n24361 , n27 , n23559 );
and ( n24362 , n1159 , n23188 );
nor ( n24363 , n24361 , n24362 );
nor ( n24364 , n24360 , n24363 );
nor ( n24365 , n1639 , n20570 , n13217 );
and ( n24366 , n1576 , n24365 );
nor ( n24367 , n24366 , n1020 );
nor ( n24368 , n20577 , n24367 );
and ( n24369 , n1609 , n24365 );
nor ( n24370 , n24369 , n1021 );
nor ( n24371 , n20582 , n24370 );
and ( n24372 , n1588 , n24365 );
nor ( n24373 , n24372 , n1032 );
nor ( n24374 , n20587 , n24373 );
and ( n24375 , n1559 , n24365 );
nor ( n24376 , n24375 , n1033 );
nor ( n24377 , n20569 , n24376 );
not ( n24378 , n2 );
not ( n24379 , n23156 );
and ( n24380 , n28 , n24379 );
and ( n24381 , n1253 , n23156 );
nor ( n24382 , n24380 , n24381 );
nor ( n24383 , n24378 , n24382 );
nor ( n24384 , n20057 , n15606 );
nand ( n24385 , n24384 , n1100 , n21349 , n15650 );
not ( n24386 , n1100 );
not ( n24387 , n15616 );
or ( n24388 , n24386 , n24387 );
nand ( n24389 , n24388 , n15617 );
not ( n24390 , n19381 );
nand ( n24391 , n24389 , n15622 , n24390 );
and ( n24392 , n1100 , n15668 );
nor ( n24393 , n24392 , n19379 );
not ( n24394 , n24393 );
nand ( n24395 , n24394 , n15676 );
and ( n24396 , n24385 , n24391 , n24395 );
nor ( n24397 , n24396 , n21342 );
nand ( n24398 , n928 , n21428 );
not ( n24399 , n24398 );
and ( n24400 , n21434 , n21679 , n24399 );
or ( n24401 , n929 , n21429 );
nand ( n24402 , n24401 , n928 );
and ( n24403 , n931 , n24402 );
nor ( n24404 , n24400 , n24403 );
not ( n24405 , n13556 );
nand ( n24406 , n21423 , n21434 , n21433 );
nand ( n24407 , n24405 , n24406 );
not ( n24408 , n24406 );
nand ( n24409 , n21432 , n24408 );
nand ( n24410 , n24407 , n24409 );
or ( n24411 , n24404 , n900 , n24410 );
not ( n24412 , n17118 );
not ( n24413 , n17122 );
or ( n24414 , n24412 , n24413 , n24409 );
nand ( n24415 , n24411 , n24414 );
not ( n24416 , n24415 );
or ( n24417 , n21675 , n928 , n930 );
and ( n24418 , n21434 , n16462 );
nor ( n24419 , n932 , n929 , n24398 );
nor ( n24420 , n24418 , n24419 );
or ( n24421 , n930 , n24420 );
nand ( n24422 , n24417 , n24421 );
not ( n24423 , n24410 );
and ( n24424 , n24422 , n24423 );
and ( n24425 , n21419 , n21669 );
nor ( n24426 , n24425 , n1623 , n24407 );
nor ( n24427 , n24424 , n24426 );
nand ( n24428 , n24416 , n24427 );
not ( n24429 , n2 );
and ( n24430 , n37 , n24350 );
and ( n24431 , n1251 , n23156 );
nor ( n24432 , n24430 , n24431 );
nor ( n24433 , n24429 , n24432 );
not ( n24434 , n940 );
not ( n24435 , n20613 );
not ( n24436 , n24435 );
or ( n24437 , n24434 , n24436 );
buf ( n24438 , n20613 );
nand ( n24439 , n964 , n24438 );
nand ( n24440 , n24437 , n24439 );
not ( n24441 , n949 );
not ( n24442 , n24435 );
or ( n24443 , n24441 , n24442 );
nand ( n24444 , n972 , n24438 );
nand ( n24445 , n24443 , n24444 );
not ( n24446 , n957 );
not ( n24447 , n24435 );
or ( n24448 , n24446 , n24447 );
nand ( n24449 , n980 , n24438 );
nand ( n24450 , n24448 , n24449 );
not ( n24451 , n966 );
not ( n24452 , n24438 );
or ( n24453 , n24451 , n24452 );
or ( n24454 , n13458 , n21778 );
nand ( n24455 , n24453 , n24454 );
not ( n24456 , n944 );
not ( n24457 , n24435 );
or ( n24458 , n24456 , n24457 );
nand ( n24459 , n967 , n24438 );
nand ( n24460 , n24458 , n24459 );
not ( n24461 , n999 );
not ( n24462 , n24435 );
or ( n24463 , n24461 , n24462 );
nand ( n24464 , n881 , n24438 );
nand ( n24465 , n24463 , n24464 );
not ( n24466 , n968 );
not ( n24467 , n24438 );
or ( n24468 , n24466 , n24467 );
not ( n24469 , n20618 );
or ( n24470 , n13441 , n24469 );
nand ( n24471 , n24468 , n24470 );
not ( n24472 , n969 );
not ( n24473 , n24438 );
or ( n24474 , n24472 , n24473 );
or ( n24475 , n12762 , n24469 );
nand ( n24476 , n24474 , n24475 );
not ( n24477 , n885 );
not ( n24478 , n24435 );
or ( n24479 , n24477 , n24478 );
nand ( n24480 , n1009 , n24438 );
nand ( n24481 , n24479 , n24480 );
not ( n24482 , n959 );
not ( n24483 , n24435 );
or ( n24484 , n24482 , n24483 );
nand ( n24485 , n983 , n24438 );
nand ( n24486 , n24484 , n24485 );
not ( n24487 , n984 );
not ( n24488 , n24438 );
or ( n24489 , n24487 , n24488 );
or ( n24490 , n14624 , n24469 );
nand ( n24491 , n24489 , n24490 );
not ( n24492 , n985 );
not ( n24493 , n24438 );
or ( n24494 , n24492 , n24493 );
or ( n24495 , n14392 , n24469 );
nand ( n24496 , n24494 , n24495 );
not ( n24497 , n1008 );
not ( n24498 , n24438 );
or ( n24499 , n24497 , n24498 );
or ( n24500 , n14403 , n21778 );
nand ( n24501 , n24499 , n24500 );
not ( n24502 , n2 );
not ( n24503 , n23156 );
and ( n24504 , n46 , n24503 );
and ( n24505 , n1250 , n23156 );
nor ( n24506 , n24504 , n24505 );
nor ( n24507 , n24502 , n24506 );
not ( n24508 , n986 );
not ( n24509 , n24438 );
or ( n24510 , n24508 , n24509 );
or ( n24511 , n14001 , n21778 );
nand ( n24512 , n24510 , n24511 );
not ( n24513 , n987 );
not ( n24514 , n24438 );
or ( n24515 , n24513 , n24514 );
or ( n24516 , n13976 , n21778 );
nand ( n24517 , n24515 , n24516 );
not ( n24518 , n887 );
not ( n24519 , n24438 );
or ( n24520 , n24518 , n24519 );
or ( n24521 , n13920 , n21778 );
nand ( n24522 , n24520 , n24521 );
not ( n24523 , n965 );
not ( n24524 , n24438 );
or ( n24525 , n24523 , n24524 );
or ( n24526 , n13934 , n21778 );
nand ( n24527 , n24525 , n24526 );
not ( n24528 , n2 );
not ( n24529 , n23156 );
and ( n24530 , n40 , n24529 );
and ( n24531 , n1249 , n23156 );
nor ( n24532 , n24530 , n24531 );
nor ( n24533 , n24528 , n24532 );
not ( n24534 , n1146 );
not ( n24535 , n17140 );
nand ( n24536 , n24535 , n17742 );
not ( n24537 , n24536 );
or ( n24538 , n24534 , n24537 );
or ( n24539 , n18385 , n24536 );
nand ( n24540 , n24538 , n24539 );
not ( n24541 , n2 );
not ( n24542 , n23156 );
and ( n24543 , n50 , n24542 );
and ( n24544 , n1151 , n23156 );
nor ( n24545 , n24543 , n24544 );
nor ( n24546 , n24541 , n24545 );
not ( n24547 , n2 );
and ( n24548 , n48 , n24542 );
and ( n24549 , n1152 , n23156 );
nor ( n24550 , n24548 , n24549 );
nor ( n24551 , n24547 , n24550 );
not ( n24552 , n2 );
not ( n24553 , n23156 );
and ( n24554 , n36 , n24553 );
and ( n24555 , n1153 , n23156 );
nor ( n24556 , n24554 , n24555 );
nor ( n24557 , n24552 , n24556 );
not ( n24558 , n2 );
and ( n24559 , n35 , n24350 );
and ( n24560 , n1154 , n23156 );
nor ( n24561 , n24559 , n24560 );
nor ( n24562 , n24558 , n24561 );
not ( n24563 , n2 );
and ( n24564 , n50 , n23189 );
and ( n24565 , n1156 , n23188 );
nor ( n24566 , n24564 , n24565 );
nor ( n24567 , n24563 , n24566 );
not ( n24568 , n2 );
and ( n24569 , n47 , n23559 );
and ( n24570 , n1157 , n23188 );
nor ( n24571 , n24569 , n24570 );
nor ( n24572 , n24568 , n24571 );
not ( n24573 , n2 );
and ( n24574 , n43 , n23565 );
and ( n24575 , n1158 , n23188 );
nor ( n24576 , n24574 , n24575 );
nor ( n24577 , n24573 , n24576 );
not ( n24578 , n2 );
and ( n24579 , n52 , n23590 );
and ( n24580 , n1160 , n23204 );
nor ( n24581 , n24579 , n24580 );
nor ( n24582 , n24578 , n24581 );
not ( n24583 , n2 );
not ( n24584 , n23204 );
and ( n24585 , n50 , n24584 );
and ( n24586 , n1161 , n23204 );
nor ( n24587 , n24585 , n24586 );
nor ( n24588 , n24583 , n24587 );
not ( n24589 , n2 );
and ( n24590 , n46 , n23590 );
and ( n24591 , n1162 , n23204 );
nor ( n24592 , n24590 , n24591 );
nor ( n24593 , n24589 , n24592 );
not ( n24594 , n1168 );
not ( n24595 , n24536 );
or ( n24596 , n24594 , n24595 );
or ( n24597 , n17967 , n24536 );
nand ( n24598 , n24596 , n24597 );
not ( n24599 , n1169 );
not ( n24600 , n24536 );
or ( n24601 , n24599 , n24600 );
or ( n24602 , n17985 , n24536 );
nand ( n24603 , n24601 , n24602 );
not ( n24604 , n1170 );
not ( n24605 , n24536 );
or ( n24606 , n24604 , n24605 );
or ( n24607 , n18483 , n24536 );
nand ( n24608 , n24606 , n24607 );
not ( n24609 , n1171 );
not ( n24610 , n24536 );
or ( n24611 , n24609 , n24610 );
or ( n24612 , n18380 , n24536 );
nand ( n24613 , n24611 , n24612 );
not ( n24614 , n1172 );
not ( n24615 , n24536 );
or ( n24616 , n24614 , n24615 );
or ( n24617 , n18473 , n24536 );
nand ( n24618 , n24616 , n24617 );
not ( n24619 , n1173 );
not ( n24620 , n24536 );
or ( n24621 , n24619 , n24620 );
or ( n24622 , n18754 , n24536 );
nand ( n24623 , n24621 , n24622 );
not ( n24624 , n1178 );
not ( n24625 , n24536 );
or ( n24626 , n24624 , n24625 );
or ( n24627 , n17954 , n24536 );
nand ( n24628 , n24626 , n24627 );
not ( n24629 , n2 );
and ( n24630 , n35 , n23129 );
and ( n24631 , n1180 , n23128 );
nor ( n24632 , n24630 , n24631 );
nor ( n24633 , n24629 , n24632 );
not ( n24634 , n2 );
not ( n24635 , n23128 );
and ( n24636 , n39 , n24635 );
and ( n24637 , n1181 , n23128 );
nor ( n24638 , n24636 , n24637 );
nor ( n24639 , n24634 , n24638 );
not ( n24640 , n2 );
and ( n24641 , n34 , n23553 );
and ( n24642 , n1183 , n23188 );
nor ( n24643 , n24641 , n24642 );
nor ( n24644 , n24640 , n24643 );
nand ( n24645 , n1184 , n23138 );
nand ( n24646 , n24645 , n2 , n22057 );
not ( n24647 , n22446 );
nand ( n24648 , n1191 , n24647 );
nand ( n24649 , n24648 , n2 , n22455 );
nand ( n24650 , n1192 , n23166 );
nand ( n24651 , n24650 , n2 , n22131 );
not ( n24652 , n21598 );
nand ( n24653 , n1193 , n24652 );
nand ( n24654 , n24653 , n2 , n24020 );
not ( n24655 , n22071 );
nand ( n24656 , n1194 , n24655 );
nand ( n24657 , n24656 , n2 , n24212 );
nand ( n24658 , n1196 , n23138 );
nand ( n24659 , n24658 , n2 , n22475 );
not ( n24660 , n2 );
and ( n24661 , n47 , n23529 );
and ( n24662 , n1197 , n23531 );
nor ( n24663 , n24661 , n24662 );
nor ( n24664 , n24660 , n24663 );
not ( n24665 , n2 );
not ( n24666 , n23128 );
and ( n24667 , n31 , n24666 );
and ( n24668 , n1199 , n23128 );
nor ( n24669 , n24667 , n24668 );
nor ( n24670 , n24665 , n24669 );
nand ( n24671 , n1200 , n24647 );
nand ( n24672 , n24671 , n2 , n22649 );
not ( n24673 , n21830 );
nand ( n24674 , n1202 , n24673 );
nand ( n24675 , n24674 , n2 , n21936 );
not ( n24676 , n2 );
and ( n24677 , n27 , n24635 );
and ( n24678 , n1203 , n23128 );
nor ( n24679 , n24677 , n24678 );
nor ( n24680 , n24676 , n24679 );
nand ( n24681 , n1204 , n22414 );
nand ( n24682 , n24681 , n2 , n21845 );
not ( n24683 , n2 );
and ( n24684 , n44 , n23553 );
and ( n24685 , n1205 , n23188 );
nor ( n24686 , n24684 , n24685 );
nor ( n24687 , n24683 , n24686 );
not ( n24688 , n2 );
and ( n24689 , n36 , n23571 );
and ( n24690 , n1207 , n23188 );
nor ( n24691 , n24689 , n24690 );
nor ( n24692 , n24688 , n24691 );
not ( n24693 , n2 );
not ( n24694 , n23128 );
and ( n24695 , n45 , n24694 );
and ( n24696 , n1210 , n23128 );
nor ( n24697 , n24695 , n24696 );
nor ( n24698 , n24693 , n24697 );
not ( n24699 , n2 );
and ( n24700 , n26 , n23571 );
and ( n24701 , n1209 , n23188 );
nor ( n24702 , n24700 , n24701 );
nor ( n24703 , n24699 , n24702 );
not ( n24704 , n2 );
and ( n24705 , n46 , n23565 );
and ( n24706 , n1212 , n23188 );
nor ( n24707 , n24705 , n24706 );
nor ( n24708 , n24704 , n24707 );
not ( n24709 , n2 );
and ( n24710 , n40 , n23571 );
and ( n24711 , n1213 , n23188 );
nor ( n24712 , n24710 , n24711 );
nor ( n24713 , n24709 , n24712 );
nand ( n24714 , n1215 , n24652 );
nand ( n24715 , n24714 , n2 , n22379 );
not ( n24716 , n2 );
and ( n24717 , n51 , n23547 );
and ( n24718 , n1221 , n23188 );
nor ( n24719 , n24717 , n24718 );
nor ( n24720 , n24716 , n24719 );
or ( n24721 , n16926 , n21830 );
nand ( n24722 , n24721 , n2 , n22021 );
not ( n24723 , n2 );
and ( n24724 , n52 , n23529 );
and ( n24725 , n1223 , n23531 );
nor ( n24726 , n24724 , n24725 );
nor ( n24727 , n24723 , n24726 );
not ( n24728 , n2 );
and ( n24729 , n51 , n23529 );
and ( n24730 , n1224 , n23531 );
nor ( n24731 , n24729 , n24730 );
nor ( n24732 , n24728 , n24731 );
not ( n24733 , n2 );
and ( n24734 , n48 , n23529 );
and ( n24735 , n1226 , n23531 );
nor ( n24736 , n24734 , n24735 );
nor ( n24737 , n24733 , n24736 );
not ( n24738 , n2 );
and ( n24739 , n46 , n23529 );
and ( n24740 , n1227 , n23531 );
nor ( n24741 , n24739 , n24740 );
nor ( n24742 , n24738 , n24741 );
not ( n24743 , n2 );
and ( n24744 , n39 , n23584 );
and ( n24745 , n1229 , n23204 );
nor ( n24746 , n24744 , n24745 );
nor ( n24747 , n24743 , n24746 );
not ( n24748 , n2 );
and ( n24749 , n42 , n24694 );
and ( n24750 , n1231 , n23128 );
nor ( n24751 , n24749 , n24750 );
nor ( n24752 , n24748 , n24751 );
not ( n24753 , n2 );
not ( n24754 , n23128 );
and ( n24755 , n51 , n24754 );
and ( n24756 , n1233 , n23128 );
nor ( n24757 , n24755 , n24756 );
nor ( n24758 , n24753 , n24757 );
not ( n24759 , n2 );
and ( n24760 , n50 , n24754 );
and ( n24761 , n1234 , n23128 );
nor ( n24762 , n24760 , n24761 );
nor ( n24763 , n24759 , n24762 );
not ( n24764 , n2 );
and ( n24765 , n48 , n24666 );
and ( n24766 , n1235 , n23128 );
nor ( n24767 , n24765 , n24766 );
nor ( n24768 , n24764 , n24767 );
not ( n24769 , n2 );
not ( n24770 , n23128 );
and ( n24771 , n46 , n24770 );
and ( n24772 , n1237 , n23128 );
nor ( n24773 , n24771 , n24772 );
nor ( n24774 , n24769 , n24773 );
not ( n24775 , n2 );
and ( n24776 , n44 , n24770 );
and ( n24777 , n1238 , n23128 );
nor ( n24778 , n24776 , n24777 );
nor ( n24779 , n24775 , n24778 );
not ( n24780 , n2 );
and ( n24781 , n43 , n23827 );
and ( n24782 , n1239 , n23128 );
nor ( n24783 , n24781 , n24782 );
nor ( n24784 , n24780 , n24783 );
not ( n24785 , n2 );
and ( n24786 , n26 , n23827 );
and ( n24787 , n1241 , n23128 );
nor ( n24788 , n24786 , n24787 );
nor ( n24789 , n24785 , n24788 );
not ( n24790 , n2 );
and ( n24791 , n25 , n24666 );
and ( n24792 , n1242 , n23128 );
nor ( n24793 , n24791 , n24792 );
nor ( n24794 , n24790 , n24793 );
not ( n24795 , n2 );
and ( n24796 , n36 , n24770 );
and ( n24797 , n1243 , n23128 );
nor ( n24798 , n24796 , n24797 );
nor ( n24799 , n24795 , n24798 );
not ( n24800 , n2 );
and ( n24801 , n33 , n24666 );
and ( n24802 , n1245 , n23128 );
nor ( n24803 , n24801 , n24802 );
nor ( n24804 , n24800 , n24803 );
not ( n24805 , n2 );
and ( n24806 , n32 , n24770 );
and ( n24807 , n1246 , n23128 );
nor ( n24808 , n24806 , n24807 );
nor ( n24809 , n24805 , n24808 );
not ( n24810 , n2 );
and ( n24811 , n28 , n24635 );
and ( n24812 , n1247 , n23128 );
nor ( n24813 , n24811 , n24812 );
nor ( n24814 , n24810 , n24813 );
not ( n24815 , n2 );
and ( n24816 , n34 , n23511 );
and ( n24817 , n1275 , n23204 );
nor ( n24818 , n24816 , n24817 );
nor ( n24819 , n24815 , n24818 );
not ( n24820 , n2 );
and ( n24821 , n32 , n23590 );
and ( n24822 , n1277 , n23204 );
nor ( n24823 , n24821 , n24822 );
nor ( n24824 , n24820 , n24823 );
not ( n24825 , n22627 );
nand ( n24826 , n1278 , n24825 );
nand ( n24827 , n24826 , n2 , n22886 );
nand ( n24828 , n1279 , n24825 );
nand ( n24829 , n24828 , n2 , n22942 );
nand ( n24830 , n1280 , n24825 );
nand ( n24831 , n24830 , n2 , n22807 );
nand ( n24832 , n1281 , n24825 );
nand ( n24833 , n24832 , n2 , n22836 );
not ( n24834 , n2 );
and ( n24835 , n36 , n23536 );
and ( n24836 , n1274 , n23204 );
nor ( n24837 , n24835 , n24836 );
nor ( n24838 , n24834 , n24837 );
not ( n24839 , n22835 );
nand ( n24840 , n1282 , n24839 );
nand ( n24841 , n24840 , n2 , n22894 );
or ( n24842 , n16853 , n22835 );
nand ( n24843 , n24842 , n2 , n22958 );
or ( n24844 , n16848 , n22835 );
nand ( n24845 , n24844 , n2 , n22628 );
or ( n24846 , n19031 , n22835 );
nand ( n24847 , n24846 , n2 , n22992 );
not ( n24848 , n22835 );
nand ( n24849 , n1290 , n24848 );
nand ( n24850 , n24849 , n2 , n23845 );
not ( n24851 , n22835 );
nand ( n24852 , n1291 , n24851 );
nand ( n24853 , n24852 , n2 , n22788 );
nand ( n24854 , n1292 , n24825 );
nand ( n24855 , n24854 , n2 , n23000 );
nand ( n24856 , n1295 , n22414 );
nand ( n24857 , n24856 , n2 , n21896 );
nand ( n24858 , n1296 , n23138 );
nand ( n24859 , n24858 , n2 , n21914 );
not ( n24860 , n21830 );
nand ( n24861 , n1297 , n24860 );
nand ( n24862 , n24861 , n2 , n23988 );
nand ( n24863 , n1299 , n23138 );
nand ( n24864 , n24863 , n2 , n23996 );
nand ( n24865 , n1300 , n24673 );
nand ( n24866 , n24865 , n2 , n21966 );
or ( n24867 , n16934 , n21830 );
nand ( n24868 , n24867 , n2 , n22002 );
nand ( n24869 , n1301 , n23138 );
nand ( n24870 , n24869 , n2 , n21984 );
not ( n24871 , n21830 );
nand ( n24872 , n1307 , n24871 );
nand ( n24873 , n24872 , n2 , n22352 );
nand ( n24874 , n1309 , n23138 );
nand ( n24875 , n24874 , n2 , n22048 );
nand ( n24876 , n1311 , n24871 );
nand ( n24877 , n24876 , n2 , n21856 );
nand ( n24878 , n1310 , n24860 );
nand ( n24879 , n24878 , n2 , n22417 );
nand ( n24880 , n1312 , n23579 );
nand ( n24881 , n24880 , n2 , n24204 );
nand ( n24882 , n1315 , n23166 );
nand ( n24883 , n24882 , n2 , n22140 );
not ( n24884 , n22071 );
nand ( n24885 , n1316 , n24884 );
nand ( n24886 , n24885 , n2 , n23008 );
nand ( n24887 , n1317 , n22239 );
nand ( n24888 , n24887 , n2 , n22114 );
nand ( n24889 , n1319 , n22239 );
nand ( n24890 , n24889 , n2 , n22232 );
nand ( n24891 , n1318 , n22239 );
nand ( n24892 , n24891 , n2 , n22148 );
not ( n24893 , n22071 );
nand ( n24894 , n1320 , n24893 );
nand ( n24895 , n24894 , n2 , n22242 );
nand ( n24896 , n1322 , n23166 );
nand ( n24897 , n24896 , n2 , n23804 );
nand ( n24898 , n1329 , n23166 );
nand ( n24899 , n24898 , n2 , n22728 );
nand ( n24900 , n1331 , n24655 );
nand ( n24901 , n24900 , n2 , n22310 );
nand ( n24902 , n1332 , n24893 );
nand ( n24903 , n24902 , n2 , n22863 );
nand ( n24904 , n1333 , n23166 );
nand ( n24905 , n24904 , n2 , n22768 );
nand ( n24906 , n1334 , n24884 );
nand ( n24907 , n24906 , n2 , n22177 );
nand ( n24908 , n1336 , n24652 );
nand ( n24909 , n24908 , n2 , n24005 );
not ( n24910 , n22446 );
nand ( n24911 , n1337 , n24910 );
nand ( n24912 , n24911 , n2 , n22438 );
nand ( n24913 , n1338 , n24652 );
nand ( n24914 , n24913 , n2 , n22463 );
nand ( n24915 , n1339 , n24910 );
nand ( n24916 , n24915 , n2 , n23874 );
not ( n24917 , n22446 );
nand ( n24918 , n1340 , n24917 );
nand ( n24919 , n24918 , n2 , n22657 );
not ( n24920 , n22446 );
nand ( n24921 , n1341 , n24920 );
nand ( n24922 , n24921 , n2 , n22666 );
or ( n24923 , n17081 , n22446 );
nand ( n24924 , n24923 , n2 , n21599 );
or ( n24925 , n17078 , n22446 );
nand ( n24926 , n24925 , n2 , n22674 );
or ( n24927 , n17075 , n22446 );
nand ( n24928 , n24927 , n2 , n23040 );
or ( n24929 , n17072 , n22446 );
nand ( n24930 , n24929 , n2 , n22683 );
or ( n24931 , n17053 , n22446 );
nand ( n24932 , n24931 , n2 , n22702 );
nand ( n24933 , n1349 , n24652 );
nand ( n24934 , n24933 , n2 , n24225 );
nand ( n24935 , n1350 , n24652 );
nand ( n24936 , n24935 , n2 , n22334 );
not ( n24937 , n22446 );
nand ( n24938 , n1351 , n24937 );
nand ( n24939 , n24938 , n2 , n23475 );
nand ( n24940 , n1352 , n24917 );
nand ( n24941 , n24940 , n2 , n23897 );
nand ( n24942 , n1353 , n24652 );
nand ( n24943 , n24942 , n2 , n23064 );
not ( n24944 , n2 );
and ( n24945 , n52 , n24379 );
and ( n24946 , n1364 , n23156 );
nor ( n24947 , n24945 , n24946 );
nor ( n24948 , n24944 , n24947 );
not ( n24949 , n2 );
and ( n24950 , n52 , n24694 );
and ( n24951 , n1366 , n23128 );
nor ( n24952 , n24950 , n24951 );
nor ( n24953 , n24949 , n24952 );
nand ( n24954 , n1367 , n22239 );
nand ( n24955 , n24954 , n2 , n22081 );
nand ( n24956 , n1368 , n22414 );
nand ( n24957 , n24956 , n2 , n21905 );
nand ( n24958 , n1369 , n23166 );
nand ( n24959 , n24958 , n2 , n23819 );
not ( n24960 , n2 );
and ( n24961 , n28 , n23205 );
and ( n24962 , n1371 , n23204 );
nor ( n24963 , n24961 , n24962 );
nor ( n24964 , n24960 , n24963 );
not ( n24965 , n22071 );
nand ( n24966 , n1373 , n24965 );
nand ( n24967 , n24966 , n2 , n22106 );
nand ( n24968 , n1374 , n23166 );
nand ( n24969 , n24968 , n2 , n22090 );
nand ( n24970 , n1375 , n23576 );
nand ( n24971 , n24970 , n2 , n21926 );
nand ( n24972 , n1376 , n23138 );
nand ( n24973 , n24972 , n2 , n22637 );
nand ( n24974 , n1377 , n24965 );
nand ( n24975 , n24974 , n2 , n23016 );
not ( n24976 , n2 );
and ( n24977 , n27 , n24379 );
and ( n24978 , n1381 , n23156 );
nor ( n24979 , n24977 , n24978 );
nor ( n24980 , n24976 , n24979 );
not ( n24981 , n2 );
and ( n24982 , n33 , n23536 );
and ( n24983 , n1382 , n23204 );
nor ( n24984 , n24982 , n24983 );
nor ( n24985 , n24981 , n24984 );
nand ( n24986 , n1383 , n22414 );
nand ( n24987 , n24986 , n2 , n21957 );
not ( n24988 , n2 );
and ( n24989 , n35 , n24584 );
and ( n24990 , n1384 , n23204 );
nor ( n24991 , n24989 , n24990 );
nor ( n24992 , n24988 , n24991 );
not ( n24993 , n2 );
and ( n24994 , n26 , n24553 );
and ( n24995 , n1385 , n23156 );
nor ( n24996 , n24994 , n24995 );
nor ( n24997 , n24993 , n24996 );
not ( n24998 , n2 );
and ( n24999 , n25 , n24542 );
and ( n25000 , n1386 , n23156 );
nor ( n25001 , n24999 , n25000 );
nor ( n25002 , n24998 , n25001 );
not ( n25003 , n2 );
and ( n25004 , n47 , n23517 );
and ( n25005 , n1387 , n23204 );
nor ( n25006 , n25004 , n25005 );
nor ( n25007 , n25003 , n25006 );
not ( n25008 , n2 );
and ( n25009 , n27 , n23536 );
and ( n25010 , n1390 , n23204 );
nor ( n25011 , n25009 , n25010 );
nor ( n25012 , n25008 , n25011 );
not ( n25013 , n2 );
and ( n25014 , n31 , n24529 );
and ( n25015 , n1391 , n23156 );
nor ( n25016 , n25014 , n25015 );
nor ( n25017 , n25013 , n25016 );
not ( n25018 , n2 );
and ( n25019 , n33 , n24503 );
and ( n25020 , n1389 , n23156 );
nor ( n25021 , n25019 , n25020 );
nor ( n25022 , n25018 , n25021 );
not ( n25023 , n2 );
and ( n25024 , n44 , n24584 );
and ( n25025 , n1394 , n23204 );
nor ( n25026 , n25024 , n25025 );
nor ( n25027 , n25023 , n25026 );
not ( n25028 , n2 );
and ( n25029 , n43 , n24542 );
and ( n25030 , n1396 , n23156 );
nor ( n25031 , n25029 , n25030 );
nor ( n25032 , n25028 , n25031 );
not ( n25033 , n2 );
and ( n25034 , n41 , n24503 );
and ( n25035 , n1397 , n23156 );
nor ( n25036 , n25034 , n25035 );
nor ( n25037 , n25033 , n25036 );
or ( n25038 , n16828 , n22835 );
nand ( n25039 , n25038 , n2 , n22749 );
not ( n25040 , n2 );
and ( n25041 , n51 , n23584 );
and ( n25042 , n1400 , n23204 );
nor ( n25043 , n25041 , n25042 );
nor ( n25044 , n25040 , n25043 );
not ( n25045 , n2 );
and ( n25046 , n47 , n24350 );
and ( n25047 , n1401 , n23156 );
nor ( n25048 , n25046 , n25047 );
nor ( n25049 , n25045 , n25048 );
not ( n25050 , n2 );
and ( n25051 , n44 , n24553 );
and ( n25052 , n1399 , n23156 );
nor ( n25053 , n25051 , n25052 );
nor ( n25054 , n25050 , n25053 );
not ( n25055 , n2 );
and ( n25056 , n45 , n24379 );
and ( n25057 , n1403 , n23156 );
nor ( n25058 , n25056 , n25057 );
nor ( n25059 , n25055 , n25058 );
not ( n25060 , n2 );
and ( n25061 , n41 , n23511 );
and ( n25062 , n1402 , n23204 );
nor ( n25063 , n25061 , n25062 );
nor ( n25064 , n25060 , n25063 );
not ( n25065 , n2 );
and ( n25066 , n49 , n23157 );
and ( n25067 , n1406 , n23156 );
nor ( n25068 , n25066 , n25067 );
nor ( n25069 , n25065 , n25068 );
not ( n25070 , n22446 );
nand ( n25071 , n1407 , n25070 );
nand ( n25072 , n25071 , n2 , n22429 );
nand ( n25073 , n1408 , n25070 );
nand ( n25074 , n25073 , n2 , n22361 );
not ( n25075 , n2 );
and ( n25076 , n51 , n24553 );
and ( n25077 , n1409 , n23156 );
nor ( n25078 , n25076 , n25077 );
nor ( n25079 , n25075 , n25078 );
nand ( n25080 , n1410 , n24652 );
nand ( n25081 , n25080 , n2 , n23032 );
nand ( n25082 , n1411 , n24920 );
nand ( n25083 , n25082 , n2 , n24028 );
or ( n25084 , n16864 , n22835 );
nand ( n25085 , n25084 , n2 , n22931 );
nand ( n25086 , n1413 , n24825 );
nand ( n25087 , n25086 , n2 , n22914 );
not ( n25088 , n22835 );
nand ( n25089 , n1421 , n25088 );
nand ( n25090 , n25089 , n2 , n24168 );
nand ( n25091 , n1434 , n24839 );
nand ( n25092 , n25091 , n2 , n22906 );
not ( n25093 , n22835 );
nand ( n25094 , n1440 , n25093 );
nand ( n25095 , n25094 , n2 , n22827 );
nand ( n25096 , n1441 , n24848 );
nand ( n25097 , n25096 , n2 , n22818 );
nand ( n25098 , n1445 , n25093 );
nand ( n25099 , n25098 , n2 , n22796 );
nand ( n25100 , n1461 , n24825 );
nand ( n25101 , n25100 , n2 , n22845 );
nand ( n25102 , n1462 , n24825 );
nand ( n25103 , n25102 , n2 , n22855 );
not ( n25104 , n2 );
and ( n25105 , n49 , n24635 );
and ( n25106 , n1467 , n23128 );
nor ( n25107 , n25105 , n25106 );
nor ( n25108 , n25104 , n25107 );
nand ( n25109 , n1472 , n24851 );
nand ( n25110 , n25109 , n2 , n22779 );
nand ( n25111 , n1473 , n25088 );
nand ( n25112 , n25111 , n2 , n24183 );
not ( n25113 , n2 );
and ( n25114 , n49 , n24584 );
and ( n25115 , n1471 , n23204 );
nor ( n25116 , n25114 , n25115 );
nor ( n25117 , n25113 , n25116 );
nand ( n25118 , n2 , n30 );
or ( n25119 , n25118 , n23130 );
not ( n25120 , n23132 );
or ( n25121 , n1490 , n25120 );
nand ( n25122 , n25121 , n23135 );
nand ( n25123 , n25119 , n25122 );
or ( n25124 , n25118 , n23158 );
not ( n25125 , n23160 );
or ( n25126 , n1489 , n25125 );
nand ( n25127 , n25126 , n23163 );
nand ( n25128 , n25124 , n25127 );
or ( n25129 , n25118 , n23190 );
not ( n25130 , n23192 );
or ( n25131 , n1498 , n25130 );
nand ( n25132 , n25131 , n23195 );
nand ( n25133 , n25129 , n25132 );
or ( n25134 , n25118 , n23206 );
not ( n25135 , n23208 );
or ( n25136 , n1542 , n25135 );
nand ( n25137 , n25136 , n23211 );
nand ( n25138 , n25134 , n25137 );
not ( n25139 , n2 );
and ( n25140 , n31 , n23511 );
and ( n25141 , n1276 , n23204 );
nor ( n25142 , n25140 , n25141 );
nor ( n25143 , n25139 , n25142 );
not ( n25144 , n2 );
and ( n25145 , n37 , n23584 );
and ( n25146 , n1272 , n23204 );
nor ( n25147 , n25145 , n25146 );
nor ( n25148 , n25144 , n25147 );
not ( n25149 , n2 );
and ( n25150 , n42 , n23517 );
and ( n25151 , n1268 , n23204 );
nor ( n25152 , n25150 , n25151 );
nor ( n25153 , n25149 , n25152 );
not ( n25154 , n2 );
and ( n25155 , n32 , n24529 );
and ( n25156 , n1252 , n23156 );
nor ( n25157 , n25155 , n25156 );
nor ( n25158 , n25154 , n25157 );
not ( n25159 , n2 );
and ( n25160 , n49 , n23559 );
and ( n25161 , n1439 , n23188 );
nor ( n25162 , n25160 , n25161 );
nor ( n25163 , n25159 , n25162 );
not ( n25164 , n2 );
and ( n25165 , n37 , n23553 );
and ( n25166 , n1260 , n23188 );
nor ( n25167 , n25165 , n25166 );
nor ( n25168 , n25164 , n25167 );
not ( n25169 , n2 );
and ( n25170 , n39 , n24503 );
and ( n25171 , n1254 , n23156 );
nor ( n25172 , n25170 , n25171 );
nor ( n25173 , n25169 , n25172 );
not ( n25174 , n2 );
and ( n25175 , n32 , n24186 );
and ( n25176 , n1264 , n23188 );
nor ( n25177 , n25175 , n25176 );
nor ( n25178 , n25174 , n25177 );
not ( n25179 , n2 );
and ( n25180 , n42 , n23547 );
and ( n25181 , n1256 , n23188 );
nor ( n25182 , n25180 , n25181 );
nor ( n25183 , n25179 , n25182 );
not ( n25184 , n2 );
and ( n25185 , n42 , n24529 );
and ( n25186 , n1248 , n23156 );
nor ( n25187 , n25185 , n25186 );
nor ( n25188 , n25184 , n25187 );
not ( n25189 , n2 );
and ( n25190 , n37 , n24694 );
and ( n25191 , n1240 , n23128 );
nor ( n25192 , n25190 , n25191 );
nor ( n25193 , n25189 , n25192 );
not ( n25194 , n2 );
and ( n25195 , n34 , n24754 );
and ( n25196 , n1244 , n23128 );
nor ( n25197 , n25195 , n25196 );
nor ( n25198 , n25194 , n25197 );
not ( n25199 , n2 );
and ( n25200 , n47 , n23827 );
and ( n25201 , n1236 , n23128 );
nor ( n25202 , n25200 , n25201 );
nor ( n25203 , n25199 , n25202 );
not ( n25204 , n2 );
and ( n25205 , n40 , n24754 );
and ( n25206 , n1232 , n23128 );
nor ( n25207 , n25205 , n25206 );
nor ( n25208 , n25204 , n25207 );
not ( n25209 , n2 );
and ( n25210 , n50 , n23529 );
and ( n25211 , n1225 , n23531 );
nor ( n25212 , n25210 , n25211 );
nor ( n25213 , n25209 , n25212 );
nand ( n25214 , n1214 , n24937 );
nand ( n25215 , n25214 , n2 , n22447 );
not ( n25216 , n17056 );
nand ( n25217 , n25216 , n17052 );
not ( n25218 , n25217 );
not ( n25219 , n19355 );
or ( n25220 , n25218 , n25219 );
or ( n25221 , n25217 , n19355 );
nand ( n25222 , n25220 , n25221 );
not ( n25223 , n15675 );
not ( n25224 , n312 );
nand ( n25225 , n25224 , n1179 , n19391 );
and ( n25226 , n25223 , n25225 );
nor ( n25227 , n25226 , n21342 );
not ( n25228 , n16915 );
nand ( n25229 , n25228 , n16911 );
not ( n25230 , n25229 );
not ( n25231 , n19223 );
or ( n25232 , n25230 , n25231 );
or ( n25233 , n25229 , n19223 );
nand ( n25234 , n25232 , n25233 );
or ( n25235 , n16844 , n16837 );
not ( n25236 , n25235 );
not ( n25237 , n19312 );
or ( n25238 , n25236 , n25237 );
or ( n25239 , n25235 , n19312 );
nand ( n25240 , n25238 , n25239 );
not ( n25241 , n16986 );
nand ( n25242 , n25241 , n16982 );
not ( n25243 , n25242 );
not ( n25244 , n19267 );
or ( n25245 , n25243 , n25244 );
or ( n25246 , n25242 , n19267 );
nand ( n25247 , n25245 , n25246 );
not ( n25248 , n2 );
and ( n25249 , n17 , n15947 );
nor ( n25250 , n14 , n21587 );
nand ( n25251 , n15961 , n25249 , n25250 , n21590 );
buf ( n25252 , n25251 );
not ( n25253 , n25252 );
and ( n25254 , n31 , n25253 );
and ( n25255 , n1457 , n25252 );
nor ( n25256 , n25254 , n25255 );
nor ( n25257 , n25248 , n25256 );
or ( n25258 , n15122 , n15097 );
and ( n25259 , n15123 , n15148 );
or ( n25260 , n25259 , n16794 );
and ( n25261 , n25259 , n16794 );
not ( n25262 , n15095 );
nor ( n25263 , n25261 , n25262 );
nand ( n25264 , n25260 , n25263 );
nand ( n25265 , n25258 , n25264 );
and ( n25266 , n15090 , n25265 );
and ( n25267 , n15193 , n15122 );
not ( n25268 , n15193 );
and ( n25269 , n25268 , n782 );
nor ( n25270 , n25267 , n25269 );
and ( n25271 , n1826 , n25270 );
nor ( n25272 , n25266 , n25271 );
nor ( n25273 , n15089 , n25272 );
or ( n25274 , n232 , n13757 );
nand ( n25275 , n25274 , n14490 );
nand ( n25276 , n353 , n20636 );
nand ( n25277 , n368 , n20638 );
not ( n25278 , n25277 );
nand ( n25279 , n25278 , n369 );
nor ( n25280 , n14543 , n19937 , n25279 );
or ( n25281 , n353 , n25280 );
and ( n25282 , n353 , n25280 );
not ( n25283 , n20633 );
nor ( n25284 , n25282 , n25283 );
nand ( n25285 , n25281 , n25284 );
and ( n25286 , n25276 , n25285 );
nor ( n25287 , n25286 , n20652 );
not ( n25288 , n1078 );
nor ( n25289 , n1109 , n1470 );
not ( n25290 , n1256 );
nand ( n25291 , n1437 , n25290 );
and ( n25292 , n1659 , n15736 );
nand ( n25293 , n1659 , n1681 );
nor ( n25294 , n1258 , n25293 );
nor ( n25295 , n25292 , n25294 );
or ( n25296 , n1157 , n1258 );
not ( n25297 , n25296 );
nand ( n25298 , n1681 , n25297 );
not ( n25299 , n1439 );
or ( n25300 , n25299 , n1687 );
not ( n25301 , n1258 );
and ( n25302 , n1659 , n25301 );
and ( n25303 , n1681 , n15736 );
nor ( n25304 , n25302 , n25303 );
and ( n25305 , n25304 , n25293 , n25296 );
and ( n25306 , n1687 , n25299 );
not ( n25307 , n1156 );
nor ( n25308 , n25306 , n25307 , n1759 );
nor ( n25309 , n25305 , n25308 );
nand ( n25310 , n25300 , n25309 );
and ( n25311 , n25295 , n25298 , n25310 );
not ( n25312 , n1259 );
and ( n25313 , n1629 , n25312 );
not ( n25314 , n1212 );
and ( n25315 , n1581 , n25314 );
nor ( n25316 , n25313 , n25315 );
nand ( n25317 , n1581 , n1629 );
or ( n25318 , n1212 , n1259 );
and ( n25319 , n25316 , n25317 , n25318 );
nor ( n25320 , n25311 , n25319 );
not ( n25321 , n1437 );
nand ( n25322 , n25321 , n1256 );
not ( n25323 , n1205 );
and ( n25324 , n1549 , n25323 );
not ( n25325 , n1158 );
and ( n25326 , n1573 , n25325 );
nor ( n25327 , n25324 , n25326 );
nand ( n25328 , n1549 , n1573 );
nor ( n25329 , n1158 , n1205 );
not ( n25330 , n25329 );
nand ( n25331 , n25327 , n25328 , n25330 );
and ( n25332 , n25320 , n25322 , n25331 );
or ( n25333 , n1212 , n25317 );
not ( n25334 , n25318 );
nand ( n25335 , n1629 , n25334 );
nand ( n25336 , n25333 , n25335 );
and ( n25337 , n25336 , n25331 );
not ( n25338 , n25328 );
and ( n25339 , n25323 , n25338 );
nor ( n25340 , n25337 , n25339 );
and ( n25341 , n1573 , n25329 );
and ( n25342 , n1549 , n25325 );
nor ( n25343 , n25341 , n25342 );
nand ( n25344 , n1581 , n25312 , n25331 );
nand ( n25345 , n25340 , n25343 , n25344 );
and ( n25346 , n25322 , n25345 );
nor ( n25347 , n25332 , n25346 );
nand ( n25348 , n25288 , n25289 , n25291 , n25347 );
not ( n25349 , n1077 );
nor ( n25350 , n1108 , n1469 );
not ( n25351 , n1248 );
nand ( n25352 , n1436 , n25351 );
not ( n25353 , n1401 );
and ( n25354 , n1658 , n25353 );
nand ( n25355 , n1658 , n1682 );
nor ( n25356 , n1152 , n25355 );
nor ( n25357 , n25354 , n25356 );
or ( n25358 , n1152 , n1401 );
not ( n25359 , n25358 );
nand ( n25360 , n1682 , n25359 );
not ( n25361 , n1406 );
or ( n25362 , n25361 , n1688 );
and ( n25363 , n1682 , n25353 );
not ( n25364 , n1152 );
and ( n25365 , n1658 , n25364 );
nor ( n25366 , n25363 , n25365 );
and ( n25367 , n25366 , n25355 , n25358 );
and ( n25368 , n1688 , n25361 );
not ( n25369 , n1151 );
nor ( n25370 , n25368 , n25369 , n1753 );
nor ( n25371 , n25367 , n25370 );
nand ( n25372 , n25362 , n25371 );
and ( n25373 , n25357 , n25360 , n25372 );
not ( n25374 , n1403 );
and ( n25375 , n1628 , n25374 );
not ( n25376 , n1250 );
and ( n25377 , n1579 , n25376 );
nor ( n25378 , n25375 , n25377 );
nand ( n25379 , n1579 , n1628 );
or ( n25380 , n1250 , n1403 );
and ( n25381 , n25378 , n25379 , n25380 );
nor ( n25382 , n25373 , n25381 );
not ( n25383 , n1436 );
nand ( n25384 , n25383 , n1248 );
and ( n25385 , n1561 , n14993 );
not ( n25386 , n1396 );
and ( n25387 , n1572 , n25386 );
nor ( n25388 , n25385 , n25387 );
nand ( n25389 , n1561 , n1572 );
nor ( n25390 , n1396 , n1399 );
not ( n25391 , n25390 );
nand ( n25392 , n25388 , n25389 , n25391 );
and ( n25393 , n25382 , n25384 , n25392 );
or ( n25394 , n1250 , n25379 );
not ( n25395 , n25380 );
nand ( n25396 , n1628 , n25395 );
nand ( n25397 , n25394 , n25396 );
and ( n25398 , n25397 , n25392 );
not ( n25399 , n25389 );
and ( n25400 , n14993 , n25399 );
nor ( n25401 , n25398 , n25400 );
and ( n25402 , n1572 , n25390 );
and ( n25403 , n1561 , n25386 );
nor ( n25404 , n25402 , n25403 );
nand ( n25405 , n1579 , n25374 , n25392 );
nand ( n25406 , n25401 , n25404 , n25405 );
and ( n25407 , n25384 , n25406 );
nor ( n25408 , n25393 , n25407 );
nand ( n25409 , n25349 , n25350 , n25352 , n25408 );
not ( n25410 , n1079 );
nor ( n25411 , n1110 , n1528 );
not ( n25412 , n1268 );
nand ( n25413 , n1438 , n25412 );
not ( n25414 , n1387 );
and ( n25415 , n1660 , n25414 );
nand ( n25416 , n1660 , n1684 );
nor ( n25417 , n1270 , n25416 );
nor ( n25418 , n25415 , n25417 );
or ( n25419 , n1270 , n1387 );
not ( n25420 , n25419 );
nand ( n25421 , n1684 , n25420 );
not ( n25422 , n1471 );
or ( n25423 , n25422 , n1686 );
and ( n25424 , n1684 , n25414 );
not ( n25425 , n1270 );
and ( n25426 , n1660 , n25425 );
nor ( n25427 , n25424 , n25426 );
and ( n25428 , n25427 , n25416 , n25419 );
and ( n25429 , n1686 , n25422 );
not ( n25430 , n1161 );
nor ( n25431 , n25429 , n25430 , n1752 );
nor ( n25432 , n25428 , n25431 );
nand ( n25433 , n25423 , n25432 );
and ( n25434 , n25418 , n25421 , n25433 );
not ( n25435 , n1271 );
and ( n25436 , n1630 , n25435 );
not ( n25437 , n1162 );
and ( n25438 , n1582 , n25437 );
nor ( n25439 , n25436 , n25438 );
nand ( n25440 , n1582 , n1630 );
or ( n25441 , n1162 , n1271 );
and ( n25442 , n25439 , n25440 , n25441 );
nor ( n25443 , n25434 , n25442 );
not ( n25444 , n1438 );
nand ( n25445 , n25444 , n1268 );
and ( n25446 , n1562 , n15110 );
not ( n25447 , n1163 );
and ( n25448 , n1575 , n25447 );
nor ( n25449 , n25446 , n25448 );
nand ( n25450 , n1562 , n1575 );
nor ( n25451 , n1163 , n1394 );
not ( n25452 , n25451 );
nand ( n25453 , n25449 , n25450 , n25452 );
and ( n25454 , n25443 , n25445 , n25453 );
or ( n25455 , n1162 , n25440 );
not ( n25456 , n25441 );
nand ( n25457 , n1630 , n25456 );
nand ( n25458 , n25455 , n25457 );
and ( n25459 , n25458 , n25453 );
not ( n25460 , n25450 );
and ( n25461 , n15110 , n25460 );
nor ( n25462 , n25459 , n25461 );
and ( n25463 , n1575 , n25451 );
and ( n25464 , n1562 , n25447 );
nor ( n25465 , n25463 , n25464 );
nand ( n25466 , n1582 , n25435 , n25453 );
nand ( n25467 , n25462 , n25465 , n25466 );
and ( n25468 , n25445 , n25467 );
nor ( n25469 , n25454 , n25468 );
nand ( n25470 , n25410 , n25411 , n25413 , n25469 );
not ( n25471 , n1076 );
nor ( n25472 , n1107 , n1527 );
nand ( n25473 , n1435 , n23081 );
not ( n25474 , n1236 );
and ( n25475 , n1657 , n25474 );
nand ( n25476 , n1657 , n1683 );
nor ( n25477 , n1235 , n25476 );
nor ( n25478 , n25475 , n25477 );
or ( n25479 , n1235 , n1236 );
not ( n25480 , n25479 );
nand ( n25481 , n1683 , n25480 );
not ( n25482 , n1467 );
or ( n25483 , n25482 , n1689 );
and ( n25484 , n1683 , n25474 );
not ( n25485 , n1235 );
and ( n25486 , n1657 , n25485 );
nor ( n25487 , n25484 , n25486 );
and ( n25488 , n25487 , n25476 , n25479 );
and ( n25489 , n1689 , n25482 );
not ( n25490 , n1234 );
nor ( n25491 , n25489 , n25490 , n1751 );
nor ( n25492 , n25488 , n25491 );
nand ( n25493 , n25483 , n25492 );
and ( n25494 , n25478 , n25481 , n25493 );
and ( n25495 , n1580 , n16273 );
not ( n25496 , n1210 );
and ( n25497 , n1627 , n25496 );
nor ( n25498 , n25495 , n25497 );
nand ( n25499 , n1580 , n1627 );
or ( n25500 , n1210 , n1237 );
and ( n25501 , n25498 , n25499 , n25500 );
nor ( n25502 , n25494 , n25501 );
not ( n25503 , n1435 );
nand ( n25504 , n25503 , n1231 );
and ( n25505 , n1571 , n16338 );
and ( n25506 , n1560 , n16300 );
nor ( n25507 , n25505 , n25506 );
nand ( n25508 , n1560 , n1571 );
nor ( n25509 , n1238 , n1239 );
not ( n25510 , n25509 );
nand ( n25511 , n25507 , n25508 , n25510 );
and ( n25512 , n25502 , n25504 , n25511 );
or ( n25513 , n1237 , n25499 );
not ( n25514 , n25500 );
nand ( n25515 , n1627 , n25514 );
nand ( n25516 , n25513 , n25515 );
and ( n25517 , n25516 , n25511 );
not ( n25518 , n25508 );
and ( n25519 , n16300 , n25518 );
nor ( n25520 , n25517 , n25519 );
and ( n25521 , n1571 , n25509 );
and ( n25522 , n1560 , n16338 );
nor ( n25523 , n25521 , n25522 );
nand ( n25524 , n1580 , n25496 , n25511 );
nand ( n25525 , n25520 , n25523 , n25524 );
and ( n25526 , n25504 , n25525 );
nor ( n25527 , n25512 , n25526 );
nand ( n25528 , n25471 , n25472 , n25473 , n25527 );
and ( n25529 , n447 , n23600 );
and ( n25530 , n140 , n23599 );
nor ( n25531 , n25529 , n25530 );
not ( n25532 , n23627 );
or ( n25533 , n25531 , n25532 );
or ( n25534 , n16029 , n23627 );
nand ( n25535 , n25533 , n25534 , n2 );
and ( n25536 , n451 , n23600 );
and ( n25537 , n145 , n23599 );
nor ( n25538 , n25536 , n25537 );
or ( n25539 , n25538 , n25532 );
or ( n25540 , n16045 , n23627 );
nand ( n25541 , n25539 , n25540 , n2 );
and ( n25542 , n452 , n23600 );
and ( n25543 , n136 , n23599 );
nor ( n25544 , n25542 , n25543 );
not ( n25545 , n23627 );
or ( n25546 , n25544 , n25545 );
or ( n25547 , n16033 , n23610 );
nand ( n25548 , n25546 , n25547 , n2 );
and ( n25549 , n454 , n23600 );
and ( n25550 , n148 , n23599 );
nor ( n25551 , n25549 , n25550 );
or ( n25552 , n25551 , n25545 );
or ( n25553 , n16041 , n23610 );
nand ( n25554 , n25552 , n25553 , n2 );
and ( n25555 , n458 , n23600 );
and ( n25556 , n157 , n23599 );
nor ( n25557 , n25555 , n25556 );
or ( n25558 , n25557 , n25545 );
or ( n25559 , n16061 , n23627 );
nand ( n25560 , n25558 , n25559 , n2 );
or ( n25561 , n15965 , n23627 );
or ( n25562 , n1795 , n23600 );
or ( n25563 , n464 , n23599 );
nand ( n25564 , n25562 , n25563 , n23627 );
nand ( n25565 , n25561 , n2 , n25564 );
and ( n25566 , n519 , n23600 );
and ( n25567 , n143 , n23599 );
nor ( n25568 , n25566 , n25567 );
or ( n25569 , n25568 , n25532 );
or ( n25570 , n16081 , n23627 );
nand ( n25571 , n25569 , n25570 , n2 );
and ( n25572 , n522 , n23600 );
and ( n25573 , n461 , n23599 );
nor ( n25574 , n25572 , n25573 );
or ( n25575 , n25574 , n25532 );
or ( n25576 , n16009 , n23627 );
nand ( n25577 , n25575 , n25576 , n2 );
and ( n25578 , n524 , n23600 );
and ( n25579 , n428 , n23599 );
nor ( n25580 , n25578 , n25579 );
or ( n25581 , n25580 , n25545 );
or ( n25582 , n16005 , n23627 );
nand ( n25583 , n25581 , n25582 , n2 );
not ( n25584 , n17331 );
and ( n25585 , n541 , n25584 );
not ( n25586 , n17332 );
nor ( n25587 , n25585 , n14974 , n25586 );
and ( n25588 , n541 , n18536 );
nand ( n25589 , n17284 , n17287 );
not ( n25590 , n17859 );
and ( n25591 , n25589 , n25590 );
or ( n25592 , n25589 , n25590 );
not ( n25593 , n14979 );
nand ( n25594 , n25592 , n25593 );
nor ( n25595 , n25591 , n25594 );
nor ( n25596 , n25588 , n1819 , n25595 );
nor ( n25597 , n14973 , n25587 , n25596 );
nand ( n25598 , n596 , n22477 );
not ( n25599 , n20234 );
or ( n25600 , n596 , n25599 );
not ( n25601 , n20235 );
nand ( n25602 , n25600 , n1800 , n25601 );
and ( n25603 , n25598 , n25602 );
nor ( n25604 , n25603 , n834 );
nand ( n25605 , n608 , n22477 );
or ( n25606 , n608 , n22481 );
and ( n25607 , n608 , n22481 );
nor ( n25608 , n25607 , n22477 );
nand ( n25609 , n25606 , n25608 );
and ( n25610 , n25605 , n25609 );
nor ( n25611 , n25610 , n834 );
not ( n25612 , n17412 );
and ( n25613 , n642 , n25612 );
not ( n25614 , n17413 );
nor ( n25615 , n25613 , n15704 , n25614 );
and ( n25616 , n642 , n16393 );
nand ( n25617 , n17365 , n17368 );
not ( n25618 , n17910 );
and ( n25619 , n25617 , n25618 );
or ( n25620 , n25617 , n25618 );
nand ( n25621 , n25620 , n15709 );
nor ( n25622 , n25619 , n25621 );
nor ( n25623 , n25616 , n1808 , n25622 );
nor ( n25624 , n15703 , n25615 , n25623 );
not ( n25625 , n2 );
and ( n25626 , n32 , n25253 );
and ( n25627 , n1456 , n25252 );
nor ( n25628 , n25626 , n25627 );
nor ( n25629 , n25625 , n25628 );
not ( n25630 , n2 );
and ( n25631 , n34 , n25253 );
and ( n25632 , n1455 , n25252 );
nor ( n25633 , n25631 , n25632 );
nor ( n25634 , n25630 , n25633 );
or ( n25635 , n15750 , n15710 );
and ( n25636 , n15751 , n15764 );
or ( n25637 , n25636 , n17169 );
and ( n25638 , n25636 , n17169 );
not ( n25639 , n15709 );
nor ( n25640 , n25638 , n25639 );
nand ( n25641 , n25637 , n25640 );
nand ( n25642 , n25635 , n25641 );
and ( n25643 , n15704 , n25642 );
and ( n25644 , n15793 , n15750 );
not ( n25645 , n15793 );
and ( n25646 , n25645 , n716 );
nor ( n25647 , n25644 , n25646 );
and ( n25648 , n1808 , n25647 );
nor ( n25649 , n25643 , n25648 );
nor ( n25650 , n15703 , n25649 );
not ( n25651 , n17676 );
and ( n25652 , n719 , n25651 );
not ( n25653 , n17677 );
nor ( n25654 , n25652 , n15090 , n25653 );
and ( n25655 , n719 , n18627 );
nand ( n25656 , n17628 , n17631 );
not ( n25657 , n17765 );
and ( n25658 , n25656 , n25657 );
or ( n25659 , n25656 , n25657 );
nand ( n25660 , n25659 , n15095 );
nor ( n25661 , n25658 , n25660 );
nor ( n25662 , n25655 , n1826 , n25661 );
nor ( n25663 , n15089 , n25654 , n25662 );
or ( n25664 , n23607 , n21760 );
buf ( n25665 , n25664 );
or ( n25666 , n16057 , n25665 );
not ( n25667 , n1125 );
not ( n25668 , n1609 );
or ( n25669 , n25667 , n25668 );
nand ( n25670 , n1609 , n1858 );
nand ( n25671 , n25669 , n25670 );
not ( n25672 , n25671 );
or ( n25673 , n159 , n25672 );
or ( n25674 , n753 , n25671 );
buf ( n25675 , n25664 );
nand ( n25676 , n25673 , n25674 , n25675 );
nand ( n25677 , n25666 , n2 , n25676 );
not ( n25678 , n25671 );
buf ( n25679 , n25678 );
and ( n25680 , n757 , n25679 );
not ( n25681 , n25678 );
and ( n25682 , n157 , n25681 );
nor ( n25683 , n25680 , n25682 );
not ( n25684 , n25675 );
or ( n25685 , n25683 , n25684 );
or ( n25686 , n16061 , n25665 );
nand ( n25687 , n25685 , n25686 , n2 );
or ( n25688 , n15901 , n25665 );
not ( n25689 , n25671 );
or ( n25690 , n152 , n25689 );
or ( n25691 , n762 , n25671 );
nand ( n25692 , n25690 , n25691 , n25675 );
nand ( n25693 , n25688 , n2 , n25692 );
or ( n25694 , n16029 , n25665 );
or ( n25695 , n140 , n25689 );
or ( n25696 , n764 , n25671 );
nand ( n25697 , n25695 , n25696 , n25675 );
nand ( n25698 , n25694 , n2 , n25697 );
and ( n25699 , n765 , n25679 );
not ( n25700 , n25671 );
not ( n25701 , n25700 );
and ( n25702 , n145 , n25701 );
nor ( n25703 , n25699 , n25702 );
not ( n25704 , n25675 );
or ( n25705 , n25703 , n25704 );
or ( n25706 , n16045 , n25665 );
nand ( n25707 , n25705 , n25706 , n2 );
and ( n25708 , n766 , n25679 );
not ( n25709 , n25700 );
and ( n25710 , n136 , n25709 );
nor ( n25711 , n25708 , n25710 );
or ( n25712 , n25711 , n25704 );
or ( n25713 , n16033 , n25665 );
nand ( n25714 , n25712 , n25713 , n2 );
and ( n25715 , n767 , n25679 );
and ( n25716 , n148 , n25709 );
nor ( n25717 , n25715 , n25716 );
not ( n25718 , n25675 );
or ( n25719 , n25717 , n25718 );
or ( n25720 , n16041 , n25665 );
nand ( n25721 , n25719 , n25720 , n2 );
and ( n25722 , n768 , n25679 );
not ( n25723 , n25700 );
and ( n25724 , n147 , n25723 );
nor ( n25725 , n25722 , n25724 );
not ( n25726 , n25675 );
or ( n25727 , n25725 , n25726 );
or ( n25728 , n16025 , n25665 );
nand ( n25729 , n25727 , n25728 , n2 );
and ( n25730 , n770 , n25679 );
and ( n25731 , n175 , n25723 );
nor ( n25732 , n25730 , n25731 );
or ( n25733 , n25732 , n25684 );
or ( n25734 , n16085 , n25665 );
nand ( n25735 , n25733 , n25734 , n2 );
and ( n25736 , n780 , n25679 );
not ( n25737 , n25700 );
and ( n25738 , n1801 , n25737 );
nor ( n25739 , n25736 , n25738 );
or ( n25740 , n25739 , n25726 );
or ( n25741 , n16065 , n25665 );
nand ( n25742 , n25740 , n25741 , n2 );
and ( n25743 , n781 , n25679 );
and ( n25744 , n1795 , n25723 );
nor ( n25745 , n25743 , n25744 );
or ( n25746 , n25745 , n25726 );
or ( n25747 , n15965 , n25665 );
nand ( n25748 , n25746 , n25747 , n2 );
and ( n25749 , n796 , n25679 );
and ( n25750 , n283 , n25681 );
nor ( n25751 , n25749 , n25750 );
not ( n25752 , n25675 );
or ( n25753 , n25751 , n25752 );
or ( n25754 , n15985 , n25665 );
nand ( n25755 , n25753 , n25754 , n2 );
and ( n25756 , n797 , n25679 );
and ( n25757 , n415 , n25737 );
nor ( n25758 , n25756 , n25757 );
or ( n25759 , n25758 , n25684 );
or ( n25760 , n16001 , n25665 );
nand ( n25761 , n25759 , n25760 , n2 );
and ( n25762 , n799 , n25679 );
and ( n25763 , n193 , n25701 );
nor ( n25764 , n25762 , n25763 );
or ( n25765 , n25764 , n25704 );
or ( n25766 , n16089 , n25665 );
nand ( n25767 , n25765 , n25766 , n2 );
and ( n25768 , n800 , n25679 );
and ( n25769 , n439 , n25701 );
nor ( n25770 , n25768 , n25769 );
or ( n25771 , n25770 , n25726 );
or ( n25772 , n16013 , n25665 );
nand ( n25773 , n25771 , n25772 , n2 );
and ( n25774 , n809 , n25679 );
and ( n25775 , n143 , n25709 );
nor ( n25776 , n25774 , n25775 );
or ( n25777 , n25776 , n25718 );
or ( n25778 , n16081 , n25665 );
nand ( n25779 , n25777 , n25778 , n2 );
or ( n25780 , n16021 , n25665 );
or ( n25781 , n144 , n25689 );
or ( n25782 , n810 , n25671 );
nand ( n25783 , n25781 , n25782 , n25675 );
nand ( n25784 , n25780 , n2 , n25783 );
and ( n25785 , n811 , n25679 );
and ( n25786 , n1082 , n25681 );
nor ( n25787 , n25785 , n25786 );
or ( n25788 , n25787 , n25752 );
or ( n25789 , n16017 , n25665 );
nand ( n25790 , n25788 , n25789 , n2 );
or ( n25791 , n16009 , n25665 );
not ( n25792 , n25671 );
or ( n25793 , n461 , n25792 );
or ( n25794 , n812 , n25671 );
nand ( n25795 , n25793 , n25794 , n25675 );
nand ( n25796 , n25791 , n2 , n25795 );
and ( n25797 , n813 , n25679 );
and ( n25798 , n186 , n25681 );
nor ( n25799 , n25797 , n25798 );
or ( n25800 , n25799 , n25752 );
or ( n25801 , n16077 , n25665 );
nand ( n25802 , n25800 , n25801 , n2 );
and ( n25803 , n814 , n25679 );
and ( n25804 , n428 , n25681 );
nor ( n25805 , n25803 , n25804 );
or ( n25806 , n25805 , n25752 );
or ( n25807 , n16005 , n25665 );
nand ( n25808 , n25806 , n25807 , n2 );
not ( n25809 , n2 );
and ( n25810 , n51 , n25253 );
and ( n25811 , n1448 , n25252 );
nor ( n25812 , n25810 , n25811 );
nor ( n25813 , n25809 , n25812 );
and ( n25814 , n815 , n25672 );
and ( n25815 , n1610 , n25701 );
nor ( n25816 , n25814 , n25815 );
or ( n25817 , n25816 , n25684 );
or ( n25818 , n15997 , n25665 );
nand ( n25819 , n25817 , n25818 , n2 );
not ( n25820 , n16 );
or ( n25821 , n25820 , n23525 );
not ( n25822 , n25821 );
not ( n25823 , n25822 );
or ( n25824 , n21585 , n23123 );
not ( n25825 , n25824 );
and ( n25826 , n315 , n25825 );
nand ( n25827 , n15951 , n22151 );
not ( n25828 , n25827 );
and ( n25829 , n1106 , n25828 );
nor ( n25830 , n25826 , n25829 );
or ( n25831 , n25823 , n25830 );
nand ( n25832 , n25820 , n23526 );
buf ( n25833 , n25832 );
or ( n25834 , n25833 , n25830 );
not ( n25835 , n21580 );
and ( n25836 , n479 , n25835 );
not ( n25837 , n21740 );
and ( n25838 , n1478 , n25837 );
nor ( n25839 , n25836 , n25838 );
not ( n25840 , n25839 );
not ( n25841 , n23124 );
and ( n25842 , n1068 , n25841 );
not ( n25843 , n22151 );
not ( n25844 , n25843 );
and ( n25845 , n535 , n25844 );
nor ( n25846 , n25842 , n25845 );
not ( n25847 , n25846 );
or ( n25848 , n25840 , n25847 );
and ( n25849 , n15952 , n21746 , n21586 );
nand ( n25850 , n25848 , n25849 );
nand ( n25851 , n25834 , n25850 );
not ( n25852 , n21581 );
and ( n25853 , n556 , n25852 );
not ( n25854 , n21740 );
not ( n25855 , n25854 );
not ( n25856 , n25855 );
and ( n25857 , n1536 , n25856 );
nor ( n25858 , n25853 , n25857 );
and ( n25859 , n1098 , n23125 );
not ( n25860 , n23604 );
and ( n25861 , n633 , n25860 );
nor ( n25862 , n25859 , n25861 );
and ( n25863 , n25858 , n25862 );
not ( n25864 , n21584 );
nand ( n25865 , n25864 , n21586 );
not ( n25866 , n25865 );
nand ( n25867 , n25820 , n25866 );
buf ( n25868 , n25867 );
nor ( n25869 , n25863 , n25868 );
not ( n25870 , n21579 );
not ( n25871 , n25870 );
and ( n25872 , n440 , n25871 );
not ( n25873 , n23604 );
and ( n25874 , n463 , n25873 );
nor ( n25875 , n25872 , n25874 );
not ( n25876 , n23153 );
and ( n25877 , n992 , n25876 );
not ( n25878 , n25855 );
and ( n25879 , n1525 , n25878 );
nor ( n25880 , n25877 , n25879 );
and ( n25881 , n25875 , n25880 );
and ( n25882 , n25820 , n21746 , n21586 );
not ( n25883 , n25882 );
nor ( n25884 , n25881 , n25883 );
nor ( n25885 , n25851 , n25869 , n25884 );
not ( n25886 , n21582 );
and ( n25887 , n644 , n25886 );
buf ( n25888 , n21741 );
not ( n25889 , n25888 );
and ( n25890 , n1482 , n25889 );
nor ( n25891 , n25887 , n25890 );
not ( n25892 , n25891 );
buf ( n25893 , n23124 );
not ( n25894 , n25893 );
buf ( n25895 , n25894 );
and ( n25896 , n1123 , n25895 );
and ( n25897 , n780 , n23606 );
nor ( n25898 , n25896 , n25897 );
not ( n25899 , n25898 );
or ( n25900 , n25892 , n25899 );
or ( n25901 , n23523 , n25865 );
not ( n25902 , n25901 );
nand ( n25903 , n25900 , n25902 );
nand ( n25904 , n25831 , n25885 , n25903 );
or ( n25905 , n15993 , n25665 );
or ( n25906 , n383 , n25689 );
or ( n25907 , n816 , n25671 );
nand ( n25908 , n25906 , n25907 , n25675 );
nand ( n25909 , n25905 , n2 , n25908 );
and ( n25910 , n817 , n25679 );
and ( n25911 , n352 , n25681 );
nor ( n25912 , n25910 , n25911 );
or ( n25913 , n25912 , n25752 );
or ( n25914 , n15989 , n25665 );
nand ( n25915 , n25913 , n25914 , n2 );
or ( n25916 , n15977 , n25665 );
or ( n25917 , n253 , n25792 );
or ( n25918 , n818 , n25671 );
nand ( n25919 , n25917 , n25918 , n25675 );
nand ( n25920 , n25916 , n2 , n25919 );
and ( n25921 , n819 , n25679 );
and ( n25922 , n284 , n25681 );
nor ( n25923 , n25921 , n25922 );
or ( n25924 , n25923 , n25704 );
or ( n25925 , n15981 , n25665 );
nand ( n25926 , n25924 , n25925 , n2 );
and ( n25927 , n820 , n25672 );
and ( n25928 , n192 , n25737 );
nor ( n25929 , n25927 , n25928 );
or ( n25930 , n25929 , n25752 );
or ( n25931 , n15969 , n25665 );
nand ( n25932 , n25930 , n25931 , n2 );
not ( n25933 , n21582 );
and ( n25934 , n450 , n25933 );
and ( n25935 , n1094 , n21742 );
nor ( n25936 , n25934 , n25935 );
and ( n25937 , n1250 , n25895 );
not ( n25938 , n25860 );
not ( n25939 , n25938 );
and ( n25940 , n456 , n25939 );
nor ( n25941 , n25937 , n25940 );
nand ( n25942 , n25936 , n25941 );
and ( n25943 , n25882 , n25942 );
buf ( n25944 , n21581 );
not ( n25945 , n25944 );
and ( n25946 , n578 , n25945 );
not ( n25947 , n23605 );
and ( n25948 , n590 , n25947 );
nor ( n25949 , n25946 , n25948 );
and ( n25950 , n1162 , n25895 );
and ( n25951 , n1177 , n21742 );
nor ( n25952 , n25950 , n25951 );
and ( n25953 , n25949 , n25952 );
nor ( n25954 , n25953 , n25868 );
nor ( n25955 , n25943 , n25954 );
nand ( n25956 , n25821 , n25832 );
nand ( n25957 , n23523 , n21579 );
not ( n25958 , n25957 );
and ( n25959 , n1451 , n25958 );
or ( n25960 , n23523 , n21738 );
not ( n25961 , n25960 );
and ( n25962 , n1822 , n25961 );
nor ( n25963 , n25959 , n25962 );
and ( n25964 , n577 , n25825 );
and ( n25965 , n1227 , n23524 );
nor ( n25966 , n25964 , n25965 );
nand ( n25967 , n25963 , n25966 );
and ( n25968 , n25956 , n25967 );
buf ( n25969 , n25870 );
not ( n25970 , n25969 );
and ( n25971 , n679 , n25970 );
and ( n25972 , n762 , n22154 );
nor ( n25973 , n25971 , n25972 );
not ( n25974 , n23124 );
buf ( n25975 , n25974 );
and ( n25976 , n1237 , n25975 );
not ( n25977 , n21741 );
and ( n25978 , n1443 , n25977 );
nor ( n25979 , n25976 , n25978 );
and ( n25980 , n25973 , n25979 );
nor ( n25981 , n25980 , n25901 );
not ( n25982 , n25969 );
and ( n25983 , n491 , n25982 );
and ( n25984 , n1119 , n25856 );
nor ( n25985 , n25983 , n25984 );
and ( n25986 , n1212 , n23125 );
and ( n25987 , n486 , n25873 );
nor ( n25988 , n25986 , n25987 );
and ( n25989 , n25985 , n25988 );
not ( n25990 , n25849 );
nor ( n25991 , n25989 , n25990 );
nor ( n25992 , n25968 , n25981 , n25991 );
nand ( n25993 , n25955 , n25992 );
and ( n25994 , n821 , n25679 );
and ( n25995 , n185 , n25681 );
nor ( n25996 , n25994 , n25995 );
or ( n25997 , n25996 , n25718 );
or ( n25998 , n16073 , n25665 );
nand ( n25999 , n25997 , n25998 , n2 );
or ( n26000 , n16049 , n25665 );
or ( n26001 , n151 , n25792 );
or ( n26002 , n822 , n25671 );
nand ( n26003 , n26001 , n26002 , n25675 );
nand ( n26004 , n26000 , n2 , n26003 );
or ( n26005 , n16053 , n25665 );
or ( n26006 , n156 , n25792 );
or ( n26007 , n823 , n25671 );
nand ( n26008 , n26006 , n26007 , n25675 );
nand ( n26009 , n26005 , n2 , n26008 );
not ( n26010 , n17596 );
and ( n26011 , n828 , n26010 );
not ( n26012 , n17597 );
nor ( n26013 , n26011 , n16258 , n26012 );
and ( n26014 , n828 , n16347 );
nand ( n26015 , n17549 , n17552 );
not ( n26016 , n17703 );
and ( n26017 , n26015 , n26016 );
or ( n26018 , n26015 , n26016 );
not ( n26019 , n16265 );
nand ( n26020 , n26018 , n26019 );
nor ( n26021 , n26017 , n26020 );
nor ( n26022 , n26014 , n1828 , n26021 );
nor ( n26023 , n16257 , n26013 , n26022 );
and ( n26024 , n832 , n25672 );
and ( n26025 , n178 , n25723 );
nor ( n26026 , n26024 , n26025 );
or ( n26027 , n26026 , n25752 );
or ( n26028 , n16069 , n25665 );
nand ( n26029 , n26027 , n26028 , n2 );
and ( n26030 , n833 , n25672 );
and ( n26031 , n323 , n25709 );
nor ( n26032 , n26030 , n26031 );
or ( n26033 , n26032 , n25718 );
or ( n26034 , n15973 , n25665 );
nand ( n26035 , n26033 , n26034 , n2 );
or ( n26036 , n16281 , n16746 );
not ( n26037 , n16282 );
nor ( n26038 , n26037 , n16316 );
or ( n26039 , n26038 , n16728 );
and ( n26040 , n26038 , n16728 );
nor ( n26041 , n26040 , n16265 );
nand ( n26042 , n26039 , n26041 );
nand ( n26043 , n26036 , n26042 );
and ( n26044 , n16258 , n26043 );
and ( n26045 , n16358 , n16281 );
not ( n26046 , n16358 );
and ( n26047 , n26046 , n848 );
nor ( n26048 , n26045 , n26047 );
and ( n26049 , n1828 , n26048 );
nor ( n26050 , n26044 , n26049 );
nor ( n26051 , n16257 , n26050 );
not ( n26052 , n25822 );
and ( n26053 , n379 , n25825 );
and ( n26054 , n857 , n25828 );
nor ( n26055 , n26053 , n26054 );
or ( n26056 , n26052 , n26055 );
or ( n26057 , n25833 , n26055 );
and ( n26058 , n561 , n25835 );
not ( n26059 , n25843 );
and ( n26060 , n627 , n26059 );
nor ( n26061 , n26058 , n26060 );
not ( n26062 , n26061 );
and ( n26063 , n1209 , n25841 );
and ( n26064 , n1519 , n25837 );
nor ( n26065 , n26063 , n26064 );
not ( n26066 , n26065 );
or ( n26067 , n26062 , n26066 );
nand ( n26068 , n26067 , n25849 );
nand ( n26069 , n26057 , n26068 );
and ( n26070 , n735 , n25852 );
not ( n26071 , n25855 );
and ( n26072 , n1511 , n26071 );
nor ( n26073 , n26070 , n26072 );
and ( n26074 , n1241 , n23125 );
not ( n26075 , n23604 );
and ( n26076 , n819 , n26075 );
nor ( n26077 , n26074 , n26076 );
and ( n26078 , n26073 , n26077 );
nor ( n26079 , n26078 , n25901 );
and ( n26080 , n475 , n25871 );
not ( n26081 , n23604 );
and ( n26082 , n530 , n26081 );
nor ( n26083 , n26080 , n26082 );
not ( n26084 , n23153 );
and ( n26085 , n1385 , n26084 );
and ( n26086 , n1513 , n25878 );
nor ( n26087 , n26085 , n26086 );
and ( n26088 , n26083 , n26087 );
nor ( n26089 , n26088 , n25883 );
nor ( n26090 , n26069 , n26079 , n26089 );
not ( n26091 , n25888 );
and ( n26092 , n1535 , n26091 );
not ( n26093 , n25873 );
not ( n26094 , n26093 );
and ( n26095 , n708 , n26094 );
nor ( n26096 , n26092 , n26095 );
not ( n26097 , n26096 );
and ( n26098 , n1273 , n25895 );
and ( n26099 , n758 , n25933 );
nor ( n26100 , n26098 , n26099 );
not ( n26101 , n26100 );
or ( n26102 , n26097 , n26101 );
not ( n26103 , n25868 );
nand ( n26104 , n26102 , n26103 );
nand ( n26105 , n26056 , n26090 , n26104 );
and ( n26106 , n384 , n25825 );
and ( n26107 , n1030 , n25828 );
nor ( n26108 , n26106 , n26107 );
or ( n26109 , n26052 , n26108 );
or ( n26110 , n25833 , n26108 );
not ( n26111 , n21580 );
and ( n26112 , n551 , n26111 );
and ( n26113 , n626 , n26059 );
nor ( n26114 , n26112 , n26113 );
not ( n26115 , n26114 );
and ( n26116 , n1159 , n25841 );
and ( n26117 , n1491 , n25837 );
nor ( n26118 , n26116 , n26117 );
not ( n26119 , n26118 );
or ( n26120 , n26115 , n26119 );
nand ( n26121 , n26120 , n25849 );
nand ( n26122 , n26110 , n26121 );
and ( n26123 , n673 , n25852 );
and ( n26124 , n1492 , n26071 );
nor ( n26125 , n26123 , n26124 );
and ( n26126 , n1203 , n23125 );
and ( n26127 , n796 , n26075 );
nor ( n26128 , n26126 , n26127 );
and ( n26129 , n26125 , n26128 );
nor ( n26130 , n26129 , n25901 );
and ( n26131 , n474 , n25871 );
and ( n26132 , n527 , n26081 );
nor ( n26133 , n26131 , n26132 );
not ( n26134 , n23153 );
and ( n26135 , n1381 , n26134 );
and ( n26136 , n1512 , n25878 );
nor ( n26137 , n26135 , n26136 );
and ( n26138 , n26133 , n26137 );
nor ( n26139 , n26138 , n25883 );
nor ( n26140 , n26122 , n26130 , n26139 );
not ( n26141 , n21582 );
and ( n26142 , n656 , n26141 );
and ( n26143 , n709 , n26094 );
nor ( n26144 , n26142 , n26143 );
not ( n26145 , n26144 );
and ( n26146 , n1390 , n25895 );
and ( n26147 , n1503 , n25889 );
nor ( n26148 , n26146 , n26147 );
not ( n26149 , n26148 );
or ( n26150 , n26145 , n26149 );
nand ( n26151 , n26150 , n26103 );
nand ( n26152 , n26109 , n26140 , n26151 );
and ( n26153 , n515 , n14993 );
and ( n26154 , n516 , n25386 );
nor ( n26155 , n26153 , n26154 );
nand ( n26156 , n26155 , n15073 , n25391 );
or ( n26157 , n1250 , n15886 );
or ( n26158 , n19789 , n25380 );
nand ( n26159 , n26157 , n26158 , n15049 );
and ( n26160 , n26156 , n26159 );
or ( n26161 , n15052 , n25391 );
or ( n26162 , n1399 , n15073 );
nand ( n26163 , n26161 , n26162 );
nor ( n26164 , n26160 , n26163 , n15059 );
or ( n26165 , n16656 , n26164 );
nand ( n26166 , n26165 , n17442 );
or ( n26167 , n26166 , n510 , n599 );
nor ( n26168 , n1248 , n1409 , n25380 );
not ( n26169 , n26168 );
nor ( n26170 , n26169 , n1151 , n1364 , n1406 );
nand ( n26171 , n26170 , n25390 , n25359 );
nand ( n26172 , n26167 , n26171 );
and ( n26173 , n613 , n25374 );
and ( n26174 , n609 , n25376 );
nor ( n26175 , n26173 , n26174 );
and ( n26176 , n26175 , n15886 , n25380 );
not ( n26177 , n26156 );
nor ( n26178 , n26176 , n26177 );
or ( n26179 , n15005 , n25358 );
or ( n26180 , n1152 , n15077 );
and ( n26181 , n637 , n25353 );
and ( n26182 , n638 , n25364 );
nor ( n26183 , n26181 , n26182 );
nand ( n26184 , n26183 , n15077 , n25358 );
and ( n26185 , n16674 , n26184 );
not ( n26186 , n15023 );
nor ( n26187 , n26185 , n26186 );
nand ( n26188 , n26179 , n26180 , n26187 );
nand ( n26189 , n26178 , n26188 , n14991 , n26171 );
nand ( n26190 , n26172 , n26189 );
not ( n26191 , n1095 );
not ( n26192 , n21349 );
or ( n26193 , n26191 , n26192 );
nand ( n26194 , n26193 , n20056 );
not ( n26195 , n15606 );
nand ( n26196 , n26194 , n15650 , n26195 );
not ( n26197 , n15601 );
nor ( n26198 , n1113 , n26197 );
and ( n26199 , n26198 , n1174 , n15584 , n15591 );
nor ( n26200 , n21635 , n15647 , n15639 );
or ( n26201 , n26199 , n26200 );
or ( n26202 , n406 , n1095 );
nand ( n26203 , n26201 , n26202 );
and ( n26204 , n26196 , n26203 );
nor ( n26205 , n26204 , n21342 );
and ( n26206 , n399 , n25825 );
and ( n26207 , n1417 , n25958 );
nor ( n26208 , n26206 , n26207 );
or ( n26209 , n26052 , n26208 );
or ( n26210 , n25833 , n26208 );
and ( n26211 , n545 , n25835 );
and ( n26212 , n1540 , n25837 );
nor ( n26213 , n26211 , n26212 );
not ( n26214 , n26213 );
and ( n26215 , n1263 , n25841 );
and ( n26216 , n621 , n25844 );
nor ( n26217 , n26215 , n26216 );
not ( n26218 , n26217 );
or ( n26219 , n26214 , n26218 );
nand ( n26220 , n26219 , n25849 );
nand ( n26221 , n26210 , n26220 );
and ( n26222 , n573 , n25852 );
and ( n26223 , n1509 , n25856 );
nor ( n26224 , n26222 , n26223 );
and ( n26225 , n1382 , n23125 );
and ( n26226 , n703 , n26075 );
nor ( n26227 , n26225 , n26226 );
and ( n26228 , n26224 , n26227 );
nor ( n26229 , n26228 , n25868 );
and ( n26230 , n468 , n25871 );
and ( n26231 , n522 , n26081 );
nor ( n26232 , n26230 , n26231 );
and ( n26233 , n1389 , n26134 );
and ( n26234 , n1518 , n25878 );
nor ( n26235 , n26233 , n26234 );
and ( n26236 , n26232 , n26235 );
nor ( n26237 , n26236 , n25883 );
nor ( n26238 , n26221 , n26229 , n26237 );
and ( n26239 , n727 , n25886 );
and ( n26240 , n1483 , n25889 );
nor ( n26241 , n26239 , n26240 );
not ( n26242 , n26241 );
and ( n26243 , n1245 , n25895 );
and ( n26244 , n812 , n23606 );
nor ( n26245 , n26243 , n26244 );
not ( n26246 , n26245 );
or ( n26247 , n26242 , n26246 );
nand ( n26248 , n26247 , n25902 );
nand ( n26249 , n26209 , n26238 , n26248 );
and ( n26250 , n1455 , n25958 );
not ( n26251 , n401 );
nor ( n26252 , n26251 , n25824 );
nor ( n26253 , n26250 , n26252 );
or ( n26254 , n25823 , n26253 );
or ( n26255 , n25833 , n26253 );
and ( n26256 , n544 , n25835 );
and ( n26257 , n1537 , n25854 );
nor ( n26258 , n26256 , n26257 );
not ( n26259 , n26258 );
and ( n26260 , n1183 , n25974 );
and ( n26261 , n620 , n25844 );
nor ( n26262 , n26260 , n26261 );
not ( n26263 , n26262 );
or ( n26264 , n26259 , n26263 );
nand ( n26265 , n26264 , n25849 );
nand ( n26266 , n26255 , n26265 );
not ( n26267 , n21581 );
and ( n26268 , n652 , n26267 );
and ( n26269 , n1534 , n25856 );
nor ( n26270 , n26268 , n26269 );
and ( n26271 , n1275 , n23125 );
and ( n26272 , n702 , n25860 );
nor ( n26273 , n26271 , n26272 );
and ( n26274 , n26270 , n26273 );
nor ( n26275 , n26274 , n25868 );
and ( n26276 , n467 , n25871 );
and ( n26277 , n1524 , n26071 );
nor ( n26278 , n26276 , n26277 );
not ( n26279 , n23153 );
and ( n26280 , n1155 , n26279 );
and ( n26281 , n559 , n26075 );
nor ( n26282 , n26280 , n26281 );
and ( n26283 , n26278 , n26282 );
nor ( n26284 , n26283 , n25883 );
nor ( n26285 , n26266 , n26275 , n26284 );
and ( n26286 , n726 , n25886 );
not ( n26287 , n25888 );
and ( n26288 , n1479 , n26287 );
nor ( n26289 , n26286 , n26288 );
not ( n26290 , n26289 );
buf ( n26291 , n23125 );
and ( n26292 , n1244 , n26291 );
not ( n26293 , n26093 );
and ( n26294 , n800 , n26293 );
nor ( n26295 , n26292 , n26294 );
not ( n26296 , n26295 );
or ( n26297 , n26290 , n26296 );
nand ( n26298 , n26297 , n25902 );
nand ( n26299 , n26254 , n26285 , n26298 );
nor ( n26300 , n391 , n15633 );
nand ( n26301 , n1148 , n26300 );
and ( n26302 , n15629 , n21349 );
nor ( n26303 , n26302 , n15606 );
nand ( n26304 , n26303 , n20056 , n15650 );
and ( n26305 , n26301 , n26304 );
nor ( n26306 , n26305 , n21342 );
and ( n26307 , n1454 , n25958 );
not ( n26308 , n400 );
nor ( n26309 , n26308 , n25824 );
nor ( n26310 , n26307 , n26309 );
or ( n26311 , n25823 , n26310 );
or ( n26312 , n25833 , n26310 );
and ( n26313 , n743 , n25835 );
and ( n26314 , n619 , n25844 );
nor ( n26315 , n26313 , n26314 );
not ( n26316 , n26315 );
and ( n26317 , n1262 , n25974 );
and ( n26318 , n1531 , n25854 );
nor ( n26319 , n26317 , n26318 );
not ( n26320 , n26319 );
or ( n26321 , n26316 , n26320 );
nand ( n26322 , n26321 , n25849 );
nand ( n26323 , n26312 , n26322 );
and ( n26324 , n725 , n26267 );
and ( n26325 , n811 , n25860 );
nor ( n26326 , n26324 , n26325 );
and ( n26327 , n1180 , n23125 );
and ( n26328 , n1484 , n25856 );
nor ( n26329 , n26327 , n26328 );
and ( n26330 , n26326 , n26329 );
nor ( n26331 , n26330 , n25901 );
and ( n26332 , n647 , n25871 );
and ( n26333 , n1516 , n26071 );
nor ( n26334 , n26332 , n26333 );
and ( n26335 , n1154 , n26279 );
and ( n26336 , n521 , n26075 );
nor ( n26337 , n26335 , n26336 );
and ( n26338 , n26334 , n26337 );
nor ( n26339 , n26338 , n25883 );
nor ( n26340 , n26323 , n26331 , n26339 );
and ( n26341 , n651 , n25886 );
and ( n26342 , n672 , n26293 );
nor ( n26343 , n26341 , n26342 );
not ( n26344 , n26343 );
and ( n26345 , n1384 , n26291 );
and ( n26346 , n1507 , n26091 );
nor ( n26347 , n26345 , n26346 );
not ( n26348 , n26347 );
or ( n26349 , n26344 , n26348 );
nand ( n26350 , n26349 , n26103 );
nand ( n26351 , n26311 , n26340 , n26350 );
not ( n26352 , n20185 );
not ( n26353 , n20182 );
or ( n26354 , n26352 , n26353 );
nand ( n26355 , n26354 , n20187 );
not ( n26356 , n20168 );
or ( n26357 , n26356 , n20194 );
and ( n26358 , n1219 , n23641 );
nand ( n26359 , n26357 , n26358 );
and ( n26360 , n26355 , n26359 );
not ( n26361 , n2 );
nor ( n26362 , n26360 , n26361 );
or ( n26363 , n20182 , n20184 );
not ( n26364 , n20186 );
nand ( n26365 , n26363 , n26364 );
and ( n26366 , n26365 , n23642 );
not ( n26367 , n2 );
and ( n26368 , n20184 , n26364 );
nor ( n26369 , n26368 , n1220 );
nor ( n26370 , n26366 , n26367 , n26369 );
and ( n26371 , n398 , n25825 );
and ( n26372 , n1453 , n25958 );
nor ( n26373 , n26371 , n26372 );
or ( n26374 , n26052 , n26373 );
or ( n26375 , n25833 , n26373 );
and ( n26376 , n543 , n26111 );
and ( n26377 , n618 , n26059 );
nor ( n26378 , n26376 , n26377 );
not ( n26379 , n26378 );
and ( n26380 , n1207 , n25841 );
and ( n26381 , n1523 , n25837 );
nor ( n26382 , n26380 , n26381 );
not ( n26383 , n26382 );
or ( n26384 , n26379 , n26383 );
nand ( n26385 , n26384 , n25849 );
nand ( n26386 , n26375 , n26385 );
and ( n26387 , n724 , n25852 );
and ( n26388 , n1486 , n26071 );
nor ( n26389 , n26387 , n26388 );
and ( n26390 , n1243 , n23125 );
and ( n26391 , n810 , n26075 );
nor ( n26392 , n26390 , n26391 );
and ( n26393 , n26389 , n26392 );
nor ( n26394 , n26393 , n25901 );
and ( n26395 , n646 , n25871 );
and ( n26396 , n520 , n26081 );
nor ( n26397 , n26395 , n26396 );
and ( n26398 , n1153 , n26134 );
and ( n26399 , n1526 , n25878 );
nor ( n26400 , n26398 , n26399 );
and ( n26401 , n26397 , n26400 );
nor ( n26402 , n26401 , n25883 );
nor ( n26403 , n26386 , n26394 , n26402 );
and ( n26404 , n650 , n26141 );
and ( n26405 , n701 , n26094 );
nor ( n26406 , n26404 , n26405 );
not ( n26407 , n26406 );
and ( n26408 , n1274 , n25895 );
and ( n26409 , n1506 , n25889 );
nor ( n26410 , n26408 , n26409 );
not ( n26411 , n26410 );
or ( n26412 , n26407 , n26411 );
nand ( n26413 , n26412 , n26103 );
nand ( n26414 , n26374 , n26403 , n26413 );
nand ( n26415 , n1066 , n24271 );
not ( n26416 , n26415 );
nand ( n26417 , n20043 , n19376 , n26416 , n20052 );
or ( n26418 , n20056 , n24279 );
nand ( n26419 , n26418 , n26415 );
nand ( n26420 , n26419 , n20043 , n20058 );
and ( n26421 , n26417 , n26420 );
nor ( n26422 , n26421 , n21342 );
not ( n26423 , n13633 );
not ( n26424 , n19960 );
and ( n26425 , n26423 , n26424 );
nor ( n26426 , n371 , n19960 );
nor ( n26427 , n26425 , n26426 );
not ( n26428 , n888 );
not ( n26429 , n19963 );
or ( n26430 , n26428 , n26429 );
nand ( n26431 , n14549 , n19963 );
nand ( n26432 , n26430 , n26431 );
not ( n26433 , n26432 );
nor ( n26434 , n26427 , n26433 );
not ( n26435 , n26434 );
or ( n26436 , n19941 , n26433 );
not ( n26437 , n26431 );
nand ( n26438 , n888 , n26437 );
nand ( n26439 , n26436 , n26438 );
not ( n26440 , n26439 );
nand ( n26441 , n938 , n26426 , n26432 );
nand ( n26442 , n26440 , n19949 , n26441 );
not ( n26443 , n26442 );
and ( n26444 , n26435 , n26443 );
not ( n26445 , n19973 );
nand ( n26446 , n26445 , n12640 );
or ( n26447 , n18835 , n26446 );
nand ( n26448 , n26447 , n19934 );
not ( n26449 , n19973 );
nand ( n26450 , n26449 , n884 );
and ( n26451 , n26450 , n26446 );
nor ( n26452 , n368 , n19969 );
and ( n26453 , n935 , n26452 );
not ( n26454 , n19927 );
nor ( n26455 , n26453 , n26454 );
nor ( n26456 , n26451 , n26455 );
nor ( n26457 , n26448 , n26456 , n26442 );
nor ( n26458 , n26444 , n26457 );
not ( n26459 , n2 );
not ( n26460 , n25251 );
and ( n26461 , n52 , n26460 );
and ( n26462 , n1420 , n25252 );
nor ( n26463 , n26461 , n26462 );
nor ( n26464 , n26459 , n26463 );
not ( n26465 , n2 );
and ( n26466 , n33 , n26460 );
and ( n26467 , n1417 , n25252 );
nor ( n26468 , n26466 , n26467 );
nor ( n26469 , n26465 , n26468 );
and ( n26470 , n671 , n26141 );
not ( n26471 , n21741 );
and ( n26472 , n1485 , n26471 );
nor ( n26473 , n26470 , n26472 );
buf ( n26474 , n25894 );
and ( n26475 , n1143 , n26474 );
and ( n26476 , n833 , n23606 );
nor ( n26477 , n26475 , n26476 );
and ( n26478 , n26473 , n26477 );
nor ( n26479 , n26478 , n25901 );
not ( n26480 , n21582 );
and ( n26481 , n745 , n26480 );
and ( n26482 , n1481 , n26471 );
nor ( n26483 , n26481 , n26482 );
and ( n26484 , n1071 , n26474 );
not ( n26485 , n25938 );
and ( n26486 , n630 , n26485 );
nor ( n26487 , n26484 , n26486 );
and ( n26488 , n26483 , n26487 );
nor ( n26489 , n26488 , n25990 );
nor ( n26490 , n26479 , n26489 );
and ( n26491 , n25825 , n25956 );
and ( n26492 , n282 , n26491 );
not ( n26493 , n25969 );
and ( n26494 , n657 , n26493 );
not ( n26495 , n25843 );
not ( n26496 , n26495 );
not ( n26497 , n26496 );
and ( n26498 , n710 , n26497 );
nor ( n26499 , n26494 , n26498 );
and ( n26500 , n1102 , n25975 );
not ( n26501 , n21741 );
and ( n26502 , n1505 , n26501 );
nor ( n26503 , n26500 , n26502 );
and ( n26504 , n26499 , n26503 );
nor ( n26505 , n26504 , n25868 );
and ( n26506 , n648 , n25970 );
not ( n26507 , n21741 );
and ( n26508 , n1515 , n26507 );
nor ( n26509 , n26506 , n26508 );
and ( n26510 , n1005 , n25975 );
not ( n26511 , n22153 );
and ( n26512 , n506 , n26511 );
nor ( n26513 , n26510 , n26512 );
and ( n26514 , n26509 , n26513 );
nor ( n26515 , n26514 , n25883 );
nor ( n26516 , n26492 , n26505 , n26515 );
nand ( n26517 , n26490 , n26516 );
not ( n26518 , n2 );
and ( n26519 , n29 , n26460 );
and ( n26520 , n1468 , n25252 );
nor ( n26521 , n26519 , n26520 );
nor ( n26522 , n26518 , n26521 );
or ( n26523 , n20606 , n15379 , n19401 );
nand ( n26524 , n26523 , n19405 );
not ( n26525 , n176 );
nor ( n26526 , n1678 , n26525 , n74 );
not ( n26527 , n12835 );
nand ( n26528 , n1821 , n26527 );
nor ( n26529 , n1821 , n14794 );
not ( n26530 , n26529 );
nand ( n26531 , n26528 , n26530 );
nor ( n26532 , n1796 , n26526 , n222 , n26531 );
not ( n26533 , n12839 );
nor ( n26534 , n26533 , n26527 , n14805 , n12846 );
and ( n26535 , n26532 , n26534 );
not ( n26536 , n2 );
nor ( n26537 , n26535 , n26536 );
not ( n26538 , n12920 );
nand ( n26539 , n14628 , n26538 );
and ( n26540 , n14661 , n26539 );
not ( n26541 , n2 );
nor ( n26542 , n26540 , n26541 );
nand ( n26543 , n371 , n20636 );
not ( n26544 , n20640 );
nor ( n26545 , n19937 , n26544 );
or ( n26546 , n371 , n26545 );
and ( n26547 , n371 , n26545 );
not ( n26548 , n20633 );
nor ( n26549 , n26547 , n26548 );
nand ( n26550 , n26546 , n26549 );
and ( n26551 , n26543 , n26550 );
nor ( n26552 , n26551 , n20652 );
not ( n26553 , n2 );
and ( n26554 , n28 , n26460 );
and ( n26555 , n1459 , n25252 );
nor ( n26556 , n26554 , n26555 );
nor ( n26557 , n26553 , n26556 );
not ( n26558 , n2 );
and ( n26559 , n30 , n26460 );
and ( n26560 , n1458 , n25252 );
nor ( n26561 , n26559 , n26560 );
nor ( n26562 , n26558 , n26561 );
not ( n26563 , n2 );
and ( n26564 , n35 , n26460 );
and ( n26565 , n1454 , n25252 );
nor ( n26566 , n26564 , n26565 );
nor ( n26567 , n26563 , n26566 );
or ( n26568 , n15754 , n15710 );
not ( n26569 , n15753 );
nand ( n26570 , n15755 , n17168 );
or ( n26571 , n26569 , n26570 );
and ( n26572 , n26569 , n26570 );
not ( n26573 , n15709 );
nor ( n26574 , n26572 , n26573 );
nand ( n26575 , n26571 , n26574 );
nand ( n26576 , n26568 , n26575 );
and ( n26577 , n15704 , n26576 );
or ( n26578 , n15752 , n747 );
or ( n26579 , n15754 , n635 );
nand ( n26580 , n26578 , n26579 );
and ( n26581 , n1808 , n26580 );
nor ( n26582 , n26577 , n26581 );
nor ( n26583 , n15703 , n26582 );
nand ( n26584 , n763 , n18895 );
nor ( n26585 , n26584 , n806 , n1530 );
not ( n26586 , n26585 );
nand ( n26587 , n18683 , n15245 , n748 , n18686 );
nand ( n26588 , n26586 , n2 , n26587 );
and ( n26589 , n755 , n26480 );
and ( n26590 , n243 , n26471 );
nor ( n26591 , n26589 , n26590 );
and ( n26592 , n1161 , n26474 );
and ( n26593 , n711 , n26485 );
nor ( n26594 , n26592 , n26593 );
and ( n26595 , n26591 , n26594 );
nor ( n26596 , n26595 , n25868 );
and ( n26597 , n564 , n26480 );
and ( n26598 , n245 , n26471 );
nor ( n26599 , n26597 , n26598 );
and ( n26600 , n1151 , n26474 );
not ( n26601 , n25938 );
and ( n26602 , n531 , n26601 );
nor ( n26603 , n26600 , n26602 );
and ( n26604 , n26599 , n26603 );
nor ( n26605 , n26604 , n25883 );
nor ( n26606 , n26596 , n26605 );
and ( n26607 , n562 , n25825 );
and ( n26608 , n1418 , n25958 );
nor ( n26609 , n26607 , n26608 );
and ( n26610 , n1811 , n25961 );
and ( n26611 , n1634 , n25828 );
nor ( n26612 , n26610 , n26611 );
nor ( n26613 , n15952 , n23124 );
and ( n26614 , n1586 , n26613 );
and ( n26615 , n1225 , n23524 );
nor ( n26616 , n26614 , n26615 );
and ( n26617 , n26609 , n26612 , n26616 );
not ( n26618 , n25956 );
nor ( n26619 , n26617 , n26618 );
and ( n26620 , n736 , n26493 );
not ( n26621 , n21741 );
and ( n26622 , n244 , n26621 );
nor ( n26623 , n26620 , n26622 );
buf ( n26624 , n25894 );
and ( n26625 , n1234 , n26624 );
not ( n26626 , n26496 );
and ( n26627 , n821 , n26626 );
nor ( n26628 , n26625 , n26627 );
and ( n26629 , n26623 , n26628 );
nor ( n26630 , n26629 , n25901 );
not ( n26631 , n25870 );
not ( n26632 , n26631 );
not ( n26633 , n26632 );
and ( n26634 , n663 , n26633 );
not ( n26635 , n22153 );
and ( n26636 , n628 , n26635 );
nor ( n26637 , n26634 , n26636 );
and ( n26638 , n1156 , n25975 );
and ( n26639 , n247 , n21742 );
nor ( n26640 , n26638 , n26639 );
and ( n26641 , n26637 , n26640 );
nor ( n26642 , n26641 , n25990 );
nor ( n26643 , n26619 , n26630 , n26642 );
nand ( n26644 , n26606 , n26643 );
and ( n26645 , n466 , n26480 );
and ( n26646 , n744 , n26471 );
nor ( n26647 , n26645 , n26646 );
and ( n26648 , n1364 , n26474 );
and ( n26649 , n518 , n26601 );
nor ( n26650 , n26648 , n26649 );
nand ( n26651 , n26647 , n26650 );
and ( n26652 , n25882 , n26651 );
and ( n26653 , n722 , n25933 );
and ( n26654 , n799 , n25939 );
nor ( n26655 , n26653 , n26654 );
and ( n26656 , n1366 , n26474 );
and ( n26657 , n664 , n26471 );
nor ( n26658 , n26656 , n26657 );
and ( n26659 , n26655 , n26658 );
nor ( n26660 , n26659 , n25901 );
nor ( n26661 , n26652 , n26660 );
and ( n26662 , n598 , n25825 );
and ( n26663 , n1420 , n25958 );
nor ( n26664 , n26662 , n26663 );
and ( n26665 , n1816 , n25961 );
and ( n26666 , n1632 , n25828 );
nor ( n26667 , n26665 , n26666 );
and ( n26668 , n1167 , n26613 );
and ( n26669 , n1223 , n23524 );
nor ( n26670 , n26668 , n26669 );
and ( n26671 , n26664 , n26667 , n26670 );
nor ( n26672 , n26671 , n26618 );
and ( n26673 , n649 , n26493 );
and ( n26674 , n721 , n26621 );
nor ( n26675 , n26673 , n26674 );
and ( n26676 , n1160 , n26624 );
and ( n26677 , n699 , n26626 );
nor ( n26678 , n26676 , n26677 );
and ( n26679 , n26675 , n26678 );
nor ( n26680 , n26679 , n25868 );
and ( n26681 , n741 , n26633 );
not ( n26682 , n21741 );
and ( n26683 , n746 , n26682 );
nor ( n26684 , n26681 , n26683 );
and ( n26685 , n1255 , n25975 );
and ( n26686 , n616 , n26497 );
nor ( n26687 , n26685 , n26686 );
and ( n26688 , n26684 , n26687 );
nor ( n26689 , n26688 , n25990 );
nor ( n26690 , n26672 , n26680 , n26689 );
nand ( n26691 , n26661 , n26690 );
nand ( n26692 , n1828 , n16283 );
or ( n26693 , n826 , n20841 );
not ( n26694 , n16284 );
and ( n26695 , n1234 , n16266 );
nor ( n26696 , n26695 , n16283 );
or ( n26697 , n26694 , n26696 );
nand ( n26698 , n26693 , n26697 , n16258 );
and ( n26699 , n26692 , n26698 );
nor ( n26700 , n26699 , n16257 );
and ( n26701 , n827 , n829 );
nor ( n26702 , n26701 , n16258 , n17596 );
and ( n26703 , n827 , n16747 );
not ( n26704 , n17554 );
nand ( n26705 , n17546 , n26704 );
and ( n26706 , n17553 , n26705 );
or ( n26707 , n17553 , n26705 );
nand ( n26708 , n26707 , n16266 );
nor ( n26709 , n26706 , n26708 );
nor ( n26710 , n26703 , n1828 , n26709 );
nor ( n26711 , n16257 , n26702 , n26710 );
or ( n26712 , n16285 , n16746 );
nand ( n26713 , n16286 , n16727 );
or ( n26714 , n26694 , n26713 );
and ( n26715 , n26694 , n26713 );
nor ( n26716 , n26715 , n16265 );
nand ( n26717 , n26714 , n26716 );
nand ( n26718 , n26712 , n26717 );
and ( n26719 , n16258 , n26718 );
or ( n26720 , n16283 , n847 );
or ( n26721 , n16285 , n826 );
nand ( n26722 , n26720 , n26721 );
and ( n26723 , n1828 , n26722 );
nor ( n26724 , n26719 , n26723 );
nor ( n26725 , n16257 , n26724 );
and ( n26726 , n1164 , n26091 );
and ( n26727 , n704 , n26601 );
nor ( n26728 , n26726 , n26727 );
and ( n26729 , n1400 , n26474 );
and ( n26730 , n658 , n25933 );
nor ( n26731 , n26729 , n26730 );
and ( n26732 , n26728 , n26731 );
nor ( n26733 , n26732 , n25868 );
and ( n26734 , n1120 , n26091 );
and ( n26735 , n523 , n26601 );
nor ( n26736 , n26734 , n26735 );
and ( n26737 , n1409 , n26474 );
not ( n26738 , n25944 );
and ( n26739 , n469 , n26738 );
nor ( n26740 , n26737 , n26739 );
and ( n26741 , n26736 , n26740 );
nor ( n26742 , n26741 , n25883 );
nor ( n26743 , n26733 , n26742 );
and ( n26744 , n603 , n25825 );
and ( n26745 , n1448 , n25958 );
nor ( n26746 , n26744 , n26745 );
and ( n26747 , n1813 , n25961 );
and ( n26748 , n1616 , n25828 );
nor ( n26749 , n26747 , n26748 );
and ( n26750 , n1608 , n26613 );
and ( n26751 , n1224 , n23524 );
nor ( n26752 , n26750 , n26751 );
and ( n26753 , n26746 , n26749 , n26752 );
nor ( n26754 , n26753 , n26618 );
and ( n26755 , n728 , n26493 );
and ( n26756 , n1294 , n26621 );
nor ( n26757 , n26755 , n26756 );
and ( n26758 , n1233 , n26624 );
and ( n26759 , n813 , n26626 );
nor ( n26760 , n26758 , n26759 );
and ( n26761 , n26757 , n26760 );
nor ( n26762 , n26761 , n25901 );
and ( n26763 , n546 , n26633 );
not ( n26764 , n26496 );
and ( n26765 , n569 , n26764 );
nor ( n26766 , n26763 , n26765 );
and ( n26767 , n1221 , n25975 );
and ( n26768 , n1166 , n21742 );
nor ( n26769 , n26767 , n26768 );
and ( n26770 , n26766 , n26769 );
nor ( n26771 , n26770 , n25990 );
nor ( n26772 , n26754 , n26762 , n26771 );
nand ( n26773 , n26743 , n26772 );
and ( n26774 , n660 , n25886 );
and ( n26775 , n1099 , n26287 );
nor ( n26776 , n26774 , n26775 );
and ( n26777 , n1471 , n26291 );
and ( n26778 , n666 , n26293 );
nor ( n26779 , n26777 , n26778 );
and ( n26780 , n26776 , n26779 );
nor ( n26781 , n26780 , n25868 );
and ( n26782 , n477 , n26141 );
not ( n26783 , n25888 );
and ( n26784 , n1087 , n26783 );
nor ( n26785 , n26782 , n26784 );
and ( n26786 , n1406 , n25895 );
and ( n26787 , n489 , n23606 );
nor ( n26788 , n26786 , n26787 );
and ( n26789 , n26785 , n26788 );
nor ( n26790 , n26789 , n25883 );
nor ( n26791 , n26781 , n26790 );
nand ( n26792 , n604 , n25825 );
nand ( n26793 , n1449 , n25958 );
and ( n26794 , n1829 , n25961 );
and ( n26795 , n1633 , n25828 );
nor ( n26796 , n26794 , n26795 );
and ( n26797 , n1860 , n26613 );
and ( n26798 , n1198 , n23524 );
nor ( n26799 , n26797 , n26798 );
nand ( n26800 , n26792 , n26793 , n26796 , n26799 );
and ( n26801 , n25956 , n26800 );
not ( n26802 , n25944 );
and ( n26803 , n738 , n26802 );
and ( n26804 , n1086 , n21742 );
nor ( n26805 , n26803 , n26804 );
and ( n26806 , n1467 , n25895 );
and ( n26807 , n832 , n25947 );
nor ( n26808 , n26806 , n26807 );
and ( n26809 , n26805 , n26808 );
nor ( n26810 , n26809 , n25901 );
not ( n26811 , n26632 );
and ( n26812 , n554 , n26811 );
and ( n26813 , n1088 , n26682 );
nor ( n26814 , n26812 , n26813 );
and ( n26815 , n1439 , n25975 );
and ( n26816 , n631 , n26764 );
nor ( n26817 , n26815 , n26816 );
and ( n26818 , n26814 , n26817 );
nor ( n26819 , n26818 , n25990 );
nor ( n26820 , n26801 , n26810 , n26819 );
nand ( n26821 , n26791 , n26820 );
not ( n26822 , n21637 );
and ( n26823 , n1104 , n1095 , n26822 );
not ( n26824 , n21625 );
not ( n26825 , n21629 );
nand ( n26826 , n1150 , n26824 , n26825 );
nor ( n26827 , n26826 , n1045 , n21658 );
nor ( n26828 , n26823 , n26827 );
and ( n26829 , n15594 , n15580 );
nand ( n26830 , n20044 , n21657 );
nor ( n26831 , n1150 , n26830 );
nand ( n26832 , n19389 , n26829 , n26831 );
nor ( n26833 , n1100 , n15674 , n26832 );
and ( n26834 , n26833 , n21517 , n15599 );
nor ( n26835 , n26834 , n21643 );
or ( n26836 , n1150 , n19389 , n21658 );
not ( n26837 , n21533 );
nand ( n26838 , n26837 , n21632 );
or ( n26839 , n26838 , n1066 , n1083 );
nand ( n26840 , n26836 , n26839 );
nand ( n26841 , n21628 , n21654 , n15585 , n26840 );
nand ( n26842 , n26841 , n1104 , n26822 );
nand ( n26843 , n26828 , n26835 , n26842 );
not ( n26844 , n405 );
nand ( n26845 , n26844 , n1124 , n21529 );
and ( n26846 , n15639 , n26845 );
nor ( n26847 , n1124 , n15647 );
nor ( n26848 , n26846 , n21342 , n26847 );
nor ( n26849 , n16505 , n20618 );
nand ( n26850 , n928 , n21679 , n24423 );
not ( n26851 , n21446 );
or ( n26852 , n26850 , n900 , n26851 );
and ( n26853 , n21675 , n21428 );
nor ( n26854 , n26853 , n21446 );
nor ( n26855 , n24410 , n929 , n26854 );
not ( n26856 , n930 );
and ( n26857 , n26855 , n928 , n26856 );
nand ( n26858 , n17121 , n17122 );
nor ( n26859 , n24409 , n26858 );
nor ( n26860 , n26857 , n26859 );
nand ( n26861 , n26852 , n26860 );
nor ( n26862 , n1799 , n24271 );
nor ( n26863 , n1799 , n21532 , n19377 );
or ( n26864 , n26862 , n26863 );
nand ( n26865 , n26864 , n20052 );
nor ( n26866 , n1799 , n21532 , n20057 );
or ( n26867 , n26862 , n26866 );
nand ( n26868 , n26867 , n20058 );
and ( n26869 , n26865 , n26868 );
nor ( n26870 , n26869 , n21342 );
nor ( n26871 , n16505 , n24438 );
and ( n26872 , n567 , n21583 );
and ( n26873 , n1489 , n26474 );
and ( n26874 , n525 , n26485 );
nor ( n26875 , n26872 , n26873 , n26874 );
or ( n26876 , n25883 , n26875 );
not ( n26877 , n25902 );
not ( n26878 , n26493 );
not ( n26879 , n26878 );
and ( n26880 , n733 , n26879 );
and ( n26881 , n1490 , n26474 );
and ( n26882 , n815 , n26485 );
nor ( n26883 , n26880 , n26881 , n26882 );
or ( n26884 , n26877 , n26883 );
nand ( n26885 , n402 , n25825 );
and ( n26886 , n1458 , n25958 );
and ( n26887 , n265 , n25828 );
nor ( n26888 , n26886 , n26887 );
and ( n26889 , n26885 , n26888 );
or ( n26890 , n25821 , n26889 );
not ( n26891 , n25893 );
and ( n26892 , n1498 , n26891 );
not ( n26893 , n25870 );
and ( n26894 , n665 , n26893 );
and ( n26895 , n624 , n22152 );
nor ( n26896 , n26892 , n26894 , n26895 );
or ( n26897 , n25990 , n26896 );
nand ( n26898 , n26890 , n26897 );
or ( n26899 , n25833 , n26889 );
not ( n26900 , n25893 );
and ( n26901 , n1542 , n26900 );
not ( n26902 , n25870 );
and ( n26903 , n654 , n26902 );
and ( n26904 , n705 , n22152 );
nor ( n26905 , n26901 , n26903 , n26904 );
or ( n26906 , n25868 , n26905 );
nand ( n26907 , n26899 , n26906 );
nor ( n26908 , n26898 , n26907 );
nand ( n26909 , n26876 , n26884 , n26908 );
and ( n26910 , n472 , n21583 );
and ( n26911 , n1313 , n26474 );
and ( n26912 , n528 , n26485 );
nor ( n26913 , n26910 , n26911 , n26912 );
or ( n26914 , n25883 , n26913 );
not ( n26915 , n23154 );
and ( n26916 , n1335 , n26915 );
and ( n26917 , n549 , n26480 );
and ( n26918 , n575 , n26094 );
nor ( n26919 , n26916 , n26917 , n26918 );
or ( n26920 , n25990 , n26919 );
nand ( n26921 , n381 , n25825 );
and ( n26922 , n1468 , n25958 );
and ( n26923 , n915 , n25828 );
nor ( n26924 , n26922 , n26923 );
and ( n26925 , n26921 , n26924 );
or ( n26926 , n25821 , n26925 );
and ( n26927 , n1354 , n26891 );
and ( n26928 , n786 , n26893 );
and ( n26929 , n706 , n22152 );
nor ( n26930 , n26927 , n26928 , n26929 );
or ( n26931 , n25868 , n26930 );
nand ( n26932 , n26926 , n26931 );
or ( n26933 , n25833 , n26925 );
and ( n26934 , n1293 , n26900 );
and ( n26935 , n731 , n26902 );
and ( n26936 , n816 , n22152 );
nor ( n26937 , n26934 , n26935 , n26936 );
or ( n26938 , n25901 , n26937 );
nand ( n26939 , n26933 , n26938 );
nor ( n26940 , n26932 , n26939 );
nand ( n26941 , n26914 , n26920 , n26940 );
and ( n26942 , n453 , n26879 );
and ( n26943 , n1403 , n25895 );
and ( n26944 , n459 , n26293 );
nor ( n26945 , n26942 , n26943 , n26944 );
or ( n26946 , n25883 , n26945 );
and ( n26947 , n687 , n26879 );
and ( n26948 , n1210 , n25895 );
and ( n26949 , n753 , n26293 );
nor ( n26950 , n26947 , n26948 , n26949 );
or ( n26951 , n26877 , n26950 );
nand ( n26952 , n1814 , n25961 );
and ( n26953 , n596 , n25825 );
and ( n26954 , n1452 , n25958 );
nor ( n26955 , n26953 , n26954 );
and ( n26956 , n26952 , n26955 );
or ( n26957 , n25821 , n26956 );
and ( n26958 , n1259 , n23125 );
and ( n26959 , n500 , n26631 );
and ( n26960 , n504 , n26495 );
nor ( n26961 , n26958 , n26959 , n26960 );
or ( n26962 , n25990 , n26961 );
nand ( n26963 , n26957 , n26962 );
or ( n26964 , n25833 , n26956 );
and ( n26965 , n1271 , n23125 );
not ( n26966 , n25870 );
and ( n26967 , n588 , n26966 );
not ( n26968 , n23604 );
and ( n26969 , n593 , n26968 );
nor ( n26970 , n26965 , n26967 , n26969 );
or ( n26971 , n25868 , n26970 );
nand ( n26972 , n26964 , n26971 );
nor ( n26973 , n26963 , n26972 );
nand ( n26974 , n26946 , n26951 , n26973 );
and ( n26975 , n372 , n18815 );
and ( n26976 , n888 , n14549 );
or ( n26977 , n14543 , n938 );
or ( n26978 , n13633 , n371 );
nand ( n26979 , n26977 , n26978 , n19941 );
nor ( n26980 , n26975 , n26976 , n26979 );
not ( n26981 , n19982 );
nor ( n26982 , n19981 , n988 );
nor ( n26983 , n19960 , n26981 , n26982 );
and ( n26984 , n26980 , n26983 , n19949 , n19963 );
and ( n26985 , n350 , n18835 );
and ( n26986 , n884 , n12640 );
or ( n26987 , n14591 , n935 );
or ( n26988 , n13660 , n368 );
and ( n26989 , n366 , n19984 );
not ( n26990 , n366 );
and ( n26991 , n26990 , n879 );
nor ( n26992 , n26989 , n26991 );
nand ( n26993 , n26987 , n26988 , n26992 );
nor ( n26994 , n26985 , n26986 , n26993 );
and ( n26995 , n14593 , n13664 );
and ( n26996 , n367 , n933 );
nor ( n26997 , n26995 , n26996 );
not ( n26998 , n19934 );
nor ( n26999 , n26997 , n26998 , n19973 );
not ( n27000 , n19969 );
and ( n27001 , n26994 , n26999 , n19927 , n27000 );
and ( n27002 , n26984 , n27001 );
not ( n27003 , n13746 );
nor ( n27004 , n27002 , n16554 , n27003 );
and ( n27005 , n587 , n26738 );
and ( n27006 , n1033 , n21742 );
nor ( n27007 , n27005 , n27006 );
and ( n27008 , n1152 , n25895 );
and ( n27009 , n457 , n25947 );
nor ( n27010 , n27008 , n27009 );
nand ( n27011 , n27007 , n27010 );
and ( n27012 , n25882 , n27011 );
and ( n27013 , n686 , n26802 );
and ( n27014 , n770 , n26626 );
nor ( n27015 , n27013 , n27014 );
and ( n27016 , n1235 , n25895 );
and ( n27017 , n1021 , n21742 );
nor ( n27018 , n27016 , n27017 );
and ( n27019 , n27015 , n27018 );
nor ( n27020 , n27019 , n25901 );
nor ( n27021 , n27012 , n27020 );
and ( n27022 , n1419 , n25958 );
and ( n27023 , n1226 , n23524 );
nor ( n27024 , n27022 , n27023 );
and ( n27025 , n605 , n25825 );
and ( n27026 , n1871 , n26613 );
and ( n27027 , n1815 , n25961 );
nor ( n27028 , n27025 , n27026 , n27027 );
and ( n27029 , n27024 , n27028 );
nor ( n27030 , n27029 , n26618 );
and ( n27031 , n688 , n25970 );
and ( n27032 , n1020 , n26507 );
nor ( n27033 , n27031 , n27032 );
and ( n27034 , n1258 , n25975 );
and ( n27035 , n503 , n26511 );
nor ( n27036 , n27034 , n27035 );
and ( n27037 , n27033 , n27036 );
nor ( n27038 , n27037 , n25990 );
not ( n27039 , n25969 );
and ( n27040 , n761 , n27039 );
and ( n27041 , n591 , n25873 );
nor ( n27042 , n27040 , n27041 );
and ( n27043 , n1270 , n23125 );
and ( n27044 , n1032 , n26507 );
nor ( n27045 , n27043 , n27044 );
and ( n27046 , n27042 , n27045 );
nor ( n27047 , n27046 , n25868 );
nor ( n27048 , n27030 , n27038 , n27047 );
nand ( n27049 , n27021 , n27048 );
not ( n27050 , n2 );
and ( n27051 , n44 , n26460 );
and ( n27052 , n1416 , n25252 );
nor ( n27053 , n27051 , n27052 );
nor ( n27054 , n27050 , n27053 );
not ( n27055 , n2 );
and ( n27056 , n48 , n26460 );
and ( n27057 , n1419 , n25252 );
nor ( n27058 , n27056 , n27057 );
nor ( n27059 , n27055 , n27058 );
not ( n27060 , n2 );
and ( n27061 , n50 , n26460 );
and ( n27062 , n1418 , n25252 );
nor ( n27063 , n27061 , n27062 );
nor ( n27064 , n27060 , n27063 );
and ( n27065 , n380 , n25825 );
and ( n27066 , n1456 , n25958 );
and ( n27067 , n773 , n25828 );
nor ( n27068 , n27065 , n27066 , n27067 );
or ( n27069 , n26618 , n27068 );
and ( n27070 , n470 , n26811 );
and ( n27071 , n1517 , n25977 );
nor ( n27072 , n27070 , n27071 );
and ( n27073 , n1252 , n25975 );
and ( n27074 , n524 , n26635 );
nor ( n27075 , n27073 , n27074 );
nand ( n27076 , n27072 , n27075 );
and ( n27077 , n25882 , n27076 );
and ( n27078 , n653 , n25970 );
and ( n27079 , n667 , n22154 );
nor ( n27080 , n27078 , n27079 );
and ( n27081 , n1277 , n25975 );
and ( n27082 , n1508 , n25977 );
nor ( n27083 , n27081 , n27082 );
and ( n27084 , n27080 , n27083 );
nor ( n27085 , n27084 , n25868 );
nor ( n27086 , n27077 , n27085 );
not ( n27087 , n26632 );
and ( n27088 , n729 , n27087 );
and ( n27089 , n814 , n26764 );
nor ( n27090 , n27088 , n27089 );
and ( n27091 , n1246 , n25975 );
and ( n27092 , n1480 , n26621 );
nor ( n27093 , n27091 , n27092 );
and ( n27094 , n27090 , n27093 );
nor ( n27095 , n27094 , n25901 );
and ( n27096 , n547 , n26811 );
and ( n27097 , n622 , n26511 );
nor ( n27098 , n27096 , n27097 );
and ( n27099 , n1264 , n25975 );
and ( n27100 , n1520 , n26682 );
nor ( n27101 , n27099 , n27100 );
and ( n27102 , n27098 , n27101 );
nor ( n27103 , n27102 , n25990 );
nor ( n27104 , n27095 , n27103 );
nand ( n27105 , n27069 , n27086 , n27104 );
and ( n27106 , n392 , n25825 );
and ( n27107 , n1457 , n25958 );
and ( n27108 , n1116 , n25828 );
nor ( n27109 , n27106 , n27107 , n27108 );
or ( n27110 , n26618 , n27109 );
and ( n27111 , n675 , n27087 );
and ( n27112 , n797 , n26764 );
nor ( n27113 , n27111 , n27112 );
and ( n27114 , n1199 , n25975 );
and ( n27115 , n1476 , n26501 );
nor ( n27116 , n27114 , n27115 );
and ( n27117 , n27113 , n27116 );
nor ( n27118 , n27117 , n25901 );
and ( n27119 , n471 , n26633 );
and ( n27120 , n507 , n26635 );
nor ( n27121 , n27119 , n27120 );
and ( n27122 , n1391 , n25975 );
and ( n27123 , n1522 , n26621 );
nor ( n27124 , n27122 , n27123 );
and ( n27125 , n27121 , n27124 );
nor ( n27126 , n27125 , n25883 );
nor ( n27127 , n27118 , n27126 );
and ( n27128 , n785 , n27087 );
and ( n27129 , n1532 , n26682 );
nor ( n27130 , n27128 , n27129 );
and ( n27131 , n1276 , n25975 );
and ( n27132 , n707 , n26497 );
nor ( n27133 , n27131 , n27132 );
and ( n27134 , n27130 , n27133 );
nor ( n27135 , n27134 , n25868 );
and ( n27136 , n548 , n26811 );
and ( n27137 , n623 , n26511 );
nor ( n27138 , n27136 , n27137 );
and ( n27139 , n1265 , n25975 );
and ( n27140 , n1541 , n21742 );
nor ( n27141 , n27139 , n27140 );
and ( n27142 , n27138 , n27141 );
nor ( n27143 , n27142 , n25990 );
nor ( n27144 , n27135 , n27143 );
nand ( n27145 , n27110 , n27127 , n27144 );
and ( n27146 , n257 , n26287 );
and ( n27147 , n592 , n26601 );
nor ( n27148 , n27146 , n27147 );
and ( n27149 , n1387 , n26474 );
and ( n27150 , n769 , n26802 );
nor ( n27151 , n27149 , n27150 );
and ( n27152 , n27148 , n27151 );
nor ( n27153 , n27152 , n25868 );
and ( n27154 , n576 , n25933 );
not ( n27155 , n23605 );
and ( n27156 , n458 , n27155 );
nor ( n27157 , n27154 , n27156 );
and ( n27158 , n1401 , n25895 );
and ( n27159 , n259 , n26471 );
nor ( n27160 , n27158 , n27159 );
and ( n27161 , n27157 , n27160 );
nor ( n27162 , n27161 , n25883 );
nor ( n27163 , n27153 , n27162 );
and ( n27164 , n1450 , n25958 );
and ( n27165 , n1810 , n25961 );
nor ( n27166 , n27164 , n27165 );
and ( n27167 , n606 , n25825 );
and ( n27168 , n1197 , n23524 );
nor ( n27169 , n27167 , n27168 );
and ( n27170 , n27166 , n27169 );
nor ( n27171 , n27170 , n26618 );
and ( n27172 , n676 , n25970 );
and ( n27173 , n757 , n26511 );
nor ( n27174 , n27172 , n27173 );
and ( n27175 , n1236 , n25975 );
and ( n27176 , n258 , n25977 );
nor ( n27177 , n27175 , n27176 );
and ( n27178 , n27174 , n27177 );
nor ( n27179 , n27178 , n25901 );
and ( n27180 , n677 , n27039 );
and ( n27181 , n505 , n22154 );
nor ( n27182 , n27180 , n27181 );
and ( n27183 , n1157 , n25975 );
and ( n27184 , n260 , n25977 );
nor ( n27185 , n27183 , n27184 );
and ( n27186 , n27182 , n27185 );
nor ( n27187 , n27186 , n25990 );
nor ( n27188 , n27171 , n27179 , n27187 );
nand ( n27189 , n27163 , n27188 );
not ( n27190 , n2 );
and ( n27191 , n49 , n26460 );
and ( n27192 , n1449 , n25252 );
nor ( n27193 , n27191 , n27192 );
nor ( n27194 , n27190 , n27193 );
not ( n27195 , n2 );
and ( n27196 , n47 , n26460 );
and ( n27197 , n1450 , n25252 );
nor ( n27198 , n27196 , n27197 );
nor ( n27199 , n27195 , n27198 );
not ( n27200 , n2 );
and ( n27201 , n45 , n26460 );
and ( n27202 , n1452 , n25252 );
nor ( n27203 , n27201 , n27202 );
nor ( n27204 , n27200 , n27203 );
not ( n27205 , n2 );
and ( n27206 , n36 , n26460 );
and ( n27207 , n1453 , n25252 );
nor ( n27208 , n27206 , n27207 );
nor ( n27209 , n27205 , n27208 );
not ( n27210 , n2 );
and ( n27211 , n46 , n26460 );
and ( n27212 , n1451 , n25252 );
nor ( n27213 , n27211 , n27212 );
nor ( n27214 , n27210 , n27213 );
and ( n27215 , n552 , n26141 );
and ( n27216 , n574 , n26094 );
nor ( n27217 , n27215 , n27216 );
and ( n27218 , n1261 , n25895 );
and ( n27219 , n1493 , n26287 );
nor ( n27220 , n27218 , n27219 );
and ( n27221 , n27217 , n27220 );
nor ( n27222 , n27221 , n25990 );
not ( n27223 , n27222 );
and ( n27224 , n734 , n26802 );
and ( n27225 , n1477 , n26501 );
nor ( n27226 , n27224 , n27225 );
and ( n27227 , n1242 , n26624 );
and ( n27228 , n818 , n25947 );
nor ( n27229 , n27227 , n27228 );
and ( n27230 , n27226 , n27229 );
nor ( n27231 , n27230 , n25901 );
not ( n27232 , n25944 );
and ( n27233 , n787 , n27232 );
and ( n27234 , n1504 , n26501 );
nor ( n27235 , n27233 , n27234 );
and ( n27236 , n1388 , n26624 );
and ( n27237 , n668 , n26626 );
nor ( n27238 , n27236 , n27237 );
and ( n27239 , n27235 , n27238 );
nor ( n27240 , n27239 , n25868 );
nor ( n27241 , n27231 , n27240 );
and ( n27242 , n1115 , n25828 , n25956 );
and ( n27243 , n443 , n27039 );
and ( n27244 , n529 , n22154 );
nor ( n27245 , n27243 , n27244 );
and ( n27246 , n1386 , n23125 );
and ( n27247 , n1514 , n26507 );
nor ( n27248 , n27246 , n27247 );
and ( n27249 , n27245 , n27248 );
nor ( n27250 , n27249 , n25883 );
nor ( n27251 , n27242 , n27250 );
nand ( n27252 , n27223 , n27241 , n27251 );
and ( n27253 , n382 , n25825 );
and ( n27254 , n1459 , n25958 );
and ( n27255 , n1044 , n25828 );
nor ( n27256 , n27253 , n27254 , n27255 );
or ( n27257 , n26618 , n27256 );
and ( n27258 , n655 , n27087 );
and ( n27259 , n669 , n26764 );
nor ( n27260 , n27258 , n27259 );
and ( n27261 , n1371 , n25975 );
and ( n27262 , n1529 , n26501 );
nor ( n27263 , n27261 , n27262 );
and ( n27264 , n27260 , n27263 );
nor ( n27265 , n27264 , n25868 );
and ( n27266 , n473 , n26633 );
and ( n27267 , n526 , n26635 );
nor ( n27268 , n27266 , n27267 );
and ( n27269 , n1253 , n25975 );
and ( n27270 , n1533 , n21742 );
nor ( n27271 , n27269 , n27270 );
and ( n27272 , n27268 , n27271 );
nor ( n27273 , n27272 , n25883 );
nor ( n27274 , n27265 , n27273 );
and ( n27275 , n732 , n27087 );
and ( n27276 , n1510 , n26682 );
nor ( n27277 , n27275 , n27276 );
and ( n27278 , n1247 , n25975 );
and ( n27279 , n817 , n26497 );
nor ( n27280 , n27278 , n27279 );
and ( n27281 , n27277 , n27280 );
nor ( n27282 , n27281 , n25901 );
and ( n27283 , n550 , n26811 );
and ( n27284 , n625 , n26635 );
nor ( n27285 , n27283 , n27284 );
and ( n27286 , n1266 , n25975 );
and ( n27287 , n1488 , n21742 );
nor ( n27288 , n27286 , n27287 );
and ( n27289 , n27285 , n27288 );
nor ( n27290 , n27289 , n25990 );
nor ( n27291 , n27282 , n27290 );
nand ( n27292 , n27257 , n27274 , n27291 );
not ( n27293 , n829 );
or ( n27294 , n27293 , n16746 );
or ( n27295 , n829 , n1234 );
nand ( n27296 , n27295 , n17553 , n16266 );
nand ( n27297 , n27294 , n27296 );
and ( n27298 , n16258 , n27297 );
and ( n27299 , n1828 , n27293 );
nor ( n27300 , n27298 , n27299 );
nor ( n27301 , n16257 , n27300 );
and ( n27302 , n478 , n21583 );
and ( n27303 , n1399 , n26624 );
and ( n27304 , n533 , n27155 );
nor ( n27305 , n27302 , n27303 , n27304 );
or ( n27306 , n25883 , n27305 );
and ( n27307 , n1394 , n26291 );
and ( n27308 , n565 , n26738 );
and ( n27309 , n713 , n25939 );
nor ( n27310 , n27307 , n27308 , n27309 );
or ( n27311 , n25868 , n27310 );
and ( n27312 , n608 , n25825 );
and ( n27313 , n1416 , n25958 );
nor ( n27314 , n27312 , n27313 );
not ( n27315 , n27314 );
not ( n27316 , n26618 );
and ( n27317 , n27315 , n27316 );
and ( n27318 , n632 , n26059 );
not ( n27319 , n23124 );
and ( n27320 , n1205 , n27319 );
and ( n27321 , n485 , n26111 );
nor ( n27322 , n27318 , n27320 , n27321 );
or ( n27323 , n25990 , n27322 );
and ( n27324 , n1238 , n25894 );
and ( n27325 , n739 , n26111 );
and ( n27326 , n823 , n25844 );
nor ( n27327 , n27324 , n27325 , n27326 );
or ( n27328 , n25901 , n27327 );
nand ( n27329 , n27323 , n27328 );
nor ( n27330 , n27317 , n27329 );
nand ( n27331 , n27306 , n27311 , n27330 );
nand ( n27332 , n1546 , n15309 , n15328 , n13535 );
nand ( n27333 , n218 , n1545 , n15336 , n13535 );
nand ( n27334 , n27332 , n27333 );
and ( n27335 , n1559 , n27334 );
nor ( n27336 , n27335 , n744 );
nor ( n27337 , n20569 , n27336 );
and ( n27338 , n1576 , n27334 );
nor ( n27339 , n27338 , n746 );
nor ( n27340 , n20577 , n27339 );
and ( n27341 , n695 , n15110 );
and ( n27342 , n698 , n25447 );
nor ( n27343 , n27341 , n27342 );
nand ( n27344 , n27343 , n15189 , n25452 );
or ( n27345 , n1162 , n15839 );
or ( n27346 , n15191 , n25441 );
nand ( n27347 , n27345 , n27346 , n15165 );
and ( n27348 , n27344 , n27347 );
or ( n27349 , n15168 , n25452 );
or ( n27350 , n1394 , n15189 );
nand ( n27351 , n27349 , n27350 );
nor ( n27352 , n27348 , n27351 , n15175 );
or ( n27353 , n16778 , n27352 );
nand ( n27354 , n27353 , n17477 );
or ( n27355 , n27354 , n750 , n774 );
nor ( n27356 , n1160 , n1471 , n25441 );
not ( n27357 , n27356 );
nor ( n27358 , n27357 , n1161 , n1268 , n1400 );
nand ( n27359 , n27358 , n25420 , n25451 );
nand ( n27360 , n27355 , n27359 );
and ( n27361 , n779 , n25435 );
and ( n27362 , n777 , n25437 );
nor ( n27363 , n27361 , n27362 );
and ( n27364 , n27363 , n15839 , n25441 );
not ( n27365 , n27344 );
nor ( n27366 , n27364 , n27365 );
or ( n27367 , n15122 , n25419 );
or ( n27368 , n1270 , n15192 );
and ( n27369 , n782 , n25414 );
and ( n27370 , n783 , n25425 );
nor ( n27371 , n27369 , n27370 );
nand ( n27372 , n27371 , n15192 , n25419 );
and ( n27373 , n16794 , n27372 );
not ( n27374 , n15139 );
nor ( n27375 , n27373 , n27374 );
nand ( n27376 , n27367 , n27368 , n27375 );
nand ( n27377 , n27366 , n27376 , n15108 , n27359 );
nand ( n27378 , n27360 , n27377 );
not ( n27379 , n2 );
and ( n27380 , n14628 , n12965 );
and ( n27381 , n1126 , n14184 );
nor ( n27382 , n27380 , n27381 );
nor ( n27383 , n27379 , n27382 );
or ( n27384 , n20634 , n20641 );
nand ( n27385 , n27384 , n19933 );
and ( n27386 , n20643 , n27385 );
and ( n27387 , n370 , n25283 );
nor ( n27388 , n27386 , n27387 );
nor ( n27389 , n20652 , n27388 );
nand ( n27390 , n372 , n20647 );
not ( n27391 , n19930 );
nand ( n27392 , n386 , n19987 , n27391 );
nor ( n27393 , n19944 , n19937 , n27392 );
or ( n27394 , n372 , n27393 );
and ( n27395 , n372 , n27393 );
not ( n27396 , n20633 );
nor ( n27397 , n27395 , n27396 );
nand ( n27398 , n27394 , n27397 );
and ( n27399 , n27390 , n27398 );
nor ( n27400 , n27399 , n20652 );
nand ( n27401 , n754 , n16462 , n15348 );
not ( n27402 , n15366 );
nor ( n27403 , n27401 , n15309 , n27402 );
or ( n27404 , n19614 , n14980 );
nand ( n27405 , n15011 , n16672 );
or ( n27406 , n15009 , n27405 );
and ( n27407 , n15009 , n27405 );
nor ( n27408 , n27407 , n14979 );
nand ( n27409 , n27406 , n27408 );
nand ( n27410 , n27404 , n27409 );
and ( n27411 , n14974 , n27410 );
or ( n27412 , n15007 , n636 );
or ( n27413 , n19614 , n537 );
nand ( n27414 , n27412 , n27413 );
and ( n27415 , n1819 , n27414 );
nor ( n27416 , n27411 , n27415 );
nor ( n27417 , n14973 , n27416 );
and ( n27418 , n1588 , n27334 );
nor ( n27419 , n27418 , n721 );
nor ( n27420 , n20587 , n27419 );
or ( n27421 , n15126 , n15828 );
not ( n27422 , n15125 );
nand ( n27423 , n15127 , n16793 );
or ( n27424 , n27422 , n27423 );
and ( n27425 , n27422 , n27423 );
nor ( n27426 , n27425 , n25262 );
nand ( n27427 , n27424 , n27426 );
nand ( n27428 , n27421 , n27427 );
and ( n27429 , n15090 , n27428 );
or ( n27430 , n15124 , n791 );
or ( n27431 , n15126 , n715 );
nand ( n27432 , n27430 , n27431 );
and ( n27433 , n1826 , n27432 );
nor ( n27434 , n27429 , n27433 );
nor ( n27435 , n15089 , n27434 );
and ( n27436 , n1609 , n27334 );
nor ( n27437 , n27436 , n664 );
nor ( n27438 , n20582 , n27437 );
and ( n27439 , n612 , n25323 );
and ( n27440 , n614 , n25325 );
nor ( n27441 , n27439 , n27440 );
nand ( n27442 , n27441 , n16400 , n25330 );
or ( n27443 , n1212 , n15792 );
or ( n27444 , n15733 , n25318 );
nand ( n27445 , n27443 , n27444 , n18572 );
and ( n27446 , n27442 , n27445 );
or ( n27447 , n15739 , n25330 );
or ( n27448 , n1205 , n16400 );
nand ( n27449 , n27447 , n27448 );
nor ( n27450 , n27446 , n27449 , n15722 );
or ( n27451 , n17215 , n27450 );
nand ( n27452 , n27451 , n17174 );
or ( n27453 , n27452 , n597 , n691 );
nor ( n27454 , n1156 , n1256 , n25318 );
not ( n27455 , n27454 );
nor ( n27456 , n27455 , n1439 , n1221 , n1255 );
nand ( n27457 , n27456 , n25329 , n25297 );
nand ( n27458 , n27453 , n27457 );
and ( n27459 , n696 , n25312 );
and ( n27460 , n678 , n25314 );
nor ( n27461 , n27459 , n27460 );
and ( n27462 , n27461 , n15792 , n25318 );
not ( n27463 , n27442 );
nor ( n27464 , n27462 , n27463 );
or ( n27465 , n15750 , n25296 );
or ( n27466 , n1258 , n16402 );
and ( n27467 , n751 , n25301 );
and ( n27468 , n716 , n15736 );
nor ( n27469 , n27467 , n27468 );
nand ( n27470 , n27469 , n16402 , n25296 );
and ( n27471 , n17169 , n27470 );
not ( n27472 , n15737 );
nor ( n27473 , n27471 , n27472 );
nand ( n27474 , n27465 , n27466 , n27473 );
nand ( n27475 , n27464 , n27474 , n15720 , n27457 );
nand ( n27476 , n27458 , n27475 );
and ( n27477 , n807 , n16338 );
and ( n27478 , n804 , n16300 );
nor ( n27479 , n27477 , n27478 );
nand ( n27480 , n27479 , n16355 , n25510 );
or ( n27481 , n1237 , n16439 );
or ( n27482 , n16357 , n25500 );
nand ( n27483 , n27481 , n27482 , n16329 );
and ( n27484 , n27480 , n27483 );
or ( n27485 , n16332 , n25510 );
or ( n27486 , n1238 , n16355 );
nand ( n27487 , n27485 , n27486 );
nor ( n27488 , n27484 , n27487 , n16339 );
or ( n27489 , n16716 , n27488 );
nand ( n27490 , n27489 , n17502 );
or ( n27491 , n27490 , n793 , n794 );
nor ( n27492 , n1231 , n1467 , n25500 );
not ( n27493 , n27492 );
nor ( n27494 , n27493 , n1234 , n1233 , n1366 );
nand ( n27495 , n27494 , n25480 , n25509 );
nand ( n27496 , n27491 , n27495 );
and ( n27497 , n843 , n16273 );
and ( n27498 , n846 , n25496 );
nor ( n27499 , n27497 , n27498 );
and ( n27500 , n27499 , n16439 , n25500 );
not ( n27501 , n27480 );
nor ( n27502 , n27500 , n27501 );
or ( n27503 , n16281 , n25479 );
or ( n27504 , n1235 , n16361 );
and ( n27505 , n848 , n25474 );
and ( n27506 , n837 , n25485 );
nor ( n27507 , n27505 , n27506 );
nand ( n27508 , n27507 , n16361 , n25479 );
and ( n27509 , n16728 , n27508 );
nor ( n27510 , n27509 , n16725 );
nand ( n27511 , n27503 , n27504 , n27510 );
nand ( n27512 , n27502 , n27511 , n16295 , n27495 );
nand ( n27513 , n27496 , n27512 );
nand ( n27514 , n1083 , n26829 , n21626 , n26831 );
nor ( n27515 , n27514 , n1124 , n1148 );
and ( n27516 , n26824 , n27515 );
nor ( n27517 , n27516 , n21622 );
and ( n27518 , n21521 , n21533 );
not ( n27519 , n21626 );
nor ( n27520 , n1066 , n1083 );
nand ( n27521 , n27520 , n21623 , n15610 , n15582 );
nor ( n27522 , n27518 , n27519 , n27521 );
and ( n27523 , n27522 , n21632 , n21628 );
and ( n27524 , n1095 , n15647 );
nor ( n27525 , n27523 , n27524 );
and ( n27526 , n1114 , n27517 , n27525 );
not ( n27527 , n13586 );
and ( n27528 , n20157 , n13583 , n27527 , n13591 );
nand ( n27529 , n27528 , n202 , n13853 );
nand ( n27530 , n1147 , n13594 , n27529 );
and ( n27531 , n13580 , n27530 );
not ( n27532 , n2 );
nor ( n27533 , n27531 , n27532 );
nand ( n27534 , n1175 , n19378 , n15668 , n15676 );
nand ( n27535 , n1175 , n15617 , n15622 );
not ( n27536 , n27535 );
not ( n27537 , n21642 );
or ( n27538 , n27536 , n27537 );
nand ( n27539 , n27538 , n24390 );
and ( n27540 , n27534 , n27539 );
nor ( n27541 , n27540 , n21342 );
not ( n27542 , n26878 );
and ( n27543 , n476 , n27542 );
and ( n27544 , n990 , n26291 );
not ( n27545 , n26093 );
and ( n27546 , n532 , n27545 );
nor ( n27547 , n27543 , n27544 , n27546 );
or ( n27548 , n25883 , n27547 );
and ( n27549 , n553 , n27542 );
and ( n27550 , n1067 , n26915 );
and ( n27551 , n629 , n22155 );
nor ( n27552 , n27549 , n27550 , n27551 );
or ( n27553 , n25990 , n27552 );
and ( n27554 , n324 , n26491 );
and ( n27555 , n737 , n26267 );
and ( n27556 , n1121 , n27319 );
not ( n27557 , n23604 );
and ( n27558 , n820 , n27557 );
nor ( n27559 , n27555 , n27556 , n27558 );
nor ( n27560 , n25901 , n27559 );
and ( n27561 , n1096 , n26900 );
not ( n27562 , n25870 );
and ( n27563 , n659 , n27562 );
and ( n27564 , n712 , n22152 );
nor ( n27565 , n27561 , n27563 , n27564 );
nor ( n27566 , n25868 , n27565 );
nor ( n27567 , n27554 , n27560 , n27566 );
nand ( n27568 , n27548 , n27553 , n27567 );
and ( n27569 , n480 , n27542 );
and ( n27570 , n1070 , n26291 );
and ( n27571 , n536 , n27545 );
nor ( n27572 , n27569 , n27570 , n27571 );
or ( n27573 , n25990 , n27572 );
and ( n27574 , n566 , n27542 );
and ( n27575 , n1122 , n26915 );
and ( n27576 , n781 , n22155 );
nor ( n27577 , n27574 , n27575 , n27576 );
or ( n27578 , n26877 , n27577 );
and ( n27579 , n314 , n26491 );
and ( n27580 , n441 , n25852 );
and ( n27581 , n991 , n27319 );
and ( n27582 , n464 , n22152 );
nor ( n27583 , n27580 , n27581 , n27582 );
nor ( n27584 , n25883 , n27583 );
and ( n27585 , n1097 , n26900 );
and ( n27586 , n557 , n26902 );
and ( n27587 , n634 , n22152 );
nor ( n27588 , n27585 , n27586 , n27587 );
nor ( n27589 , n25868 , n27588 );
nor ( n27590 , n27579 , n27584 , n27589 );
nand ( n27591 , n27573 , n27578 , n27590 );
and ( n27592 , n1256 , n26915 );
and ( n27593 , n493 , n21583 );
and ( n27594 , n498 , n27545 );
nor ( n27595 , n27592 , n27593 , n27594 );
or ( n27596 , n25990 , n27595 );
and ( n27597 , n680 , n27542 );
and ( n27598 , n1231 , n26915 );
and ( n27599 , n765 , n22155 );
nor ( n27600 , n27597 , n27598 , n27599 );
or ( n27601 , n26877 , n27600 );
and ( n27602 , n602 , n26491 );
and ( n27603 , n580 , n26267 );
and ( n27604 , n1268 , n27319 );
and ( n27605 , n585 , n27557 );
nor ( n27606 , n27603 , n27604 , n27605 );
nor ( n27607 , n25868 , n27606 );
and ( n27608 , n1248 , n26900 );
and ( n27609 , n445 , n27562 );
and ( n27610 , n451 , n22152 );
nor ( n27611 , n27608 , n27609 , n27610 );
nor ( n27612 , n25883 , n27611 );
nor ( n27613 , n27602 , n27607 , n27612 );
nand ( n27614 , n27596 , n27601 , n27613 );
and ( n27615 , n1402 , n26915 );
and ( n27616 , n579 , n21583 );
and ( n27617 , n589 , n27545 );
nor ( n27618 , n27615 , n27616 , n27617 );
or ( n27619 , n25868 , n27618 );
and ( n27620 , n496 , n27542 );
and ( n27621 , n1257 , n26915 );
and ( n27622 , n501 , n22155 );
nor ( n27623 , n27620 , n27621 , n27622 );
or ( n27624 , n25990 , n27623 );
and ( n27625 , n594 , n26491 );
and ( n27626 , n684 , n26267 );
and ( n27627 , n1372 , n27319 );
and ( n27628 , n767 , n26968 );
nor ( n27629 , n27626 , n27627 , n27628 );
nor ( n27630 , n25901 , n27629 );
and ( n27631 , n1397 , n26900 );
and ( n27632 , n448 , n27562 );
and ( n27633 , n454 , n22152 );
nor ( n27634 , n27631 , n27632 , n27633 );
nor ( n27635 , n25883 , n27634 );
nor ( n27636 , n27625 , n27630 , n27635 );
nand ( n27637 , n27619 , n27624 , n27636 );
and ( n27638 , n1158 , n26915 );
and ( n27639 , n555 , n21583 );
and ( n27640 , n572 , n27545 );
nor ( n27641 , n27638 , n27639 , n27640 );
or ( n27642 , n25990 , n27641 );
and ( n27643 , n740 , n27542 );
and ( n27644 , n1239 , n26915 );
and ( n27645 , n822 , n22155 );
nor ( n27646 , n27643 , n27644 , n27645 );
or ( n27647 , n26877 , n27646 );
and ( n27648 , n607 , n26491 );
and ( n27649 , n1163 , n26279 );
and ( n27650 , n788 , n26893 );
and ( n27651 , n714 , n22152 );
nor ( n27652 , n27649 , n27650 , n27651 );
nor ( n27653 , n25868 , n27652 );
and ( n27654 , n1396 , n26900 );
and ( n27655 , n442 , n27562 );
and ( n27656 , n534 , n22152 );
nor ( n27657 , n27654 , n27655 , n27656 );
nor ( n27658 , n25883 , n27657 );
nor ( n27659 , n27648 , n27653 , n27658 );
nand ( n27660 , n27642 , n27647 , n27659 );
and ( n27661 , n16885 , n16856 );
not ( n27662 , n27661 );
not ( n27663 , n16881 );
not ( n27664 , n27663 );
or ( n27665 , n27662 , n27664 );
or ( n27666 , n27661 , n27663 );
nand ( n27667 , n27665 , n27666 );
not ( n27668 , n895 );
not ( n27669 , n917 );
nor ( n27670 , n27669 , n19915 );
nand ( n27671 , n912 , n27670 );
not ( n27672 , n27671 );
and ( n27673 , n893 , n27672 );
nand ( n27674 , n919 , n894 , n27673 );
not ( n27675 , n27674 );
or ( n27676 , n27668 , n27675 );
or ( n27677 , n895 , n27674 );
nand ( n27678 , n27676 , n27677 );
and ( n27679 , n1249 , n25895 );
and ( n27680 , n645 , n25945 );
and ( n27681 , n519 , n27155 );
nor ( n27682 , n27679 , n27680 , n27681 );
or ( n27683 , n25883 , n27682 );
and ( n27684 , n1232 , n26291 );
and ( n27685 , n730 , n26738 );
and ( n27686 , n809 , n25939 );
nor ( n27687 , n27684 , n27685 , n27686 );
or ( n27688 , n25901 , n27687 );
not ( n27689 , n25990 );
and ( n27690 , n1213 , n23125 );
and ( n27691 , n742 , n26631 );
and ( n27692 , n617 , n26495 );
nor ( n27693 , n27690 , n27691 , n27692 );
not ( n27694 , n27693 );
and ( n27695 , n27689 , n27694 );
and ( n27696 , n1269 , n26891 );
and ( n27697 , n568 , n26893 );
and ( n27698 , n700 , n22152 );
nor ( n27699 , n27696 , n27697 , n27698 );
nor ( n27700 , n25868 , n27699 );
nor ( n27701 , n27695 , n27700 );
nand ( n27702 , n27683 , n27688 , n27701 );
and ( n27703 , n718 , n723 );
nor ( n27704 , n27703 , n15090 , n17676 );
and ( n27705 , n718 , n18627 );
not ( n27706 , n17633 );
nand ( n27707 , n17625 , n27706 );
and ( n27708 , n17632 , n27707 );
or ( n27709 , n17632 , n27707 );
nand ( n27710 , n27709 , n15095 );
nor ( n27711 , n27708 , n27710 );
nor ( n27712 , n27705 , n1826 , n27711 );
nor ( n27713 , n15089 , n27704 , n27712 );
buf ( n27714 , n13198 );
not ( n27715 , n14803 );
nand ( n27716 , n27715 , n14800 );
nor ( n27717 , n27714 , n27716 );
or ( n27718 , n27717 , n12836 );
nand ( n27719 , n27718 , n188 );
or ( n27720 , n188 , n1821 );
not ( n27721 , n14794 );
nand ( n27722 , n27720 , n27721 );
nand ( n27723 , n27719 , n2 , n27722 );
nor ( n27724 , n1711 , n1697 , n12493 );
not ( n27725 , n27724 );
not ( n27726 , n1711 );
not ( n27727 , n1697 );
nand ( n27728 , n27726 , n27727 , n13557 );
or ( n27729 , n27728 , n1699 , n1709 );
or ( n27730 , n1699 , n12512 );
nand ( n27731 , n27729 , n27730 );
not ( n27732 , n27731 );
and ( n27733 , n27725 , n27732 );
nor ( n27734 , n27733 , n13551 );
not ( n27735 , n2 );
not ( n27736 , n12903 );
and ( n27737 , n14628 , n27736 );
and ( n27738 , n1127 , n14184 );
nor ( n27739 , n27737 , n27738 );
nor ( n27740 , n27735 , n27739 );
not ( n27741 , n539 );
or ( n27742 , n27741 , n14980 );
or ( n27743 , n539 , n1151 );
nand ( n27744 , n27743 , n17288 , n25593 );
nand ( n27745 , n27742 , n27744 );
and ( n27746 , n14974 , n27745 );
and ( n27747 , n1819 , n27741 );
nor ( n27748 , n27746 , n27747 );
nor ( n27749 , n14973 , n27748 );
nand ( n27750 , n1819 , n15007 );
or ( n27751 , n537 , n15874 );
and ( n27752 , n1151 , n25593 );
nor ( n27753 , n27752 , n15007 );
or ( n27754 , n15009 , n27753 );
nand ( n27755 , n27751 , n27754 , n14974 );
and ( n27756 , n27750 , n27755 );
nor ( n27757 , n27756 , n14973 );
and ( n27758 , n539 , n540 );
nor ( n27759 , n27758 , n14974 , n17331 );
and ( n27760 , n540 , n18536 );
not ( n27761 , n17289 );
nand ( n27762 , n17281 , n27761 );
and ( n27763 , n17288 , n27762 );
or ( n27764 , n17288 , n27762 );
nand ( n27765 , n27764 , n25593 );
nor ( n27766 , n27763 , n27765 );
nor ( n27767 , n27760 , n1819 , n27766 );
nor ( n27768 , n14973 , n27759 , n27767 );
nand ( n27769 , n577 , n22477 );
or ( n27770 , n577 , n20233 );
nand ( n27771 , n27770 , n1800 , n20234 );
and ( n27772 , n27769 , n27771 );
nor ( n27773 , n27772 , n834 );
nand ( n27774 , n606 , n22477 );
or ( n27775 , n606 , n22500 );
nand ( n27776 , n27775 , n1800 , n22501 );
and ( n27777 , n27774 , n27776 );
nor ( n27778 , n27777 , n834 );
and ( n27779 , n640 , n641 );
nor ( n27780 , n27779 , n15704 , n17412 );
and ( n27781 , n641 , n16393 );
not ( n27782 , n17370 );
nand ( n27783 , n17362 , n27782 );
and ( n27784 , n17369 , n27783 );
or ( n27785 , n17369 , n27783 );
nand ( n27786 , n27785 , n15709 );
nor ( n27787 , n27784 , n27786 );
nor ( n27788 , n27781 , n1808 , n27787 );
nor ( n27789 , n15703 , n27780 , n27788 );
not ( n27790 , n1105 );
not ( n27791 , n27525 );
or ( n27792 , n27790 , n27791 );
nand ( n27793 , n27792 , n27517 );
and ( n27794 , n15611 , n19379 );
and ( n27795 , n15624 , n19384 );
nor ( n27796 , n27794 , n27795 , n1167 );
not ( n27797 , n15630 );
not ( n27798 , n15638 );
and ( n27799 , n27797 , n27798 );
nor ( n27800 , n27799 , n1806 );
not ( n27801 , n21658 );
and ( n27802 , n21532 , n15601 , n21627 , n27801 );
nand ( n27803 , n27800 , n21647 , n27802 );
nand ( n27804 , n1100 , n15651 );
not ( n27805 , n15674 );
nand ( n27806 , n27805 , n15631 , n27802 , n21624 );
nand ( n27807 , n27803 , n27804 , n27806 );
nor ( n27808 , n27796 , n27807 );
or ( n27809 , n15217 , n267 );
nand ( n27810 , n27809 , n24239 );
nand ( n27811 , n27810 , n15216 );
nand ( n27812 , n1217 , n23641 , n15221 );
not ( n27813 , n15217 );
not ( n27814 , n20158 );
or ( n27815 , n27813 , n27814 );
and ( n27816 , n20161 , n20163 );
nand ( n27817 , n27815 , n27816 );
and ( n27818 , n27811 , n27812 , n27817 );
not ( n27819 , n2 );
nor ( n27820 , n27818 , n27819 );
not ( n27821 , n2 );
and ( n27822 , n1499 , n20158 , n27816 );
or ( n27823 , n15207 , n267 );
nand ( n27824 , n27823 , n24239 );
and ( n27825 , n27824 , n15221 );
nor ( n27826 , n27822 , n27825 );
nor ( n27827 , n27821 , n27826 );
and ( n27828 , n1254 , n25895 );
and ( n27829 , n446 , n25945 );
and ( n27830 , n452 , n27155 );
nor ( n27831 , n27828 , n27829 , n27830 );
or ( n27832 , n25883 , n27831 );
and ( n27833 , n1229 , n26291 );
and ( n27834 , n582 , n26738 );
and ( n27835 , n586 , n25939 );
nor ( n27836 , n27833 , n27834 , n27835 );
or ( n27837 , n25868 , n27836 );
not ( n27838 , n25990 );
and ( n27839 , n1267 , n23125 );
and ( n27840 , n494 , n26966 );
and ( n27841 , n499 , n26495 );
nor ( n27842 , n27839 , n27840 , n27841 );
not ( n27843 , n27842 );
and ( n27844 , n27838 , n27843 );
and ( n27845 , n1181 , n26891 );
and ( n27846 , n683 , n26893 );
and ( n27847 , n766 , n22152 );
nor ( n27848 , n27845 , n27846 , n27847 );
nor ( n27849 , n25901 , n27848 );
nor ( n27850 , n27844 , n27849 );
nand ( n27851 , n27832 , n27837 , n27850 );
and ( n27852 , n1251 , n25895 );
and ( n27853 , n449 , n25945 );
and ( n27854 , n455 , n25947 );
nor ( n27855 , n27852 , n27853 , n27854 );
or ( n27856 , n25883 , n27855 );
and ( n27857 , n1240 , n25895 );
and ( n27858 , n685 , n25945 );
and ( n27859 , n768 , n27155 );
nor ( n27860 , n27857 , n27858 , n27859 );
or ( n27861 , n25901 , n27860 );
not ( n27862 , n25990 );
and ( n27863 , n1260 , n23125 );
and ( n27864 , n497 , n26966 );
and ( n27865 , n502 , n26968 );
nor ( n27866 , n27863 , n27864 , n27865 );
not ( n27867 , n27866 );
and ( n27868 , n27862 , n27867 );
and ( n27869 , n1272 , n26891 );
and ( n27870 , n584 , n26902 );
and ( n27871 , n661 , n22152 );
nor ( n27872 , n27869 , n27870 , n27871 );
nor ( n27873 , n25868 , n27872 );
nor ( n27874 , n27868 , n27873 );
nand ( n27875 , n27856 , n27861 , n27874 );
not ( n27876 , n1548 );
or ( n27877 , n25960 , n23527 );
not ( n27878 , n27877 );
or ( n27879 , n27876 , n27878 );
or ( n27880 , n16073 , n27877 );
nand ( n27881 , n27879 , n27880 );
nand ( n27882 , n16981 , n19826 );
nand ( n27883 , n1321 , n1405 );
nand ( n27884 , n17005 , n27883 );
not ( n27885 , n27884 );
and ( n27886 , n17002 , n27885 );
nand ( n27887 , n16983 , n19843 , n27886 );
nor ( n27888 , n1330 , n27882 , n27887 );
and ( n27889 , n27888 , n1165 );
not ( n27890 , n27888 );
and ( n27891 , n27890 , n19230 );
nor ( n27892 , n27889 , n27891 );
not ( n27893 , n1552 );
not ( n27894 , n27877 );
or ( n27895 , n27893 , n27894 );
or ( n27896 , n16077 , n27877 );
nand ( n27897 , n27895 , n27896 );
not ( n27898 , n1554 );
not ( n27899 , n27877 );
or ( n27900 , n27898 , n27899 );
or ( n27901 , n16089 , n27877 );
nand ( n27902 , n27900 , n27901 );
not ( n27903 , n1555 );
not ( n27904 , n27877 );
or ( n27905 , n27903 , n27904 );
or ( n27906 , n16069 , n27877 );
nand ( n27907 , n27905 , n27906 );
not ( n27908 , n1836 );
nand ( n27909 , n27908 , n1557 );
and ( n27910 , n27909 , n27877 );
not ( n27911 , n2 );
nor ( n27912 , n27910 , n27911 );
nand ( n27913 , n16910 , n19743 );
nand ( n27914 , n1206 , n1370 );
nand ( n27915 , n16934 , n27914 );
not ( n27916 , n27915 );
and ( n27917 , n16931 , n27916 );
nand ( n27918 , n16912 , n19760 , n27917 );
nor ( n27919 , n1306 , n27913 , n27918 );
and ( n27920 , n27919 , n1308 );
not ( n27921 , n27919 );
and ( n27922 , n27921 , n19186 );
nor ( n27923 , n27920 , n27922 );
nand ( n27924 , n17051 , n18958 );
nand ( n27925 , n1342 , n1343 );
nand ( n27926 , n17075 , n27925 );
not ( n27927 , n27926 );
and ( n27928 , n17072 , n27927 );
nand ( n27929 , n17053 , n18975 , n27928 );
nor ( n27930 , n1361 , n27924 , n27929 );
and ( n27931 , n27930 , n1395 );
not ( n27932 , n27930 );
and ( n27933 , n27932 , n18949 );
nor ( n27934 , n27931 , n27933 );
not ( n27935 , n16927 );
nor ( n27936 , n27935 , n16961 );
not ( n27937 , n27936 );
nor ( n27938 , n21371 , n21362 );
not ( n27939 , n27938 );
or ( n27940 , n27937 , n27939 );
or ( n27941 , n27936 , n27938 );
nand ( n27942 , n27940 , n27941 );
not ( n27943 , n16854 );
nor ( n27944 , n27943 , n16888 );
not ( n27945 , n27944 );
nor ( n27946 , n21615 , n21603 );
not ( n27947 , n27946 );
or ( n27948 , n27945 , n27947 );
or ( n27949 , n27944 , n27946 );
nand ( n27950 , n27948 , n27949 );
not ( n27951 , n16998 );
nor ( n27952 , n27951 , n17032 );
not ( n27953 , n27952 );
nor ( n27954 , n21390 , n21381 );
not ( n27955 , n27954 );
or ( n27956 , n27953 , n27955 );
or ( n27957 , n27952 , n27954 );
nand ( n27958 , n27956 , n27957 );
not ( n27959 , n17068 );
nor ( n27960 , n27959 , n17102 );
not ( n27961 , n27960 );
nor ( n27962 , n21409 , n21400 );
not ( n27963 , n27962 );
or ( n27964 , n27961 , n27963 );
or ( n27965 , n27960 , n27962 );
nand ( n27966 , n27964 , n27965 );
not ( n27967 , n407 );
nand ( n27968 , n27967 , n1113 , n24277 );
and ( n27969 , n15678 , n27968 );
nor ( n27970 , n406 , n1113 );
nor ( n27971 , n27969 , n21342 , n27970 );
nand ( n27972 , n17099 , n17070 );
not ( n27973 , n27972 );
not ( n27974 , n17095 );
or ( n27975 , n27973 , n27974 );
or ( n27976 , n27972 , n17095 );
nand ( n27977 , n27975 , n27976 );
nand ( n27978 , n16836 , n19038 );
nand ( n27979 , n1412 , n1460 );
nand ( n27980 , n16861 , n27979 );
not ( n27981 , n27980 );
and ( n27982 , n16858 , n27981 );
nand ( n27983 , n16839 , n19055 , n27982 );
nor ( n27984 , n1398 , n27978 , n27983 );
and ( n27985 , n27984 , n1289 );
not ( n27986 , n27984 );
and ( n27987 , n27986 , n19031 );
nor ( n27988 , n27985 , n27987 );
not ( n27989 , n26534 );
not ( n27990 , n723 );
or ( n27991 , n27990 , n15828 );
or ( n27992 , n723 , n1161 );
nand ( n27993 , n27992 , n17632 , n15095 );
nand ( n27994 , n27991 , n27993 );
and ( n27995 , n15090 , n27994 );
and ( n27996 , n1826 , n27990 );
nor ( n27997 , n27995 , n27996 );
nor ( n27998 , n15089 , n27997 );
and ( n27999 , n1609 , n15365 );
nor ( n28000 , n27999 , n1294 );
nor ( n28001 , n20582 , n28000 );
not ( n28002 , n153 );
not ( n28003 , n13880 );
or ( n28004 , n28002 , n28003 );
not ( n28005 , n13880 );
nand ( n28006 , n158 , n28005 );
nand ( n28007 , n28004 , n28006 );
not ( n28008 , n2 );
and ( n28009 , n223 , n13199 );
and ( n28010 , n195 , n13200 );
nor ( n28011 , n28009 , n28010 );
nor ( n28012 , n28008 , n28011 , n26531 );
not ( n28013 , n116 );
not ( n28014 , n1708 );
or ( n28015 , n28013 , n28014 );
not ( n28016 , n20633 );
and ( n28017 , n326 , n28016 );
not ( n28018 , n326 );
not ( n28019 , n12880 );
not ( n28020 , n28019 );
not ( n28021 , n28020 );
not ( n28022 , n28021 );
and ( n28023 , n28018 , n28022 );
not ( n28024 , n28019 );
or ( n28025 , n1838 , n28024 );
nand ( n28026 , n28025 , n20633 );
nor ( n28027 , n28023 , n28026 );
nor ( n28028 , n28017 , n28027 );
or ( n28029 , n1708 , n28028 );
nand ( n28030 , n28015 , n28029 );
not ( n28031 , n118 );
not ( n28032 , n1708 );
or ( n28033 , n28031 , n28032 );
and ( n28034 , n330 , n28016 );
not ( n28035 , n330 );
not ( n28036 , n28021 );
and ( n28037 , n28035 , n28036 );
not ( n28038 , n28019 );
or ( n28039 , n1842 , n28038 );
buf ( n28040 , n20632 );
nand ( n28041 , n28039 , n28040 );
nor ( n28042 , n28037 , n28041 );
nor ( n28043 , n28034 , n28042 );
or ( n28044 , n1708 , n28043 );
nand ( n28045 , n28033 , n28044 );
not ( n28046 , n117 );
not ( n28047 , n1708 );
or ( n28048 , n28046 , n28047 );
and ( n28049 , n331 , n28016 );
not ( n28050 , n331 );
not ( n28051 , n28020 );
not ( n28052 , n28051 );
and ( n28053 , n28050 , n28052 );
or ( n28054 , n1843 , n28024 );
nand ( n28055 , n28054 , n20633 );
nor ( n28056 , n28053 , n28055 );
nor ( n28057 , n28049 , n28056 );
or ( n28058 , n1708 , n28057 );
nand ( n28059 , n28048 , n28058 );
not ( n28060 , n115 );
not ( n28061 , n1708 );
or ( n28062 , n28060 , n28061 );
and ( n28063 , n332 , n28016 );
not ( n28064 , n332 );
not ( n28065 , n28021 );
and ( n28066 , n28064 , n28065 );
or ( n28067 , n1846 , n28038 );
nand ( n28068 , n28067 , n20633 );
nor ( n28069 , n28066 , n28068 );
nor ( n28070 , n28063 , n28069 );
or ( n28071 , n1708 , n28070 );
nand ( n28072 , n28062 , n28071 );
not ( n28073 , n114 );
not ( n28074 , n1708 );
or ( n28075 , n28073 , n28074 );
and ( n28076 , n333 , n28016 );
not ( n28077 , n333 );
not ( n28078 , n28051 );
and ( n28079 , n28077 , n28078 );
or ( n28080 , n1847 , n28038 );
nand ( n28081 , n28080 , n20633 );
nor ( n28082 , n28079 , n28081 );
nor ( n28083 , n28076 , n28082 );
or ( n28084 , n1708 , n28083 );
nand ( n28085 , n28075 , n28084 );
not ( n28086 , n113 );
not ( n28087 , n1708 );
or ( n28088 , n28086 , n28087 );
and ( n28089 , n334 , n28016 );
not ( n28090 , n334 );
not ( n28091 , n28021 );
and ( n28092 , n28090 , n28091 );
or ( n28093 , n1840 , n28024 );
nand ( n28094 , n28093 , n28040 );
nor ( n28095 , n28092 , n28094 );
nor ( n28096 , n28089 , n28095 );
or ( n28097 , n1708 , n28096 );
nand ( n28098 , n28088 , n28097 );
not ( n28099 , n111 );
not ( n28100 , n1708 );
or ( n28101 , n28099 , n28100 );
and ( n28102 , n335 , n28016 );
not ( n28103 , n335 );
not ( n28104 , n12878 );
not ( n28105 , n28104 );
not ( n28106 , n28105 );
not ( n28107 , n28106 );
and ( n28108 , n28103 , n28107 );
not ( n28109 , n28104 );
or ( n28110 , n1845 , n28109 );
nand ( n28111 , n28110 , n28040 );
nor ( n28112 , n28108 , n28111 );
nor ( n28113 , n28102 , n28112 );
or ( n28114 , n1708 , n28113 );
nand ( n28115 , n28101 , n28114 );
not ( n28116 , n105 );
not ( n28117 , n1708 );
or ( n28118 , n28116 , n28117 );
and ( n28119 , n336 , n28016 );
not ( n28120 , n336 );
not ( n28121 , n28106 );
and ( n28122 , n28120 , n28121 );
not ( n28123 , n28104 );
or ( n28124 , n1840 , n28123 );
nand ( n28125 , n28124 , n20633 );
nor ( n28126 , n28122 , n28125 );
nor ( n28127 , n28119 , n28126 );
or ( n28128 , n1708 , n28127 );
nand ( n28129 , n28118 , n28128 );
not ( n28130 , n109 );
not ( n28131 , n1708 );
or ( n28132 , n28130 , n28131 );
and ( n28133 , n348 , n28016 );
not ( n28134 , n348 );
not ( n28135 , n28105 );
not ( n28136 , n28135 );
and ( n28137 , n28134 , n28136 );
or ( n28138 , n1843 , n28109 );
nand ( n28139 , n28138 , n28040 );
nor ( n28140 , n28137 , n28139 );
nor ( n28141 , n28133 , n28140 );
or ( n28142 , n1708 , n28141 );
nand ( n28143 , n28132 , n28142 );
not ( n28144 , n112 );
not ( n28145 , n1708 );
or ( n28146 , n28144 , n28145 );
and ( n28147 , n349 , n28016 );
not ( n28148 , n349 );
not ( n28149 , n28135 );
and ( n28150 , n28148 , n28149 );
or ( n28151 , n1841 , n28123 );
nand ( n28152 , n28151 , n28040 );
nor ( n28153 , n28150 , n28152 );
nor ( n28154 , n28147 , n28153 );
or ( n28155 , n1708 , n28154 );
nand ( n28156 , n28146 , n28155 );
not ( n28157 , n20633 );
nand ( n28158 , n350 , n28157 );
not ( n28159 , n27392 );
or ( n28160 , n350 , n28159 );
and ( n28161 , n350 , n28159 );
not ( n28162 , n20632 );
nor ( n28163 , n28161 , n28162 );
nand ( n28164 , n28160 , n28163 );
and ( n28165 , n28158 , n28164 );
nor ( n28166 , n28165 , n20652 );
not ( n28167 , n110 );
not ( n28168 , n1708 );
or ( n28169 , n28167 , n28168 );
and ( n28170 , n354 , n28016 );
not ( n28171 , n354 );
not ( n28172 , n28135 );
and ( n28173 , n28171 , n28172 );
or ( n28174 , n1842 , n28109 );
nand ( n28175 , n28174 , n28040 );
nor ( n28176 , n28173 , n28175 );
nor ( n28177 , n28170 , n28176 );
or ( n28178 , n1708 , n28177 );
nand ( n28179 , n28169 , n28178 );
not ( n28180 , n108 );
not ( n28181 , n1708 );
or ( n28182 , n28180 , n28181 );
and ( n28183 , n355 , n28157 );
not ( n28184 , n355 );
not ( n28185 , n28106 );
and ( n28186 , n28184 , n28185 );
or ( n28187 , n1838 , n28109 );
nand ( n28188 , n28187 , n20633 );
nor ( n28189 , n28186 , n28188 );
nor ( n28190 , n28183 , n28189 );
or ( n28191 , n1708 , n28190 );
nand ( n28192 , n28182 , n28191 );
not ( n28193 , n107 );
not ( n28194 , n1708 );
or ( n28195 , n28193 , n28194 );
and ( n28196 , n356 , n28016 );
not ( n28197 , n356 );
not ( n28198 , n28106 );
and ( n28199 , n28197 , n28198 );
or ( n28200 , n1846 , n28123 );
nand ( n28201 , n28200 , n20633 );
nor ( n28202 , n28199 , n28201 );
nor ( n28203 , n28196 , n28202 );
or ( n28204 , n1708 , n28203 );
nand ( n28205 , n28195 , n28204 );
not ( n28206 , n119 );
not ( n28207 , n1708 );
or ( n28208 , n28206 , n28207 );
and ( n28209 , n357 , n28016 );
not ( n28210 , n357 );
not ( n28211 , n28051 );
and ( n28212 , n28210 , n28211 );
or ( n28213 , n1845 , n28038 );
nand ( n28214 , n28213 , n20633 );
nor ( n28215 , n28212 , n28214 );
nor ( n28216 , n28209 , n28215 );
or ( n28217 , n1708 , n28216 );
nand ( n28218 , n28208 , n28217 );
not ( n28219 , n106 );
not ( n28220 , n1708 );
or ( n28221 , n28219 , n28220 );
and ( n28222 , n375 , n28016 );
not ( n28223 , n375 );
not ( n28224 , n28135 );
and ( n28225 , n28223 , n28224 );
or ( n28226 , n1847 , n28123 );
nand ( n28227 , n28226 , n28040 );
nor ( n28228 , n28225 , n28227 );
nor ( n28229 , n28222 , n28228 );
or ( n28230 , n1708 , n28229 );
nand ( n28231 , n28221 , n28230 );
not ( n28232 , n120 );
not ( n28233 , n1708 );
or ( n28234 , n28232 , n28233 );
and ( n28235 , n377 , n28016 );
not ( n28236 , n377 );
not ( n28237 , n28051 );
and ( n28238 , n28236 , n28237 );
or ( n28239 , n1841 , n28024 );
nand ( n28240 , n28239 , n28040 );
nor ( n28241 , n28238 , n28240 );
nor ( n28242 , n28235 , n28241 );
or ( n28243 , n1708 , n28242 );
nand ( n28244 , n28234 , n28243 );
not ( n28245 , n20203 );
nand ( n28246 , n28245 , n20175 );
and ( n28247 , n23646 , n28246 );
not ( n28248 , n20636 );
or ( n28249 , n281 , n328 );
not ( n28250 , n28249 );
nor ( n28251 , n28247 , n28248 , n28250 );
and ( n28252 , n605 , n22477 );
and ( n28253 , n22499 , n20232 );
nor ( n28254 , n28253 , n22477 , n22500 );
nor ( n28255 , n28252 , n28254 );
nor ( n28256 , n834 , n28255 );
nand ( n28257 , n1808 , n15752 );
or ( n28258 , n635 , n17197 );
and ( n28259 , n1156 , n15709 );
nor ( n28260 , n28259 , n15752 );
or ( n28261 , n26569 , n28260 );
nand ( n28262 , n28258 , n28261 , n15704 );
and ( n28263 , n28257 , n28262 );
nor ( n28264 , n28263 , n15703 );
and ( n28265 , n640 , n1808 );
and ( n28266 , n640 , n15711 );
or ( n28267 , n15704 , n640 );
or ( n28268 , n640 , n1156 );
nand ( n28269 , n28268 , n17369 , n15709 );
nand ( n28270 , n28267 , n28269 );
nor ( n28271 , n28266 , n28270 );
nor ( n28272 , n28265 , n15703 , n28271 );
nand ( n28273 , n1826 , n15124 );
or ( n28274 , n715 , n15097 );
and ( n28275 , n1161 , n15095 );
nor ( n28276 , n28275 , n15124 );
or ( n28277 , n27422 , n28276 );
nand ( n28278 , n28274 , n28277 , n15090 );
and ( n28279 , n28273 , n28278 );
nor ( n28280 , n28279 , n15089 );
and ( n28281 , n1576 , n15365 );
nor ( n28282 , n28281 , n1166 );
nor ( n28283 , n20577 , n28282 );
and ( n28284 , n1559 , n15365 );
nor ( n28285 , n28284 , n1120 );
nor ( n28286 , n20569 , n28285 );
and ( n28287 , n1588 , n15365 );
nor ( n28288 , n28287 , n1164 );
nor ( n28289 , n20587 , n28288 );
not ( n28290 , n406 );
nand ( n28291 , n1174 , n28290 , n26199 );
and ( n28292 , n15633 , n28291 );
nor ( n28293 , n391 , n1174 );
nor ( n28294 , n28292 , n21342 , n28293 );
not ( n28295 , n919 );
not ( n28296 , n27673 );
not ( n28297 , n28296 );
or ( n28298 , n28295 , n28297 );
or ( n28299 , n919 , n28296 );
nand ( n28300 , n28298 , n28299 );
not ( n28301 , n16621 );
not ( n28302 , n28301 );
nand ( n28303 , n1622 , n28302 );
and ( n28304 , n28303 , n15395 );
not ( n28305 , n2 );
nor ( n28306 , n28304 , n28305 );
not ( n28307 , n1398 );
not ( n28308 , n27978 );
and ( n28309 , n16855 , n27979 , n19071 );
and ( n28310 , n16853 , n28309 );
nand ( n28311 , n16839 , n28310 );
not ( n28312 , n28311 );
nand ( n28313 , n28308 , n28312 );
not ( n28314 , n28313 );
or ( n28315 , n28307 , n28314 );
or ( n28316 , n1398 , n28313 );
nand ( n28317 , n28315 , n28316 );
not ( n28318 , n1589 );
not ( n28319 , n1593 );
nand ( n28320 , n1594 , n1595 );
nor ( n28321 , n28319 , n28320 );
nand ( n28322 , n1601 , n28321 );
nor ( n28323 , n28318 , n28322 );
nand ( n28324 , n1607 , n28323 );
xor ( n28325 , n1592 , n28324 );
nor ( n28326 , n1755 , n28325 );
not ( n28327 , n1306 );
not ( n28328 , n27913 );
and ( n28329 , n16928 , n27914 , n19774 );
and ( n28330 , n16926 , n28329 );
nand ( n28331 , n16912 , n28330 );
not ( n28332 , n28331 );
nand ( n28333 , n28328 , n28332 );
not ( n28334 , n28333 );
or ( n28335 , n28327 , n28334 );
or ( n28336 , n1306 , n28333 );
nand ( n28337 , n28335 , n28336 );
not ( n28338 , n1361 );
not ( n28339 , n27924 );
and ( n28340 , n17098 , n27925 , n18986 );
and ( n28341 , n17067 , n28340 );
nand ( n28342 , n17053 , n28341 );
not ( n28343 , n28342 );
nand ( n28344 , n28339 , n28343 );
not ( n28345 , n28344 );
or ( n28346 , n28338 , n28345 );
or ( n28347 , n1361 , n28344 );
nand ( n28348 , n28346 , n28347 );
and ( n28349 , n444 , n26879 );
and ( n28350 , n447 , n22155 );
nor ( n28351 , n28349 , n28350 );
or ( n28352 , n25883 , n28351 );
and ( n28353 , n492 , n26879 );
and ( n28354 , n495 , n22155 );
nor ( n28355 , n28353 , n28354 );
or ( n28356 , n25990 , n28355 );
not ( n28357 , n25868 );
and ( n28358 , n581 , n26493 );
and ( n28359 , n583 , n26497 );
nor ( n28360 , n28358 , n28359 );
not ( n28361 , n28360 );
and ( n28362 , n28357 , n28361 );
and ( n28363 , n682 , n27039 );
and ( n28364 , n764 , n22154 );
nor ( n28365 , n28363 , n28364 );
nor ( n28366 , n25901 , n28365 );
nor ( n28367 , n28362 , n28366 );
nand ( n28368 , n28352 , n28356 , n28367 );
not ( n28369 , n1330 );
not ( n28370 , n27882 );
and ( n28371 , n16999 , n27883 , n19857 );
and ( n28372 , n16997 , n28371 );
nand ( n28373 , n16983 , n28372 );
not ( n28374 , n28373 );
nand ( n28375 , n28370 , n28374 );
not ( n28376 , n28375 );
or ( n28377 , n28369 , n28376 );
or ( n28378 , n1330 , n28375 );
nand ( n28379 , n28377 , n28378 );
and ( n28380 , n935 , n27000 );
nor ( n28381 , n28380 , n26452 );
not ( n28382 , n26434 );
nor ( n28383 , n28381 , n26451 , n28382 );
or ( n28384 , n27396 , n25277 );
nand ( n28385 , n28384 , n19926 );
and ( n28386 , n25279 , n28385 );
and ( n28387 , n369 , n20634 );
nor ( n28388 , n28386 , n28387 );
nor ( n28389 , n20652 , n28388 );
not ( n28390 , n100 );
not ( n28391 , n1708 );
or ( n28392 , n28390 , n28391 );
not ( n28393 , n346 );
not ( n28394 , n28162 );
not ( n28395 , n28394 );
not ( n28396 , n28395 );
or ( n28397 , n28393 , n28396 );
not ( n28398 , n20155 );
or ( n28399 , n346 , n28398 );
or ( n28400 , n1838 , n20155 );
nand ( n28401 , n28399 , n28400 , n28394 );
nand ( n28402 , n28397 , n28401 );
nand ( n28403 , n14176 , n28402 );
nand ( n28404 , n28392 , n28403 );
not ( n28405 , n97 );
not ( n28406 , n1708 );
or ( n28407 , n28405 , n28406 );
not ( n28408 , n343 );
not ( n28409 , n28394 );
not ( n28410 , n28409 );
or ( n28411 , n28408 , n28410 );
not ( n28412 , n20155 );
or ( n28413 , n343 , n28412 );
or ( n28414 , n1840 , n20155 );
not ( n28415 , n28162 );
nand ( n28416 , n28413 , n28414 , n28415 );
nand ( n28417 , n28411 , n28416 );
nand ( n28418 , n14176 , n28417 );
nand ( n28419 , n28407 , n28418 );
not ( n28420 , n98 );
not ( n28421 , n1708 );
or ( n28422 , n28420 , n28421 );
not ( n28423 , n342 );
not ( n28424 , n28395 );
or ( n28425 , n28423 , n28424 );
or ( n28426 , n342 , n28412 );
or ( n28427 , n1847 , n20155 );
nand ( n28428 , n28426 , n28427 , n28415 );
nand ( n28429 , n28425 , n28428 );
nand ( n28430 , n14176 , n28429 );
nand ( n28431 , n28422 , n28430 );
not ( n28432 , n99 );
not ( n28433 , n1708 );
or ( n28434 , n28432 , n28433 );
not ( n28435 , n341 );
not ( n28436 , n28409 );
or ( n28437 , n28435 , n28436 );
or ( n28438 , n341 , n28412 );
or ( n28439 , n1846 , n20155 );
nand ( n28440 , n28438 , n28439 , n28415 );
nand ( n28441 , n28437 , n28440 );
nand ( n28442 , n14176 , n28441 );
nand ( n28443 , n28434 , n28442 );
not ( n28444 , n101 );
not ( n28445 , n1708 );
or ( n28446 , n28444 , n28445 );
not ( n28447 , n340 );
not ( n28448 , n28409 );
or ( n28449 , n28447 , n28448 );
or ( n28450 , n340 , n28398 );
or ( n28451 , n1843 , n20155 );
nand ( n28452 , n28450 , n28451 , n28415 );
nand ( n28453 , n28449 , n28452 );
nand ( n28454 , n14176 , n28453 );
nand ( n28455 , n28446 , n28454 );
not ( n28456 , n104 );
not ( n28457 , n1708 );
or ( n28458 , n28456 , n28457 );
not ( n28459 , n338 );
not ( n28460 , n28409 );
or ( n28461 , n28459 , n28460 );
or ( n28462 , n338 , n20156 );
or ( n28463 , n1841 , n20155 );
nand ( n28464 , n28462 , n28463 , n28415 );
nand ( n28465 , n28461 , n28464 );
nand ( n28466 , n14176 , n28465 );
nand ( n28467 , n28458 , n28466 );
not ( n28468 , n102 );
not ( n28469 , n1708 );
or ( n28470 , n28468 , n28469 );
not ( n28471 , n339 );
not ( n28472 , n28395 );
or ( n28473 , n28471 , n28472 );
or ( n28474 , n339 , n28412 );
or ( n28475 , n1842 , n20155 );
nand ( n28476 , n28474 , n28475 , n28415 );
nand ( n28477 , n28473 , n28476 );
nand ( n28478 , n14176 , n28477 );
nand ( n28479 , n28470 , n28478 );
not ( n28480 , n26832 );
and ( n28481 , n15599 , n21647 , n28480 );
and ( n28482 , n312 , n1179 );
nor ( n28483 , n28482 , n1586 );
nor ( n28484 , n28481 , n28483 );
not ( n28485 , n2 );
and ( n28486 , n1623 , n16621 , n13560 );
not ( n28487 , n15394 );
nor ( n28488 , n28486 , n28487 );
nor ( n28489 , n28485 , n28488 );
not ( n28490 , n103 );
not ( n28491 , n1708 );
or ( n28492 , n28490 , n28491 );
not ( n28493 , n337 );
not ( n28494 , n28395 );
or ( n28495 , n28493 , n28494 );
or ( n28496 , n337 , n28398 );
or ( n28497 , n1845 , n20155 );
nand ( n28498 , n28496 , n28497 , n28415 );
nand ( n28499 , n28495 , n28498 );
nand ( n28500 , n14176 , n28499 );
nand ( n28501 , n28492 , n28500 );
nand ( n28502 , n1551 , n12836 );
and ( n28503 , n28502 , n12839 , n12847 );
not ( n28504 , n2 );
nor ( n28505 , n28503 , n28504 );
or ( n28506 , n26527 , n26529 );
nand ( n28507 , n28506 , n1558 );
and ( n28508 , n26528 , n28507 );
not ( n28509 , n2 );
nor ( n28510 , n28508 , n28509 );
not ( n28511 , n2 );
and ( n28512 , n1530 , n15245 );
nor ( n28513 , n28512 , n18682 , n18685 );
nor ( n28514 , n28511 , n15253 , n28513 );
not ( n28515 , n1547 );
nand ( n28516 , n28515 , n13594 );
or ( n28517 , n28162 , n20639 );
nand ( n28518 , n28517 , n14591 );
and ( n28519 , n25277 , n28518 );
and ( n28520 , n368 , n27396 );
nor ( n28521 , n28519 , n28520 );
nor ( n28522 , n20652 , n28521 );
not ( n28523 , n18928 );
or ( n28524 , n18385 , n28523 );
nand ( n28525 , n1414 , n28523 );
nand ( n28526 , n28524 , n28525 );
not ( n28527 , n18685 );
nor ( n28528 , n28527 , n15274 );
nand ( n28529 , n21743 , n28528 );
nor ( n28530 , n21796 , n28529 );
not ( n28531 , n27886 );
nor ( n28532 , n1326 , n1327 );
nand ( n28533 , n28532 , n19843 );
nor ( n28534 , n28531 , n28533 );
and ( n28535 , n28534 , n1328 );
not ( n28536 , n28534 );
and ( n28537 , n28536 , n16979 );
nor ( n28538 , n28535 , n28537 );
or ( n28539 , n18483 , n28523 );
nand ( n28540 , n1463 , n28523 );
nand ( n28541 , n28539 , n28540 );
or ( n28542 , n18380 , n28523 );
nand ( n28543 , n1464 , n28523 );
nand ( n28544 , n28542 , n28543 );
or ( n28545 , n18473 , n28523 );
nand ( n28546 , n1465 , n28523 );
nand ( n28547 , n28545 , n28546 );
or ( n28548 , n18754 , n28523 );
nand ( n28549 , n1466 , n28523 );
nand ( n28550 , n28548 , n28549 );
not ( n28551 , n1211 );
nor ( n28552 , n1218 , n1304 );
nand ( n28553 , n16908 , n28552 , n28330 );
not ( n28554 , n28553 );
or ( n28555 , n28551 , n28554 );
or ( n28556 , n1211 , n28553 );
nand ( n28557 , n28555 , n28556 );
not ( n28558 , n1186 );
nor ( n28559 , n1347 , n1348 );
nand ( n28560 , n17047 , n28559 , n28341 );
not ( n28561 , n28560 );
or ( n28562 , n28558 , n28561 );
or ( n28563 , n1186 , n28560 );
nand ( n28564 , n28562 , n28563 );
nor ( n28565 , n21747 , n28529 );
not ( n28566 , n21588 );
nor ( n28567 , n28566 , n28529 );
not ( n28568 , n2 );
and ( n28569 , n1587 , n15395 );
nor ( n28570 , n28569 , n28301 );
nor ( n28571 , n28568 , n28570 );
not ( n28572 , n1218 );
not ( n28573 , n27918 );
or ( n28574 , n28572 , n28573 );
or ( n28575 , n1218 , n27918 );
nand ( n28576 , n28574 , n28575 );
not ( n28577 , n27917 );
nand ( n28578 , n19760 , n28552 );
nor ( n28579 , n28577 , n28578 );
and ( n28580 , n28579 , n1305 );
not ( n28581 , n28579 );
and ( n28582 , n28581 , n16908 );
nor ( n28583 , n28580 , n28582 );
not ( n28584 , n1288 );
nor ( n28585 , n1287 , n1404 );
nand ( n28586 , n16832 , n28585 , n28310 );
not ( n28587 , n28586 );
or ( n28588 , n28584 , n28587 );
or ( n28589 , n1288 , n28586 );
nand ( n28590 , n28588 , n28589 );
not ( n28591 , n1378 );
nand ( n28592 , n16979 , n28532 , n28372 );
not ( n28593 , n28592 );
or ( n28594 , n28591 , n28593 );
or ( n28595 , n1378 , n28592 );
nand ( n28596 , n28594 , n28595 );
not ( n28597 , n21759 );
nor ( n28598 , n28597 , n28529 );
not ( n28599 , n1287 );
not ( n28600 , n27983 );
or ( n28601 , n28599 , n28600 );
or ( n28602 , n1287 , n27983 );
nand ( n28603 , n28601 , n28602 );
not ( n28604 , n1348 );
not ( n28605 , n27929 );
or ( n28606 , n28604 , n28605 );
or ( n28607 , n1348 , n27929 );
nand ( n28608 , n28606 , n28607 );
nand ( n28609 , n16880 , n16859 );
not ( n28610 , n28609 );
not ( n28611 , n19301 );
or ( n28612 , n28610 , n28611 );
or ( n28613 , n28609 , n19301 );
nand ( n28614 , n28612 , n28613 );
nand ( n28615 , n16953 , n16932 );
not ( n28616 , n28615 );
not ( n28617 , n19213 );
or ( n28618 , n28616 , n28617 );
or ( n28619 , n28615 , n19213 );
nand ( n28620 , n28618 , n28619 );
nand ( n28621 , n17024 , n17003 );
not ( n28622 , n28621 );
not ( n28623 , n19257 );
or ( n28624 , n28622 , n28623 );
or ( n28625 , n28621 , n19257 );
nand ( n28626 , n28624 , n28625 );
nand ( n28627 , n17094 , n17073 );
not ( n28628 , n28627 );
not ( n28629 , n19345 );
or ( n28630 , n28628 , n28629 );
or ( n28631 , n28627 , n19345 );
nand ( n28632 , n28630 , n28631 );
not ( n28633 , n14911 );
not ( n28634 , n17119 );
and ( n28635 , n28633 , n28634 );
not ( n28636 , n14911 );
not ( n28637 , n17121 );
or ( n28638 , n28636 , n28637 );
nand ( n28639 , n28638 , n1111 );
nor ( n28640 , n28635 , n28639 );
and ( n28641 , n1145 , n17118 );
nor ( n28642 , n1145 , n24413 );
nor ( n28643 , n28641 , n1111 , n28642 );
nor ( n28644 , n28640 , n28643 );
not ( n28645 , n1327 );
not ( n28646 , n27887 );
or ( n28647 , n28645 , n28646 );
or ( n28648 , n1327 , n27887 );
nand ( n28649 , n28647 , n28648 );
or ( n28650 , n17985 , n28523 );
or ( n28651 , n17811 , n18928 );
nand ( n28652 , n28650 , n28651 );
nand ( n28653 , n2 , n850 );
or ( n28654 , n1733 , n28653 );
not ( n28655 , n2 );
not ( n28656 , n19099 );
and ( n28657 , n1668 , n216 , n28656 );
and ( n28658 , n313 , n1649 , n216 , n19099 );
nor ( n28659 , n28657 , n28658 );
or ( n28660 , n28655 , n28659 );
not ( n28661 , n68 );
nand ( n28662 , n28661 , n216 , n2 );
nand ( n28663 , n28654 , n28660 , n28662 );
nand ( n28664 , n2 , n805 );
or ( n28665 , n1736 , n28664 );
not ( n28666 , n2 );
not ( n28667 , n19807 );
and ( n28668 , n1669 , n214 , n28667 );
and ( n28669 , n272 , n1606 , n214 , n19807 );
nor ( n28670 , n28668 , n28669 );
or ( n28671 , n28666 , n28670 );
not ( n28672 , n71 );
nand ( n28673 , n28672 , n214 , n2 );
nand ( n28674 , n28665 , n28671 , n28673 );
nand ( n28675 , n2 , n842 );
or ( n28676 , n1712 , n28675 );
not ( n28677 , n2 );
not ( n28678 , n19017 );
and ( n28679 , n1667 , n213 , n28678 );
and ( n28680 , n271 , n1620 , n213 , n19017 );
nor ( n28681 , n28679 , n28680 );
or ( n28682 , n28677 , n28681 );
not ( n28683 , n69 );
nand ( n28684 , n28683 , n213 , n2 );
nand ( n28685 , n28676 , n28682 , n28684 );
nand ( n28686 , n2 , n840 );
or ( n28687 , n1737 , n28686 );
not ( n28688 , n2 );
not ( n28689 , n19889 );
and ( n28690 , n1670 , n201 , n28689 );
and ( n28691 , n266 , n1621 , n201 , n19889 );
nor ( n28692 , n28690 , n28691 );
or ( n28693 , n28688 , n28692 );
not ( n28694 , n70 );
nand ( n28695 , n28694 , n201 , n2 );
nand ( n28696 , n28687 , n28693 , n28695 );
nand ( n28697 , n184 , n12842 , n12846 );
and ( n28698 , n27716 , n28697 );
not ( n28699 , n2 );
nor ( n28700 , n184 , n27714 );
nor ( n28701 , n28698 , n28699 , n28700 );
not ( n28702 , n1475 );
and ( n28703 , n19055 , n28585 );
nand ( n28704 , n27982 , n28703 );
not ( n28705 , n28704 );
or ( n28706 , n28702 , n28705 );
or ( n28707 , n1475 , n28704 );
nand ( n28708 , n28706 , n28707 );
not ( n28709 , n13594 );
not ( n28710 , n558 );
nand ( n28711 , n314 , n28710 );
not ( n28712 , n324 );
nand ( n28713 , n282 , n315 );
nor ( n28714 , n28712 , n28713 );
or ( n28715 , n314 , n28714 );
and ( n28716 , n314 , n28714 );
nor ( n28717 , n28716 , n28710 );
nand ( n28718 , n28715 , n28717 );
and ( n28719 , n28711 , n28718 );
not ( n28720 , n835 );
not ( n28721 , n28710 );
or ( n28722 , n28720 , n28721 );
nand ( n28723 , n28722 , n2 );
nor ( n28724 , n28719 , n28723 );
not ( n28725 , n128 );
not ( n28726 , n1708 );
or ( n28727 , n28725 , n28726 );
and ( n28728 , n358 , n25283 );
not ( n28729 , n358 );
not ( n28730 , n28250 );
and ( n28731 , n28729 , n28730 );
or ( n28732 , n1841 , n28249 );
buf ( n28733 , n20632 );
nand ( n28734 , n28732 , n28733 );
nor ( n28735 , n28731 , n28734 );
nor ( n28736 , n28728 , n28735 );
or ( n28737 , n1708 , n28736 );
nand ( n28738 , n28727 , n28737 );
not ( n28739 , n127 );
not ( n28740 , n1708 );
or ( n28741 , n28739 , n28740 );
and ( n28742 , n359 , n28157 );
not ( n28743 , n359 );
not ( n28744 , n28250 );
and ( n28745 , n28743 , n28744 );
or ( n28746 , n1845 , n28249 );
nand ( n28747 , n28746 , n28733 );
nor ( n28748 , n28745 , n28747 );
nor ( n28749 , n28742 , n28748 );
or ( n28750 , n1708 , n28749 );
nand ( n28751 , n28741 , n28750 );
not ( n28752 , n124 );
not ( n28753 , n1708 );
or ( n28754 , n28752 , n28753 );
and ( n28755 , n360 , n28157 );
not ( n28756 , n360 );
not ( n28757 , n28250 );
and ( n28758 , n28756 , n28757 );
or ( n28759 , n1838 , n28249 );
nand ( n28760 , n28759 , n28733 );
nor ( n28761 , n28758 , n28760 );
nor ( n28762 , n28755 , n28761 );
or ( n28763 , n1708 , n28762 );
nand ( n28764 , n28754 , n28763 );
not ( n28765 , n123 );
not ( n28766 , n1708 );
or ( n28767 , n28765 , n28766 );
and ( n28768 , n361 , n28157 );
not ( n28769 , n361 );
not ( n28770 , n28250 );
and ( n28771 , n28769 , n28770 );
or ( n28772 , n1846 , n28249 );
nand ( n28773 , n28772 , n28733 );
nor ( n28774 , n28771 , n28773 );
nor ( n28775 , n28768 , n28774 );
or ( n28776 , n1708 , n28775 );
nand ( n28777 , n28767 , n28776 );
not ( n28778 , n121 );
not ( n28779 , n1708 );
or ( n28780 , n28778 , n28779 );
and ( n28781 , n363 , n25283 );
not ( n28782 , n363 );
not ( n28783 , n28250 );
and ( n28784 , n28782 , n28783 );
or ( n28785 , n1840 , n28249 );
nand ( n28786 , n28785 , n28733 );
nor ( n28787 , n28784 , n28786 );
nor ( n28788 , n28781 , n28787 );
or ( n28789 , n1708 , n28788 );
nand ( n28790 , n28780 , n28789 );
not ( n28791 , n125 );
not ( n28792 , n1708 );
or ( n28793 , n28791 , n28792 );
and ( n28794 , n364 , n28157 );
not ( n28795 , n364 );
not ( n28796 , n28250 );
and ( n28797 , n28795 , n28796 );
or ( n28798 , n1843 , n28249 );
nand ( n28799 , n28798 , n28733 );
nor ( n28800 , n28797 , n28799 );
nor ( n28801 , n28794 , n28800 );
or ( n28802 , n1708 , n28801 );
nand ( n28803 , n28793 , n28802 );
not ( n28804 , n126 );
not ( n28805 , n1708 );
or ( n28806 , n28804 , n28805 );
and ( n28807 , n376 , n25283 );
not ( n28808 , n376 );
not ( n28809 , n28250 );
and ( n28810 , n28808 , n28809 );
or ( n28811 , n1842 , n28249 );
nand ( n28812 , n28811 , n28733 );
nor ( n28813 , n28810 , n28812 );
nor ( n28814 , n28807 , n28813 );
or ( n28815 , n1708 , n28814 );
nand ( n28816 , n28806 , n28815 );
not ( n28817 , n835 );
nand ( n28818 , n22477 , n2 , n28817 );
nand ( n28819 , n397 , n460 );
not ( n28820 , n28819 );
nand ( n28821 , n28820 , n403 );
not ( n28822 , n28821 );
nand ( n28823 , n404 , n28822 );
xor ( n28824 , n414 , n28823 );
nor ( n28825 , n28818 , n28824 );
nand ( n28826 , n604 , n22477 );
or ( n28827 , n604 , n20231 );
nand ( n28828 , n28827 , n1800 , n20232 );
and ( n28829 , n28826 , n28828 );
nor ( n28830 , n28829 , n834 );
not ( n28831 , n122 );
not ( n28832 , n1708 );
or ( n28833 , n28831 , n28832 );
and ( n28834 , n362 , n25283 );
not ( n28835 , n362 );
not ( n28836 , n28250 );
and ( n28837 , n28835 , n28836 );
or ( n28838 , n1847 , n28249 );
nand ( n28839 , n28838 , n28733 );
nor ( n28840 , n28837 , n28839 );
nor ( n28841 , n28834 , n28840 );
or ( n28842 , n1708 , n28841 );
nand ( n28843 , n28833 , n28842 );
not ( n28844 , n2 );
nand ( n28845 , n17150 , n17155 );
or ( n28846 , n17133 , n28845 );
not ( n28847 , n28846 );
and ( n28848 , n1856 , n28847 );
and ( n28849 , n1365 , n28846 );
nor ( n28850 , n28848 , n28849 );
nor ( n28851 , n28844 , n28850 );
not ( n28852 , n2 );
and ( n28853 , n1862 , n28847 );
and ( n28854 , n1356 , n28846 );
nor ( n28855 , n28853 , n28854 );
nor ( n28856 , n28852 , n28855 );
not ( n28857 , n2 );
and ( n28858 , n1870 , n28847 );
and ( n28859 , n1357 , n28846 );
nor ( n28860 , n28858 , n28859 );
nor ( n28861 , n28857 , n28860 );
or ( n28862 , n17967 , n28523 );
or ( n28863 , n15522 , n18928 );
nand ( n28864 , n28862 , n28863 );
or ( n28865 , n17954 , n28523 );
or ( n28866 , n15467 , n18928 );
nand ( n28867 , n28865 , n28866 );
and ( n28868 , n18 , n25250 , n25249 , n28528 );
not ( n28869 , n1185 );
and ( n28870 , n18975 , n28559 );
nand ( n28871 , n27928 , n28870 );
not ( n28872 , n28871 );
or ( n28873 , n28869 , n28872 );
or ( n28874 , n1185 , n28871 );
nand ( n28875 , n28873 , n28874 );
not ( n28876 , n19101 );
and ( n28877 , n18308 , n28876 );
nor ( n28878 , n28877 , n19099 );
not ( n28879 , n2 );
and ( n28880 , n1851 , n28847 );
and ( n28881 , n1358 , n28846 );
nor ( n28882 , n28880 , n28881 );
nor ( n28883 , n28879 , n28882 );
not ( n28884 , n28324 );
nand ( n28885 , n28884 , n1592 );
not ( n28886 , n1631 );
not ( n28887 , n1637 );
nand ( n28888 , n1646 , n1647 );
nor ( n28889 , n28887 , n28888 );
nand ( n28890 , n1635 , n28889 );
nor ( n28891 , n28886 , n28890 );
nand ( n28892 , n1650 , n28891 );
not ( n28893 , n28892 );
nand ( n28894 , n28893 , n1645 );
xor ( n28895 , n893 , n27672 );
nand ( n28896 , n1474 , n1624 );
or ( n28897 , n1474 , n1624 );
not ( n28898 , n13539 );
not ( n28899 , n19375 );
or ( n28900 , n28898 , n28899 );
nand ( n28901 , n28900 , n21636 );
nand ( n28902 , n28897 , n28901 );
and ( n28903 , n28896 , n28902 );
not ( n28904 , n2 );
nor ( n28905 , n28903 , n28904 );
not ( n28906 , n2 );
nor ( n28907 , n28906 , n14804 );
nand ( n28908 , n562 , n22477 );
not ( n28909 , n20230 );
or ( n28910 , n562 , n28909 );
nor ( n28911 , n22477 , n20231 );
nand ( n28912 , n28910 , n28911 );
and ( n28913 , n28908 , n28912 );
nor ( n28914 , n28913 , n834 );
nand ( n28915 , n324 , n28710 );
not ( n28916 , n28713 );
or ( n28917 , n324 , n28916 );
not ( n28918 , n28714 );
nand ( n28919 , n28917 , n558 , n28918 );
and ( n28920 , n28915 , n28919 );
nor ( n28921 , n28920 , n28723 );
xor ( n28922 , n1589 , n28322 );
nor ( n28923 , n1755 , n28922 );
or ( n28924 , n16912 , n28330 );
nand ( n28925 , n28924 , n28331 );
or ( n28926 , n17053 , n28341 );
nand ( n28927 , n28926 , n28342 );
or ( n28928 , n16983 , n28372 );
nand ( n28929 , n28928 , n28373 );
xor ( n28930 , n1631 , n28890 );
nor ( n28931 , n1710 , n28930 );
or ( n28932 , n16839 , n28310 );
nand ( n28933 , n28932 , n28311 );
nor ( n28934 , n20456 , n27671 );
and ( n28935 , n28934 , n894 );
not ( n28936 , n28934 );
and ( n28937 , n28936 , n21305 );
nor ( n28938 , n28935 , n28937 );
not ( n28939 , n19019 );
and ( n28940 , n18195 , n28939 );
nor ( n28941 , n28940 , n19017 );
not ( n28942 , n19809 );
and ( n28943 , n18058 , n28942 );
nor ( n28944 , n28943 , n19807 );
not ( n28945 , n19891 );
and ( n28946 , n18111 , n28945 );
nor ( n28947 , n28946 , n19889 );
or ( n28948 , n1556 , n17145 );
or ( n28949 , n18754 , n28846 );
nand ( n28950 , n1208 , n28846 );
nand ( n28951 , n28949 , n28950 , n2 );
nand ( n28952 , n17089 , n17076 );
not ( n28953 , n28952 );
not ( n28954 , n17085 );
or ( n28955 , n28953 , n28954 );
or ( n28956 , n28952 , n17085 );
nand ( n28957 , n28955 , n28956 );
nand ( n28958 , n17019 , n17006 );
not ( n28959 , n28958 );
not ( n28960 , n17015 );
or ( n28961 , n28959 , n28960 );
or ( n28962 , n28958 , n17015 );
nand ( n28963 , n28961 , n28962 );
or ( n28964 , n16853 , n28309 );
not ( n28965 , n28310 );
nand ( n28966 , n28964 , n28965 );
and ( n28967 , n27928 , n1195 );
not ( n28968 , n27928 );
and ( n28969 , n28968 , n17098 );
nor ( n28970 , n28967 , n28969 );
or ( n28971 , n17072 , n27927 );
not ( n28972 , n27928 );
nand ( n28973 , n28971 , n28972 );
or ( n28974 , n16858 , n27981 );
not ( n28975 , n27982 );
nand ( n28976 , n28974 , n28975 );
or ( n28977 , n17067 , n28340 );
not ( n28978 , n28341 );
nand ( n28979 , n28977 , n28978 );
or ( n28980 , n16997 , n28371 );
not ( n28981 , n28372 );
nand ( n28982 , n28980 , n28981 );
or ( n28983 , n16926 , n28329 );
not ( n28984 , n28330 );
nand ( n28985 , n28983 , n28984 );
and ( n28986 , n27917 , n1303 );
not ( n28987 , n27917 );
and ( n28988 , n28987 , n16928 );
nor ( n28989 , n28986 , n28988 );
and ( n28990 , n27886 , n1325 );
not ( n28991 , n27886 );
and ( n28992 , n28991 , n16999 );
nor ( n28993 , n28990 , n28992 );
or ( n28994 , n17002 , n27885 );
not ( n28995 , n27886 );
nand ( n28996 , n28994 , n28995 );
not ( n28997 , n21647 );
nor ( n28998 , n26830 , n28997 );
and ( n28999 , n28998 , n15599 , n26829 );
nor ( n29000 , n889 , n1608 );
nor ( n29001 , n28999 , n29000 );
and ( n29002 , n941 , n942 , n943 , n949 );
and ( n29003 , n945 , n885 , n959 );
nand ( n29004 , n29002 , n29003 , n957 , n963 );
nand ( n29005 , n960 , n961 , n940 , n962 );
nand ( n29006 , n886 , n946 , n944 , n999 );
nor ( n29007 , n29004 , n29005 , n29006 );
or ( n29008 , n958 , n29007 );
and ( n29009 , n887 , n965 , n966 , n972 );
and ( n29010 , n1008 , n983 , n987 );
nand ( n29011 , n29009 , n29010 , n980 , n1009 );
nand ( n29012 , n881 , n967 , n964 , n969 );
nand ( n29013 , n984 , n985 , n968 , n986 );
nor ( n29014 , n29011 , n29012 , n29013 );
or ( n29015 , n982 , n29014 );
or ( n29016 , n18385 , n28846 );
nand ( n29017 , n1187 , n28846 );
nand ( n29018 , n29016 , n29017 , n2 );
nor ( n29019 , n1747 , n1748 );
and ( n29020 , n1044 , n1419 );
nor ( n29021 , n29020 , n1746 );
and ( n29022 , n1030 , n1450 );
and ( n29023 , n1116 , n1448 );
nor ( n29024 , n29022 , n29023 );
nand ( n29025 , n29021 , n29024 );
nor ( n29026 , n1745 , n29025 );
and ( n29027 , n857 , n1451 );
and ( n29028 , n773 , n1420 );
and ( n29029 , n1106 , n1416 );
nor ( n29030 , n29027 , n29028 , n29029 );
and ( n29031 , n1115 , n1452 );
and ( n29032 , n915 , n1449 );
and ( n29033 , n265 , n1418 );
nor ( n29034 , n29031 , n29032 , n29033 );
nand ( n29035 , n29019 , n29026 , n29030 , n29034 );
nor ( n29036 , n1742 , n1749 );
and ( n29037 , n1116 , n1454 );
nor ( n29038 , n29037 , n1740 );
and ( n29039 , n1030 , n1457 );
and ( n29040 , n1044 , n1456 );
nor ( n29041 , n29039 , n29040 );
nand ( n29042 , n29038 , n29041 );
nor ( n29043 , n1741 , n29042 );
and ( n29044 , n1106 , n1459 );
and ( n29045 , n857 , n1458 );
and ( n29046 , n773 , n1453 );
nor ( n29047 , n29044 , n29045 , n29046 );
and ( n29048 , n1115 , n1468 );
and ( n29049 , n265 , n1455 );
and ( n29050 , n915 , n1417 );
nor ( n29051 , n29048 , n29049 , n29050 );
nand ( n29052 , n29036 , n29043 , n29047 , n29051 );
or ( n29053 , n18380 , n28846 );
nand ( n29054 , n1359 , n28846 );
nand ( n29055 , n29053 , n29054 , n2 );
not ( n29056 , n18830 );
nor ( n29057 , n855 , n1487 );
not ( n29058 , n749 );
nand ( n29059 , n29057 , n29058 , n18845 );
nor ( n29060 , n29056 , n29059 , n462 , n674 );
not ( n29061 , n29060 );
not ( n29062 , n409 );
not ( n29063 , n482 );
not ( n29064 , n484 );
nand ( n29065 , n29062 , n29063 , n29064 , n18819 );
nor ( n29066 , n29061 , n29065 , n329 , n347 );
and ( n29067 , n27982 , n1285 );
not ( n29068 , n27982 );
and ( n29069 , n29068 , n16855 );
nor ( n29070 , n29067 , n29069 );
not ( n29071 , n20632 );
or ( n29072 , n29071 , n14572 );
nand ( n29073 , n29072 , n14593 );
and ( n29074 , n20639 , n29073 );
not ( n29075 , n20633 );
and ( n29076 , n367 , n29075 );
nor ( n29077 , n29074 , n29076 );
nor ( n29078 , n20652 , n29077 );
or ( n29079 , n18473 , n28846 );
nand ( n29080 , n1360 , n28846 );
nand ( n29081 , n29079 , n29080 , n2 );
or ( n29082 , n16931 , n27916 );
not ( n29083 , n27917 );
nand ( n29084 , n29082 , n29083 );
not ( n29085 , n19995 );
nand ( n29086 , n29085 , n879 );
or ( n29087 , n366 , n19995 );
and ( n29088 , n29086 , n29087 );
or ( n29089 , n26982 , n29088 );
or ( n29090 , n19984 , n29087 );
or ( n29091 , n13664 , n367 );
nand ( n29092 , n29089 , n29090 , n29091 );
not ( n29093 , n1771 );
or ( n29094 , n15203 , n167 );
buf ( n29095 , n29094 );
not ( n29096 , n29095 );
or ( n29097 , n29093 , n29096 );
buf ( n29098 , n29094 );
not ( n29099 , n29098 );
nand ( n29100 , n124 , n29099 );
nand ( n29101 , n29097 , n29100 );
nand ( n29102 , n19071 , n19038 , n19025 , n28703 );
and ( n29103 , n19063 , n29102 );
not ( n29104 , n1772 );
not ( n29105 , n29095 );
or ( n29106 , n29104 , n29105 );
not ( n29107 , n29098 );
nand ( n29108 , n98 , n29107 );
nand ( n29109 , n29106 , n29108 );
not ( n29110 , n1793 );
not ( n29111 , n29095 );
or ( n29112 , n29110 , n29111 );
nand ( n29113 , n117 , n29107 );
nand ( n29114 , n29112 , n29113 );
not ( n29115 , n1792 );
not ( n29116 , n29095 );
or ( n29117 , n29115 , n29116 );
not ( n29118 , n29098 );
nand ( n29119 , n113 , n29118 );
nand ( n29120 , n29117 , n29119 );
not ( n29121 , n1791 );
not ( n29122 , n29095 );
or ( n29123 , n29121 , n29122 );
not ( n29124 , n29098 );
nand ( n29125 , n116 , n29124 );
nand ( n29126 , n29123 , n29125 );
not ( n29127 , n1790 );
not ( n29128 , n29095 );
or ( n29129 , n29127 , n29128 );
nand ( n29130 , n103 , n29118 );
nand ( n29131 , n29129 , n29130 );
not ( n29132 , n1789 );
not ( n29133 , n29095 );
or ( n29134 , n29132 , n29133 );
nand ( n29135 , n115 , n29118 );
nand ( n29136 , n29134 , n29135 );
not ( n29137 , n1788 );
not ( n29138 , n29095 );
or ( n29139 , n29137 , n29138 );
nand ( n29140 , n106 , n29124 );
nand ( n29141 , n29139 , n29140 );
not ( n29142 , n1787 );
not ( n29143 , n29095 );
or ( n29144 , n29142 , n29143 );
nand ( n29145 , n121 , n29118 );
nand ( n29146 , n29144 , n29145 );
not ( n29147 , n1786 );
not ( n29148 , n29095 );
or ( n29149 , n29147 , n29148 );
nand ( n29150 , n111 , n29124 );
nand ( n29151 , n29149 , n29150 );
not ( n29152 , n1785 );
not ( n29153 , n29095 );
or ( n29154 , n29152 , n29153 );
nand ( n29155 , n112 , n29118 );
nand ( n29156 , n29154 , n29155 );
not ( n29157 , n1784 );
not ( n29158 , n29095 );
or ( n29159 , n29157 , n29158 );
nand ( n29160 , n108 , n29118 );
nand ( n29161 , n29159 , n29160 );
not ( n29162 , n1783 );
not ( n29163 , n29095 );
or ( n29164 , n29162 , n29163 );
nand ( n29165 , n107 , n29118 );
nand ( n29166 , n29164 , n29165 );
xor ( n29167 , n404 , n28821 );
nor ( n29168 , n28818 , n29167 );
nand ( n29169 , n366 , n27396 );
not ( n29170 , n14574 );
nand ( n29171 , n29170 , n14572 , n28394 );
and ( n29172 , n29169 , n29171 );
nor ( n29173 , n29172 , n20652 );
not ( n29174 , n1782 );
not ( n29175 , n29095 );
or ( n29176 , n29174 , n29175 );
nand ( n29177 , n119 , n29107 );
nand ( n29178 , n29176 , n29177 );
not ( n29179 , n1781 );
not ( n29180 , n29095 );
or ( n29181 , n29179 , n29180 );
nand ( n29182 , n99 , n29124 );
nand ( n29183 , n29181 , n29182 );
not ( n29184 , n1780 );
not ( n29185 , n29095 );
or ( n29186 , n29184 , n29185 );
nand ( n29187 , n127 , n29118 );
nand ( n29188 , n29186 , n29187 );
not ( n29189 , n1779 );
not ( n29190 , n29095 );
or ( n29191 , n29189 , n29190 );
nand ( n29192 , n128 , n29099 );
nand ( n29193 , n29191 , n29192 );
not ( n29194 , n28578 );
nand ( n29195 , n29194 , n19743 , n19801 , n19774 );
and ( n29196 , n19772 , n29195 );
not ( n29197 , n28533 );
nand ( n29198 , n29197 , n19883 , n19826 , n19857 );
and ( n29199 , n19855 , n29198 );
nor ( n29200 , n20570 , n20617 );
not ( n29201 , n20456 );
not ( n29202 , n916 );
nand ( n29203 , n890 , n29202 );
not ( n29204 , n29203 );
nand ( n29205 , n29201 , n894 , n895 , n29204 );
not ( n29206 , n912 );
nor ( n29207 , n29205 , n29206 , n917 );
not ( n29208 , n17082 );
nand ( n29209 , n17080 , n17083 );
not ( n29210 , n29209 );
or ( n29211 , n29208 , n29210 );
or ( n29212 , n17082 , n29209 );
nand ( n29213 , n29211 , n29212 );
not ( n29214 , n17012 );
nand ( n29215 , n17010 , n17013 );
not ( n29216 , n29215 );
or ( n29217 , n29214 , n29216 );
or ( n29218 , n17012 , n29215 );
nand ( n29219 , n29217 , n29218 );
not ( n29220 , n16942 );
nand ( n29221 , n16939 , n16940 );
not ( n29222 , n29221 );
or ( n29223 , n29220 , n29222 );
or ( n29224 , n16942 , n29221 );
nand ( n29225 , n29223 , n29224 );
not ( n29226 , n16869 );
nand ( n29227 , n16866 , n16867 );
not ( n29228 , n29227 );
or ( n29229 , n29226 , n29228 );
or ( n29230 , n16869 , n29227 );
nand ( n29231 , n29229 , n29230 );
not ( n29232 , n1761 );
not ( n29233 , n29095 );
or ( n29234 , n29232 , n29233 );
nand ( n29235 , n126 , n29107 );
nand ( n29236 , n29234 , n29235 );
not ( n29237 , n1762 );
not ( n29238 , n29095 );
or ( n29239 , n29237 , n29238 );
nand ( n29240 , n97 , n29107 );
nand ( n29241 , n29239 , n29240 );
not ( n29242 , n1763 );
not ( n29243 , n29095 );
or ( n29244 , n29242 , n29243 );
nand ( n29245 , n100 , n29099 );
nand ( n29246 , n29244 , n29245 );
not ( n29247 , n1764 );
not ( n29248 , n29095 );
or ( n29249 , n29247 , n29248 );
nand ( n29250 , n122 , n29099 );
nand ( n29251 , n29249 , n29250 );
not ( n29252 , n1765 );
not ( n29253 , n29095 );
or ( n29254 , n29252 , n29253 );
nand ( n29255 , n105 , n29124 );
nand ( n29256 , n29254 , n29255 );
not ( n29257 , n1767 );
not ( n29258 , n29095 );
or ( n29259 , n29257 , n29258 );
nand ( n29260 , n109 , n29107 );
nand ( n29261 , n29259 , n29260 );
not ( n29262 , n1768 );
not ( n29263 , n29095 );
or ( n29264 , n29262 , n29263 );
nand ( n29265 , n104 , n29107 );
nand ( n29266 , n29264 , n29265 );
not ( n29267 , n1769 );
not ( n29268 , n29095 );
or ( n29269 , n29267 , n29268 );
nand ( n29270 , n110 , n29099 );
nand ( n29271 , n29269 , n29270 );
not ( n29272 , n1770 );
not ( n29273 , n29095 );
or ( n29274 , n29272 , n29273 );
nand ( n29275 , n118 , n29124 );
nand ( n29276 , n29274 , n29275 );
not ( n29277 , n1773 );
not ( n29278 , n29095 );
or ( n29279 , n29277 , n29278 );
nand ( n29280 , n101 , n29099 );
nand ( n29281 , n29279 , n29280 );
not ( n29282 , n1774 );
not ( n29283 , n29095 );
or ( n29284 , n29282 , n29283 );
nand ( n29285 , n125 , n29124 );
nand ( n29286 , n29284 , n29285 );
not ( n29287 , n1775 );
not ( n29288 , n29095 );
or ( n29289 , n29287 , n29288 );
nand ( n29290 , n123 , n29107 );
nand ( n29291 , n29289 , n29290 );
not ( n29292 , n1776 );
not ( n29293 , n29095 );
or ( n29294 , n29292 , n29293 );
nand ( n29295 , n120 , n29099 );
nand ( n29296 , n29294 , n29295 );
not ( n29297 , n1777 );
not ( n29298 , n29095 );
or ( n29299 , n29297 , n29298 );
nand ( n29300 , n102 , n29124 );
nand ( n29301 , n29299 , n29300 );
not ( n29302 , n1778 );
not ( n29303 , n29095 );
or ( n29304 , n29302 , n29303 );
nand ( n29305 , n114 , n29099 );
nand ( n29306 , n29304 , n29305 );
not ( n29307 , n18954 );
nand ( n29308 , n18986 , n29307 , n18958 , n28870 );
and ( n29309 , n18983 , n29308 );
not ( n29310 , n28891 );
not ( n29311 , n1593 );
or ( n29312 , n1595 , n1601 );
nor ( n29313 , n29311 , n29312 , n1605 , n1592 );
not ( n29314 , n29313 );
and ( n29315 , n28318 , n13539 );
and ( n29316 , n1589 , n1608 );
nor ( n29317 , n29315 , n29316 );
and ( n29318 , n1594 , n1608 );
nor ( n29319 , n1594 , n1608 );
nor ( n29320 , n29318 , n29319 );
and ( n29321 , n1607 , n13539 );
not ( n29322 , n1607 );
and ( n29323 , n1608 , n29322 );
nor ( n29324 , n29321 , n29323 );
nor ( n29325 , n29314 , n29317 , n29320 , n29324 );
and ( n29326 , n920 , n20028 );
and ( n29327 , n922 , n892 , n29326 );
nor ( n29328 , n412 , n420 );
not ( n29329 , n29328 );
nand ( n29330 , n419 , n421 , n422 , n16135 );
nor ( n29331 , n29329 , n29330 , n418 , n1663 );
not ( n29332 , n20156 );
or ( n29333 , n20634 , n29332 );
not ( n29334 , n387 );
nand ( n29335 , n29333 , n29334 );
and ( n29336 , n20633 , n19981 );
not ( n29337 , n20633 );
and ( n29338 , n29337 , n386 );
nor ( n29339 , n29336 , n29338 );
nor ( n29340 , n20652 , n29339 );
not ( n29341 , n1637 );
nor ( n29342 , n29341 , n1635 );
not ( n29343 , n29342 );
nor ( n29344 , n29343 , n1645 , n1646 , n1648 );
not ( n29345 , n29344 );
and ( n29346 , n1650 , n13539 );
not ( n29347 , n1650 );
and ( n29348 , n29347 , n1608 );
nor ( n29349 , n29346 , n29348 );
and ( n29350 , n13539 , n28886 );
and ( n29351 , n1608 , n1631 );
nor ( n29352 , n29350 , n29351 );
and ( n29353 , n1608 , n1647 );
nor ( n29354 , n1608 , n1647 );
nor ( n29355 , n29353 , n29354 );
nor ( n29356 , n29345 , n29349 , n29352 , n29355 );
not ( n29357 , n912 );
not ( n29358 , n27670 );
not ( n29359 , n29358 );
or ( n29360 , n29357 , n29359 );
or ( n29361 , n912 , n29358 );
nand ( n29362 , n29360 , n29361 );
nand ( n29363 , n603 , n22477 );
or ( n29364 , n598 , n603 );
nand ( n29365 , n29364 , n20230 , n1800 );
and ( n29366 , n29363 , n29365 );
nor ( n29367 , n29366 , n834 );
not ( n29368 , n123 );
nand ( n29369 , n167 , n1230 );
not ( n29370 , n29369 );
not ( n29371 , n29370 );
or ( n29372 , n29368 , n29371 );
buf ( n29373 , n29369 );
nand ( n29374 , n1725 , n29373 );
nand ( n29375 , n29372 , n29374 );
not ( n29376 , n2 );
nand ( n29377 , n1559 , n1824 );
and ( n29378 , n29377 , n1005 );
not ( n29379 , n29377 );
and ( n29380 , n29379 , n178 );
nor ( n29381 , n29378 , n29380 );
nor ( n29382 , n29376 , n29381 );
not ( n29383 , n2 );
nand ( n29384 , n1588 , n1824 );
and ( n29385 , n29384 , n1102 );
not ( n29386 , n29384 );
and ( n29387 , n29386 , n178 );
nor ( n29388 , n29385 , n29387 );
nor ( n29389 , n29383 , n29388 );
and ( n29390 , n1187 , n1358 );
not ( n29391 , n1187 );
not ( n29392 , n1358 );
and ( n29393 , n29391 , n29392 );
nor ( n29394 , n29390 , n29393 );
and ( n29395 , n1359 , n1356 );
not ( n29396 , n1359 );
and ( n29397 , n29396 , n15319 );
nor ( n29398 , n29395 , n29397 );
and ( n29399 , n1360 , n1357 );
not ( n29400 , n1360 );
and ( n29401 , n29400 , n13518 );
nor ( n29402 , n29399 , n29401 );
xor ( n29403 , n1208 , n1365 );
nand ( n29404 , n29394 , n29398 , n29402 , n29403 );
not ( n29405 , n2 );
nand ( n29406 , n1588 , n1827 );
and ( n29407 , n29406 , n1097 );
not ( n29408 , n29406 );
and ( n29409 , n29408 , n186 );
nor ( n29410 , n29407 , n29409 );
nor ( n29411 , n29405 , n29410 );
not ( n29412 , n2 );
and ( n29413 , n29406 , n1096 );
not ( n29414 , n29406 );
and ( n29415 , n29414 , n193 );
nor ( n29416 , n29413 , n29415 );
nor ( n29417 , n29412 , n29416 );
nand ( n29418 , n282 , n28710 );
or ( n29419 , n282 , n315 );
nand ( n29420 , n29419 , n28713 , n558 );
and ( n29421 , n29418 , n29420 );
nor ( n29422 , n29421 , n28723 );
xor ( n29423 , n403 , n28819 );
nor ( n29424 , n28818 , n29423 );
not ( n29425 , n2 );
nand ( n29426 , n1559 , n1827 );
and ( n29427 , n29426 , n991 );
not ( n29428 , n29426 );
and ( n29429 , n29428 , n186 );
nor ( n29430 , n29427 , n29429 );
nor ( n29431 , n29425 , n29430 );
not ( n29432 , n2 );
nand ( n29433 , n1576 , n1824 );
and ( n29434 , n29433 , n1068 );
not ( n29435 , n29433 );
and ( n29436 , n29435 , n185 );
nor ( n29437 , n29434 , n29436 );
nor ( n29438 , n29432 , n29437 );
not ( n29439 , n2 );
and ( n29440 , n29433 , n1071 );
not ( n29441 , n29433 );
and ( n29442 , n29441 , n178 );
nor ( n29443 , n29440 , n29442 );
nor ( n29444 , n29439 , n29443 );
not ( n29445 , n2 );
and ( n29446 , n29384 , n1098 );
not ( n29447 , n29384 );
and ( n29448 , n29447 , n185 );
nor ( n29449 , n29446 , n29448 );
nor ( n29450 , n29445 , n29449 );
not ( n29451 , n2 );
nand ( n29452 , n1609 , n1827 );
and ( n29453 , n29452 , n1122 );
not ( n29454 , n29452 );
and ( n29455 , n29454 , n186 );
nor ( n29456 , n29453 , n29455 );
nor ( n29457 , n29451 , n29456 );
not ( n29458 , n2 );
nand ( n29459 , n1609 , n1824 );
and ( n29460 , n29459 , n1143 );
not ( n29461 , n29459 );
and ( n29462 , n29461 , n178 );
nor ( n29463 , n29460 , n29462 );
nor ( n29464 , n29458 , n29463 );
not ( n29465 , n2 );
and ( n29466 , n29377 , n992 );
not ( n29467 , n29377 );
and ( n29468 , n29467 , n185 );
nor ( n29469 , n29466 , n29468 );
nor ( n29470 , n29465 , n29469 );
not ( n29471 , n109 );
not ( n29472 , n29370 );
or ( n29473 , n29471 , n29472 );
nand ( n29474 , n1692 , n29373 );
nand ( n29475 , n29473 , n29474 );
not ( n29476 , n127 );
not ( n29477 , n29370 );
or ( n29478 , n29476 , n29477 );
nand ( n29479 , n1693 , n29373 );
nand ( n29480 , n29478 , n29479 );
not ( n29481 , n121 );
not ( n29482 , n29370 );
or ( n29483 , n29481 , n29482 );
nand ( n29484 , n1704 , n29373 );
nand ( n29485 , n29483 , n29484 );
not ( n29486 , n101 );
not ( n29487 , n29370 );
or ( n29488 , n29486 , n29487 );
nand ( n29489 , n1714 , n29373 );
nand ( n29490 , n29488 , n29489 );
not ( n29491 , n125 );
not ( n29492 , n29370 );
or ( n29493 , n29491 , n29492 );
nand ( n29494 , n1715 , n29373 );
nand ( n29495 , n29493 , n29494 );
not ( n29496 , n128 );
not ( n29497 , n29370 );
or ( n29498 , n29496 , n29497 );
nand ( n29499 , n1716 , n29373 );
nand ( n29500 , n29498 , n29499 );
not ( n29501 , n116 );
not ( n29502 , n29370 );
or ( n29503 , n29501 , n29502 );
nand ( n29504 , n1717 , n29373 );
nand ( n29505 , n29503 , n29504 );
not ( n29506 , n126 );
not ( n29507 , n29370 );
or ( n29508 , n29506 , n29507 );
nand ( n29509 , n1718 , n29373 );
nand ( n29510 , n29508 , n29509 );
not ( n29511 , n120 );
not ( n29512 , n29370 );
or ( n29513 , n29511 , n29512 );
nand ( n29514 , n1719 , n29373 );
nand ( n29515 , n29513 , n29514 );
not ( n29516 , n110 );
not ( n29517 , n29370 );
or ( n29518 , n29516 , n29517 );
nand ( n29519 , n1720 , n29373 );
nand ( n29520 , n29518 , n29519 );
not ( n29521 , n100 );
not ( n29522 , n29370 );
or ( n29523 , n29521 , n29522 );
nand ( n29524 , n1721 , n29373 );
nand ( n29525 , n29523 , n29524 );
not ( n29526 , n114 );
not ( n29527 , n29370 );
or ( n29528 , n29526 , n29527 );
nand ( n29529 , n1722 , n29373 );
nand ( n29530 , n29528 , n29529 );
not ( n29531 , n122 );
not ( n29532 , n29370 );
or ( n29533 , n29531 , n29532 );
nand ( n29534 , n1724 , n29373 );
nand ( n29535 , n29533 , n29534 );
not ( n29536 , n119 );
not ( n29537 , n29370 );
or ( n29538 , n29536 , n29537 );
nand ( n29539 , n1726 , n29373 );
nand ( n29540 , n29538 , n29539 );
not ( n29541 , n108 );
not ( n29542 , n29370 );
or ( n29543 , n29541 , n29542 );
nand ( n29544 , n1727 , n29373 );
nand ( n29545 , n29543 , n29544 );
not ( n29546 , n113 );
not ( n29547 , n29370 );
or ( n29548 , n29546 , n29547 );
nand ( n29549 , n1729 , n29373 );
nand ( n29550 , n29548 , n29549 );
not ( n29551 , n105 );
not ( n29552 , n29370 );
or ( n29553 , n29551 , n29552 );
nand ( n29554 , n1730 , n29373 );
nand ( n29555 , n29553 , n29554 );
not ( n29556 , n111 );
not ( n29557 , n29370 );
or ( n29558 , n29556 , n29557 );
nand ( n29559 , n1732 , n29373 );
nand ( n29560 , n29558 , n29559 );
not ( n29561 , n124 );
not ( n29562 , n29370 );
or ( n29563 , n29561 , n29562 );
nand ( n29564 , n1735 , n29373 );
nand ( n29565 , n29563 , n29564 );
not ( n29566 , n99 );
not ( n29567 , n29370 );
or ( n29568 , n29566 , n29567 );
nand ( n29569 , n1738 , n29373 );
nand ( n29570 , n29568 , n29569 );
not ( n29571 , n118 );
not ( n29572 , n29370 );
or ( n29573 , n29571 , n29572 );
nand ( n29574 , n1739 , n29373 );
nand ( n29575 , n29573 , n29574 );
not ( n29576 , n117 );
not ( n29577 , n29370 );
or ( n29578 , n29576 , n29577 );
nand ( n29579 , n1743 , n29373 );
nand ( n29580 , n29578 , n29579 );
not ( n29581 , n115 );
not ( n29582 , n29370 );
or ( n29583 , n29581 , n29582 );
nand ( n29584 , n1744 , n29373 );
nand ( n29585 , n29583 , n29584 );
not ( n29586 , n2 );
and ( n29587 , n29426 , n990 );
not ( n29588 , n29426 );
and ( n29589 , n29588 , n193 );
nor ( n29590 , n29587 , n29589 );
nor ( n29591 , n29586 , n29590 );
not ( n29592 , n1593 );
not ( n29593 , n28320 );
and ( n29594 , n29592 , n29593 );
and ( n29595 , n1593 , n28320 );
nor ( n29596 , n29594 , n29595 );
nor ( n29597 , n1755 , n29596 );
not ( n29598 , n107 );
not ( n29599 , n29370 );
or ( n29600 , n29598 , n29599 );
nand ( n29601 , n1706 , n29373 );
nand ( n29602 , n29600 , n29601 );
not ( n29603 , n102 );
not ( n29604 , n29370 );
or ( n29605 , n29603 , n29604 );
nand ( n29606 , n1713 , n29373 );
nand ( n29607 , n29605 , n29606 );
not ( n29608 , n1637 );
not ( n29609 , n28888 );
and ( n29610 , n29608 , n29609 );
and ( n29611 , n1637 , n28888 );
nor ( n29612 , n29610 , n29611 );
nor ( n29613 , n1710 , n29612 );
not ( n29614 , n112 );
not ( n29615 , n29370 );
or ( n29616 , n29614 , n29615 );
nand ( n29617 , n1734 , n29373 );
nand ( n29618 , n29616 , n29617 );
nor ( n29619 , n408 , n426 );
not ( n29620 , n424 );
nor ( n29621 , n29620 , n436 );
nand ( n29622 , n29619 , n29621 , n425 , n437 );
nor ( n29623 , n29622 , n423 , n427 );
not ( n29624 , n2 );
nand ( n29625 , n1576 , n1827 );
and ( n29626 , n29625 , n1070 );
not ( n29627 , n29625 );
and ( n29628 , n29627 , n186 );
nor ( n29629 , n29626 , n29628 );
nor ( n29630 , n29624 , n29629 );
not ( n29631 , n106 );
not ( n29632 , n29370 );
or ( n29633 , n29631 , n29632 );
nand ( n29634 , n1728 , n29373 );
nand ( n29635 , n29633 , n29634 );
not ( n29636 , n2 );
and ( n29637 , n29459 , n1123 );
not ( n29638 , n29459 );
and ( n29639 , n29638 , n185 );
nor ( n29640 , n29637 , n29639 );
nor ( n29641 , n29636 , n29640 );
not ( n29642 , n2 );
and ( n29643 , n29452 , n1121 );
not ( n29644 , n29452 );
and ( n29645 , n29644 , n193 );
nor ( n29646 , n29643 , n29645 );
nor ( n29647 , n29642 , n29646 );
not ( n29648 , n2 );
and ( n29649 , n29625 , n1067 );
not ( n29650 , n29625 );
and ( n29651 , n29650 , n193 );
nor ( n29652 , n29649 , n29651 );
nor ( n29653 , n29648 , n29652 );
not ( n29654 , n97 );
not ( n29655 , n29370 );
or ( n29656 , n29654 , n29655 );
nand ( n29657 , n1702 , n29373 );
nand ( n29658 , n29656 , n29657 );
not ( n29659 , n98 );
not ( n29660 , n29370 );
or ( n29661 , n29659 , n29660 );
nand ( n29662 , n1703 , n29373 );
nand ( n29663 , n29661 , n29662 );
not ( n29664 , n103 );
not ( n29665 , n29370 );
or ( n29666 , n29664 , n29665 );
nand ( n29667 , n1731 , n29373 );
nand ( n29668 , n29666 , n29667 );
not ( n29669 , n104 );
not ( n29670 , n29370 );
or ( n29671 , n29669 , n29670 );
or ( n29672 , n13168 , n29370 );
nand ( n29673 , n29671 , n29672 );
and ( n29674 , n598 , n22477 );
not ( n29675 , n598 );
and ( n29676 , n29675 , n1800 );
nor ( n29677 , n29674 , n29676 );
nor ( n29678 , n834 , n29677 );
not ( n29679 , n2 );
not ( n29680 , n1825 );
and ( n29681 , n1691 , n29680 );
nor ( n29682 , n29681 , n68 );
nor ( n29683 , n29679 , n29682 );
not ( n29684 , n2 );
not ( n29685 , n1821 );
and ( n29686 , n194 , n29685 );
nor ( n29687 , n29686 , n222 );
nor ( n29688 , n29684 , n29687 );
and ( n29689 , n257 , n1536 );
and ( n29690 , n1177 , n1505 );
and ( n29691 , n1032 , n1504 );
nor ( n29692 , n29689 , n29690 , n29691 );
and ( n29693 , n721 , n1529 );
and ( n29694 , n1164 , n1503 );
nor ( n29695 , n29693 , n29694 );
and ( n29696 , n243 , n1535 );
and ( n29697 , n1099 , n1504 );
nor ( n29698 , n29696 , n29697 );
nand ( n29699 , n29692 , n29695 , n29698 );
not ( n29700 , n2 );
not ( n29701 , n1859 );
and ( n29702 , n1737 , n29701 );
nor ( n29703 , n29702 , n840 );
nor ( n29704 , n29700 , n29703 );
and ( n29705 , n1119 , n1481 );
and ( n29706 , n260 , n1478 );
and ( n29707 , n1020 , n1493 );
nor ( n29708 , n29705 , n29706 , n29707 );
and ( n29709 , n1166 , n1491 );
and ( n29710 , n746 , n1488 );
nor ( n29711 , n29709 , n29710 );
and ( n29712 , n247 , n1519 );
and ( n29713 , n1088 , n1493 );
nor ( n29714 , n29712 , n29713 );
nand ( n29715 , n29708 , n29711 , n29714 );
and ( n29716 , n259 , n1525 );
and ( n29717 , n1094 , n1515 );
and ( n29718 , n1033 , n1514 );
nor ( n29719 , n29716 , n29717 , n29718 );
and ( n29720 , n1087 , n1514 );
and ( n29721 , n245 , n1513 );
nor ( n29722 , n29720 , n29721 );
and ( n29723 , n744 , n1533 );
and ( n29724 , n1120 , n1512 );
nor ( n29725 , n29723 , n29724 );
nand ( n29726 , n29719 , n29722 , n29725 );
not ( n29727 , n2 );
not ( n29728 , n1818 );
and ( n29729 , n1685 , n29728 );
nor ( n29730 , n29729 , n70 );
nor ( n29731 , n29727 , n29730 );
not ( n29732 , n2 );
and ( n29733 , n381 , n28817 );
and ( n29734 , n835 , n1173 );
nor ( n29735 , n29733 , n29734 );
nor ( n29736 , n29732 , n29735 );
not ( n29737 , n2 );
and ( n29738 , n384 , n28817 );
and ( n29739 , n835 , n1446 );
nor ( n29740 , n29738 , n29739 );
nor ( n29741 , n29737 , n29740 );
xnor ( n29742 , n397 , n460 );
nor ( n29743 , n28818 , n29742 );
not ( n29744 , n2 );
and ( n29745 , n399 , n28817 );
and ( n29746 , n835 , n1170 );
nor ( n29747 , n29745 , n29746 );
nor ( n29748 , n29744 , n29747 );
nor ( n29749 , n460 , n28818 );
not ( n29750 , n2 );
and ( n29751 , n402 , n28817 );
and ( n29752 , n835 , n1146 );
nor ( n29753 , n29751 , n29752 );
nor ( n29754 , n29750 , n29753 );
not ( n29755 , n2 );
and ( n29756 , n400 , n28817 );
and ( n29757 , n835 , n1169 );
nor ( n29758 , n29756 , n29757 );
nor ( n29759 , n29755 , n29758 );
not ( n29760 , n2 );
and ( n29761 , n401 , n28817 );
and ( n29762 , n835 , n1178 );
nor ( n29763 , n29761 , n29762 );
nor ( n29764 , n29760 , n29763 );
not ( n29765 , n2 );
and ( n29766 , n398 , n28817 );
and ( n29767 , n835 , n1168 );
nor ( n29768 , n29766 , n29767 );
nor ( n29769 , n29765 , n29768 );
not ( n29770 , n2 );
and ( n29771 , n392 , n28817 );
and ( n29772 , n835 , n1172 );
nor ( n29773 , n29771 , n29772 );
nor ( n29774 , n29770 , n29773 );
not ( n29775 , n2 );
and ( n29776 , n382 , n28817 );
and ( n29777 , n835 , n1442 );
nor ( n29778 , n29776 , n29777 );
nor ( n29779 , n29775 , n29778 );
not ( n29780 , n2 );
and ( n29781 , n380 , n28817 );
and ( n29782 , n835 , n1171 );
nor ( n29783 , n29781 , n29782 );
nor ( n29784 , n29780 , n29783 );
not ( n29785 , n2 );
and ( n29786 , n379 , n28817 );
and ( n29787 , n835 , n1447 );
nor ( n29788 , n29786 , n29787 );
nor ( n29789 , n29785 , n29788 );
or ( n29790 , n16861 , n27979 );
nand ( n29791 , n29790 , n27980 );
not ( n29792 , n2 );
not ( n29793 , n1820 );
and ( n29794 , n1690 , n29793 );
nor ( n29795 , n29794 , n71 );
nor ( n29796 , n29792 , n29795 );
not ( n29797 , n2 );
not ( n29798 , n1863 );
and ( n29799 , n1736 , n29798 );
nor ( n29800 , n29799 , n805 );
nor ( n29801 , n29797 , n29800 );
and ( n29802 , n1020 , n1540 );
and ( n29803 , n260 , n1520 );
and ( n29804 , n1119 , n1541 );
nor ( n29805 , n29802 , n29803 , n29804 );
and ( n29806 , n1166 , n1531 );
and ( n29807 , n746 , n1523 );
nor ( n29808 , n29806 , n29807 );
and ( n29809 , n1088 , n1540 );
and ( n29810 , n247 , n1537 );
nor ( n29811 , n29809 , n29810 );
nand ( n29812 , n29805 , n29808 , n29811 );
and ( n29813 , n1032 , n1509 );
and ( n29814 , n257 , n1508 );
and ( n29815 , n1177 , n1532 );
nor ( n29816 , n29813 , n29814 , n29815 );
and ( n29817 , n1164 , n1507 );
and ( n29818 , n721 , n1506 );
nor ( n29819 , n29817 , n29818 );
and ( n29820 , n243 , n1534 );
and ( n29821 , n1099 , n1509 );
nor ( n29822 , n29820 , n29821 );
nand ( n29823 , n29816 , n29819 , n29822 );
and ( n29824 , n245 , n1524 );
and ( n29825 , n1087 , n1518 );
and ( n29826 , n1094 , n1522 );
nor ( n29827 , n29824 , n29825 , n29826 );
and ( n29828 , n1033 , n1518 );
and ( n29829 , n259 , n1517 );
nor ( n29830 , n29828 , n29829 );
and ( n29831 , n744 , n1526 );
and ( n29832 , n1120 , n1516 );
nor ( n29833 , n29831 , n29832 );
nand ( n29834 , n29827 , n29830 , n29833 );
and ( n29835 , n1443 , n1485 );
and ( n29836 , n258 , n1482 );
and ( n29837 , n1021 , n1477 );
nor ( n29838 , n29835 , n29836 , n29837 );
and ( n29839 , n664 , n1510 );
and ( n29840 , n1294 , n1492 );
nor ( n29841 , n29839 , n29840 );
and ( n29842 , n244 , n1511 );
and ( n29843 , n1086 , n1477 );
nor ( n29844 , n29842 , n29843 );
nand ( n29845 , n29838 , n29841 , n29844 );
and ( n29846 , n1021 , n1483 );
and ( n29847 , n258 , n1480 );
and ( n29848 , n1443 , n1476 );
nor ( n29849 , n29846 , n29847 , n29848 );
and ( n29850 , n1086 , n1483 );
and ( n29851 , n244 , n1479 );
nor ( n29852 , n29850 , n29851 );
and ( n29853 , n664 , n1486 );
and ( n29854 , n1294 , n1484 );
nor ( n29855 , n29853 , n29854 );
nand ( n29856 , n29849 , n29852 , n29855 );
not ( n29857 , n20041 );
and ( n29858 , n1050 , n29857 );
and ( n29859 , n315 , n28710 );
not ( n29860 , n315 );
and ( n29861 , n29860 , n558 );
nor ( n29862 , n29859 , n29861 );
nor ( n29863 , n28723 , n29862 );
not ( n29864 , n2 );
not ( n29865 , n1872 );
and ( n29866 , n1712 , n29865 );
nor ( n29867 , n29866 , n842 );
nor ( n29868 , n29864 , n29867 );
not ( n29869 , n2 );
not ( n29870 , n1857 );
and ( n29871 , n1733 , n29870 );
nor ( n29872 , n29871 , n850 );
nor ( n29873 , n29869 , n29872 );
not ( n29874 , n2 );
not ( n29875 , n1823 );
and ( n29876 , n1680 , n29875 );
nor ( n29877 , n29876 , n69 );
nor ( n29878 , n29874 , n29877 );
or ( n29879 , n16934 , n27914 );
nand ( n29880 , n29879 , n27915 );
or ( n29881 , n17005 , n27883 );
nand ( n29882 , n29881 , n27884 );
or ( n29883 , n17075 , n27925 );
nand ( n29884 , n29883 , n27926 );
not ( n29885 , n13544 );
not ( n29886 , n14785 );
not ( n29887 , n2 );
nor ( n29888 , n72 , n923 );
nor ( n29889 , n1444 , n29887 , n29888 );
not ( n29890 , n915 );
not ( n29891 , n1809 );
nor ( n29892 , n29891 , n1804 );
not ( n29893 , n29892 );
and ( n29894 , n29890 , n29893 );
not ( n29895 , n2 );
or ( n29896 , n29895 , n1553 );
nor ( n29897 , n29894 , n29896 );
not ( n29898 , n1443 );
and ( n29899 , n29898 , n25670 );
nor ( n29900 , n29899 , n20582 );
and ( n29901 , n327 , n1609 );
nor ( n29902 , n29901 , n244 );
nor ( n29903 , n20582 , n29902 );
not ( n29904 , n265 );
not ( n29905 , n351 );
and ( n29906 , n29904 , n29905 );
nor ( n29907 , n29906 , n29896 );
not ( n29908 , n1044 );
not ( n29909 , n1804 );
nor ( n29910 , n29909 , n1809 );
not ( n29911 , n29910 );
and ( n29912 , n29908 , n29911 );
nor ( n29913 , n29912 , n29896 );
not ( n29914 , n1094 );
and ( n29915 , n29914 , n23598 );
nor ( n29916 , n29915 , n20569 );
not ( n29917 , n1177 );
and ( n29918 , n29917 , n23860 );
nor ( n29919 , n29918 , n20587 );
not ( n29920 , n773 );
not ( n29921 , n1022 );
and ( n29922 , n29920 , n29921 );
nor ( n29923 , n29922 , n29896 );
or ( n29924 , n17011 , n640 );
nand ( n29925 , n29924 , n17012 );
not ( n29926 , n917 );
not ( n29927 , n19915 );
or ( n29928 , n29926 , n29927 );
or ( n29929 , n917 , n19915 );
nand ( n29930 , n29928 , n29929 );
not ( n29931 , n403 );
nand ( n29932 , n404 , n414 );
nor ( n29933 , n29931 , n29932 , n460 , n397 );
or ( n29934 , n29202 , n890 );
nand ( n29935 , n29934 , n29203 );
xnor ( n29936 , n1646 , n1647 );
nor ( n29937 , n1710 , n29936 );
not ( n29938 , n857 );
not ( n29939 , n1805 );
nor ( n29940 , n29939 , n1855 );
not ( n29941 , n29940 );
and ( n29942 , n29938 , n29941 );
nor ( n29943 , n29942 , n29896 );
xnor ( n29944 , n1594 , n1595 );
nor ( n29945 , n1755 , n29944 );
or ( n29946 , n17081 , n723 );
nand ( n29947 , n29946 , n17082 );
or ( n29948 , n16941 , n539 );
nand ( n29949 , n29948 , n16942 );
not ( n29950 , n1106 );
not ( n29951 , n1672 );
and ( n29952 , n29950 , n29951 );
nor ( n29953 , n29952 , n29896 );
not ( n29954 , n1115 );
not ( n29955 , n1677 );
and ( n29956 , n29954 , n29955 );
nor ( n29957 , n29956 , n29896 );
not ( n29958 , n1116 );
not ( n29959 , n1652 );
and ( n29960 , n29958 , n29959 );
nor ( n29961 , n29960 , n29896 );
not ( n29962 , n1119 );
and ( n29963 , n29962 , n22163 );
nor ( n29964 , n29963 , n20577 );
and ( n29965 , n388 , n1609 );
nor ( n29966 , n29965 , n258 );
nor ( n29967 , n20582 , n29966 );
and ( n29968 , n388 , n1559 );
nor ( n29969 , n29968 , n259 );
nor ( n29970 , n20569 , n29969 );
and ( n29971 , n388 , n1576 );
nor ( n29972 , n29971 , n260 );
nor ( n29973 , n20577 , n29972 );
and ( n29974 , n388 , n1588 );
nor ( n29975 , n29974 , n257 );
nor ( n29976 , n20587 , n29975 );
or ( n29977 , n16868 , n829 );
nand ( n29978 , n29977 , n16869 );
and ( n29979 , n327 , n1576 );
nor ( n29980 , n29979 , n247 );
nor ( n29981 , n20577 , n29980 );
not ( n29982 , n1030 );
not ( n29983 , n1855 );
nor ( n29984 , n29983 , n1805 );
not ( n29985 , n29984 );
and ( n29986 , n29982 , n29985 );
nor ( n29987 , n29986 , n29896 );
and ( n29988 , n327 , n1559 );
nor ( n29989 , n29988 , n245 );
nor ( n29990 , n20569 , n29989 );
and ( n29991 , n327 , n1588 );
nor ( n29992 , n29991 , n243 );
nor ( n29993 , n20587 , n29992 );
nand ( n29994 , n16948 , n16935 );
and ( n29995 , n17029 , n17000 );
and ( n29996 , n16958 , n16929 );
not ( n29997 , n28889 );
nand ( n29998 , n16875 , n16862 );
not ( n29999 , n367 );
not ( n30000 , n1228 );
or ( n30001 , n29999 , n30000 );
or ( n30002 , n18845 , n1228 );
nand ( n30003 , n30001 , n30002 );
nor ( n30004 , n1176 , n1655 );
nor ( n30005 , n16258 , n30004 );
not ( n30006 , n368 );
not ( n30007 , n1228 );
or ( n30008 , n30006 , n30007 );
or ( n30009 , n18849 , n1228 );
nand ( n30010 , n30008 , n30009 );
not ( n30011 , n371 );
not ( n30012 , n1228 );
or ( n30013 , n30011 , n30012 );
or ( n30014 , n29064 , n1228 );
nand ( n30015 , n30013 , n30014 );
not ( n30016 , n370 );
not ( n30017 , n1228 );
or ( n30018 , n30016 , n30017 );
or ( n30019 , n18819 , n1228 );
nand ( n30020 , n30018 , n30019 );
not ( n30021 , n1167 );
or ( n30022 , n30021 , n1812 );
not ( n30023 , n86 );
or ( n30024 , n30023 , n87 );
nand ( n30025 , n30022 , n30024 );
or ( n30026 , n16937 , n1370 );
or ( n30027 , n16941 , n1206 );
nand ( n30028 , n30026 , n30027 );
or ( n30029 , n16864 , n1460 );
or ( n30030 , n16868 , n1412 );
nand ( n30031 , n30029 , n30030 );
nor ( n30032 , n15090 , n30004 );
nor ( n30033 , n14974 , n30004 );
or ( n30034 , n17011 , n1405 );
or ( n30035 , n17008 , n1321 );
nand ( n30036 , n30034 , n30035 );
nor ( n30037 , n15704 , n30004 );
nand ( n30038 , n15219 , n15214 );
or ( n30039 , n17081 , n1343 );
or ( n30040 , n17078 , n1342 );
nand ( n30041 , n30039 , n30040 );
and ( n30042 , n390 , n335 );
not ( n30043 , n390 );
and ( n30044 , n30043 , n292 );
or ( n30045 , n30042 , n30044 );
and ( n30046 , n3 , n122 );
not ( n30047 , n3 );
and ( n30048 , n30047 , n1433 );
or ( n30049 , n30046 , n30048 );
and ( n30050 , n3 , n124 );
not ( n30051 , n3 );
and ( n30052 , n30051 , n1415 );
or ( n30053 , n30050 , n30052 );
and ( n30054 , n390 , n360 );
not ( n30055 , n390 );
and ( n30056 , n30055 , n307 );
or ( n30057 , n30054 , n30056 );
and ( n30058 , n390 , n336 );
not ( n30059 , n390 );
and ( n30060 , n30059 , n298 );
or ( n30061 , n30058 , n30060 );
and ( n30062 , n3 , n99 );
not ( n30063 , n3 );
and ( n30064 , n30063 , n1494 );
or ( n30065 , n30062 , n30064 );
and ( n30066 , n3 , n125 );
not ( n30067 , n3 );
and ( n30068 , n30067 , n1015 );
or ( n30069 , n30066 , n30068 );
and ( n30070 , n390 , n359 );
not ( n30071 , n390 );
and ( n30072 , n30071 , n275 );
or ( n30073 , n30070 , n30072 );
and ( n30074 , n3 , n103 );
not ( n30075 , n3 );
and ( n30076 , n30075 , n1429 );
or ( n30077 , n30074 , n30076 );
and ( n30078 , n3 , n115 );
not ( n30079 , n3 );
and ( n30080 , n30079 , n1543 );
or ( n30081 , n30078 , n30080 );
and ( n30082 , n3 , n128 );
not ( n30083 , n3 );
and ( n30084 , n30083 , n1012 );
or ( n30085 , n30082 , n30084 );
and ( n30086 , n3 , n112 );
not ( n30087 , n3 );
and ( n30088 , n30087 , n1423 );
or ( n30089 , n30086 , n30088 );
and ( n30090 , n3 , n121 );
not ( n30091 , n3 );
and ( n30092 , n30091 , n1190 );
or ( n30093 , n30090 , n30092 );
and ( n30094 , n3 , n126 );
not ( n30095 , n3 );
and ( n30096 , n30095 , n1014 );
or ( n30097 , n30094 , n30096 );
and ( n30098 , n3 , n117 );
not ( n30099 , n3 );
and ( n30100 , n30099 , n1501 );
or ( n30101 , n30098 , n30100 );
not ( n30102 , n759 );
nor ( n30103 , n30102 , n385 , n483 );
and ( n30104 , n3 , n123 );
not ( n30105 , n3 );
and ( n30106 , n30105 , n1432 );
or ( n30107 , n30104 , n30106 );
not ( n30108 , n15580 );
and ( n30109 , n390 , n377 );
not ( n30110 , n390 );
and ( n30111 , n30110 , n310 );
or ( n30112 , n30109 , n30111 );
and ( n30113 , n1228 , n350 );
not ( n30114 , n1228 );
and ( n30115 , n30114 , n462 );
or ( n30116 , n30113 , n30115 );
and ( n30117 , n390 , n376 );
not ( n30118 , n390 );
and ( n30119 , n30118 , n304 );
or ( n30120 , n30117 , n30119 );
and ( n30121 , n1228 , n369 );
not ( n30122 , n1228 );
and ( n30123 , n30122 , n749 );
or ( n30124 , n30121 , n30123 );
and ( n30125 , n390 , n337 );
not ( n30126 , n390 );
and ( n30127 , n30126 , n300 );
or ( n30128 , n30125 , n30127 );
and ( n30129 , n390 , n364 );
not ( n30130 , n390 );
and ( n30131 , n30130 , n306 );
or ( n30132 , n30129 , n30131 );
and ( n30133 , n3 , n120 );
not ( n30134 , n3 );
and ( n30135 , n30134 , n1201 );
or ( n30136 , n30133 , n30135 );
and ( n30137 , n390 , n375 );
not ( n30138 , n390 );
and ( n30139 , n30138 , n297 );
or ( n30140 , n30137 , n30139 );
and ( n30141 , n3 , n108 );
not ( n30142 , n3 );
and ( n30143 , n30142 , n1422 );
or ( n30144 , n30141 , n30143 );
and ( n30145 , n3 , n109 );
not ( n30146 , n3 );
and ( n30147 , n30146 , n1426 );
or ( n30148 , n30145 , n30147 );
and ( n30149 , n390 , n356 );
not ( n30150 , n390 );
and ( n30151 , n30150 , n296 );
or ( n30152 , n30149 , n30151 );
and ( n30153 , n3 , n110 );
not ( n30154 , n3 );
and ( n30155 , n30154 , n1425 );
or ( n30156 , n30153 , n30155 );
and ( n30157 , n1228 , n372 );
not ( n30158 , n1228 );
and ( n30159 , n30158 , n409 );
or ( n30160 , n30157 , n30159 );
and ( n30161 , n390 , n348 );
not ( n30162 , n390 );
and ( n30163 , n30162 , n294 );
or ( n30164 , n30161 , n30163 );
and ( n30165 , n1228 , n365 );
not ( n30166 , n1228 );
and ( n30167 , n30166 , n347 );
or ( n30168 , n30165 , n30167 );
and ( n30169 , n3 , n101 );
not ( n30170 , n3 );
and ( n30171 , n30170 , n1497 );
or ( n30172 , n30169 , n30171 );
and ( n30173 , n390 , n331 );
not ( n30174 , n390 );
and ( n30175 , n30174 , n288 );
or ( n30176 , n30173 , n30175 );
and ( n30177 , n390 , n354 );
not ( n30178 , n390 );
and ( n30179 , n30178 , n293 );
or ( n30180 , n30177 , n30179 );
and ( n30181 , n3 , n100 );
not ( n30182 , n3 );
and ( n30183 , n30182 , n1431 );
or ( n30184 , n30181 , n30183 );
and ( n30185 , n3 , n118 );
not ( n30186 , n3 );
and ( n30187 , n30186 , n1500 );
or ( n30188 , n30185 , n30187 );
and ( n30189 , n3 , n106 );
not ( n30190 , n3 );
and ( n30191 , n30190 , n1188 );
or ( n30192 , n30189 , n30191 );
and ( n30193 , n3 , n104 );
not ( n30194 , n3 );
and ( n30195 , n30194 , n1428 );
or ( n30196 , n30193 , n30195 );
and ( n30197 , n3 , n119 );
not ( n30198 , n3 );
and ( n30199 , n30198 , n1502 );
or ( n30200 , n30197 , n30199 );
and ( n30201 , n390 , n343 );
not ( n30202 , n390 );
and ( n30203 , n30202 , n305 );
or ( n30204 , n30201 , n30203 );
and ( n30205 , n3 , n127 );
not ( n30206 , n3 );
and ( n30207 , n30206 , n882 );
or ( n30208 , n30205 , n30207 );
and ( n30209 , n3 , n116 );
not ( n30210 , n3 );
and ( n30211 , n30210 , n1521 );
or ( n30212 , n30209 , n30211 );
and ( n30213 , n390 , n340 );
not ( n30214 , n390 );
and ( n30215 , n30214 , n274 );
or ( n30216 , n30213 , n30215 );
and ( n30217 , n390 , n349 );
not ( n30218 , n390 );
and ( n30219 , n30218 , n276 );
or ( n30220 , n30217 , n30219 );
and ( n30221 , n1228 , n353 );
not ( n30222 , n1228 );
and ( n30223 , n30222 , n482 );
or ( n30224 , n30221 , n30223 );
and ( n30225 , n390 , n358 );
not ( n30226 , n390 );
and ( n30227 , n30226 , n285 );
or ( n30228 , n30225 , n30227 );
and ( n30229 , n390 , n330 );
not ( n30230 , n390 );
and ( n30231 , n30230 , n286 );
or ( n30232 , n30229 , n30231 );
and ( n30233 , n390 , n333 );
not ( n30234 , n390 );
and ( n30235 , n30234 , n290 );
or ( n30236 , n30233 , n30235 );
and ( n30237 , n1228 , n386 );
not ( n30238 , n1228 );
and ( n30239 , n30238 , n1487 );
or ( n30240 , n30237 , n30239 );
and ( n30241 , n3 , n105 );
not ( n30242 , n3 );
and ( n30243 , n30242 , n1189 );
or ( n30244 , n30241 , n30243 );
and ( n30245 , n390 , n326 );
not ( n30246 , n390 );
and ( n30247 , n30246 , n287 );
or ( n30248 , n30245 , n30247 );
and ( n30249 , n3 , n114 );
not ( n30250 , n3 );
and ( n30251 , n30250 , n1574 );
or ( n30252 , n30249 , n30251 );
and ( n30253 , n3 , n111 );
not ( n30254 , n3 );
and ( n30255 , n30254 , n1424 );
or ( n30256 , n30253 , n30255 );
and ( n30257 , n3 , n102 );
not ( n30258 , n3 );
and ( n30259 , n30258 , n1430 );
or ( n30260 , n30257 , n30259 );
not ( n30261 , n390 );
nor ( n30262 , n30261 , n325 );
and ( n30263 , n3 , n97 );
not ( n30264 , n3 );
and ( n30265 , n30264 , n1496 );
or ( n30266 , n30263 , n30265 );
and ( n30267 , n390 , n362 );
not ( n30268 , n390 );
and ( n30269 , n30268 , n308 );
or ( n30270 , n30267 , n30269 );
and ( n30271 , n390 , n363 );
not ( n30272 , n390 );
and ( n30273 , n30272 , n309 );
or ( n30274 , n30271 , n30273 );
and ( n30275 , n3 , n98 );
not ( n30276 , n3 );
and ( n30277 , n30276 , n1495 );
or ( n30278 , n30275 , n30277 );
and ( n30279 , n390 , n357 );
not ( n30280 , n390 );
and ( n30281 , n30280 , n311 );
or ( n30282 , n30279 , n30281 );
and ( n30283 , n1228 , n366 );
not ( n30284 , n1228 );
and ( n30285 , n30284 , n855 );
or ( n30286 , n30283 , n30285 );
and ( n30287 , n390 , n346 );
not ( n30288 , n390 );
and ( n30289 , n30288 , n302 );
or ( n30290 , n30287 , n30289 );
and ( n30291 , n390 , n341 );
not ( n30292 , n390 );
and ( n30293 , n30292 , n303 );
or ( n30294 , n30291 , n30293 );
and ( n30295 , n390 , n339 );
not ( n30296 , n390 );
and ( n30297 , n30296 , n301 );
or ( n30298 , n30295 , n30297 );
and ( n30299 , n3 , n107 );
not ( n30300 , n3 );
and ( n30301 , n30300 , n1427 );
or ( n30302 , n30299 , n30301 );
nor ( n30303 , n18004 , n1228 );
and ( n30304 , n390 , n338 );
not ( n30305 , n390 );
and ( n30306 , n30305 , n299 );
or ( n30307 , n30304 , n30306 );
and ( n30308 , n390 , n355 );
not ( n30309 , n390 );
and ( n30310 , n30309 , n295 );
or ( n30311 , n30308 , n30310 );
and ( n30312 , n390 , n334 );
not ( n30313 , n390 );
and ( n30314 , n30313 , n291 );
or ( n30315 , n30312 , n30314 );
and ( n30316 , n390 , n332 );
not ( n30317 , n390 );
and ( n30318 , n30317 , n289 );
or ( n30319 , n30316 , n30318 );
and ( n30320 , n390 , n361 );
not ( n30321 , n390 );
and ( n30322 , n30321 , n273 );
or ( n30323 , n30320 , n30322 );
or ( n30324 , n221 , n237 );
nand ( n30325 , n30324 , n26525 );
and ( n30326 , n390 , n342 );
not ( n30327 , n390 );
and ( n30328 , n30327 , n270 );
or ( n30329 , n30326 , n30328 );
and ( n30330 , n3 , n113 );
not ( n30331 , n3 );
and ( n30332 , n30331 , n1544 );
or ( n30333 , n30330 , n30332 );
or ( n30334 , n1742 , n1745 );
not ( n30335 , n215 );
nor ( n30336 , n30335 , n1228 );
and ( n30337 , n2 , n77 );
and ( n30338 , n54 , n55 );
buf ( n30339 , n73 );
buf ( n30340 , n30339 );
buf ( n30341 , n73 );
buf ( n30342 , n30341 );
buf ( n30343 , n30341 );
buf ( n30344 , n73 );
buf ( n30345 , n30344 );
buf ( n30346 , n30344 );
buf ( n30347 , n30339 );
buf ( n30348 , n30339 );
buf ( n30349 , n30341 );
buf ( n30350 , n73 );
buf ( n30351 , n30350 );
buf ( n30352 , n30350 );
buf ( n30353 , n30350 );
buf ( n30354 , n30339 );
buf ( n30355 , n30339 );
buf ( n30356 , n30339 );
buf ( n30357 , n30341 );
buf ( n30358 , n30344 );
or ( n30359 , n1748 , n1749 );
nor ( n30360 , n1646 , n1710 );
and ( n30361 , n2 , n76 );
not ( n30362 , n329 );
nor ( n30363 , n30362 , n1228 );
and ( n30364 , n2 , n75 );
or ( n30365 , n1741 , n1747 );
or ( n30366 , n1740 , n1746 );
not ( n30367 , n410 );
nor ( n30368 , n30367 , n1228 );
nor ( n30369 , n1595 , n1755 );
buf ( n30370 , n73 );
buf ( n30371 , n30370 );
buf ( n30372 , n30339 );
buf ( n30373 , n30370 );
buf ( n30374 , n30339 );
buf ( n30375 , n30344 );
buf ( n30376 , n30350 );
buf ( n30377 , n30370 );
buf ( n30378 , n30370 );
and ( n30379 , n29092 , n28383 );
nor ( n30380 , n30379 , n926 , n26458 );
and ( n30381 , n1126 , n13756 );
not ( n30382 , n1126 );
and ( n30383 , n30382 , n13757 );
nor ( n30384 , n30381 , n30383 );
xor ( n30385 , n1605 , n28885 );
nor ( n30386 , n30385 , n1755 );
xor ( n30387 , n29996 , n16954 );
xor ( n30388 , n29995 , n17025 );
xor ( n30389 , n1648 , n28894 );
nor ( n30390 , n30389 , n1710 );
xor ( n30391 , n1645 , n28892 );
nor ( n30392 , n30391 , n1710 );
xnor ( n30393 , n1607 , n28323 );
nor ( n30394 , n30393 , n1755 );
xor ( n30395 , n1650 , n29310 );
nor ( n30396 , n30395 , n1710 );
xnor ( n30397 , n29998 , n16871 );
xnor ( n30398 , n29994 , n16944 );
xor ( n30399 , n1635 , n29997 );
nor ( n30400 , n30399 , n1710 );
xnor ( n30401 , n1601 , n28321 );
nor ( n30402 , n30401 , n1755 );
endmodule

