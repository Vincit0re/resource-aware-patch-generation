module top (g98, g97, g96, g95, g94, g93, g92, g91, g90, g9, g89, g88, g87, g86, g85, g84, g83, g82, g81, g80, g8, g79, g78, g77, g76, g75, g74, g73, g72, g71, g70, g7, g69, g68, g67, g66, g65, g64, g63, g62, g61, g60, g6, g59, g58, g57, g56, g55, g54, g53, g52, g51, g50, g5, g49, g48, g47, g46, g45, g44, g43, g42, g41, g40, g4, g39, g38, g37, g36, g35, g34, g33, g32, g31, g30, g3, g29, g28, g27, g26, g25, g24, g23, g22, g21, g20, g2, g19, g18, g17, g16, g15, g14, g13, g12, g11, g10, g1, g0, g99, g100, g101, g102, g103, g104, g105, g106, g107, g108, g109, g110, g111, g112, g113, g114, g115, g116, g117, g118, g119, g120, g121, g122, g123, g124, g125, g126, g127, g128, g129, g130, g131, g132, g133, g134, g135, g136, g137, g138, g139, g140, g141, g142, g143, g144, g145, g146, g147, g148, g149, g150, g151, g152, g153, g154, g155, g156, g157, g158, g159, g160, g161, g162, g163, g164, g165, g166, g167, g168, g169, g170, g171, g172, g173, g174, g175, g176, g177, g178, g179, g180, g181, g182, g183, g184, g185, g186, g187, g188, g189, g190, g191, g192, g193, g194, g195, g196, g197, g198, g199, g200, g201, g202, g203, g204, g205, g206, g207, g208, g209, g210, g211, g212, g213, g214, g215, g216, g217, g218, g219, g220, g221, g222, g223, g224, g225, g226);
   input g98, g97, g96, g95, g94, g93, g92, g91, g90, g9, g89, g88, g87, g86, g85, g84, g83, g82, g81, g80, g8, g79, g78, g77, g76, g75, g74, g73, g72, g71, g70, g7, g69, g68, g67, g66, g65, g64, g63, g62, g61, g60, g6, g59, g58, g57, g56, g55, g54, g53, g52, g51, g50, g5, g49, g48, g47, g46, g45, g44, g43, g42, g41, g40, g4, g39, g38, g37, g36, g35, g34, g33, g32, g31, g30, g3, g29, g28, g27, g26, g25, g24, g23, g22, g21, g20, g2, g19, g18, g17, g16, g15, g14, g13, g12, g11, g10, g1, g0;
   output g99, g100, g101, g102, g103, g104, g105, g106, g107, g108, g109, g110, g111, g112, g113, g114, g115, g116, g117, g118, g119, g120, g121, g122, g123, g124, g125, g126, g127, g128, g129, g130, g131, g132, g133, g134, g135, g136, g137, g138, g139, g140, g141, g142, g143, g144, g145, g146, g147, g148, g149, g150, g151, g152, g153, g154, g155, g156, g157, g158, g159, g160, g161, g162, g163, g164, g165, g166, g167, g168, g169, g170, g171, g172, g173, g174, g175, g176, g177, g178, g179, g180, g181, g182, g183, g184, g185, g186, g187, g188, g189, g190, g191, g192, g193, g194, g195, g196, g197, g198, g199, g200, g201, g202, g203, g204, g205, g206, g207, g208, g209, g210, g211, g212, g213, g214, g215, g216, g217, g218, g219, g220, g221, g222, g223, g224, g225, g226;
   wire n1, n10, n100, n1000, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009, n1001, n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019, n1002, n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029, n1003, n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039, n1004, n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049, n1005, n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059, n1006, n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069, n1007, n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079, n1008, n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089, n1009, n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099, n101, n1010, n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109, n1011, n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119, n1012, n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129, n1013, n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139, n1014, n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149, n1015, n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159, n1016, n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169, n1017, n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179, n1018, n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189, n1019, n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199, n102, n1020, n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209, n1021, n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219, n1022, n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229, n1023, n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239, n1024, n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249, n1025, n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259, n1026, n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269, n1027, n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279, n1028, n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289, n1029, n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299, n103, n1030, n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309, n1031, n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319, n1032, n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329, n1033, n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339, n1034, n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349, n1035, n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359, n1036, n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369, n1037, n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379, n1038, n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389, n1039, n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399, n104, n1040, n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409, n1041, n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419, n1042, n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429, n1043, n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439, n1044, n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449, n1045, n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459, n1046, n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469, n1047, n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479, n1048, n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489, n1049, n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499, n105, n1050, n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509, n1051, n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519, n1052, n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529, n1053, n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539, n1054, n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549, n1055, n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559, n1056, n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569, n1057, n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579, n1058, n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589, n1059, n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599, n106, n1060, n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609, n1061, n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619, n1062, n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629, n1063, n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639, n1064, n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649, n1065, n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659, n1066, n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669, n1067, n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679, n1068, n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689, n1069, n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699, n107, n1070, n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709, n1071, n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719, n1072, n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729, n1073, n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739, n1074, n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749, n1075, n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759, n1076, n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769, n1077, n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779, n1078, n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789, n1079, n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799, n108, n1080, n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809, n1081, n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819, n1082, n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829, n1083, n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839, n1084, n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849, n1085, n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859, n1086, n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869, n1087, n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879, n1088, n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889, n1089, n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899, n109, n1090, n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909, n1091, n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919, n1092, n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929, n1093, n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939, n1094, n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949, n1095, n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959, n1096, n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969, n1097, n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979, n1098, n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989, n1099, n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11, n110, n1100, n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009, n1101, n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019, n1102, n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029, n1103, n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039, n1104, n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049, n1105, n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059, n1106, n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069, n1107, n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079, n1108, n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089, n1109, n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099, n111, n1110, n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109, n1111, n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119, n1112, n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129, n1113, n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139, n1114, n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149, n1115, n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159, n1116, n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169, n1117, n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179, n1118, n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189, n1119, n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199, n112, n1120, n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209, n1121, n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219, n1122, n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229, n1123, n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239, n1124, n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249, n1125, n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259, n1126, n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269, n1127, n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279, n1128, n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289, n1129, n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299, n113, n1130, n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309, n1131, n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319, n1132, n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329, n1133, n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339, n1134, n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349, n1135, n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359, n1136, n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369, n1137, n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379, n1138, n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389, n1139, n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399, n114, n1140, n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409, n1141, n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419, n1142, n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429, n1143, n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439, n1144, n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449, n1145, n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459, n1146, n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469, n1147, n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479, n1148, n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489, n1149, n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499, n115, n1150, n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509, n1151, n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519, n1152, n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529, n1153, n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539, n1154, n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549, n1155, n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559, n1156, n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569, n1157, n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579, n1158, n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589, n1159, n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599, n116, n1160, n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609, n1161, n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619, n1162, n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629, n1163, n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639, n1164, n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649, n1165, n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659, n1166, n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669, n1167, n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679, n1168, n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689, n1169, n11690, n11691, n11692, n117, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n118, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n119, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n12, n120, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n121, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n122, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n123, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n124, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n125, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n126, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n127, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n128, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n129, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n13, n130, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n131, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n132, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n133, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n134, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n135, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n136, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n137, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n138, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n139, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n14, n140, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n141, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n142, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n143, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n144, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n145, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n146, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n147, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n148, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n149, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n15, n150, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n151, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n152, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n153, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n154, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n155, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n156, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n157, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n158, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n159, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n16, n160, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n161, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n162, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n163, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n164, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n165, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n166, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n167, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n168, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n169, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n17, n170, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n171, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n172, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n173, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n174, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n175, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n176, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n177, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n178, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n179, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n18, n180, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n181, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n182, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n183, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n184, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n185, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n186, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n187, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n188, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n189, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n19, n190, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n191, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n192, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n193, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n194, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n195, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n196, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n197, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n198, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n199, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2, n20, n200, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n201, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n202, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n203, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n204, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n205, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n206, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n207, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n208, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n209, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n21, n210, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n211, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n212, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n213, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n214, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n215, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n216, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n217, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n218, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n219, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n22, n220, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n221, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n222, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n223, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n224, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n225, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n226, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n227, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n23, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n237, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n238, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n239, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n24, n240, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n241, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n242, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n243, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n244, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n245, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n246, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n247, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n248, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n249, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n25, n250, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n251, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n252, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n253, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n254, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n255, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n256, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n257, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n258, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n259, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n26, n260, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n261, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n262, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n263, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n264, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n265, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n266, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n267, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n268, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n269, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n27, n270, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n271, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n272, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n273, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n274, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n275, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n276, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n277, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n278, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n279, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n28, n280, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n281, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n282, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n283, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n284, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n285, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n286, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n287, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n288, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n289, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n29, n290, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n291, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n292, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n293, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n294, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n295, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n296, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n297, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n298, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n299, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3, n30, n300, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n301, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n302, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n303, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n304, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n305, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n306, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n307, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n308, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n309, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n31, n310, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n311, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n312, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n313, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n314, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n315, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n316, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n317, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n318, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n319, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n32, n320, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n321, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n322, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n323, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n324, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n325, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n326, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n327, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n328, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n329, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n33, n330, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n331, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n332, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n333, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n334, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n335, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n336, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n337, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n338, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n339, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n34, n340, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n341, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n342, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n343, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n344, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n345, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n346, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n347, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n348, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n349, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n35, n350, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n351, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n352, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n353, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n354, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n355, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n356, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n357, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n358, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n359, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n36, n360, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n361, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n362, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n363, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n364, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n365, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n366, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n367, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n368, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n369, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n37, n370, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n371, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n372, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n373, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n374, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n375, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n376, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n377, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n378, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n379, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n38, n380, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n381, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n382, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n383, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n384, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n385, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n386, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n387, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n388, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n389, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n39, n390, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n391, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n392, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n393, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n394, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n395, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n396, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n397, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n398, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n399, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4, n40, n400, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n401, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n402, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n403, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n404, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n405, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n406, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n407, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n408, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n409, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n41, n410, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n411, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n412, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n413, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n414, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n415, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n416, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n417, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n418, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n419, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n42, n420, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n421, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n422, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n423, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n424, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n425, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n426, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n427, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n428, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n429, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n43, n430, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n431, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n432, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n433, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n434, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n435, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n436, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n437, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n438, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n439, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n44, n440, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n441, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n442, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n443, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n444, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n445, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n446, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n447, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n448, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n449, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n45, n450, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n451, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n452, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n453, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n454, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n455, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n456, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n457, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n458, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n459, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n46, n460, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n461, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n462, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n463, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n464, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n465, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n466, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n467, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n468, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n469, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n47, n470, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n471, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n472, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n473, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n474, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n475, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n476, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n477, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n478, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n479, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n48, n480, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n481, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n482, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n483, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n484, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n485, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n486, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n487, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n488, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n489, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n49, n490, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n491, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n492, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n493, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n494, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n495, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n496, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n497, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n498, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n499, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5, n50, n500, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n501, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n502, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n503, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n504, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n505, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n506, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n507, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n508, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n509, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n51, n510, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n511, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n512, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n513, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n514, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n515, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n516, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n517, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n518, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n519, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n52, n520, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n521, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n522, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n523, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n524, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n525, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n526, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n527, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n528, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n529, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n53, n530, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n531, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n532, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n533, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n534, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n535, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n536, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n537, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n538, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n539, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n54, n540, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n541, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n542, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n543, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n544, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n545, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n546, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n547, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n548, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n549, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n55, n550, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n551, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n552, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n553, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n554, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n555, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n556, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n557, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n558, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n559, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n56, n560, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n561, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n562, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n563, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n564, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n565, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n566, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n567, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n568, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n569, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n57, n570, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n571, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n572, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n573, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n574, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n575, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n576, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n577, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n578, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n579, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n58, n580, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n581, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n582, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n583, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n584, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n585, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n586, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n587, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n588, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n589, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n59, n590, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n591, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n592, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n593, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n594, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n595, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n596, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n597, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n598, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n599, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6, n60, n600, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n601, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n602, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n603, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n604, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n605, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n606, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n607, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n608, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n609, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n61, n610, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n611, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n612, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n613, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n614, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n615, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n616, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n617, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n618, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n619, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n62, n620, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n621, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n622, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n623, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n624, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n625, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n626, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n627, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n628, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n629, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n63, n630, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n631, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n632, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n633, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n634, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n635, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n636, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n637, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n638, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n639, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n64, n640, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n641, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n642, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n643, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n644, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n645, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n646, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n647, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n648, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n649, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n65, n650, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n651, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n652, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n653, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n654, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n655, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n656, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n657, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n658, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n659, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n66, n660, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n661, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n662, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n663, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n664, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n665, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n666, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n667, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n668, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n669, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n67, n670, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n671, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n672, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n673, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n674, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n675, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n676, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n677, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n678, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n679, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n68, n680, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n681, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n682, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n683, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n684, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n685, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n686, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n687, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n688, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n689, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n69, n690, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n691, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n692, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n693, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n694, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n695, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n696, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n697, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n698, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n699, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7, n70, n700, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n701, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n702, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n703, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n704, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n705, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n706, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n707, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n708, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n709, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n71, n710, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n711, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n712, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n713, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n714, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n715, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n716, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n717, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n718, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n719, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n72, n720, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n721, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n722, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n723, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n724, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n725, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n726, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n727, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n728, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n729, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n73, n730, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n731, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n732, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n733, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n734, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n735, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n736, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n737, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n738, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n739, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n74, n740, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n741, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n742, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n743, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n744, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n745, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n746, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n747, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n748, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n749, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n75, n750, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n751, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n752, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n753, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n754, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n755, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n756, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n757, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n758, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n759, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n76, n760, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n761, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n762, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n763, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n764, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n765, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n766, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n767, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n768, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n769, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n77, n770, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n771, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n772, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n773, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n774, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n775, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n776, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n777, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n778, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n779, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n78, n780, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n781, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n782, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n783, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n784, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n785, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n786, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n787, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n788, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n789, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n79, n790, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n791, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n792, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n793, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n794, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n795, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n796, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n797, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n798, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n799, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8, n80, n800, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n801, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n802, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n803, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n804, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n805, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n806, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n807, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n808, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n809, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n81, n810, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n811, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n812, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n813, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n814, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n815, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n816, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n817, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n818, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n819, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n82, n820, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n821, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n822, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n823, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n824, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n825, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n826, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n827, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n828, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n829, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n83, n830, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n831, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n832, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n833, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n834, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n835, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n836, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n837, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n838, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n839, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n84, n840, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n841, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n842, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n843, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n844, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n845, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n846, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n847, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n848, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n849, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n85, n850, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n851, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n852, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n853, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n854, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n855, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n856, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n857, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n858, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n859, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n86, n860, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n861, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n862, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n863, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n864, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n865, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n866, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n867, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n868, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n869, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n87, n870, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n871, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n872, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n873, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n874, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n875, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n876, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n877, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n878, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n879, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n88, n880, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n881, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n882, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n883, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n884, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n885, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n886, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n887, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n888, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n89, n890, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n891, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n892, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n893, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n894, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n895, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n896, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n897, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n898, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n899, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9, n90, n900, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n901, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n902, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n903, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n904, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n905, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n906, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n907, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n908, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n909, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n91, n910, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n911, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n912, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n913, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n914, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n915, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n916, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n917, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n918, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n919, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n92, n920, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n921, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n922, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n923, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n924, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n925, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n926, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n927, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n928, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n929, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n93, n930, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n931, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n932, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n933, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n934, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n935, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n936, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n937, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n938, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n939, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n94, n940, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n941, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n942, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n943, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n944, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n945, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n946, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n947, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n948, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n949, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n95, n950, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n951, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n952, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n953, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n954, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n955, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n956, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n957, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n958, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n959, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n96, n960, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n961, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n962, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n963, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n964, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n965, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n966, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n967, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n968, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n969, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n97, n970, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n971, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n972, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n973, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n974, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n975, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n976, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n977, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n978, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n979, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n98, n980, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n981, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n982, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n983, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n984, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n985, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n986, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n987, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n988, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n989, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n99, n990, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n991, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n992, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n993, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n994, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n995, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n996, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n997, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n998, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n999, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999;
   buf (g100, n101);
   buf (g101, n102);
   buf (g102, n103);
   buf (g103, n104);
   buf (g104, n105);
   buf (g105, n106);
   buf (g106, n107);
   buf (g107, n108);
   buf (g108, n109);
   buf (g109, n110);
   buf (g110, n111);
   buf (g111, n112);
   buf (g112, n113);
   buf (g113, n114);
   buf (g114, n115);
   buf (g115, n116);
   buf (g116, n117);
   buf (g117, n118);
   buf (g118, n119);
   buf (g119, n120);
   buf (g120, n121);
   buf (g121, n122);
   buf (g122, n123);
   buf (g123, n124);
   buf (g124, n125);
   buf (g125, n126);
   buf (g126, n127);
   buf (g127, n128);
   buf (g128, n129);
   buf (g129, n130);
   buf (g130, n131);
   buf (g131, n132);
   buf (g132, n133);
   buf (g133, n134);
   buf (g134, n135);
   buf (g135, n136);
   buf (g136, n137);
   buf (g137, n138);
   buf (g138, n139);
   buf (g139, n140);
   buf (g140, n141);
   buf (g141, n142);
   buf (g142, n143);
   buf (g143, n144);
   buf (g144, n145);
   buf (g145, n146);
   buf (g146, n147);
   buf (g147, n148);
   buf (g148, n149);
   buf (g149, n150);
   buf (g150, n151);
   buf (g151, n152);
   buf (g152, n153);
   buf (g153, n154);
   buf (g154, n155);
   buf (g155, n156);
   buf (g156, n157);
   buf (g157, n158);
   buf (g158, n159);
   buf (g159, n160);
   buf (g160, n161);
   buf (g161, n162);
   buf (g162, n163);
   buf (g163, n164);
   buf (g164, n165);
   buf (g165, n166);
   buf (g166, n167);
   buf (g167, n168);
   buf (g168, n169);
   buf (g169, n170);
   buf (g170, n171);
   buf (g171, n172);
   buf (g172, n173);
   buf (g173, n174);
   buf (g174, n175);
   buf (g175, n176);
   buf (g176, n177);
   buf (g177, n178);
   buf (g178, n179);
   buf (g179, n180);
   buf (g180, n181);
   buf (g181, n182);
   buf (g182, n183);
   buf (g183, n184);
   buf (g184, n185);
   buf (g185, n186);
   buf (g186, n187);
   buf (g187, n188);
   buf (g188, n189);
   buf (g189, n190);
   buf (g190, n191);
   buf (g191, n192);
   buf (g192, n193);
   buf (g193, n194);
   buf (g194, n195);
   buf (g195, n196);
   buf (g196, n197);
   buf (g197, n198);
   buf (g198, n199);
   buf (g199, n200);
   buf (g200, n201);
   buf (g201, n202);
   buf (g202, n203);
   buf (g203, n204);
   buf (g204, n205);
   buf (g205, n206);
   buf (g206, n207);
   buf (g207, n208);
   buf (g208, n209);
   buf (g209, n210);
   buf (g210, n211);
   buf (g211, n212);
   buf (g212, n213);
   buf (g213, n214);
   buf (g214, n215);
   buf (g215, n216);
   buf (g216, n217);
   buf (g217, n218);
   buf (g218, n219);
   buf (g219, n220);
   buf (g220, n221);
   buf (g221, n222);
   buf (g222, n223);
   buf (g223, n224);
   buf (g224, n225);
   buf (g225, n226);
   buf (g226, n227);
   buf (g99, n100);
   buf (n1, g0);
   buf (n10, g9);
   buf (n100, n11417);
   nand (n1000, n996, n999);
   and (n10000, n43, n2925);
   not (n10001, n43);
   and (n10002, n10001, n2928);
   nor (n10003, n10000, n10002);
   or (n10004, n9679, n10003);
   or (n10005, n9646, n5307);
   nand (n10006, n10004, n10005);
   and (n10007, n9999, n10006);
   and (n10008, n9997, n9998);
   nor (n10009, n10007, n10008);
   not (n1001, n1000);
   or (n10010, n9948, n5427);
   not (n10011, n5248);
   or (n10012, n9957, n10011);
   nand (n10013, n10010, n10012);
   nor (n10014, n10013, n4924);
   and (n10015, n10014, n9961);
   not (n10016, n10014);
   and (n10017, n10016, n9962);
   nor (n10018, n10015, n10017);
   or (n10019, n10009, n10018);
   nand (n1002, n36, n66);
   or (n10020, n10014, n9962);
   nand (n10021, n10019, n10020);
   xor (n10022, n9990, n10021);
   xor (n10023, n9932, n9935);
   xor (n10024, n10023, n9939);
   not (n10025, n10024);
   xnor (n10026, n9918, n9919);
   and (n10027, n3386, n4580);
   not (n10028, n3386);
   and (n10029, n10028, n45);
   and (n1003, n1002, n50);
   nor (n10030, n10027, n10029);
   or (n10031, n9578, n10030);
   or (n10032, n9582, n5275);
   nand (n10033, n10031, n10032);
   and (n10034, n39, n3127);
   not (n10035, n39);
   and (n10036, n10035, n3826);
   nor (n10037, n10034, n10036);
   or (n10038, n9928, n10037);
   or (n10039, n9885, n9929);
   not (n1004, n1002);
   nand (n10040, n10038, n10039);
   xor (n10041, n10033, n10040);
   and (n10042, n2832, n3564);
   nor (n10043, n10042, n9919);
   not (n10044, n10043);
   or (n10045, n9596, n10044);
   or (n10046, n9603, n5318);
   nand (n10047, n10045, n10046);
   and (n10048, n10041, n10047);
   and (n10049, n10033, n10040);
   not (n1005, n50);
   nor (n10050, n10048, n10049);
   xor (n10051, n10026, n10050);
   not (n10052, n10051);
   or (n10053, n10025, n10052);
   or (n10054, n10050, n10026);
   nand (n10055, n10053, n10054);
   and (n10056, n10022, n10055);
   and (n10057, n9990, n10021);
   nor (n10058, n10056, n10057);
   xor (n10059, n9989, n10058);
   and (n1006, n1004, n1005);
   not (n10060, n10059);
   xor (n10061, n10022, n10055);
   xnor (n10062, n9923, n9924);
   xor (n10063, n10061, n10062);
   xor (n10064, n10009, n10018);
   not (n10065, n10064);
   not (n10066, n3919);
   not (n10067, n9994);
   not (n10068, n10067);
   not (n10069, n9752);
   nor (n1007, n1003, n1006);
   or (n10070, n10068, n10069);
   or (n10071, n9910, n3906);
   nand (n10072, n10070, n10071);
   not (n10073, n10072);
   or (n10074, n10066, n10073);
   or (n10075, n10072, n3919);
   nand (n10076, n10074, n10075);
   or (n10077, n9679, n3848);
   or (n10078, n9645, n10003);
   nand (n10079, n10077, n10078);
   not (n1008, n1007);
   and (n10080, n10076, n10079);
   not (n10081, n3919);
   and (n10082, n10072, n10081);
   nor (n10083, n10080, n10082);
   not (n10084, n3842);
   not (n10085, n9947);
   or (n10086, n10084, n10085);
   not (n10087, n5427);
   nand (n10088, n10087, n9958);
   nand (n10089, n10086, n10088);
   or (n1009, n1001, n1008);
   not (n10090, n2762);
   not (n10091, n3768);
   or (n10092, n10090, n10091);
   buf (n10093, n3363);
   nor (n10094, n3351, n10093);
   not (n10095, n10094);
   nand (n10096, n10092, n10095);
   nand (n10097, n10089, n10096);
   xor (n10098, n10083, n10097);
   not (n10099, n9596);
   buf (n101, n11417);
   or (n1010, n1002, n50);
   not (n10100, n3807);
   and (n10101, n10099, n10100);
   and (n10102, n9602, n10043);
   nor (n10103, n10101, n10102);
   buf (n10104, n9883);
   not (n10105, n10104);
   not (n10106, n10037);
   and (n10107, n10105, n10106);
   not (n10108, n3830);
   nor (n10109, n10108, n9928);
   nand (n1011, n1009, n1010);
   nor (n10110, n10107, n10109);
   xor (n10111, n10103, n10110);
   not (n10112, n3792);
   not (n10113, n10112);
   not (n10114, n9577);
   or (n10115, n10113, n10114);
   or (n10116, n9582, n10030);
   nand (n10117, n10115, n10116);
   not (n10118, n10117);
   and (n10119, n10111, n10118);
   and (n1012, n46, n55);
   and (n10120, n10103, n10110);
   or (n10121, n10119, n10120);
   and (n10122, n10098, n10121);
   and (n10123, n10083, n10097);
   nor (n10124, n10122, n10123);
   not (n10125, n10124);
   or (n10126, n10065, n10125);
   xnor (n10127, n10124, n10064);
   xor (n10128, n10041, n10047);
   not (n10129, n10014);
   not (n1013, n46);
   nand (n10130, n10013, n4924);
   nand (n10131, n10129, n10130);
   xor (n10132, n10128, n10131);
   xor (n10133, n9999, n10006);
   and (n10134, n10132, n10133);
   and (n10135, n10128, n10131);
   nor (n10136, n10134, n10135);
   or (n10137, n10127, n10136);
   nand (n10138, n10126, n10137);
   and (n10139, n10063, n10138);
   and (n1014, n1013, n377);
   and (n10140, n10061, n10062);
   nor (n10141, n10139, n10140);
   not (n10142, n10141);
   or (n10143, n10060, n10142);
   not (n10144, n3372);
   not (n10145, n9621);
   or (n10146, n10144, n10145);
   not (n10147, n3650);
   nand (n10148, n10147, n9644);
   nand (n10149, n10146, n10148);
   nor (n1015, n1012, n1014);
   not (n10150, n39);
   not (n10151, n10094);
   or (n10152, n10150, n10151);
   nand (n10153, n3351, n3363);
   not (n10154, n10153);
   or (n10155, n3768, n39);
   nand (n10156, n3739, n40);
   nand (n10157, n10155, n10156);
   nor (n10158, n10154, n10157);
   nand (n10159, n10152, n10158);
   not (n1016, n1015);
   xor (n10160, n10149, n10159);
   not (n10161, n10160);
   not (n10162, n4040);
   not (n10163, n9577);
   or (n10164, n10162, n10163);
   and (n10165, n2845, n610);
   not (n10166, n2845);
   and (n10167, n10166, n49);
   nor (n10168, n10165, n10167);
   not (n10169, n10168);
   not (n1017, n535);
   or (n10170, n9582, n10169);
   nand (n10171, n10164, n10170);
   and (n10172, n10161, n10171);
   not (n10173, n10159);
   and (n10174, n10149, n10173);
   nor (n10175, n10172, n10174);
   not (n10176, n10175);
   nand (n10177, n9602, n51);
   not (n10178, n9589);
   nand (n10179, n10178, n2833);
   or (n1018, n1016, n1017);
   not (n10180, n10179);
   and (n10181, n10177, n10180);
   not (n10182, n3356);
   not (n10183, n10093);
   and (n10184, n10182, n10183);
   not (n10185, n39);
   not (n10186, n3739);
   or (n10187, n10185, n10186);
   nand (n10188, n10187, n10153);
   nor (n10189, n10184, n10188);
   not (n1019, n815);
   or (n10190, n10181, n10189);
   nand (n10191, n10181, n10189);
   nand (n10192, n10190, n10191);
   not (n10193, n10192);
   or (n10194, n9749, n4127);
   and (n10195, n3071, n4580);
   not (n10196, n3071);
   and (n10197, n10196, n45);
   nor (n10198, n10195, n10197);
   not (n10199, n10198);
   buf (n102, n11417);
   nand (n1020, n1019, n917);
   or (n10200, n9753, n10199);
   nand (n10201, n10194, n10200);
   not (n10202, n10201);
   not (n10203, n10177);
   not (n10204, n3577);
   not (n10205, n9946);
   not (n10206, n10205);
   or (n10207, n10204, n10206);
   not (n10208, n335);
   not (n10209, n9959);
   nand (n1021, n1018, n1020);
   or (n10210, n10208, n10209);
   nand (n10211, n4570, n41);
   nand (n10212, n10210, n10211);
   nand (n10213, n9958, n10212);
   nand (n10214, n10207, n10213);
   not (n10215, n10214);
   or (n10216, n10203, n10215);
   or (n10217, n10214, n10177);
   nand (n10218, n10216, n10217);
   not (n10219, n10218);
   not (n1022, n1021);
   or (n10220, n10202, n10219);
   not (n10221, n10177);
   nand (n10222, n10221, n10214);
   nand (n10223, n10220, n10222);
   not (n10224, n10223);
   or (n10225, n10193, n10224);
   or (n10226, n10223, n10192);
   nand (n10227, n10225, n10226);
   nand (n10228, n10176, n10227);
   not (n10229, n10192);
   and (n1023, n909, n430);
   nand (n10230, n10229, n10223);
   nand (n10231, n10228, n10230);
   not (n10232, n3538);
   not (n10233, n9577);
   or (n10234, n10232, n10233);
   not (n10235, n3890);
   and (n10236, n9574, n9580);
   nand (n10237, n10235, n10236);
   nand (n10238, n10234, n10237);
   not (n10239, n3331);
   and (n1024, n42, n59);
   not (n10240, n10239);
   not (n10241, n9595);
   or (n10242, n10240, n10241);
   not (n10243, n3920);
   nand (n10244, n10243, n9602);
   nand (n10245, n10242, n10244);
   xor (n10246, n10238, n10245);
   not (n10247, n10191);
   and (n10248, n10246, n10247);
   not (n10249, n10246);
   not (n1025, n42);
   and (n10250, n10249, n10191);
   nor (n10251, n10248, n10250);
   not (n10252, n3477);
   not (n10253, n10252);
   not (n10254, n9621);
   or (n10255, n10253, n10254);
   and (n10256, n2925, n4580);
   not (n10257, n2925);
   and (n10258, n10257, n45);
   nor (n10259, n10256, n10258);
   and (n1026, n1025, n578);
   nand (n10260, n9644, n10259);
   nand (n10261, n10255, n10260);
   not (n10262, n3527);
   not (n10263, n9697);
   or (n10264, n10262, n10263);
   not (n10265, n3562);
   not (n10266, n43);
   and (n10267, n10265, n10266);
   and (n10268, n3071, n43);
   nor (n10269, n10267, n10268);
   nor (n1027, n1024, n1026);
   not (n10270, n10269);
   nand (n10271, n10270, n9752);
   nand (n10272, n10264, n10271);
   xor (n10273, n10261, n10272);
   not (n10274, n3444);
   or (n10275, n9880, n10274);
   and (n10276, n3127, n335);
   not (n10277, n3127);
   and (n10278, n10277, n41);
   nor (n10279, n10276, n10278);
   and (n1028, n421, n1027);
   not (n10280, n10279);
   or (n10281, n9885, n10280);
   nand (n10282, n10275, n10281);
   xor (n10283, n10273, n10282);
   xnor (n10284, n10251, n10283);
   xor (n10285, n10231, n10284);
   or (n10286, n9679, n3650);
   or (n10287, n9645, n3477);
   nand (n10288, n10286, n10287);
   not (n10289, n10288);
   nor (n1029, n1023, n1028);
   not (n10290, n10198);
   not (n10291, n9697);
   or (n10292, n10290, n10291);
   nand (n10293, n9752, n3527);
   nand (n10294, n10292, n10293);
   not (n10295, n10294);
   not (n10296, n9957);
   not (n10297, n3424);
   not (n10298, n10297);
   and (n10299, n10296, n10298);
   buf (n103, n11417);
   not (n1030, n1029);
   and (n10300, n9947, n10212);
   nor (n10301, n10299, n10300);
   not (n10302, n10301);
   or (n10303, n10295, n10302);
   or (n10304, n10301, n10294);
   nand (n10305, n10303, n10304);
   not (n10306, n10305);
   or (n10307, n10289, n10306);
   not (n10308, n10301);
   nand (n10309, n10308, n10294);
   and (n1031, n1022, n1030);
   nand (n10310, n10307, n10309);
   not (n10311, n10310);
   and (n10312, n2845, n3334);
   not (n10313, n2845);
   and (n10314, n10313, n51);
   nor (n10315, n10312, n10314);
   not (n10316, n10315);
   and (n10317, n9597, n10316);
   and (n10318, n9602, n10239);
   nor (n10319, n10317, n10318);
   and (n1032, n1029, n1021);
   not (n10320, n10319);
   not (n10321, n10168);
   not (n10322, n9577);
   or (n10323, n10321, n10322);
   nand (n10324, n9581, n3538);
   nand (n10325, n10323, n10324);
   xnor (n10326, n3127, n43);
   not (n10327, n10326);
   not (n10328, n9811);
   or (n10329, n10327, n10328);
   nor (n1033, n1031, n1032);
   not (n10330, n10104);
   nand (n10331, n10330, n3444);
   nand (n10332, n10329, n10331);
   xor (n10333, n10325, n10332);
   nand (n10334, n10320, n10333);
   nand (n10335, n10332, n10325);
   and (n10336, n10334, n10335);
   not (n10337, n10336);
   and (n10338, n10311, n10337);
   buf (n10339, n10336);
   and (n1034, n48, n53);
   and (n10340, n10310, n10339);
   nor (n10341, n10338, n10340);
   nand (n10342, n2833, n51);
   not (n10343, n10342);
   not (n10344, n3073);
   not (n10345, n10094);
   or (n10346, n10344, n10345);
   nand (n10347, n3768, n3363);
   not (n10348, n10347);
   not (n10349, n38);
   nor (n1035, n48, n53);
   and (n10350, n10348, n10349);
   not (n10351, n3363);
   and (n10352, n3351, n10351, n37);
   nor (n10353, n10350, n10352);
   nand (n10354, n10346, n10353);
   not (n10355, n10354);
   not (n10356, n10355);
   or (n10357, n10343, n10356);
   not (n10358, n10342);
   nand (n10359, n10358, n10354);
   nor (n1036, n1034, n1035);
   nand (n10360, n10357, n10359);
   not (n10361, n9957);
   not (n10362, n39);
   not (n10363, n4570);
   or (n10364, n10362, n10363);
   or (n10365, n4570, n39);
   nand (n10366, n10364, n10365);
   not (n10367, n10366);
   not (n10368, n10367);
   and (n10369, n10361, n10368);
   and (n1037, n712, n1036);
   and (n10370, n9949, n3424);
   nor (n10371, n10369, n10370);
   xnor (n10372, n10360, n10371);
   xnor (n10373, n10341, n10372);
   xor (n10374, n10285, n10373);
   xor (n10375, n10305, n10288);
   not (n10376, n10319);
   not (n10377, n10333);
   or (n10378, n10376, n10377);
   or (n10379, n10333, n10319);
   not (n1038, n614);
   nand (n10380, n10378, n10379);
   xor (n10381, n10375, n10380);
   not (n10382, n3567);
   not (n10383, n10382);
   not (n10384, n9697);
   or (n10385, n10383, n10384);
   or (n10386, n9751, n4127);
   nand (n10387, n10385, n10386);
   and (n10388, n2907, n610);
   not (n10389, n2907);
   not (n1039, n1038);
   and (n10390, n10389, n49);
   nor (n10391, n10388, n10390);
   not (n10392, n10391);
   not (n10393, n9620);
   not (n10394, n10393);
   or (n10395, n10392, n10394);
   not (n10396, n3372);
   or (n10397, n9645, n10396);
   nand (n10398, n10395, n10397);
   xor (n10399, n10387, n10398);
   buf (n104, n11417);
   and (n1040, n1039, n703);
   not (n10400, n10093);
   and (n10401, n4078, n10400);
   not (n10402, n41);
   not (n10403, n10093);
   or (n10404, n10402, n10403);
   nand (n10405, n10404, n10153);
   nor (n10406, n10401, n10405);
   and (n10407, n10399, n10406);
   and (n10408, n10387, n10398);
   nor (n10409, n10407, n10408);
   nor (n1041, n1037, n1040);
   and (n10410, n4570, n4944);
   not (n10411, n4570);
   and (n10412, n10411, n43);
   nor (n10413, n10410, n10412);
   not (n10414, n10413);
   not (n10415, n9947);
   or (n10416, n10414, n10415);
   nand (n10417, n9958, n3577);
   nand (n10418, n10416, n10417);
   nand (n10419, n10236, n51);
   or (n1042, n1033, n1041);
   and (n10420, n9580, n2846);
   and (n10421, n10419, n10420);
   nand (n10422, n10418, n10421);
   or (n10423, n9880, n3589);
   not (n10424, n10326);
   or (n10425, n9885, n10424);
   nand (n10426, n10423, n10425);
   and (n10427, n10422, n10426);
   not (n10428, n10422);
   not (n10429, n10426);
   not (n1043, n1021);
   and (n10430, n10428, n10429);
   nor (n10431, n10427, n10430);
   or (n10432, n10409, n10431);
   or (n10433, n10422, n10429);
   nand (n10434, n10432, n10433);
   and (n10435, n10381, n10434);
   and (n10436, n10375, n10380);
   nor (n10437, n10435, n10436);
   xnor (n10438, n10374, n10437);
   not (n10439, n10175);
   or (n1044, n1043, n1029);
   not (n10440, n10227);
   or (n10441, n10439, n10440);
   or (n10442, n10227, n10175);
   nand (n10443, n10441, n10442);
   buf (n10444, n10443);
   not (n10445, n10444);
   xnor (n10446, n10218, n10201);
   not (n10447, n10171);
   not (n10448, n10160);
   or (n10449, n10447, n10448);
   nand (n1045, n1042, n1044);
   or (n10450, n10160, n10171);
   nand (n10451, n10449, n10450);
   not (n10452, n10451);
   and (n10453, n10446, n10452);
   not (n10454, n10446);
   and (n10455, n10454, n10451);
   nor (n10456, n10453, n10455);
   or (n10457, n10418, n10421);
   nand (n10458, n10457, n10422);
   not (n10459, n10458);
   xor (n1046, n1011, n1045);
   and (n10460, n3127, n45);
   not (n10461, n3127);
   and (n10462, n10461, n4580);
   nor (n10463, n10460, n10462);
   or (n10464, n9880, n10463);
   or (n10465, n10104, n3589);
   nand (n10466, n10464, n10465);
   and (n10467, n9577, n10315);
   and (n10468, n9581, n4040);
   nor (n10469, n10467, n10468);
   and (n1047, n953, n931);
   not (n10470, n10469);
   and (n10471, n10466, n10470);
   not (n10472, n10466);
   and (n10473, n10472, n10469);
   nor (n10474, n10471, n10473);
   and (n10475, n10459, n10474);
   and (n10476, n10466, n10470);
   nor (n10477, n10475, n10476);
   and (n10478, n10456, n10477);
   and (n10479, n10452, n10446);
   not (n1048, n953);
   nor (n10480, n10478, n10479);
   not (n10481, n10480);
   and (n10482, n10445, n10481);
   xor (n10483, n10480, n10444);
   xnor (n10484, n10381, n10434);
   and (n10485, n10483, n10484);
   nor (n10486, n10482, n10485);
   and (n10487, n10438, n10486);
   not (n10488, n3330);
   not (n10489, n10366);
   and (n1049, n1048, n932);
   not (n10490, n9947);
   or (n10491, n10489, n10490);
   nand (n10492, n9958, n3842);
   nand (n10493, n10491, n10492);
   not (n10494, n10493);
   or (n10495, n10488, n10494);
   or (n10496, n10493, n3330);
   nand (n10497, n10495, n10496);
   not (n10498, n10497);
   not (n10499, n3783);
   buf (n105, n11417);
   nor (n1050, n1047, n1049);
   not (n10500, n9752);
   or (n10501, n10499, n10500);
   or (n10502, n9749, n10269);
   nand (n10503, n10501, n10502);
   not (n10504, n10503);
   and (n10505, n10498, n10504);
   and (n10506, n10497, n10503);
   nor (n10507, n10505, n10506);
   not (n10508, n10507);
   xor (n10509, n10261, n10272);
   not (n1051, n1050);
   and (n10510, n10509, n10282);
   and (n10511, n10261, n10272);
   nor (n10512, n10510, n10511);
   not (n10513, n10512);
   not (n10514, n10279);
   not (n10515, n9811);
   or (n10516, n10514, n10515);
   not (n10517, n10104);
   nand (n10518, n10517, n3830);
   nand (n10519, n10516, n10518);
   and (n1052, n1046, n1051);
   not (n10520, n10259);
   not (n10521, n9621);
   or (n10522, n10520, n10521);
   nand (n10523, n9644, n3957);
   nand (n10524, n10522, n10523);
   xor (n10525, n10519, n10524);
   or (n10526, n9578, n3890);
   or (n10527, n9582, n3792);
   nand (n10528, n10526, n10527);
   xor (n10529, n10525, n10528);
   and (n1053, n1011, n1045);
   not (n10530, n10529);
   or (n10531, n10513, n10530);
   or (n10532, n10512, n10529);
   nand (n10533, n10531, n10532);
   not (n10534, n10533);
   or (n10535, n10508, n10534);
   not (n10536, n10512);
   nand (n10537, n10536, n10529);
   nand (n10538, n10535, n10537);
   not (n10539, n10503);
   nor (n1054, n1052, n1053);
   nand (n10540, n10539, n10497);
   not (n10541, n10493);
   nand (n10542, n10541, n3330);
   nand (n10543, n10540, n10542);
   or (n10544, n10089, n10096);
   nand (n10545, n10544, n10097);
   and (n10546, n10543, n10545);
   nor (n10547, n10543, n10545);
   nor (n10548, n10546, n10547);
   not (n10549, n10548);
   xnor (n1055, n993, n1054);
   or (n10550, n10360, n10371);
   nand (n10551, n10550, n10359);
   or (n10552, n9596, n3920);
   or (n10553, n9601, n3807);
   nand (n10554, n10552, n10553);
   not (n10555, n10554);
   not (n10556, n10351);
   not (n10557, n3770);
   or (n10558, n10556, n10557);
   nor (n10559, n10351, n3073);
   nand (n1056, n36, n67);
   nor (n10560, n10154, n10559);
   nand (n10561, n10558, n10560);
   not (n10562, n10561);
   or (n10563, n10555, n10562);
   or (n10564, n10561, n10554);
   nand (n10565, n10563, n10564);
   and (n10566, n10551, n10565);
   not (n10567, n10561);
   and (n10568, n10567, n10554);
   nor (n10569, n10566, n10568);
   not (n1057, n1056);
   not (n10570, n10569);
   and (n10571, n10549, n10570);
   and (n10572, n10548, n10569);
   nor (n10573, n10571, n10572);
   and (n10574, n10538, n10573);
   not (n10575, n10538);
   not (n10576, n10573);
   and (n10577, n10575, n10576);
   or (n10578, n10574, n10577);
   xnor (n10579, n10076, n10079);
   not (n1058, n50);
   xor (n10580, n10519, n10524);
   and (n10581, n10580, n10528);
   and (n10582, n10519, n10524);
   nor (n10583, n10581, n10582);
   xor (n10584, n10103, n10110);
   not (n10585, n10117);
   xor (n10586, n10584, n10585);
   xnor (n10587, n10583, n10586);
   xor (n10588, n10579, n10587);
   xnor (n10589, n10578, n10588);
   not (n1059, n267);
   xnor (n10590, n10551, n10565);
   not (n10591, n10590);
   and (n10592, n10246, n10247);
   and (n10593, n10238, n10245);
   nor (n10594, n10592, n10593);
   not (n10595, n10594);
   and (n10596, n10591, n10595);
   xor (n10597, n10590, n10594);
   or (n10598, n10341, n10372);
   not (n10599, n10310);
   buf (n106, n11417);
   or (n1060, n1058, n1059);
   or (n10600, n10599, n10339);
   nand (n10601, n10598, n10600);
   and (n10602, n10597, n10601);
   nor (n10603, n10596, n10602);
   xnor (n10604, n10589, n10603);
   not (n10605, n10604);
   or (n10606, n10231, n10284);
   or (n10607, n10251, n10283);
   nand (n10608, n10606, n10607);
   xnor (n10609, n10533, n10507);
   nand (n1061, n50, n51);
   xor (n10610, n10608, n10609);
   xnor (n10611, n10601, n10597);
   and (n10612, n10610, n10611);
   and (n10613, n10608, n10609);
   nor (n10614, n10612, n10613);
   nand (n10615, n10605, n10614);
   xor (n10616, n10608, n10609);
   xor (n10617, n10616, n10611);
   not (n10618, n10617);
   xor (n10619, n10285, n10373);
   nand (n1062, n1060, n1061);
   and (n10620, n10619, n10437);
   and (n10621, n10285, n10373);
   nor (n10622, n10620, n10621);
   nand (n10623, n10618, n10622);
   nand (n10624, n10615, n10623);
   nor (n10625, n10487, n10624);
   not (n10626, n10625);
   xnor (n10627, n10399, n10406);
   nand (n10628, n10094, n41);
   and (n10629, n4924, n335);
   not (n1063, n1062);
   nor (n10630, n3737, n423);
   nor (n10631, n10629, n10630);
   nand (n10632, n10628, n10153, n10631);
   not (n10633, n10632);
   not (n10634, n4328);
   not (n10635, n10634);
   not (n10636, n10393);
   or (n10637, n10635, n10636);
   nand (n10638, n9644, n10391);
   nand (n10639, n10637, n10638);
   not (n1064, n1063);
   not (n10640, n10639);
   or (n10641, n10633, n10640);
   or (n10642, n10632, n10639);
   nand (n10643, n10641, n10642);
   not (n10644, n4462);
   or (n10645, n9928, n10644);
   or (n10646, n9885, n10463);
   nand (n10647, n10645, n10646);
   and (n10648, n10643, n10647);
   not (n10649, n10632);
   or (n1065, n1057, n1064);
   and (n10650, n10649, n10639);
   nor (n10651, n10648, n10650);
   not (n10652, n10651);
   not (n10653, n4365);
   or (n10654, n9749, n10653);
   or (n10655, n9753, n3567);
   nand (n10656, n10654, n10655);
   not (n10657, n10656);
   not (n10658, n10419);
   not (n10659, n4215);
   not (n1066, n1056);
   not (n10660, n9947);
   or (n10661, n10659, n10660);
   nand (n10662, n9958, n10413);
   nand (n10663, n10661, n10662);
   not (n10664, n10663);
   or (n10665, n10658, n10664);
   or (n10666, n10663, n10419);
   nand (n10667, n10665, n10666);
   not (n10668, n10667);
   or (n10669, n10657, n10668);
   nand (n1067, n1066, n1062);
   not (n10670, n10419);
   nand (n10671, n10670, n10663);
   nand (n10672, n10669, n10671);
   not (n10673, n10672);
   or (n10674, n10652, n10673);
   or (n10675, n10672, n10651);
   nand (n10676, n10674, n10675);
   and (n10677, n10627, n10676);
   not (n10678, n10672);
   and (n10679, n10678, n10651);
   nand (n1068, n1065, n1067);
   nor (n10680, n10677, n10679);
   xor (n10681, n10409, n10431);
   xor (n10682, n10680, n10681);
   xnor (n10683, n10456, n10477);
   and (n10684, n10682, n10683);
   and (n10685, n10680, n10681);
   nor (n10686, n10684, n10685);
   not (n10687, n10686);
   xor (n10688, n10480, n10444);
   xnor (n10689, n10688, n10484);
   and (n1069, n48, n54);
   not (n10690, n10689);
   or (n10691, n10687, n10690);
   or (n10692, n10689, n10686);
   nand (n10693, n10691, n10692);
   not (n10694, n10693);
   xnor (n10695, n10682, n10683);
   not (n10696, n10695);
   xor (n10697, n10676, n10627);
   not (n10698, n10458);
   not (n10699, n10474);
   buf (n107, n11417);
   not (n1070, n48);
   and (n10700, n10698, n10699);
   and (n10701, n10458, n10474);
   nor (n10702, n10700, n10701);
   and (n10703, n10697, n10702);
   not (n10704, n10697);
   not (n10705, n10702);
   and (n10706, n10704, n10705);
   nor (n10707, n10703, n10706);
   not (n10708, n4226);
   not (n10709, n9697);
   and (n1071, n1070, n299);
   or (n10710, n10708, n10709);
   or (n10711, n9751, n10653);
   nand (n10712, n10710, n10711);
   not (n10713, n3204);
   not (n10714, n3334);
   and (n10715, n10713, n10714);
   and (n10716, n3071, n3334);
   nor (n10717, n10715, n10716);
   not (n10718, n10717);
   not (n10719, n10718);
   nor (n1072, n1069, n1071);
   not (n10720, n10393);
   or (n10721, n10719, n10720);
   nand (n10722, n9644, n10634);
   nand (n10723, n10721, n10722);
   xor (n10724, n10712, n10723);
   or (n10725, n4254, n10093);
   and (n10726, n3739, n43);
   nor (n10727, n10726, n10154);
   nand (n10728, n10725, n10727);
   not (n10729, n10728);
   not (n1073, n705);
   and (n10730, n10724, n10729);
   and (n10731, n10712, n10723);
   nor (n10732, n10730, n10731);
   nand (n10733, n9644, n51);
   nand (n10734, n10733, n9624);
   not (n10735, n10734);
   not (n10736, n10205);
   not (n10737, n45);
   not (n10738, n4570);
   or (n10739, n10737, n10738);
   nor (n1074, n1073, n710);
   or (n10740, n4570, n45);
   nand (n10741, n10739, n10740);
   not (n10742, n10741);
   or (n10743, n10736, n10742);
   nand (n10744, n9958, n4215);
   nand (n10745, n10743, n10744);
   nand (n10746, n10735, n10745);
   buf (n10747, n10746);
   not (n10748, n10747);
   and (n10749, n10732, n10748);
   buf (n1075, n1074);
   not (n10750, n10732);
   and (n10751, n10750, n10747);
   nor (n10752, n10749, n10751);
   xnor (n10753, n10667, n10656);
   or (n10754, n10752, n10753);
   or (n10755, n10732, n10747);
   nand (n10756, n10754, n10755);
   not (n10757, n10756);
   and (n10758, n10707, n10757);
   and (n10759, n10697, n10702);
   and (n1076, n1072, n1075);
   nor (n10760, n10758, n10759);
   not (n10761, n10760);
   or (n10762, n10696, n10761);
   or (n10763, n10760, n10695);
   nand (n10764, n10762, n10763);
   not (n10765, n10764);
   and (n10766, n10707, n10756);
   not (n10767, n10707);
   and (n10768, n10767, n10757);
   nor (n10769, n10766, n10768);
   and (n1077, n1039, n1036);
   not (n10770, n10769);
   not (n10771, n10733);
   nor (n10772, n4924, n3363);
   nand (n10773, n10772, n43);
   not (n10774, n4944);
   not (n10775, n4924);
   or (n10776, n10774, n10775);
   nand (n10777, n10776, n4661);
   not (n10778, n10777);
   and (n10779, n10773, n10153, n10778);
   nor (n1078, n1076, n1077);
   not (n10780, n10779);
   or (n10781, n10771, n10780);
   or (n10782, n10779, n10733);
   nand (n10783, n10781, n10782);
   not (n10784, n10783);
   or (n10785, n9910, n4937);
   not (n10786, n4226);
   or (n10787, n9753, n10786);
   nand (n10788, n10785, n10787);
   or (n10789, n10784, n10788);
   or (n1079, n1068, n1078);
   not (n10790, n10733);
   or (n10791, n10779, n10790);
   nand (n10792, n10789, n10791);
   not (n10793, n10745);
   nand (n10794, n10793, n10734);
   nand (n10795, n10746, n10794);
   or (n10796, n9880, n4383);
   or (n10797, n9885, n10644);
   nand (n10798, n10796, n10797);
   xor (n10799, n10795, n10798);
   buf (n108, n11417);
   nand (n1080, n1079, n1067);
   or (n10800, n10792, n10799);
   not (n10801, n10798);
   or (n10802, n10795, n10801);
   nand (n10803, n10800, n10802);
   xor (n10804, n10643, n10647);
   xor (n10805, n10803, n10804);
   xor (n10806, n10752, n10753);
   and (n10807, n10805, n10806);
   and (n10808, n10803, n10804);
   nor (n10809, n10807, n10808);
   and (n1081, n423, n647);
   not (n10810, n10809);
   or (n10811, n10770, n10810);
   or (n10812, n10809, n10769);
   nand (n10813, n10811, n10812);
   not (n10814, n10813);
   not (n10815, n10792);
   and (n10816, n10799, n10815);
   not (n10817, n10799);
   and (n10818, n10817, n10792);
   nor (n10819, n10816, n10818);
   and (n1082, n42, n60);
   not (n10820, n4983);
   not (n10821, n9811);
   or (n10822, n10820, n10821);
   or (n10823, n10104, n4383);
   nand (n10824, n10822, n10823);
   not (n10825, n4972);
   not (n10826, n10205);
   or (n10827, n10825, n10826);
   nand (n10828, n9958, n10741);
   nand (n10829, n10827, n10828);
   nor (n1083, n1081, n1082);
   xor (n10830, n10824, n10829);
   not (n10831, n9751);
   nand (n10832, n10831, n51);
   nand (n10833, n10832, n9652);
   not (n10834, n10351);
   nand (n10835, n10834, n45);
   and (n10836, n10153, n10835);
   not (n10837, n4926);
   nand (n10838, n10837, n10351);
   nand (n10839, n10836, n10838);
   and (n1084, n421, n1083);
   nor (n10840, n10833, n10839);
   and (n10841, n10830, n10840);
   and (n10842, n10824, n10829);
   nor (n10843, n10841, n10842);
   not (n10844, n10724);
   not (n10845, n10728);
   and (n10846, n10844, n10845);
   and (n10847, n10724, n10728);
   nor (n10848, n10846, n10847);
   xor (n10849, n10843, n10848);
   and (n1085, n513, n1027);
   and (n10850, n10819, n10849);
   and (n10851, n10843, n10848);
   nor (n10852, n10850, n10851);
   not (n10853, n10852);
   xor (n10854, n10803, n10804);
   xor (n10855, n10854, n10806);
   not (n10856, n10855);
   or (n10857, n10853, n10856);
   not (n10858, n4572);
   or (n10859, n9948, n10858);
   nor (n1086, n1084, n1085);
   and (n10860, n4213, n47);
   not (n10861, n4213);
   and (n10862, n10861, n3564);
   nor (n10863, n10860, n10862);
   or (n10864, n9957, n10863);
   nand (n10865, n10859, n10864);
   not (n10866, n10865);
   and (n10867, n10772, n45);
   not (n10868, n4580);
   not (n10869, n4924);
   not (n1087, n1086);
   or (n10870, n10868, n10869);
   nand (n10871, n10870, n4608);
   not (n10872, n10871);
   nand (n10873, n10872, n10153);
   nor (n10874, n10867, n10873);
   not (n10875, n10874);
   not (n10876, n10832);
   and (n10877, n10875, n10876);
   and (n10878, n10874, n10832);
   nor (n10879, n10877, n10878);
   not (n1088, n1087);
   not (n10880, n10879);
   not (n10881, n10880);
   or (n10882, n10866, n10881);
   not (n10883, n10832);
   nand (n10884, n10883, n10874);
   nand (n10885, n10882, n10884);
   not (n10886, n10885);
   nand (n10887, n10833, n10839);
   not (n10888, n10887);
   nor (n10889, n10888, n10840);
   or (n1089, n36, n66);
   not (n10890, n10889);
   and (n10891, n10886, n10890);
   xnor (n10892, n10885, n10889);
   not (n10893, n10892);
   not (n10894, n10863);
   not (n10895, n10894);
   not (n10896, n10205);
   or (n10897, n10895, n10896);
   nand (n10898, n9956, n4972);
   nand (n10899, n10897, n10898);
   buf (n109, n11417);
   nand (n1090, n1089, n1002);
   not (n10900, n9751);
   not (n10901, n4937);
   and (n10902, n10900, n10901);
   and (n10903, n9697, n10717);
   nor (n10904, n10902, n10903);
   xnor (n10905, n10899, n10904);
   and (n10906, n3239, n49);
   not (n10907, n3239);
   and (n10908, n10907, n610);
   nor (n10909, n10906, n10908);
   or (n1091, n245, n1090);
   or (n10910, n9880, n10909);
   not (n10911, n4983);
   or (n10912, n10104, n10911);
   nand (n10913, n10910, n10912);
   not (n10914, n10913);
   and (n10915, n10905, n10914);
   not (n10916, n10905);
   and (n10917, n10916, n10913);
   nor (n10918, n10915, n10917);
   and (n10919, n10893, n10918);
   or (n1092, n400, n995);
   nor (n10920, n10891, n10919);
   not (n10921, n10920);
   not (n10922, n10899);
   not (n10923, n10922);
   not (n10924, n10904);
   and (n10925, n10923, n10924);
   and (n10926, n10905, n10913);
   nor (n10927, n10925, n10926);
   and (n10928, n10788, n10783);
   not (n10929, n10788);
   nand (n1093, n1091, n1092);
   and (n10930, n10929, n10784);
   or (n10931, n10928, n10930);
   xor (n10932, n10927, n10931);
   xor (n10933, n10824, n10829);
   xor (n10934, n10933, n10840);
   xor (n10935, n10932, n10934);
   not (n10936, n10935);
   or (n10937, n10921, n10936);
   not (n10938, n4642);
   not (n10939, n10938);
   not (n1094, n1093);
   not (n10940, n9947);
   or (n10941, n10939, n10940);
   nand (n10942, n9958, n4572);
   nand (n10943, n10941, n10942);
   not (n10944, n10943);
   or (n10945, n3238, n3334);
   nand (n10946, n10945, n4680);
   and (n10947, n10946, n9810);
   nor (n10948, n9883, n4518);
   nor (n10949, n10947, n10948);
   not (n1095, n1094);
   not (n10950, n10949);
   or (n10951, n10944, n10950);
   or (n10952, n10949, n10943);
   nand (n10953, n10951, n10952);
   not (n10954, n10953);
   not (n10955, n9883);
   nand (n10956, n10955, n51);
   nand (n10957, n10956, n9763);
   not (n10958, n10957);
   not (n10959, n4602);
   and (n1096, n44, n58);
   not (n10960, n10959);
   not (n10961, n3737);
   or (n10962, n10960, n10961);
   nand (n10963, n10093, n47);
   and (n10964, n10153, n10963);
   nand (n10965, n10962, n10964);
   not (n10966, n10965);
   or (n10967, n10958, n10966);
   or (n10968, n10957, n10965);
   nand (n10969, n10967, n10968);
   not (n1097, n44);
   not (n10970, n10969);
   or (n10971, n10954, n10970);
   or (n10972, n10969, n10953);
   nand (n10973, n10971, n10972);
   not (n10974, n10973);
   not (n10975, n10974);
   not (n10976, n4760);
   not (n10977, n10976);
   not (n10978, n9947);
   or (n10979, n10977, n10978);
   and (n1098, n1097, n769);
   nand (n10980, n10938, n9956);
   nand (n10981, n10979, n10980);
   not (n10982, n10981);
   not (n10983, n10982);
   not (n10984, n10956);
   and (n10985, n10983, n10984);
   not (n10986, n10956);
   not (n10987, n10981);
   or (n10988, n10986, n10987);
   or (n10989, n10981, n10956);
   nor (n1099, n1096, n1098);
   nand (n10990, n10988, n10989);
   not (n10991, n47);
   not (n10992, n10094);
   or (n10993, n10991, n10992);
   or (n10994, n3768, n47);
   nand (n10995, n10994, n4713);
   nor (n10996, n10154, n10995);
   nand (n10997, n10993, n10996);
   not (n10998, n10997);
   and (n10999, n10990, n10998);
   buf (n11, g10);
   buf (n110, n11417);
   and (n1100, n798, n1099);
   nor (n11000, n10985, n10999);
   not (n11001, n11000);
   and (n11002, n10975, n11001);
   not (n11003, n10976);
   not (n11004, n9958);
   or (n11005, n11003, n11004);
   not (n11006, n9945);
   and (n11007, n11006, n51);
   not (n11008, n9943);
   and (n11009, n11008, n3334);
   and (n1101, n44, n57);
   nor (n11010, n11007, n11009);
   nand (n11011, n11005, n11010);
   nand (n11012, n9956, n51);
   nand (n11013, n9890, n11012);
   and (n11014, n3363, n49);
   not (n11015, n3363);
   not (n11016, n4791);
   and (n11017, n11015, n11016);
   nor (n11018, n11014, n11017);
   nand (n11019, n11018, n10153);
   not (n1102, n44);
   nor (n11020, n11013, n11019);
   not (n11021, n11020);
   not (n11022, n11018);
   not (n11023, n10153);
   or (n11024, n11022, n11023);
   nand (n11025, n11024, n11013);
   nand (n11026, n11021, n11025);
   xnor (n11027, n11011, n11026);
   and (n11028, n4549, n10400);
   nand (n11029, n3768, n1005);
   and (n1103, n1102, n498);
   and (n11030, n11029, n10093);
   nor (n11031, n11028, n11030);
   not (n11032, n11031);
   not (n11033, n11012);
   and (n11034, n11029, n10347);
   nor (n11035, n11034, n51);
   nor (n11036, n11033, n11035);
   nor (n11037, n11032, n11036);
   and (n11038, n11027, n11037);
   not (n11039, n11026);
   nor (n1104, n1101, n1103);
   and (n11040, n11039, n11011);
   nor (n11041, n11038, n11040);
   not (n11042, n10990);
   not (n11043, n10997);
   and (n11044, n11042, n11043);
   and (n11045, n10990, n10997);
   nor (n11046, n11044, n11045);
   xor (n11047, n11046, n11020);
   or (n11048, n11041, n11047);
   not (n11049, n11046);
   and (n1105, n1104, n556);
   nand (n11050, n11049, n11020);
   nand (n11051, n11048, n11050);
   not (n11052, n11000);
   not (n11053, n10973);
   or (n11054, n11052, n11053);
   or (n11055, n11000, n10973);
   nand (n11056, n11054, n11055);
   and (n11057, n11051, n11056);
   nor (n11058, n11002, n11057);
   not (n11059, n10943);
   nor (n1106, n1100, n1105);
   not (n11060, n11059);
   not (n11061, n10949);
   and (n11062, n11060, n11061);
   not (n11063, n10969);
   and (n11064, n11063, n10953);
   nor (n11065, n11062, n11064);
   not (n11066, n9885);
   not (n11067, n10909);
   and (n11068, n11066, n11067);
   not (n11069, n4518);
   not (n1107, n1106);
   and (n11070, n9811, n11069);
   nor (n11071, n11068, n11070);
   xor (n11072, n11071, n10968);
   not (n11073, n11072);
   not (n11074, n10865);
   not (n11075, n10879);
   or (n11076, n11074, n11075);
   or (n11077, n10865, n10879);
   nand (n11078, n11076, n11077);
   not (n11079, n11078);
   not (n1108, n1107);
   and (n11080, n11073, n11079);
   and (n11081, n11078, n11072);
   nor (n11082, n11080, n11081);
   and (n11083, n11065, n11082);
   not (n11084, n11065);
   not (n11085, n11082);
   and (n11086, n11084, n11085);
   nor (n11087, n11083, n11086);
   or (n11088, n11058, n11087);
   or (n11089, n11085, n11065);
   or (n1109, n1095, n1108);
   nand (n11090, n11088, n11089);
   not (n11091, n11090);
   not (n11092, n11072);
   not (n11093, n11092);
   not (n11094, n11078);
   and (n11095, n11093, n11094);
   and (n11096, n10968, n11071);
   nor (n11097, n11095, n11096);
   not (n11098, n11097);
   xnor (n11099, n10918, n10892);
   buf (n111, n11417);
   nand (n1110, n1106, n1093);
   not (n11100, n11099);
   or (n11101, n11098, n11100);
   or (n11102, n11097, n11099);
   nand (n11103, n11101, n11102);
   not (n11104, n11103);
   or (n11105, n11091, n11104);
   not (n11106, n11099);
   nand (n11107, n11106, n11097);
   nand (n11108, n11105, n11107);
   xor (n11109, n10935, n10920);
   nand (n1111, n1109, n1110);
   nand (n11110, n11108, n11109);
   nand (n11111, n10937, n11110);
   xnor (n11112, n10819, n10849);
   not (n11113, n10934);
   not (n11114, n10932);
   or (n11115, n11113, n11114);
   or (n11116, n10927, n10931);
   nand (n11117, n11115, n11116);
   xor (n11118, n11112, n11117);
   and (n11119, n11111, n11118);
   not (n1112, n1111);
   and (n11120, n11112, n11117);
   nor (n11121, n11119, n11120);
   xnor (n11122, n10855, n10852);
   or (n11123, n11121, n11122);
   nand (n11124, n10857, n11123);
   not (n11125, n11124);
   or (n11126, n10814, n11125);
   not (n11127, n10809);
   nand (n11128, n11127, n10769);
   nand (n11129, n11126, n11128);
   or (n1113, n1088, n1112);
   not (n11130, n11129);
   or (n11131, n10765, n11130);
   not (n11132, n10695);
   nand (n11133, n11132, n10760);
   nand (n11134, n11131, n11133);
   not (n11135, n11134);
   or (n11136, n10694, n11135);
   not (n11137, n10686);
   nand (n11138, n11137, n10689);
   nand (n11139, n11136, n11138);
   nand (n1114, n1107, n1093);
   not (n11140, n11139);
   not (n11141, n11140);
   or (n11142, n10626, n11141);
   not (n11143, n10624);
   or (n11144, n10438, n10486);
   not (n11145, n10622);
   not (n11146, n10617);
   or (n11147, n11145, n11146);
   or (n11148, n10617, n10622);
   nand (n11149, n11147, n11148);
   nand (n1115, n1113, n1114);
   nand (n11150, n11144, n11149);
   and (n11151, n11143, n11150);
   not (n11152, n10604);
   not (n11153, n10614);
   and (n11154, n11152, n11153);
   and (n11155, n10604, n10614);
   nor (n11156, n11154, n11155);
   and (n11157, n11156, n10615);
   nor (n11158, n11151, n11157);
   nand (n11159, n11142, n11158);
   xor (n1116, n1080, n1115);
   not (n11160, n10589);
   not (n11161, n10603);
   and (n11162, n11160, n11161);
   and (n11163, n10578, n10588);
   nor (n11164, n11162, n11163);
   and (n11165, n10576, n10538);
   not (n11166, n10569);
   and (n11167, n10548, n11166);
   nor (n11168, n11165, n11167);
   xnor (n11169, n10132, n10133);
   not (n1117, n40);
   xor (n11170, n11168, n11169);
   xor (n11171, n10083, n10097);
   xor (n11172, n11171, n10121);
   not (n11173, n11172);
   xor (n11174, n11173, n10547);
   or (n11175, n10587, n10579);
   or (n11176, n10586, n10583);
   nand (n11177, n11175, n11176);
   xnor (n11178, n11174, n11177);
   xor (n11179, n11170, n11178);
   not (n1118, n62);
   xnor (n11180, n11164, n11179);
   or (n11181, n11159, n11180);
   or (n11182, n11179, n11164);
   nand (n11183, n11181, n11182);
   xnor (n11184, n10127, n10136);
   and (n11185, n11174, n11177);
   and (n11186, n11173, n10547);
   nor (n11187, n11185, n11186);
   xnor (n11188, n10051, n10024);
   xnor (n11189, n11187, n11188);
   and (n1119, n1117, n1118);
   xor (n11190, n11184, n11189);
   xor (n11191, n11168, n11169);
   and (n11192, n11191, n11178);
   and (n11193, n11168, n11169);
   nor (n11194, n11192, n11193);
   xor (n11195, n11190, n11194);
   and (n11196, n11183, n11195);
   and (n11197, n11190, n11194);
   nor (n11198, n11196, n11197);
   xor (n11199, n10022, n10055);
   buf (n112, n11417);
   and (n1120, n40, n62);
   xor (n11200, n11199, n10062);
   or (n11201, n11189, n11184);
   or (n11202, n11187, n11188);
   nand (n11203, n11201, n11202);
   xor (n11204, n10138, n11203);
   xor (n11205, n11200, n11204);
   nand (n11206, n11198, n11205);
   xor (n11207, n10061, n10062);
   xor (n11208, n11207, n10138);
   or (n11209, n11203, n11208);
   nor (n1121, n1119, n1120);
   nand (n11210, n11206, n11209);
   xor (n11211, n10059, n10141);
   nand (n11212, n11210, n11211);
   nand (n11213, n10143, n11212);
   xor (n11214, n9860, n9907);
   xor (n11215, n11214, n9978);
   not (n11216, n11215);
   xor (n11217, n9987, n9988);
   and (n11218, n11217, n10058);
   and (n11219, n9987, n9988);
   and (n1122, n857, n1121);
   nor (n11220, n11218, n11219);
   not (n11221, n11220);
   and (n11222, n11216, n11221);
   and (n11223, n11220, n11215);
   nor (n11224, n11222, n11223);
   or (n11225, n11213, n11224);
   not (n11226, n11215);
   nand (n11227, n11226, n11220);
   nand (n11228, n11225, n11227);
   not (n11229, n11228);
   and (n1123, n40, n61);
   or (n11230, n9986, n11229);
   not (n11231, n9858);
   nand (n11232, n11231, n9981);
   nand (n11233, n11230, n11232);
   not (n11234, n11233);
   or (n11235, n9856, n11234);
   not (n11236, n9789);
   nand (n11237, n11236, n9851);
   nand (n11238, n11235, n11237);
   not (n11239, n11238);
   not (n1124, n40);
   or (n11240, n9788, n11239);
   not (n11241, n9783);
   nand (n11242, n11241, n9717);
   nand (n11243, n11240, n11242);
   not (n11244, n11243);
   or (n11245, n9716, n11244);
   not (n11246, n9667);
   nand (n11247, n11246, n9711);
   nand (n11248, n11245, n11247);
   not (n11249, n11248);
   and (n1125, n1124, n692);
   not (n11250, n11249);
   xor (n11251, n9632, n9638);
   and (n11252, n11251, n9666);
   and (n11253, n9632, n9638);
   nor (n11254, n11252, n11253);
   not (n11255, n11254);
   not (n11256, n2837);
   not (n11257, n9597);
   or (n11258, n11256, n11257);
   or (n11259, n9603, n5781);
   nor (n1126, n1123, n1125);
   nand (n11260, n11258, n11259);
   xor (n11261, n11260, n9605);
   and (n11262, n9577, n2953);
   and (n11263, n10420, n9574);
   nor (n11264, n11262, n11263);
   xor (n11265, n11261, n11264);
   xor (n11266, n9636, n9624);
   and (n11267, n11266, n2956);
   and (n11268, n9636, n9624);
   nor (n11269, n11267, n11268);
   and (n1127, n273, n1126);
   xor (n11270, n11265, n11269);
   or (n11271, n9612, n9631);
   or (n11272, n9626, n9630);
   nand (n11273, n11271, n11272);
   xnor (n11274, n11270, n11273);
   not (n11275, n11274);
   and (n11276, n11255, n11275);
   and (n11277, n11254, n11274);
   nor (n11278, n11276, n11277);
   not (n11279, n11278);
   nor (n1128, n1122, n1127);
   not (n11280, n11279);
   and (n11281, n11250, n11280);
   nor (n11282, n11248, n11278);
   nor (n11283, n11281, n11282);
   not (n11284, n11283);
   nand (n11285, n11284, n9565);
   nand (n11286, n9537, n9567, n9569, n11285);
   not (n11287, n9561);
   not (n11288, n9524);
   or (n11289, n11287, n11288);
   and (n1129, n38, n64);
   and (n11290, n9534, n9062);
   nand (n11291, n11289, n11290);
   nor (n11292, n9534, n9565);
   nand (n11293, n9561, n11292, n9524);
   xor (n11294, n11243, n9715);
   nand (n11295, n11294, n9565);
   nand (n11296, n11291, n11293, n11295);
   nor (n11297, n9557, n9554);
   nand (n11298, n6575, n11297);
   not (n11299, n11298);
   buf (n113, n11417);
   not (n1130, n38);
   not (n11300, n11299);
   nor (n11301, n9521, n9499);
   and (n11302, n9546, n9549, n1);
   nor (n11303, n11302, n9540);
   nand (n11304, n9550, n11303);
   nand (n11305, n11301, n11304);
   not (n11306, n11305);
   or (n11307, n11300, n11306);
   nand (n11308, n11307, n9062);
   nor (n11309, n9560, n9523);
   not (n1131, n64);
   or (n11310, n11308, n11309);
   buf (n11311, n11238);
   xnor (n11312, n9787, n11311);
   or (n11313, n11312, n9062);
   nand (n11314, n11310, n11313);
   xnor (n11315, n11233, n9855);
   or (n11316, n11315, n9062);
   buf (n11317, n9499);
   not (n11318, n11317);
   and (n11319, n11318, n9522);
   and (n1132, n1130, n1131);
   nor (n11320, n11319, n11304);
   nand (n11321, n9062, n11305);
   or (n11322, n11320, n11321);
   nand (n11323, n11316, n11322);
   not (n11324, n9565);
   or (n11325, n9596, n5781);
   or (n11326, n9603, n2878);
   nand (n11327, n11325, n11326);
   or (n11328, n11327, n10420);
   nand (n11329, n11327, n10420);
   nor (n1133, n1129, n1132);
   nand (n11330, n11328, n11329);
   xnor (n11331, n11330, n2836);
   xnor (n11332, n11331, n11264);
   xor (n11333, n11260, n9605);
   and (n11334, n11333, n11264);
   and (n11335, n11260, n9605);
   nor (n11336, n11334, n11335);
   or (n11337, n11332, n11336);
   or (n11338, n11331, n11264);
   nand (n11339, n11337, n11338);
   not (n1134, n1133);
   not (n11340, n11339);
   or (n11341, n9596, n2878);
   not (n11342, n9593);
   or (n11343, n10179, n11342);
   nand (n11344, n11341, n11343);
   xor (n11345, n11344, n5780);
   and (n11346, n11330, n2836);
   not (n11347, n10420);
   and (n11348, n11327, n11347);
   nor (n11349, n11346, n11348);
   not (n1135, n376);
   and (n11350, n11345, n11349);
   not (n11351, n11345);
   not (n11352, n11349);
   and (n11353, n11351, n11352);
   nor (n11354, n11350, n11353);
   not (n11355, n11354);
   and (n11356, n11340, n11355);
   and (n11357, n11339, n11354);
   nor (n11358, n11356, n11357);
   xor (n11359, n11332, n11336);
   or (n1136, n1134, n1135);
   not (n11360, n11359);
   and (n11361, n11270, n11273);
   and (n11362, n11265, n11269);
   nor (n11363, n11361, n11362);
   not (n11364, n11363);
   or (n11365, n11360, n11364);
   or (n11366, n11363, n11359);
   nand (n11367, n11365, n11366);
   not (n11368, n11367);
   not (n11369, n11274);
   not (n1137, n38);
   nor (n11370, n11369, n11254);
   nor (n11371, n11282, n11370);
   not (n11372, n11371);
   or (n11373, n11368, n11372);
   not (n11374, n11363);
   nand (n11375, n11374, n11359);
   nand (n11376, n11373, n11375);
   xnor (n11377, n11358, n11376);
   not (n11378, n11377);
   or (n11379, n11324, n11378);
   not (n1138, n63);
   buf (n11380, n6575);
   not (n11381, n11380);
   nand (n11382, n11305, n11381, n9062);
   nand (n11383, n11379, n11382);
   not (n11384, n9565);
   xor (n11385, n11367, n11371);
   not (n11386, n11385);
   or (n11387, n11384, n11386);
   nand (n11388, n11387, n11382);
   not (n11389, n9565);
   and (n1139, n1137, n1138);
   and (n11390, n10178, n244);
   nor (n11391, n10178, n244);
   nor (n11392, n11390, n11391, n2834);
   not (n11393, n11392);
   and (n11394, n11352, n11345);
   and (n11395, n11344, n5780);
   nor (n11396, n11394, n11395);
   not (n11397, n11396);
   or (n11398, n11393, n11397);
   or (n11399, n11396, n11392);
   buf (n114, n11417);
   and (n1140, n38, n63);
   nand (n11400, n11398, n11399);
   not (n11401, n11400);
   not (n11402, n11358);
   not (n11403, n11402);
   not (n11404, n11376);
   or (n11405, n11403, n11404);
   not (n11406, n11354);
   nand (n11407, n11406, n11339);
   nand (n11408, n11405, n11407);
   not (n11409, n11408);
   nor (n1141, n1139, n1140);
   or (n11410, n11401, n11409);
   or (n11411, n11408, n11400);
   nand (n11412, n11410, n11411);
   not (n11413, n11412);
   or (n11414, n11389, n11413);
   nand (n11415, n11414, n11382);
   not (n11416, n11382);
   not (n11417, n11380);
   nand (n11418, n11417, n9062);
   nor (n11419, n11418, n11305);
   nand (n1142, n310, n1141);
   not (n11420, n11317);
   not (n11421, n9521);
   or (n11422, n11420, n11421);
   nand (n11423, n11422, n9062);
   not (n11424, n11423);
   buf (n11425, n9478);
   or (n11426, n11425, n9498);
   nand (n11427, n11426, n9062);
   or (n11428, n11427, n11318);
   xnor (n11429, n11213, n11224);
   nand (n1143, n1136, n1142);
   or (n11430, n11429, n9062);
   nand (n11431, n11428, n11430);
   not (n11432, n9451);
   not (n11433, n9477);
   or (n11434, n11432, n11433);
   nand (n11435, n11434, n9062);
   or (n11436, n11435, n11425);
   not (n11437, n11210);
   not (n11438, n11211);
   and (n11439, n11437, n11438);
   xnor (n1144, n1128, n1143);
   not (n11440, n11212);
   nor (n11441, n11439, n11440);
   or (n11442, n11441, n9062);
   nand (n11443, n11436, n11442);
   not (n11444, n11301);
   not (n11445, n9449);
   not (n11446, n11445);
   buf (n11447, n9389);
   not (n11448, n9417);
   nand (n11449, n11447, n11448);
   not (n1145, n1144);
   nand (n11450, n11446, n11449);
   nand (n11451, n11450, n9451, n9062);
   or (n11452, n11205, n11198);
   nand (n11453, n11452, n11206);
   nand (n11454, n11453, n9565);
   nand (n11455, n11451, n11454);
   not (n11456, n11447);
   nand (n11457, n11456, n9417);
   nand (n11458, n11457, n11449, n9062);
   xor (n11459, n11195, n11183);
   and (n1146, n46, n56);
   nand (n11460, n11459, n9565);
   nand (n11461, n11458, n11460);
   not (n11462, n9565);
   xor (n11463, n11180, n11159);
   not (n11464, n11463);
   or (n11465, n11462, n11464);
   nand (n11466, n9382, n1);
   nand (n11467, n11466, n9386);
   nand (n11468, n11467, n9375);
   not (n11469, n9126);
   not (n1147, n46);
   not (n11470, n11469);
   and (n11471, n11468, n11470);
   nor (n11472, n11471, n9565);
   nand (n11473, n11472, n11456);
   nand (n11474, n11465, n11473);
   not (n11475, n11467);
   not (n11476, n11475);
   buf (n11477, n9349);
   buf (n11478, n9374);
   and (n11479, n11477, n11478);
   and (n1148, n1147, n479);
   buf (n11480, n9358);
   nand (n11481, n11479, n11480);
   not (n11482, n11481);
   or (n11483, n11476, n11482);
   nand (n11484, n11483, n9062);
   not (n11485, n11468);
   or (n11486, n11484, n11485);
   buf (n11487, n11139);
   or (n11488, n11487, n10486);
   xnor (n11489, n10486, n11487);
   nor (n1149, n1146, n1148);
   nor (n11490, n11489, n10438);
   not (n11491, n11490);
   nand (n11492, n11488, n11491);
   not (n11493, n11149);
   or (n11494, n11492, n11493);
   nand (n11495, n11494, n10623);
   not (n11496, n11495);
   not (n11497, n11156);
   and (n11498, n11496, n11497);
   and (n11499, n11495, n11156);
   buf (n115, n11417);
   and (n1150, n913, n1149);
   nor (n11500, n11498, n11499);
   or (n11501, n11500, n9062);
   nand (n11502, n11486, n11501);
   or (n11503, n11479, n11480);
   nand (n11504, n11503, n9062);
   not (n11505, n11481);
   or (n11506, n11504, n11505);
   xnor (n11507, n11492, n11493);
   or (n11508, n11507, n9062);
   nand (n11509, n11506, n11508);
   not (n1151, n627);
   or (n11510, n11478, n11477);
   nand (n11511, n11510, n9062);
   or (n11512, n11511, n11479);
   and (n11513, n11489, n10438);
   nor (n11514, n11513, n11490);
   or (n11515, n11514, n9062);
   nand (n11516, n11512, n11515);
   buf (n11517, n9322);
   not (n11518, n9335);
   nor (n11519, n11517, n11518);
   and (n1152, n1151, n1015);
   or (n11520, n11519, n9347);
   nand (n11521, n11520, n9062);
   or (n11522, n11477, n11521);
   xnor (n11523, n11134, n10693);
   or (n11524, n11523, n9062);
   nand (n11525, n11522, n11524);
   not (n11526, n11518);
   not (n11527, n11517);
   or (n11528, n11526, n11527);
   nand (n11529, n11528, n9062);
   nor (n1153, n1150, n1152);
   or (n11530, n11529, n11519);
   xnor (n11531, n11129, n10764);
   or (n11532, n11531, n9062);
   nand (n11533, n11530, n11532);
   buf (n11534, n9309);
   or (n11535, n11534, n9321);
   nand (n11536, n11535, n9062);
   not (n11537, n11517);
   or (n11538, n11536, n11537);
   xnor (n11539, n11124, n10813);
   or (n1154, n1145, n1153);
   or (n11540, n11539, n9062);
   nand (n11541, n11538, n11540);
   not (n11542, n9565);
   xor (n11543, n11121, n11122);
   not (n11544, n11543);
   or (n11545, n11542, n11544);
   not (n11546, n9307);
   not (n11547, n11546);
   not (n11548, n9273);
   nand (n11549, n11548, n9293);
   not (n1155, n1143);
   not (n11550, n11549);
   or (n11551, n11547, n11550);
   nor (n11552, n11534, n9565);
   nand (n11553, n11551, n11552);
   nand (n11554, n11545, n11553);
   not (n11555, n9293);
   not (n11556, n11555);
   not (n11557, n9273);
   or (n11558, n11556, n11557);
   nand (n11559, n11558, n9062);
   or (n1156, n1155, n1128);
   not (n11560, n11559);
   nand (n11561, n11560, n11549);
   xor (n11562, n11111, n11118);
   nand (n11563, n11562, n9565);
   nand (n11564, n11561, n11563);
   xnor (n11565, n11108, n11109);
   or (n11566, n11565, n9062);
   not (n11567, n9271);
   not (n11568, n11567);
   buf (n11569, n9241);
   nand (n1157, n1154, n1156);
   not (n11570, n9255);
   nand (n11571, n11569, n11570);
   nand (n11572, n11568, n11571);
   nand (n11573, n11572, n9273, n9062);
   nand (n11574, n11566, n11573);
   not (n11575, n9225);
   nand (n11576, n9213, n9240);
   nand (n11577, n11575, n11576);
   nand (n11578, n11577, n9062);
   or (n11579, n11578, n11569);
   and (n1158, n1116, n1157);
   xnor (n11580, n11058, n11087);
   or (n11581, n11580, n9062);
   nand (n11582, n11579, n11581);
   not (n11583, n11571);
   or (n11584, n11569, n11570);
   nand (n11585, n11584, n9062);
   or (n11586, n11583, n11585);
   xnor (n11587, n11090, n11103);
   or (n11588, n11587, n9062);
   nand (n11589, n11586, n11588);
   and (n1159, n1080, n1115);
   not (n11590, n11576);
   or (n11591, n9213, n9240);
   nand (n11592, n11591, n9062);
   or (n11593, n11590, n11592);
   xnor (n11594, n11051, n11056);
   or (n11595, n11594, n9062);
   nand (n11596, n11593, n11595);
   not (n11597, n9985);
   not (n11598, n11228);
   not (n11599, n11598);
   buf (n116, n11417);
   nor (n1160, n1158, n1159);
   or (n11600, n11597, n11599);
   or (n11601, n11598, n9985);
   nand (n11602, n11600, n11601);
   nand (n11603, n11602, n9565);
   not (n11604, n9209);
   and (n11605, n9191, n11604);
   not (n11606, n9191);
   and (n11607, n11606, n9209);
   nor (n11608, n11605, n11607);
   or (n11609, n11608, n9565);
   not (n1161, n245);
   xnor (n11610, n11041, n11047);
   or (n11611, n11610, n9062);
   nand (n11612, n11609, n11611);
   xnor (n11613, n9141, n9187);
   or (n11614, n11613, n9565);
   xnor (n11615, n11027, n11037);
   or (n11616, n11615, n9062);
   nand (n11617, n11614, n11616);
   and (n11618, n17, n9184);
   not (n11619, n17);
   not (n1162, n998);
   not (n11620, n9184);
   and (n11621, n11619, n11620);
   nor (n11622, n11618, n11621);
   and (n11623, n11622, n9176);
   nor (n11624, n11622, n9176);
   nor (n11625, n11623, n11624);
   or (n11626, n11625, n9565);
   not (n11627, n11036);
   not (n11628, n11031);
   and (n11629, n11627, n11628);
   and (n1163, n1161, n1162);
   and (n11630, n11036, n11031);
   nor (n11631, n11629, n11630);
   or (n11632, n11631, n9062);
   nand (n11633, n11626, n11632);
   or (n11634, n3768, n1005);
   nand (n11635, n11634, n11029);
   and (n11636, n11635, n10400);
   and (n11637, n4875, n3768);
   nor (n11638, n11636, n11637);
   or (n11639, n11638, n11035, n9062);
   nor (n1164, n253, n719);
   and (n11640, n9174, n3489);
   not (n11641, n9174);
   and (n11642, n11641, n18);
   nor (n11643, n11640, n11642);
   and (n11644, n11643, n9157);
   nor (n11645, n11643, n9157);
   nor (n11646, n11644, n11645);
   or (n11647, n11646, n9565);
   nand (n11648, n11639, n11647);
   or (n11649, n9155, n19);
   nor (n1165, n1163, n1164);
   nand (n11650, n11649, n9062);
   or (n11651, n11650, n9157);
   or (n11652, n4875, n9062);
   nand (n11653, n11651, n11652);
   not (n11654, n6279);
   not (n11655, n6219);
   and (n11656, n11654, n11655);
   not (n11657, n6280);
   nor (n11658, n11656, n11657);
   or (n11659, n11658, n6569);
   not (n1166, n1165);
   and (n11660, n8861, n8903);
   not (n11661, n8904);
   nor (n11662, n11660, n11661);
   or (n11663, n11662, n1);
   nand (n11664, n11659, n11663);
   xnor (n11665, n6264, n6276);
   or (n11666, n11665, n6569);
   xnor (n11667, n8898, n8888);
   or (n11668, n11667, n1);
   nand (n11669, n11666, n11668);
   not (n1167, n928);
   not (n11670, n1);
   xor (n11671, n97, n6233);
   xor (n11672, n11671, n6261);
   not (n11673, n11672);
   or (n11674, n11670, n11673);
   xnor (n11675, n8870, n8885);
   or (n11676, n11675, n1);
   nand (n11677, n11674, n11676);
   xnor (n11678, n6248, n6257);
   or (n11679, n11678, n6569);
   not (n1168, n556);
   xnor (n11680, n8878, n8881);
   or (n11681, n11680, n1);
   nand (n11682, n11679, n11681);
   and (n11683, n83, n99);
   nor (n11684, n11683, n19);
   or (n11685, n11684, n8872, n1);
   or (n11686, n99, n6256);
   nand (n11687, n11686, n6257, n1);
   nand (n11688, n11685, n11687);
   not (n11689, n11424);
   or (n1169, n1167, n1168);
   not (n11690, n11444);
   or (n11691, n11689, n11690);
   nand (n11692, n11691, n11603);
   buf (n117, n11417);
   nand (n1170, n566, n1104);
   nand (n1171, n1169, n1170);
   not (n1172, n1171);
   or (n1173, n1166, n1172);
   or (n1174, n1171, n1165);
   nand (n1175, n1173, n1174);
   not (n1176, n1175);
   not (n1177, n715);
   and (n1178, n1176, n1177);
   and (n1179, n1175, n715);
   buf (n118, n11417);
   nor (n1180, n1178, n1179);
   xor (n1181, n905, n911);
   xor (n1182, n1181, n920);
   not (n1183, n1182);
   and (n1184, n1180, n1183);
   not (n1185, n1180);
   and (n1186, n1185, n1182);
   nor (n1187, n1184, n1186);
   or (n1188, n1160, n1187);
   or (n1189, n1180, n1182);
   buf (n119, n11417);
   nand (n1190, n1188, n1189);
   nand (n1191, n1055, n1190);
   not (n1192, n1054);
   nand (n1193, n1192, n993);
   and (n1194, n1191, n1193);
   not (n1195, n1194);
   not (n1196, n1195);
   not (n1197, n715);
   not (n1198, n1197);
   not (n1199, n1175);
   buf (n12, g11);
   buf (n120, n11417);
   or (n1200, n1198, n1199);
   not (n1201, n1165);
   nand (n1202, n1201, n1171);
   nand (n1203, n1200, n1202);
   xor (n1204, n699, n715);
   xor (n1205, n1204, n724);
   xor (n1206, n1203, n1205);
   and (n1207, n574, n586);
   not (n1208, n574);
   and (n1209, n1208, n587);
   buf (n121, n11417);
   nor (n1210, n1207, n1209);
   not (n1211, n1210);
   and (n1212, n1206, n1211);
   and (n1213, n1203, n1205);
   or (n1214, n1212, n1213);
   not (n1215, n1214);
   and (n1216, n1196, n1215);
   not (n1217, n1214);
   and (n1218, n1194, n1217);
   not (n1219, n1194);
   buf (n122, n11417);
   and (n1220, n1219, n1214);
   nor (n1221, n1218, n1220);
   not (n1222, n972);
   and (n1223, n971, n1222);
   not (n1224, n971);
   and (n1225, n1224, n972);
   nor (n1226, n1223, n1225);
   and (n1227, n1221, n1226);
   nor (n1228, n1216, n1227);
   buf (n1229, n1228);
   buf (n123, n11417);
   not (n1230, n1229);
   or (n1231, n986, n1230);
   xnor (n1232, n1226, n1221);
   xor (n1233, n1190, n1055);
   not (n1234, n1233);
   xnor (n1235, n1000, n1007);
   and (n1236, n1033, n1041);
   not (n1237, n1033);
   not (n1238, n1041);
   and (n1239, n1237, n1238);
   buf (n124, n11417);
   nor (n1240, n1236, n1239);
   xnor (n1241, n1235, n1240);
   not (n1242, n1241);
   and (n1243, n46, n57);
   not (n1244, n46);
   and (n1245, n1244, n498);
   nor (n1246, n1243, n1245);
   and (n1247, n535, n1246);
   and (n1248, n627, n1149);
   nor (n1249, n1247, n1248);
   buf (n125, n11417);
   xor (n1250, n40, n63);
   and (n1251, n857, n1250);
   and (n1252, n274, n1121);
   nor (n1253, n1251, n1252);
   xor (n1254, n1249, n1253);
   and (n1255, n423, n692);
   and (n1256, n42, n61);
   nor (n1257, n1255, n1256);
   and (n1258, n421, n1257);
   buf (n1259, n513);
   buf (n126, n11417);
   and (n1260, n1259, n1083);
   nor (n1261, n1258, n1260);
   and (n1262, n1254, n1261);
   and (n1263, n1249, n1253);
   nor (n1264, n1262, n1263);
   not (n1265, n1264);
   nand (n1266, n252, n67);
   and (n1267, n242, n36);
   nand (n1268, n1266, n1267);
   not (n1269, n52);
   buf (n127, n11417);
   not (n1270, n1061);
   not (n1271, n1270);
   or (n1272, n1269, n1271);
   nor (n1273, n50, n51);
   buf (n1274, n1273);
   or (n1275, n50, n52);
   or (n1276, n312, n51);
   nand (n1277, n1275, n1276);
   nor (n1278, n1274, n1277);
   nand (n1279, n1272, n1278);
   buf (n128, n11417);
   or (n1280, n1268, n1279);
   buf (n1281, n1280);
   not (n1282, n1281);
   and (n1283, n44, n59);
   not (n1284, n44);
   and (n1285, n1284, n578);
   nor (n1286, n1283, n1285);
   and (n1287, n566, n1286);
   and (n1288, n556, n1099);
   nor (n1289, n1287, n1288);
   buf (n129, n11417);
   not (n1290, n1289);
   not (n1291, n1290);
   not (n1292, n1038);
   not (n1293, n1072);
   not (n1294, n1293);
   and (n1295, n1292, n1294);
   and (n1296, n48, n55);
   not (n1297, n48);
   and (n1298, n1297, n377);
   nor (n1299, n1296, n1298);
   buf (n13, g12);
   buf (n130, n11417);
   and (n1300, n1075, n1299);
   nor (n1301, n1295, n1300);
   and (n1302, n38, n67);
   nor (n1303, n38, n67);
   nor (n1304, n1302, n1303);
   not (n1305, n1304);
   nand (n1306, n1305, n747);
   not (n1307, n1090);
   nand (n1308, n1307, n252);
   nand (n1309, n1306, n1308);
   buf (n131, n11417);
   not (n1310, n1309);
   and (n1311, n1301, n1310);
   not (n1312, n1301);
   and (n1313, n1312, n1309);
   nor (n1314, n1311, n1313);
   not (n1315, n1314);
   or (n1316, n1291, n1315);
   or (n1317, n1301, n1310);
   nand (n1318, n1316, n1317);
   not (n1319, n1318);
   buf (n132, n9564);
   or (n1320, n1282, n1319);
   or (n1321, n1318, n1281);
   nand (n1322, n1320, n1321);
   not (n1323, n1322);
   or (n1324, n1265, n1323);
   not (n1325, n1281);
   nand (n1326, n1325, n1318);
   nand (n1327, n1324, n1326);
   not (n1328, n1327);
   or (n1329, n1242, n1328);
   buf (n133, n9535);
   not (n1330, n1235);
   nand (n1331, n1330, n1240);
   nand (n1332, n1329, n1331);
   and (n1333, n857, n1126);
   and (n1334, n274, n937);
   nor (n1335, n1333, n1334);
   not (n1336, n1335);
   not (n1337, n1336);
   and (n1338, n376, n1141);
   and (n1339, n382, n947);
   buf (n134, n11298);
   nor (n1340, n1338, n1339);
   and (n1341, n1340, n1171);
   not (n1342, n1340);
   not (n1343, n1171);
   and (n1344, n1342, n1343);
   nor (n1345, n1341, n1344);
   not (n1346, n1345);
   or (n1347, n1337, n1346);
   not (n1348, n1340);
   nand (n1349, n1348, n1343);
   buf (n135, n11304);
   nand (n1350, n1347, n1349);
   xor (n1351, n1050, n1350);
   xnor (n1352, n1351, n1046);
   and (n1353, n1332, n1352);
   and (n1354, n1046, n1051);
   not (n1355, n1046);
   and (n1356, n1355, n1050);
   nor (n1357, n1354, n1356);
   and (n1358, n1357, n1350);
   nor (n1359, n1353, n1358);
   buf (n136, n9522);
   not (n1360, n1359);
   xor (n1361, n1203, n1205);
   not (n1362, n1210);
   xor (n1363, n1361, n1362);
   not (n1364, n1363);
   or (n1365, n1360, n1364);
   or (n1366, n1359, n1363);
   nand (n1367, n1365, n1366);
   not (n1368, n1367);
   or (n1369, n1234, n1368);
   buf (n137, n9498);
   not (n1370, n1359);
   nand (n1371, n1370, n1363);
   nand (n1372, n1369, n1371);
   nand (n1373, n1232, n1372);
   not (n1374, n1352);
   not (n1375, n1374);
   not (n1376, n1332);
   or (n1377, n1375, n1376);
   or (n1378, n1332, n1374);
   nand (n1379, n1377, n1378);
   buf (n138, n11433);
   not (n1380, n1379);
   not (n1381, n1153);
   not (n1382, n1144);
   or (n1383, n1381, n1382);
   or (n1384, n1144, n1153);
   nand (n1385, n1383, n1384);
   not (n1386, n1385);
   xor (n1387, n1086, n1111);
   xor (n1388, n1068, n1078);
   xnor (n1389, n1387, n1388);
   buf (n139, n11445);
   not (n1390, n1389);
   or (n1391, n1386, n1390);
   xor (n1392, n1111, n1087);
   nand (n1393, n1392, n1388);
   nand (n1394, n1391, n1393);
   not (n1395, n1394);
   not (n1396, n1395);
   and (n1397, n1345, n1336);
   not (n1398, n1345);
   and (n1399, n1398, n1335);
   buf (n14, g13);
   buf (n140, n11448);
   nor (n1400, n1397, n1399);
   not (n1401, n1400);
   not (n1402, n1401);
   and (n1403, n1396, n1402);
   not (n1404, n1400);
   not (n1405, n1395);
   or (n1406, n1404, n1405);
   or (n1407, n1395, n1400);
   nand (n1408, n1406, n1407);
   xor (n1409, n1080, n1115);
   buf (n141, n11469);
   xor (n1410, n1409, n1157);
   and (n1411, n1408, n1410);
   nor (n1412, n1403, n1411);
   xor (n1413, n1160, n1187);
   not (n1414, n1413);
   and (n1415, n1412, n1414);
   not (n1416, n1412);
   and (n1417, n1416, n1413);
   nor (n1418, n1415, n1417);
   not (n1419, n1418);
   buf (n142, n11467);
   or (n1420, n1380, n1419);
   or (n1421, n1412, n1414);
   nand (n1422, n1420, n1421);
   buf (n1423, n1367);
   and (n1424, n1423, n1233);
   not (n1425, n1423);
   not (n1426, n1233);
   and (n1427, n1425, n1426);
   nor (n1428, n1424, n1427);
   nand (n1429, n1422, n1428);
   buf (n143, n11480);
   xor (n1430, n1241, n1327);
   not (n1431, n1430);
   xor (n1432, n1410, n1408);
   not (n1433, n1432);
   not (n1434, n1433);
   or (n1435, n1431, n1434);
   not (n1436, n1430);
   nand (n1437, n1436, n1432);
   nand (n1438, n1435, n1437);
   not (n1439, n1438);
   buf (n144, n11478);
   not (n1440, n1264);
   not (n1441, n1440);
   not (n1442, n1322);
   or (n1443, n1441, n1442);
   or (n1444, n1440, n1322);
   nand (n1445, n1443, n1444);
   not (n1446, n1445);
   not (n1447, n65);
   and (n1448, n298, n1447);
   and (n1449, n38, n65);
   buf (n145, n9347);
   nor (n1450, n1448, n1449);
   and (n1451, n495, n1450);
   and (n1452, n311, n1133);
   nor (n1453, n1451, n1452);
   not (n1454, n1268);
   not (n1455, n1279);
   or (n1456, n1454, n1455);
   nand (n1457, n1456, n1280);
   xor (n1458, n1453, n1457);
   not (n1459, n1458);
   buf (n146, n9335);
   and (n1460, n48, n56);
   not (n1461, n48);
   and (n1462, n1461, n479);
   nor (n1463, n1460, n1462);
   and (n1464, n712, n1463);
   and (n1465, n1039, n1299);
   nor (n1466, n1464, n1465);
   not (n1467, n1466);
   not (n1468, n1467);
   not (n1469, n1266);
   buf (n147, n9321);
   not (n1470, n299);
   not (n1471, n51);
   nand (n1472, n1471, n50);
   not (n1473, n1472);
   not (n1474, n1473);
   or (n1475, n1470, n1474);
   not (n1476, n51);
   nor (n1477, n1476, n50);
   nand (n1478, n1477, n53);
   nand (n1479, n1475, n1478);
   buf (n148, n9307);
   buf (n1480, n1061);
   nor (n1481, n1480, n53);
   nor (n1482, n1479, n1481);
   not (n1483, n1482);
   not (n1484, n1483);
   or (n1485, n1469, n1484);
   not (n1486, n1266);
   nand (n1487, n1486, n1482);
   nand (n1488, n1485, n1487);
   not (n1489, n1488);
   buf (n149, n9293);
   or (n1490, n1468, n1489);
   not (n1491, n1266);
   nand (n1492, n1491, n1483);
   nand (n1493, n1490, n1492);
   not (n1494, n1493);
   or (n1495, n1459, n1494);
   or (n1496, n1457, n1453);
   nand (n1497, n1495, n1496);
   not (n1498, n1497);
   and (n1499, n1446, n1498);
   buf (n15, g14);
   buf (n150, n11567);
   xor (n1500, n1445, n1497);
   and (n1501, n1314, n1290);
   not (n1502, n1314);
   and (n1503, n1502, n1289);
   nor (n1504, n1501, n1503);
   not (n1505, n1504);
   and (n1506, n42, n62);
   nor (n1507, n42, n62);
   nor (n1508, n1506, n1507);
   and (n1509, n421, n1508);
   buf (n151, n11570);
   and (n1510, n513, n1257);
   nor (n1511, n1509, n1510);
   not (n1512, n1511);
   not (n1513, n1512);
   not (n1514, n1246);
   not (n1515, n815);
   or (n1516, n1514, n1515);
   and (n1517, n46, n58);
   not (n1518, n46);
   and (n1519, n1518, n769);
   buf (n152, n9225);
   nor (n1520, n1517, n1519);
   nand (n1521, n535, n1520);
   nand (n1522, n1516, n1521);
   not (n1523, n1522);
   not (n1524, n1523);
   not (n1525, n797);
   and (n1526, n44, n60);
   not (n1527, n44);
   and (n1528, n1527, n647);
   nor (n1529, n1526, n1528);
   buf (n153, n9240);
   not (n1530, n1529);
   not (n1531, n1530);
   and (n1532, n1525, n1531);
   and (n1533, n556, n1286);
   nor (n1534, n1532, n1533);
   not (n1535, n1534);
   not (n1536, n1535);
   or (n1537, n1524, n1536);
   nand (n1538, n1534, n1522);
   nand (n1539, n1537, n1538);
   buf (n154, n9204);
   not (n1540, n1539);
   or (n1541, n1513, n1540);
   not (n1542, n1523);
   nand (n1543, n1542, n1535);
   nand (n1544, n1541, n1543);
   not (n1545, n1544);
   not (n1546, n1545);
   and (n1547, n1505, n1546);
   and (n1548, n1545, n1504);
   nor (n1549, n1547, n1548);
   buf (n155, n9137);
   xor (n1550, n1249, n1253);
   xor (n1551, n1550, n1261);
   not (n1552, n1551);
   or (n1553, n1549, n1552);
   or (n1554, n1544, n1504);
   nand (n1555, n1553, n1554);
   and (n1556, n1500, n1555);
   nor (n1557, n1499, n1556);
   not (n1558, n1557);
   or (n1559, n1439, n1558);
   buf (n156, n11620);
   not (n1560, n1433);
   nand (n1561, n1560, n1430);
   nand (n1562, n1559, n1561);
   xor (n1563, n1418, n1379);
   and (n1564, n1562, n1563);
   not (n1565, n1564);
   and (n1566, n1373, n1429, n1565);
   not (n1567, n1566);
   not (n1568, n67);
   not (n1569, n295);
   buf (n157, n9174);
   or (n1570, n1568, n1569);
   and (n1571, n308, n38);
   nand (n1572, n1570, n1571);
   not (n1573, n1572);
   not (n1574, n1480);
   nand (n1575, n1574, n299);
   not (n1576, n1472);
   nand (n1577, n377, n1576);
   nand (n1578, n1477, n54);
   nand (n1579, n1575, n1577, n1578);
   buf (n158, n9155);
   nand (n1580, n1573, n1579);
   and (n1581, n274, n1250);
   not (n1582, n265);
   not (n1583, n1582);
   not (n1584, n40);
   not (n1585, n64);
   and (n1586, n1584, n1585);
   and (n1587, n40, n64);
   nor (n1588, n1586, n1587);
   and (n1589, n1583, n1588);
   buf (n159, n11664);
   nor (n1590, n1581, n1589);
   not (n1591, n1590);
   and (n1592, n1580, n1591);
   not (n1593, n1580);
   and (n1594, n1593, n1590);
   or (n1595, n1592, n1594);
   not (n1596, n1595);
   xor (n1597, n66, n38);
   and (n1598, n651, n1597);
   and (n1599, n311, n1450);
   buf (n16, g15);
   buf (n160, n11669);
   nor (n1600, n1598, n1599);
   or (n1601, n1596, n1600);
   or (n1602, n1580, n1590);
   nand (n1603, n1601, n1602);
   not (n1604, n1603);
   xnor (n1605, n1493, n1458);
   not (n1606, n1605);
   or (n1607, n1604, n1606);
   or (n1608, n1605, n1603);
   nand (n1609, n1607, n1608);
   buf (n161, n11677);
   and (n1610, n42, n63);
   not (n1611, n42);
   not (n1612, n63);
   and (n1613, n1611, n1612);
   nor (n1614, n1610, n1613);
   and (n1615, n421, n1614);
   and (n1616, n513, n1508);
   nor (n1617, n1615, n1616);
   not (n1618, n1617);
   not (n1619, n1618);
   buf (n162, n11682);
   and (n1620, n48, n57);
   not (n1621, n48);
   and (n1622, n1621, n498);
   nor (n1623, n1620, n1622);
   not (n1624, n1623);
   not (n1625, n1075);
   or (n1626, n1624, n1625);
   buf (n1627, n614);
   nand (n1628, n1627, n1463);
   nand (n1629, n1626, n1628);
   buf (n163, n11688);
   not (n1630, n1629);
   not (n1631, n1630);
   or (n1632, n1619, n1631);
   nand (n1633, n1617, n1629);
   nand (n1634, n1632, n1633);
   not (n1635, n1634);
   and (n1636, n44, n61);
   not (n1637, n44);
   and (n1638, n1637, n692);
   nor (n1639, n1636, n1638);
   buf (n164, 1'b0);
   and (n1640, n798, n1639);
   and (n1641, n556, n1529);
   nor (n1642, n1640, n1641);
   or (n1643, n1635, n1642);
   or (n1644, n1630, n1617);
   nand (n1645, n1643, n1644);
   not (n1646, n1645);
   nand (n1647, n542, n1520);
   not (n1648, n59);
   not (n1649, n46);
   buf (n165, 1'b0);
   or (n1650, n1648, n1649);
   or (n1651, n46, n59);
   nand (n1652, n1650, n1651);
   not (n1653, n1652);
   nand (n1654, n1653, n535);
   and (n1655, n1647, n1654);
   not (n1656, n1655);
   not (n1657, n1656);
   and (n1658, n40, n65);
   nor (n1659, n40, n65);
   buf (n166, 1'b0);
   nor (n1660, n1658, n1659);
   and (n1661, n1583, n1660);
   and (n1662, n274, n1588);
   nor (n1663, n1661, n1662);
   not (n1664, n1663);
   not (n1665, n1664);
   not (n1666, n1304);
   not (n1667, n376);
   or (n1668, n1666, n1667);
   nand (n1669, n310, n1597);
   buf (n167, 1'b0);
   nand (n1670, n1668, n1669);
   not (n1671, n1670);
   not (n1672, n1671);
   or (n1673, n1665, n1672);
   nand (n1674, n1670, n1663);
   nand (n1675, n1673, n1674);
   not (n1676, n1675);
   or (n1677, n1657, n1676);
   nand (n1678, n1670, n1664);
   nand (n1679, n1677, n1678);
   buf (n168, 1'b0);
   not (n1680, n1679);
   and (n1681, n1488, n1467);
   not (n1682, n1488);
   and (n1683, n1682, n1466);
   nor (n1684, n1681, n1683);
   not (n1685, n1684);
   not (n1686, n1685);
   or (n1687, n1680, n1686);
   not (n1688, n1679);
   nand (n1689, n1688, n1684);
   buf (n169, 1'b0);
   nand (n1690, n1687, n1689);
   not (n1691, n1690);
   or (n1692, n1646, n1691);
   not (n1693, n1685);
   nand (n1694, n1693, n1679);
   nand (n1695, n1692, n1694);
   nand (n1696, n1609, n1695);
   not (n1697, n1605);
   nand (n1698, n1697, n1603);
   and (n1699, n1696, n1698);
   buf (n17, g16);
   buf (n170, 1'b0);
   xnor (n1700, n1389, n1385);
   buf (n1701, n1700);
   xor (n1702, n1699, n1701);
   xor (n1703, n1555, n1500);
   and (n1704, n1702, n1703);
   and (n1705, n1699, n1701);
   nor (n1706, n1704, n1705);
   not (n1707, n1706);
   not (n1708, n1438);
   and (n1709, n1557, n1708);
   buf (n171, n11419);
   not (n1710, n1557);
   and (n1711, n1710, n1438);
   nor (n1712, n1709, n1711);
   not (n1713, n1712);
   not (n1714, n1713);
   or (n1715, n1707, n1714);
   not (n1716, n1706);
   not (n1717, n1716);
   not (n1718, n1713);
   or (n1719, n1717, n1718);
   buf (n172, n11416);
   nand (n1720, n1712, n1706);
   nand (n1721, n1719, n1720);
   not (n1722, n797);
   and (n1723, n44, n63);
   not (n1724, n44);
   and (n1725, n1724, n1612);
   nor (n1726, n1723, n1725);
   not (n1727, n1726);
   not (n1728, n1727);
   and (n1729, n1722, n1728);
   buf (n173, n11416);
   xor (n1730, n44, n62);
   and (n1731, n1730, n556);
   nor (n1732, n1729, n1731);
   not (n1733, n1732);
   not (n1734, n429);
   not (n1735, n42);
   not (n1736, n64);
   and (n1737, n1735, n1736);
   and (n1738, n42, n64);
   nor (n1739, n1737, n1738);
   buf (n174, n11416);
   not (n1740, n1739);
   not (n1741, n1740);
   and (n1742, n1734, n1741);
   not (n1743, n415);
   not (n1744, n412);
   or (n1745, n1743, n1744);
   nand (n1746, n1745, n419);
   not (n1747, n42);
   not (n1748, n65);
   and (n1749, n1747, n1748);
   buf (n175, n11416);
   and (n1750, n42, n65);
   nor (n1751, n1749, n1750);
   and (n1752, n1746, n1751);
   nor (n1753, n1742, n1752);
   not (n1754, n1753);
   not (n1755, n1754);
   nand (n1756, n1473, n498);
   nand (n1757, n1270, n479);
   nand (n1758, n1477, n56);
   nand (n1759, n1756, n1757, n1758);
   buf (n176, n11416);
   not (n1760, n1759);
   not (n1761, n1760);
   or (n1762, n1755, n1761);
   nand (n1763, n1759, n1753);
   nand (n1764, n1762, n1763);
   not (n1765, n1764);
   or (n1766, n1733, n1765);
   or (n1767, n1764, n1732);
   nand (n1768, n1766, n1767);
   not (n1769, n1768);
   buf (n177, n11416);
   not (n1770, n1769);
   nand (n1771, n273, n67);
   not (n1772, n1771);
   and (n1773, n48, n60);
   not (n1774, n48);
   and (n1775, n1774, n647);
   nor (n1776, n1773, n1775);
   not (n1777, n1776);
   not (n1778, n1074);
   not (n1779, n1778);
   buf (n178, n11416);
   not (n1780, n1779);
   or (n1781, n1777, n1780);
   and (n1782, n48, n59);
   not (n1783, n48);
   and (n1784, n1783, n578);
   nor (n1785, n1782, n1784);
   nand (n1786, n614, n1785);
   nand (n1787, n1781, n1786);
   not (n1788, n1787);
   not (n1789, n1788);
   buf (n179, n11416);
   or (n1790, n1772, n1789);
   not (n1791, n1771);
   not (n1792, n1791);
   not (n1793, n1787);
   or (n1794, n1792, n1793);
   not (n1795, n797);
   not (n1796, n44);
   not (n1797, n64);
   and (n1798, n1796, n1797);
   and (n1799, n44, n64);
   buf (n18, g17);
   buf (n180, n11416);
   nor (n1800, n1798, n1799);
   not (n1801, n1800);
   not (n1802, n1801);
   and (n1803, n1795, n1802);
   and (n1804, n556, n1726);
   nor (n1805, n1803, n1804);
   nand (n1806, n1794, n1805);
   nand (n1807, n1790, n1806);
   not (n1808, n1807);
   not (n1809, n534);
   buf (n181, n11416);
   and (n1810, n46, n62);
   not (n1811, n46);
   not (n1812, n62);
   and (n1813, n1811, n1812);
   nor (n1814, n1810, n1813);
   not (n1815, n1814);
   not (n1816, n1815);
   and (n1817, n1809, n1816);
   and (n1818, n46, n61);
   not (n1819, n46);
   buf (n182, n11416);
   and (n1820, n1819, n692);
   nor (n1821, n1818, n1820);
   and (n1822, n815, n1821);
   nor (n1823, n1817, n1822);
   not (n1824, n1823);
   not (n1825, n1824);
   not (n1826, n1472);
   nand (n1827, n1826, n769);
   nand (n1828, n50, n51);
   not (n1829, n1828);
   buf (n183, n11416);
   nand (n1830, n1829, n498);
   not (n1831, n51);
   nor (n1832, n1831, n50);
   nand (n1833, n57, n1832);
   nand (n1834, n1827, n1830, n1833);
   not (n1835, n1834);
   not (n1836, n512);
   not (n1837, n1751);
   not (n1838, n1837);
   and (n1839, n1836, n1838);
   buf (n184, n11416);
   and (n1840, n42, n66);
   not (n1841, n42);
   not (n1842, n66);
   and (n1843, n1841, n1842);
   nor (n1844, n1840, n1843);
   and (n1845, n1746, n1844);
   nor (n1846, n1839, n1845);
   not (n1847, n1846);
   or (n1848, n1835, n1847);
   or (n1849, n1834, n1846);
   buf (n185, n11416);
   nand (n1850, n1848, n1849);
   not (n1851, n1850);
   or (n1852, n1825, n1851);
   not (n1853, n1846);
   nand (n1854, n1853, n1834);
   nand (n1855, n1852, n1854);
   not (n1856, n1855);
   or (n1857, n1808, n1856);
   or (n1858, n1855, n1807);
   nand (n1859, n1857, n1858);
   buf (n186, n11416);
   not (n1860, n1859);
   or (n1861, n1770, n1860);
   not (n1862, n1855);
   nand (n1863, n1862, n1807);
   nand (n1864, n1861, n1863);
   not (n1865, n1864);
   not (n1866, n543);
   not (n1867, n1652);
   and (n1868, n1866, n1867);
   and (n1869, n46, n60);
   buf (n187, n11416);
   not (n1870, n46);
   and (n1871, n1870, n647);
   nor (n1872, n1869, n1871);
   and (n1873, n913, n1872);
   nor (n1874, n1868, n1873);
   not (n1875, n1874);
   not (n1876, n1785);
   not (n1877, n711);
   or (n1878, n1876, n1877);
   and (n1879, n48, n58);
   buf (n188, n11416);
   not (n1880, n48);
   and (n1881, n1880, n769);
   nor (n1882, n1879, n1881);
   nand (n1883, n1627, n1882);
   nand (n1884, n1878, n1883);
   not (n1885, n67);
   not (n1886, n1885);
   not (n1887, n260);
   and (n1888, n1886, n1887);
   nor (n1889, n1888, n337);
   buf (n189, n11416);
   nand (n1890, n1884, n1889);
   not (n1891, n1890);
   not (n1892, n1891);
   or (n1893, n1875, n1892);
   or (n1894, n1891, n1874);
   nand (n1895, n1893, n1894);
   not (n1896, n1759);
   not (n1897, n1754);
   or (n1898, n1896, n1897);
   not (n1899, n1732);
   buf (n19, g18);
   buf (n190, n11416);
   nand (n1900, n1899, n1764);
   nand (n1901, n1898, n1900);
   xor (n1902, n1895, n1901);
   xor (n1903, n1865, n1902);
   not (n1904, n1903);
   not (n1905, n1821);
   not (n1906, n1905);
   not (n1907, n534);
   and (n1908, n1906, n1907);
   and (n1909, n541, n1872);
   buf (n191, n11416);
   nor (n1910, n1908, n1909);
   xor (n1911, n66, n40);
   not (n1912, n1911);
   not (n1913, n274);
   or (n1914, n1912, n1913);
   and (n1915, n1885, n335);
   and (n1916, n41, n67);
   nor (n1917, n1915, n1916);
   or (n1918, n1582, n1917);
   nand (n1919, n1914, n1918);
   buf (n192, n11416);
   not (n1920, n1919);
   and (n1921, n1910, n1920);
   not (n1922, n1910);
   and (n1923, n1922, n1919);
   nor (n1924, n1921, n1923);
   not (n1925, n1924);
   not (n1926, n1890);
   nor (n1927, n1884, n1889);
   nor (n1928, n1926, n1927);
   not (n1929, n1928);
   buf (n193, n11416);
   or (n1930, n1925, n1929);
   not (n1931, n1910);
   nand (n1932, n1931, n1919);
   nand (n1933, n1930, n1932);
   and (n1934, n556, n1639);
   and (n1935, n565, n1730);
   nor (n1936, n1934, n1935);
   nand (n1937, n310, n67);
   nor (n1938, n1936, n1937);
   not (n1939, n1938);
   buf (n194, n11416);
   nand (n1940, n1936, n1937);
   nand (n1941, n1939, n1940);
   not (n1942, n1941);
   and (n1943, n1075, n1882);
   not (n1944, n1038);
   and (n1945, n1944, n1623);
   nor (n1946, n1943, n1945);
   not (n1947, n1946);
   and (n1948, n1942, n1947);
   and (n1949, n1941, n1946);
   buf (n195, n11416);
   nor (n1950, n1948, n1949);
   xor (n1951, n1933, n1950);
   and (n1952, n465, n1911);
   and (n1953, n274, n1660);
   nor (n1954, n1952, n1953);
   nand (n1955, n1574, n377);
   buf (n1956, n1576);
   nand (n1957, n1956, n479);
   nand (n1958, n1477, n55);
   nand (n1959, n1955, n1957, n1958);
   buf (n196, n11416);
   and (n1960, n867, n1739);
   and (n1961, n1259, n1614);
   nor (n1962, n1960, n1961);
   xor (n1963, n1959, n1962);
   xor (n1964, n1954, n1963);
   xor (n1965, n1951, n1964);
   not (n1966, n1965);
   and (n1967, n1904, n1966);
   and (n1968, n1903, n1965);
   nor (n1969, n1967, n1968);
   buf (n197, n11416);
   not (n1970, n1969);
   not (n1971, n1970);
   xor (n1972, n1771, n1787);
   xor (n1973, n1972, n1805);
   not (n1974, n1973);
   not (n1975, n1974);
   and (n1976, n48, n61);
   not (n1977, n48);
   and (n1978, n1977, n692);
   nor (n1979, n1976, n1978);
   buf (n198, n11415);
   not (n1980, n1979);
   not (n1981, n1075);
   or (n1982, n1980, n1981);
   nand (n1983, n614, n1776);
   nand (n1984, n1982, n1983);
   nand (n1985, n428, n67);
   and (n1986, n1985, n352);
   nand (n1987, n1984, n1986);
   buf (n1988, n1987);
   not (n1989, n1988);
   buf (n199, n11383);
   and (n1990, n1975, n1989);
   and (n1991, n1259, n1844);
   and (n1992, n421, n1885);
   nor (n1993, n1991, n1992);
   not (n1994, n1993);
   not (n1995, n1994);
   nand (n1996, n1473, n578);
   nand (n1997, n1270, n769);
   nand (n1998, n1477, n58);
   nand (n1999, n1996, n1997, n1998);
   buf (n2, g1);
   buf (n20, g19);
   buf (n200, n11388);
   not (n2000, n1999);
   not (n2001, n2000);
   and (n2002, n44, n65);
   not (n2003, n44);
   and (n2004, n2003, n1447);
   nor (n2005, n2002, n2004);
   and (n2006, n566, n2005);
   and (n2007, n556, n1800);
   nor (n2008, n2006, n2007);
   not (n2009, n2008);
   buf (n201, n11286);
   not (n2010, n2009);
   or (n2011, n2001, n2010);
   nand (n2012, n2008, n1999);
   nand (n2013, n2011, n2012);
   not (n2014, n2013);
   or (n2015, n1995, n2014);
   or (n2016, n2008, n2000);
   nand (n2017, n2015, n2016);
   not (n2018, n1988);
   not (n2019, n2018);
   buf (n202, n11296);
   not (n2020, n1974);
   or (n2021, n2019, n2020);
   nand (n2022, n1973, n1988);
   nand (n2023, n2021, n2022);
   and (n2024, n2017, n2023);
   nor (n2025, n1990, n2024);
   not (n2026, n2025);
   xor (n2027, n1924, n1928);
   not (n2028, n2027);
   not (n2029, n1771);
   buf (n203, n11314);
   not (n2030, n1788);
   or (n2031, n2029, n2030);
   nand (n2032, n2031, n1806);
   xor (n2033, n2032, n1855);
   xnor (n2034, n2033, n1768);
   not (n2035, n2034);
   not (n2036, n2035);
   or (n2037, n2028, n2036);
   not (n2038, n2027);
   nand (n2039, n2038, n2034);
   buf (n204, n11323);
   nand (n2040, n2037, n2039);
   not (n2041, n2040);
   or (n2042, n2026, n2041);
   not (n2043, n2027);
   nand (n2044, n2043, n2035);
   nand (n2045, n2042, n2044);
   not (n2046, n2045);
   not (n2047, n2046);
   or (n2048, n1971, n2047);
   nand (n2049, n2045, n1969);
   buf (n205, n11692);
   nand (n2050, n2048, n2049);
   and (n2051, n2023, n2017);
   not (n2052, n2023);
   not (n2053, n2017);
   and (n2054, n2052, n2053);
   nor (n2055, n2051, n2054);
   not (n2056, n1814);
   not (n2057, n815);
   or (n2058, n2056, n2057);
   and (n2059, n504, n1612);
   buf (n206, n11431);
   and (n2060, n46, n63);
   nor (n2061, n2059, n2060);
   nand (n2062, n913, n2061);
   nand (n2063, n2058, n2062);
   not (n2064, n1987);
   nor (n2065, n1984, n1986);
   nor (n2066, n2064, n2065);
   xor (n2067, n2063, n2066);
   not (n2068, n1985);
   not (n2069, n2068);
   buf (n207, n11443);
   nand (n2070, n1576, n647);
   nand (n2071, n59, n1832);
   nand (n2072, n1270, n578);
   and (n2073, n2070, n2071, n2072);
   not (n2074, n2073);
   not (n2075, n2074);
   or (n2076, n2069, n2075);
   and (n2077, n44, n66);
   not (n2078, n44);
   and (n2079, n2078, n1842);
   buf (n208, n11455);
   nor (n2080, n2077, n2079);
   and (n2081, n2080, n566);
   and (n2082, n556, n2005);
   nor (n2083, n2081, n2082);
   not (n2084, n2083);
   and (n2085, n2073, n1985);
   not (n2086, n2073);
   and (n2087, n2086, n2068);
   nor (n2088, n2085, n2087);
   nand (n2089, n2084, n2088);
   buf (n209, n11461);
   nand (n2090, n2076, n2089);
   and (n2091, n2067, n2090);
   and (n2092, n2063, n2066);
   or (n2093, n2091, n2092);
   and (n2094, n1850, n1824);
   not (n2095, n1850);
   and (n2096, n2095, n1823);
   nor (n2097, n2094, n2096);
   and (n2098, n2093, n2097);
   not (n2099, n2093);
   buf (n21, g20);
   buf (n210, n11474);
   not (n2100, n2097);
   and (n2101, n2099, n2100);
   nor (n2102, n2098, n2101);
   and (n2103, n2055, n2102);
   and (n2104, n2093, n2097);
   nor (n2105, n2103, n2104);
   not (n2106, n2105);
   and (n2107, n2040, n2025);
   not (n2108, n2040);
   not (n2109, n2025);
   buf (n211, n11502);
   and (n2110, n2108, n2109);
   nor (n2111, n2107, n2110);
   not (n2112, n2111);
   not (n2113, n2112);
   or (n2114, n2106, n2113);
   not (n2115, n2105);
   nand (n2116, n2115, n2111);
   nand (n2117, n2114, n2116);
   not (n2118, n2117);
   xor (n2119, n2055, n2102);
   buf (n212, n11509);
   not (n2120, n2119);
   and (n2121, n2013, n1993);
   not (n2122, n2013);
   and (n2123, n2122, n1994);
   nor (n2124, n2121, n2123);
   not (n2125, n2124);
   not (n2126, n2125);
   xor (n2127, n46, n64);
   and (n2128, n913, n2127);
   and (n2129, n815, n2061);
   buf (n213, n11516);
   nor (n2130, n2128, n2129);
   not (n2131, n2130);
   and (n2132, n48, n62);
   not (n2133, n48);
   and (n2134, n2133, n1812);
   nor (n2135, n2132, n2134);
   not (n2136, n2135);
   not (n2137, n1075);
   or (n2138, n2136, n2137);
   nand (n2139, n1627, n1979);
   buf (n214, n11525);
   nand (n2140, n2138, n2139);
   not (n2141, n801);
   not (n2142, n1885);
   or (n2143, n2141, n2142);
   not (n2144, n803);
   nand (n2145, n2143, n2144);
   nand (n2146, n2145, n44);
   not (n2147, n2146);
   nand (n2148, n1576, n692);
   nand (n2149, n1832, n60);
   buf (n215, n11533);
   nand (n2150, n1270, n647);
   nand (n2151, n2148, n2149, n2150);
   nand (n2152, n2147, n2151);
   nor (n2153, n2140, n2152);
   not (n2154, n2153);
   nand (n2155, n2140, n2152);
   nand (n2156, n2154, n2155);
   nand (n2157, n2131, n2156);
   not (n2158, n2152);
   nand (n2159, n2158, n2140);
   buf (n216, n11541);
   nand (n2160, n2157, n2159);
   not (n2161, n2160);
   not (n2162, n2161);
   or (n2163, n2126, n2162);
   nand (n2164, n2160, n2124);
   nand (n2165, n2163, n2164);
   xor (n2166, n2063, n2066);
   xor (n2167, n2166, n2090);
   and (n2168, n2165, n2167);
   and (n2169, n2160, n2125);
   buf (n217, n11554);
   nor (n2170, n2168, n2169);
   not (n2171, n2170);
   and (n2172, n2120, n2171);
   and (n2173, n2119, n2170);
   nor (n2174, n2172, n2173);
   not (n2175, n2170);
   nand (n2176, n2175, n2119);
   nand (n2177, n2174, n2176);
   not (n2178, n2177);
   or (n2179, n2118, n2178);
   buf (n218, n11564);
   not (n2180, n2105);
   nand (n2181, n2180, n2112);
   nand (n2182, n2179, n2181);
   nand (n2183, n2050, n2182);
   not (n2184, n1903);
   not (n2185, n1965);
   not (n2186, n2185);
   or (n2187, n2184, n2186);
   or (n2188, n1865, n1902);
   nand (n2189, n2187, n2188);
   buf (n219, n11574);
   not (n2190, n2189);
   not (n2191, n1655);
   not (n2192, n1675);
   or (n2193, n2191, n2192);
   or (n2194, n1675, n1655);
   nand (n2195, n2193, n2194);
   not (n2196, n2195);
   xnor (n2197, n1642, n1634);
   not (n2198, n2197);
   not (n2199, n2198);
   buf (n22, g21);
   buf (n220, n11589);
   or (n2200, n2196, n2199);
   not (n2201, n2195);
   nand (n2202, n2201, n2197);
   nand (n2203, n2200, n2202);
   not (n2204, n1901);
   not (n2205, n1895);
   or (n2206, n2204, n2205);
   not (n2207, n1874);
   nand (n2208, n2207, n1891);
   nand (n2209, n2206, n2208);
   buf (n221, n11582);
   xor (n2210, n2203, n2209);
   not (n2211, n2210);
   and (n2212, n1951, n1964);
   and (n2213, n1933, n1950);
   nor (n2214, n2212, n2213);
   or (n2215, n1963, n1954);
   and (n2216, n1955, n1957, n1958);
   or (n2217, n2216, n1962);
   nand (n2218, n2215, n2217);
   not (n2219, n1572);
   buf (n222, n11596);
   not (n2220, n1579);
   not (n2221, n2220);
   or (n2222, n2219, n2221);
   nand (n2223, n2222, n1580);
   not (n2224, n2223);
   not (n2225, n1938);
   nand (n2226, n2225, n1946);
   nand (n2227, n2226, n1940);
   not (n2228, n2227);
   not (n2229, n2228);
   buf (n223, n11612);
   or (n2230, n2224, n2229);
   not (n2231, n2223);
   nand (n2232, n2231, n2227);
   nand (n2233, n2230, n2232);
   xor (n2234, n2218, n2233);
   xor (n2235, n2214, n2234);
   not (n2236, n2235);
   or (n2237, n2211, n2236);
   or (n2238, n2235, n2210);
   nand (n2239, n2237, n2238);
   buf (n224, n11617);
   nand (n2240, n2190, n2239);
   not (n2241, n1970);
   nand (n2242, n2241, n2046);
   nand (n2243, n2183, n2240, n2242);
   not (n2244, n805);
   not (n2245, n2080);
   not (n2246, n2245);
   and (n2247, n2244, n2246);
   and (n2248, n46, n67);
   not (n2249, n46);
   buf (n225, n11633);
   and (n2250, n2249, n1885);
   nor (n2251, n2248, n2250);
   and (n2252, n566, n2251);
   nor (n2253, n2247, n2252);
   not (n2254, n2253);
   not (n2255, n2254);
   and (n2256, n48, n63);
   not (n2257, n48);
   and (n2258, n2257, n1612);
   nor (n2259, n2256, n2258);
   buf (n226, n11648);
   and (n2260, n1075, n2259);
   and (n2261, n1627, n2135);
   nor (n2262, n2260, n2261);
   not (n2263, n46);
   not (n2264, n65);
   and (n2265, n2263, n2264);
   and (n2266, n46, n65);
   nor (n2267, n2265, n2266);
   and (n2268, n535, n2267);
   and (n2269, n541, n2127);
   buf (n227, n11653);
   nor (n2270, n2268, n2269);
   xor (n2271, n2262, n2270);
   not (n2272, n2271);
   or (n2273, n2255, n2272);
   or (n2274, n2262, n2270);
   nand (n2275, n2273, n2274);
   not (n2276, n2275);
   xnor (n2277, n2083, n2088);
   not (n2278, n2277);
   and (n2279, n2276, n2278);
   not (n2280, n2276);
   and (n2281, n2280, n2277);
   nor (n2282, n2279, n2281);
   not (n2283, n2282);
   not (n2284, n2130);
   not (n2285, n2156);
   or (n2286, n2284, n2285);
   or (n2287, n2156, n2130);
   nand (n2288, n2286, n2287);
   or (n2289, n2283, n2288);
   or (n2290, n2275, n2277);
   nand (n2291, n2289, n2290);
   not (n2292, n2291);
   and (n2293, n2165, n2167);
   not (n2294, n2165);
   not (n2295, n2167);
   and (n2296, n2294, n2295);
   nor (n2297, n2293, n2296);
   nand (n2298, n2292, n2297);
   and (n2299, n2181, n2176, n2298);
   buf (n23, g22);
   not (n2300, n2288);
   not (n2301, n2282);
   or (n2302, n2300, n2301);
   or (n2303, n2288, n2282);
   nand (n2304, n2302, n2303);
   not (n2305, n2304);
   not (n2306, n2146);
   not (n2307, n2151);
   not (n2308, n2307);
   or (n2309, n2306, n2308);
   nand (n2310, n2309, n2152);
   not (n2311, n2310);
   not (n2312, n2311);
   nand (n2313, n556, n67);
   not (n2314, n2313);
   nand (n2315, n1576, n1812);
   nand (n2316, n1832, n61);
   nand (n2317, n1829, n692);
   nand (n2318, n2315, n2316, n2317);
   not (n2319, n2318);
   not (n2320, n2319);
   or (n2321, n2314, n2320);
   nand (n2322, n2318, n556, n67);
   nand (n2323, n2321, n2322);
   and (n2324, n48, n64);
   not (n2325, n48);
   and (n2326, n2325, n1131);
   nor (n2327, n2324, n2326);
   and (n2328, n1075, n2327);
   and (n2329, n1627, n2259);
   nor (n2330, n2328, n2329);
   or (n2331, n2323, n2330);
   buf (n2332, n2322);
   nand (n2333, n2331, n2332);
   not (n2334, n2333);
   and (n2335, n2312, n2334);
   xor (n2336, n2333, n2310);
   not (n2337, n2336);
   not (n2338, n2271);
   not (n2339, n2253);
   and (n2340, n2338, n2339);
   and (n2341, n2271, n2253);
   nor (n2342, n2340, n2341);
   and (n2343, n2337, n2342);
   nor (n2344, n2335, n2343);
   nand (n2345, n2305, n2344);
   not (n2346, n2345);
   xnor (n2347, n2344, n2304);
   not (n2348, n2342);
   not (n2349, n2336);
   or (n2350, n2348, n2349);
   or (n2351, n2342, n2336);
   nand (n2352, n2350, n2351);
   not (n2353, n2352);
   not (n2354, n2353);
   not (n2355, n627);
   not (n2356, n2267);
   not (n2357, n2356);
   and (n2358, n2355, n2357);
   and (n2359, n46, n66);
   not (n2360, n46);
   and (n2361, n2360, n1842);
   nor (n2362, n2359, n2361);
   and (n2363, n535, n2362);
   nor (n2364, n2358, n2363);
   not (n2365, n2364);
   not (n2366, n2365);
   nand (n2367, n541, n67);
   nand (n2368, n47, n48);
   and (n2369, n2368, n46);
   not (n237, n2);
   nand (n2370, n2367, n2369);
   not (n2371, n2370);
   nand (n2372, n1473, n1612);
   nand (n2373, n1477, n62);
   nand (n2374, n1829, n1812);
   nand (n2375, n2372, n2373, n2374);
   nand (n2376, n2371, n2375);
   not (n2377, n2376);
   not (n2378, n2377);
   or (n2379, n2366, n2378);
   not (n238, n237);
   nand (n2380, n2376, n2364);
   nand (n2381, n2379, n2380);
   not (n2382, n2381);
   not (n2383, n2330);
   and (n2384, n2323, n2383);
   not (n2385, n2323);
   and (n2386, n2385, n2330);
   nor (n2387, n2384, n2386);
   or (n2388, n2382, n2387);
   or (n2389, n2377, n2364);
   not (n239, n37);
   nand (n2390, n2388, n2389);
   not (n2391, n2390);
   and (n2392, n2354, n2391);
   not (n2393, n2367);
   not (n2394, n1828);
   not (n2395, n1612);
   and (n2396, n2394, n2395);
   not (n2397, n1273);
   not (n2398, n50);
   nand (n2399, n2398, n1612);
   buf (n24, g23);
   not (n240, n38);
   not (n2400, n51);
   nand (n2401, n2400, n64);
   nand (n2402, n2397, n2399, n2401);
   nor (n2403, n2396, n2402);
   not (n2404, n2403);
   or (n2405, n2393, n2404);
   or (n2406, n2367, n2403);
   nand (n2407, n2405, n2406);
   not (n2408, n2407);
   and (n2409, n48, n66);
   nand (n241, n239, n240);
   not (n2410, n48);
   and (n2411, n2410, n1842);
   nor (n2412, n2409, n2411);
   and (n2413, n1779, n2412);
   and (n2414, n48, n65);
   not (n2415, n48);
   and (n2416, n2415, n1447);
   nor (n2417, n2414, n2416);
   and (n2418, n614, n2417);
   nor (n2419, n2413, n2418);
   nand (n242, n37, n38);
   or (n2420, n2408, n2419);
   not (n2421, n2403);
   or (n2422, n2367, n2421);
   nand (n2423, n2420, n2422);
   not (n2424, n2417);
   not (n2425, n1779);
   or (n2426, n2424, n2425);
   nand (n2427, n614, n2327);
   nand (n2428, n2426, n2427);
   not (n2429, n541);
   nand (n243, n241, n242);
   not (n2430, n2362);
   or (n2431, n2429, n2430);
   nand (n2432, n535, n2251);
   nand (n2433, n2431, n2432);
   xor (n2434, n2428, n2433);
   not (n2435, n2370);
   nor (n2436, n2435, n2375);
   not (n2437, n2436);
   nand (n2438, n2437, n2376);
   xnor (n2439, n2434, n2438);
   xor (n244, n36, n37);
   xor (n2440, n2423, n2439);
   not (n2441, n67);
   nand (n2442, n610, n1005);
   not (n2443, n2442);
   or (n2444, n2441, n2443);
   nand (n2445, n2444, n616);
   not (n2446, n1480);
   not (n2447, n64);
   and (n2448, n2446, n2447);
   not (n2449, n1447);
   nand (n245, n243, n244);
   not (n2450, n1576);
   or (n2451, n2449, n2450);
   nand (n2452, n1832, n64);
   nand (n2453, n2451, n2452);
   nor (n2454, n2448, n2453);
   nor (n2455, n2445, n2454);
   not (n2456, n2455);
   nand (n2457, n2445, n2454);
   nand (n2458, n2456, n2457);
   not (n2459, n1885);
   not (n246, n245);
   not (n2460, n711);
   or (n2461, n2459, n2460);
   nand (n2462, n614, n2412);
   nand (n2463, n2461, n2462);
   nand (n2464, n51, n65);
   nand (n2465, n1842, n2464);
   and (n2466, n1038, n2465);
   not (n2467, n2464);
   or (n2468, n2467, n50);
   nand (n2469, n50, n66);
   not (n247, n246);
   nor (n2470, n2464, n2469);
   nor (n2471, n2470, n1885);
   nand (n2472, n2468, n2471);
   nor (n2473, n2466, n2472);
   nand (n2474, n2463, n2473);
   and (n2475, n2458, n2474);
   nor (n2476, n2463, n2473);
   nor (n2477, n2475, n2476);
   not (n2478, n2477);
   not (n2479, n2455);
   or (n248, n36, n55);
   not (n2480, n2479);
   not (n2481, n2419);
   not (n2482, n2481);
   not (n2483, n2408);
   or (n2484, n2482, n2483);
   nand (n2485, n2407, n2419);
   nand (n2486, n2484, n2485);
   not (n2487, n2486);
   or (n2488, n2480, n2487);
   or (n2489, n2486, n2479);
   nand (n249, n36, n55);
   nand (n2490, n2488, n2489);
   not (n2491, n2490);
   or (n2492, n2478, n2491);
   not (n2493, n2479);
   nand (n2494, n2493, n2486);
   nand (n2495, n2492, n2494);
   and (n2496, n2440, n2495);
   and (n2497, n2423, n2439);
   or (n2498, n2496, n2497);
   not (n2499, n2428);
   buf (n25, g24);
   nand (n250, n248, n249);
   not (n2500, n2433);
   or (n2501, n2499, n2500);
   not (n2502, n2438);
   nand (n2503, n2502, n2434);
   nand (n2504, n2501, n2503);
   not (n2505, n2504);
   not (n2506, n2505);
   not (n2507, n2381);
   not (n2508, n2387);
   and (n2509, n2507, n2508);
   or (n251, n247, n250);
   and (n2510, n2381, n2387);
   nor (n2511, n2509, n2510);
   not (n2512, n2511);
   or (n2513, n2506, n2512);
   or (n2514, n2511, n2505);
   nand (n2515, n2513, n2514);
   nand (n2516, n2498, n2515);
   and (n2517, n2353, n2390);
   nand (n2518, n2511, n2504);
   not (n2519, n2518);
   not (n252, n243);
   nor (n2520, n2517, n2519);
   and (n2521, n2516, n2520);
   nor (n2522, n2392, n2521);
   nand (n2523, n2347, n2522);
   not (n2524, n2523);
   or (n2525, n2346, n2524);
   xnor (n2526, n2291, n2297);
   nand (n2527, n2525, n2526);
   nand (n2528, n2299, n2527, n2240, n2242);
   not (n2529, n2218);
   not (n253, n252);
   not (n2530, n2233);
   or (n2531, n2529, n2530);
   not (n2532, n2223);
   nand (n2533, n2532, n2228);
   nand (n2534, n2531, n2533);
   not (n2535, n2534);
   not (n2536, n1600);
   not (n2537, n1595);
   or (n2538, n2536, n2537);
   or (n2539, n1595, n1600);
   or (n254, n36, n54);
   nand (n2540, n2538, n2539);
   not (n2541, n2540);
   and (n2542, n1539, n1512);
   not (n2543, n1539);
   and (n2544, n2543, n1511);
   or (n2545, n2542, n2544);
   not (n2546, n2545);
   and (n2547, n2541, n2546);
   and (n2548, n2540, n2545);
   nor (n2549, n2547, n2548);
   nand (n255, n36, n54);
   not (n2550, n2549);
   or (n2551, n2535, n2550);
   or (n2552, n2534, n2549);
   nand (n2553, n2551, n2552);
   and (n2554, n1690, n1645);
   not (n2555, n1690);
   not (n2556, n1645);
   and (n2557, n2555, n2556);
   or (n2558, n2554, n2557);
   not (n2559, n2558);
   nand (n256, n254, n255);
   not (n2560, n2209);
   not (n2561, n2203);
   or (n2562, n2560, n2561);
   not (n2563, n2198);
   nand (n2564, n2563, n2195);
   nand (n2565, n2562, n2564);
   not (n2566, n2565);
   or (n2567, n2559, n2566);
   or (n2568, n2558, n2565);
   nand (n2569, n2567, n2568);
   or (n257, n253, n256);
   xor (n2570, n2553, n2569);
   not (n2571, n2234);
   not (n2572, n2571);
   not (n2573, n2214);
   and (n2574, n2572, n2573);
   not (n2575, n2235);
   and (n2576, n2575, n2210);
   nor (n2577, n2574, n2576);
   xor (n2578, n2570, n2577);
   not (n2579, n2239);
   nand (n258, n251, n257);
   and (n2580, n2189, n2579);
   nor (n2581, n2578, n2580);
   nand (n2582, n2243, n2528, n2581);
   xor (n2583, n1609, n1695);
   not (n2584, n2583);
   xor (n2585, n1552, n1549);
   not (n2586, n2585);
   not (n2587, n2549);
   not (n2588, n2587);
   not (n2589, n2534);
   not (n259, n40);
   or (n2590, n2588, n2589);
   not (n2591, n2545);
   nand (n2592, n2591, n2540);
   nand (n2593, n2590, n2592);
   not (n2594, n2593);
   and (n2595, n2586, n2594);
   and (n2596, n2593, n2585);
   nor (n2597, n2595, n2596);
   not (n2598, n2597);
   not (n2599, n2598);
   buf (n26, g25);
   nor (n260, n41, n42);
   or (n2600, n2584, n2599);
   not (n2601, n2585);
   nand (n2602, n2601, n2593);
   nand (n2603, n2600, n2602);
   not (n2604, n1703);
   and (n2605, n1702, n2604);
   not (n2606, n1702);
   and (n2607, n2606, n1703);
   nor (n2608, n2605, n2607);
   and (n2609, n2603, n2608);
   not (n261, n260);
   not (n2610, n2577);
   nand (n2611, n2610, n2570);
   not (n2612, n2558);
   not (n2613, n2565);
   not (n2614, n2613);
   and (n2615, n2612, n2614);
   and (n2616, n2569, n2553);
   nor (n2617, n2615, n2616);
   not (n2618, n2617);
   xnor (n2619, n2597, n2583);
   or (n262, n259, n261);
   nand (n2620, n2618, n2619);
   nand (n2621, n2611, n2620);
   nor (n2622, n2609, n2621);
   nand (n2623, n2582, n2622);
   not (n2624, n2620);
   not (n2625, n2619);
   not (n2626, n2617);
   and (n2627, n2625, n2626);
   and (n2628, n2619, n2617);
   nor (n2629, n2627, n2628);
   not (n263, n40);
   not (n2630, n2629);
   or (n2631, n2624, n2630);
   xor (n2632, n2603, n2608);
   nand (n2633, n2631, n2632);
   not (n2634, n2609);
   nand (n2635, n2633, n2634);
   nand (n2636, n1721, n2623, n2635);
   nand (n2637, n1715, n2636);
   not (n2638, n2637);
   not (n2639, n2638);
   nand (n264, n263, n41, n42);
   or (n2640, n1567, n2639);
   and (n2641, n1373, n1429);
   xor (n2642, n1562, n1563);
   or (n2643, n2642, n1564);
   xor (n2644, n1422, n1428);
   nand (n2645, n2643, n2644);
   and (n2646, n2641, n2645);
   not (n2647, n1373);
   xnor (n2648, n1232, n1372);
   not (n2649, n2648);
   nand (n265, n262, n264);
   or (n2650, n2647, n2649);
   xor (n2651, n1229, n985);
   nand (n2652, n2650, n2651);
   nor (n2653, n2646, n2652);
   nand (n2654, n2640, n2653);
   nand (n2655, n1231, n2654);
   xor (n2656, n892, n978);
   nand (n2657, n2655, n2656);
   nand (n2658, n980, n2657);
   xor (n2659, n766, n849);
   not (n266, n265);
   and (n2660, n2659, n891);
   and (n2661, n766, n849);
   nor (n2662, n2660, n2661);
   not (n2663, n2662);
   and (n2664, n876, n890);
   and (n2665, n855, n875);
   nor (n2666, n2664, n2665);
   xnor (n2667, n472, n462);
   not (n2668, n807);
   not (n2669, n791);
   not (n267, n52);
   or (n2670, n2668, n2669);
   nand (n2671, n776, n786);
   nand (n2672, n2670, n2671);
   and (n2673, n2672, n870);
   not (n2674, n2672);
   and (n2675, n2674, n871);
   or (n2676, n2673, n2675);
   xnor (n2677, n2667, n2676);
   xor (n2678, n503, n506);
   xor (n2679, n2678, n517);
   and (n268, n40, n267);
   not (n2680, n2679);
   or (n2681, n866, n871);
   not (n2682, n861);
   or (n2683, n2682, n751);
   nand (n2684, n2681, n2683);
   xor (n2685, n2680, n2684);
   xor (n2686, n2677, n2685);
   and (n2687, n828, n848);
   and (n2688, n808, n827);
   nor (n2689, n2687, n2688);
   not (n269, n40);
   xor (n2690, n2686, n2689);
   xor (n2691, n2666, n2690);
   nand (n2692, n2663, n2691);
   xnor (n2693, n522, n523);
   not (n2694, n2667);
   and (n2695, n2676, n2694);
   and (n2696, n2672, n871);
   nor (n2697, n2695, n2696);
   xor (n2698, n2693, n2697);
   not (n2699, n2667);
   buf (n27, g26);
   and (n270, n269, n52);
   not (n2700, n2676);
   or (n2701, n2699, n2700);
   or (n2702, n2676, n2667);
   nand (n2703, n2701, n2702);
   and (n2704, n2703, n2685);
   and (n2705, n2680, n2684);
   nor (n2706, n2704, n2705);
   xor (n2707, n2698, n2706);
   not (n2708, n2707);
   or (n2709, n2690, n2666);
   nor (n271, n268, n270);
   xnor (n2710, n2703, n2685);
   or (n2711, n2710, n2689);
   nand (n2712, n2709, n2711);
   nand (n2713, n2708, n2712);
   nand (n2714, n2692, n2713);
   nor (n2715, n2658, n2714);
   not (n2716, n2692);
   not (n2717, n2662);
   not (n2718, n2691);
   and (n2719, n2717, n2718);
   or (n272, n266, n271);
   and (n2720, n2662, n2691);
   nor (n2721, n2719, n2720);
   not (n2722, n2721);
   or (n2723, n2716, n2722);
   not (n2724, n2707);
   not (n2725, n2712);
   or (n2726, n2724, n2725);
   or (n2727, n2712, n2707);
   nand (n2728, n2726, n2727);
   nand (n2729, n2723, n2728);
   xor (n273, n41, n42);
   nand (n2730, n2729, n2713);
   xor (n2731, n494, n526);
   not (n2732, n2731);
   xor (n2733, n2693, n2697);
   and (n2734, n2733, n2706);
   and (n2735, n2693, n2697);
   nor (n2736, n2734, n2735);
   not (n2737, n2736);
   or (n2738, n2732, n2737);
   or (n2739, n2736, n2731);
   buf (n274, n273);
   nand (n2740, n2738, n2739);
   nand (n2741, n2730, n2740);
   or (n2742, n2715, n2741);
   not (n2743, n2731);
   nand (n2744, n2743, n2736);
   nand (n2745, n2742, n2744);
   xnor (n2746, n454, n529);
   nand (n2747, n2745, n2746);
   not (n2748, n2747);
   or (n2749, n531, n2748);
   not (n275, n274);
   and (n2750, n373, n450);
   not (n2751, n373);
   and (n2752, n2751, n451);
   nor (n2753, n2750, n2752);
   not (n2754, n2753);
   nand (n2755, n2749, n2754);
   nand (n2756, n453, n2755);
   and (n2757, n334, n337);
   and (n2758, n332, n333);
   nor (n2759, n2757, n2758);
   not (n276, n40);
   or (n2760, n247, n256);
   and (n2761, n312, n36);
   not (n2762, n36);
   and (n2763, n2762, n53);
   nor (n2764, n2761, n2763);
   or (n2765, n253, n2764);
   nand (n2766, n2760, n2765);
   or (n2767, n2766, n249);
   nand (n2768, n2766, n249);
   nand (n2769, n2767, n2768);
   nor (n277, n275, n276);
   not (n2770, n2769);
   or (n2771, n296, n330);
   nand (n2772, n311, n38);
   nand (n2773, n2771, n2772);
   not (n2774, n2773);
   and (n2775, n2770, n2774);
   and (n2776, n2769, n2773);
   nor (n2777, n2775, n2776);
   xnor (n2778, n2759, n2777);
   and (n2779, n321, n280);
   not (n278, n277);
   and (n2780, n258, n279);
   nor (n2781, n2779, n2780);
   xor (n2782, n2778, n2781);
   and (n2783, n343, n372);
   and (n2784, n322, n342);
   nor (n2785, n2783, n2784);
   xnor (n2786, n2782, n2785);
   and (n2787, n2756, n2786);
   not (n2788, n249);
   or (n2789, n2766, n2773, n2788);
   nand (n279, n272, n278);
   nand (n2790, n2766, n2773, n2788);
   nand (n2791, n2789, n2790);
   or (n2792, n247, n2764);
   and (n2793, n267, n36);
   and (n2794, n2762, n52);
   nor (n2795, n2793, n2794);
   or (n2796, n253, n2795);
   nand (n2797, n2792, n2796);
   not (n2798, n255);
   not (n2799, n1571);
   buf (n28, g27);
   xor (n280, n258, n279);
   and (n2800, n2798, n2799);
   not (n2801, n2798);
   and (n2802, n2801, n1571);
   nor (n2803, n2800, n2802);
   xnor (n2804, n2797, n2803);
   xnor (n2805, n2791, n2804);
   not (n2806, n2805);
   or (n2807, n2781, n2778);
   or (n2808, n2759, n2777);
   nand (n2809, n2807, n2808);
   or (n281, n36, n56);
   not (n2810, n2809);
   or (n2811, n2806, n2810);
   or (n2812, n2809, n2805);
   nand (n2813, n2811, n2812);
   not (n2814, n2813);
   not (n2815, n2785);
   nand (n2816, n2815, n2782);
   nand (n2817, n2814, n2816);
   nor (n2818, n2787, n2817);
   not (n2819, n2818);
   nand (n282, n36, n56);
   not (n2820, n2816);
   nand (n2821, n2756, n2786);
   not (n2822, n2821);
   or (n2823, n2820, n2822);
   nand (n2824, n2823, n2813);
   nand (n2825, n2819, n2824);
   not (n2826, n2825);
   or (n2827, n238, n2826);
   and (n2828, n3, n4);
   not (n2829, n3);
   nand (n283, n281, n282);
   and (n2830, n2829, n20);
   nor (n2831, n2828, n2830);
   buf (n2832, n2831);
   not (n2833, n2832);
   not (n2834, n2833);
   and (n2835, n2834, n298);
   nor (n2836, n2834, n298);
   nor (n2837, n2835, n2836);
   and (n2838, n2837, n297);
   not (n2839, n2772);
   or (n284, n247, n283);
   nor (n2840, n2838, n2839);
   and (n2841, n3, n6);
   not (n2842, n3);
   and (n2843, n2842, n22);
   nor (n2844, n2841, n2843);
   buf (n2845, n2844);
   not (n2846, n2845);
   xnor (n2847, n2846, n37);
   buf (n2848, n747);
   buf (n2849, n2848);
   or (n285, n253, n250);
   and (n2850, n2847, n2849);
   and (n2851, n3, n5);
   not (n2852, n3);
   and (n2853, n2852, n21);
   nor (n2854, n2851, n2853);
   not (n2855, n2854);
   and (n2856, n2855, n2762);
   not (n2857, n2855);
   and (n2858, n2857, n36);
   nor (n2859, n2856, n2858);
   nand (n286, n284, n285);
   not (n2860, n2859);
   not (n2861, n253);
   and (n2862, n2860, n2861);
   nor (n2863, n2850, n2862);
   and (n2864, n3, n7);
   not (n2865, n3);
   and (n2866, n2865, n23);
   nor (n2867, n2864, n2866);
   not (n2868, n2867);
   and (n2869, n2868, n36);
   not (n287, n286);
   not (n2870, n2869);
   and (n2871, n2840, n2863, n2870);
   nor (n2872, n2840, n2863, n2870);
   nor (n2873, n2871, n2872);
   or (n2874, n2859, n247);
   and (n2875, n2834, n36);
   not (n2876, n2834);
   and (n2877, n2876, n2762);
   nor (n2878, n2875, n2877);
   or (n2879, n2878, n253);
   nand (n288, n36, n57);
   nand (n2880, n2874, n2879);
   nor (n2881, n2845, n2762);
   or (n2882, n2881, n1571);
   nand (n2883, n2881, n1571);
   nand (n2884, n2882, n2883);
   xor (n2885, n2880, n2884);
   xor (n2886, n2873, n2885);
   not (n2887, n2886);
   or (n2888, n2840, n2869);
   nand (n2889, n2840, n2869);
   not (n289, n288);
   nand (n2890, n2888, n2889);
   not (n2891, n2890);
   not (n2892, n2863);
   and (n2893, n2891, n2892);
   and (n2894, n2890, n2863);
   nor (n2895, n2893, n2894);
   and (n2896, n2855, n38);
   not (n2897, n2855);
   and (n2898, n2897, n298);
   nor (n2899, n2896, n2898);
   buf (n29, g28);
   and (n290, n287, n289);
   and (n2900, n297, n2899);
   and (n2901, n2837, n311);
   nor (n2902, n2900, n2901);
   and (n2903, n3, n8);
   not (n2904, n3);
   and (n2905, n2904, n24);
   nor (n2906, n2903, n2905);
   buf (n2907, n2906);
   not (n2908, n2907);
   nand (n2909, n2908, n36);
   and (n291, n286, n288);
   and (n2910, n2909, n340);
   not (n2911, n2909);
   and (n2912, n2911, n337);
   nor (n2913, n2910, n2912);
   and (n2914, n2902, n2913);
   and (n2915, n2909, n340);
   nor (n2916, n2914, n2915);
   xor (n2917, n2895, n2916);
   not (n2918, n9);
   and (n2919, n3, n2918);
   nor (n292, n290, n291);
   not (n2920, n3);
   not (n2921, n25);
   and (n2922, n2920, n2921);
   nor (n2923, n2919, n2922);
   and (n2924, n2923, n36);
   buf (n2925, n2907);
   and (n2926, n37, n2925);
   not (n2927, n37);
   not (n2928, n2925);
   and (n2929, n2927, n2928);
   xor (n293, n38, n39);
   nor (n2930, n2926, n2929);
   and (n2931, n2930, n2849);
   not (n2932, n2868);
   and (n2933, n2932, n2762);
   nor (n2934, n2933, n2869);
   and (n2935, n2934, n2861);
   nor (n2936, n2931, n2935);
   not (n2937, n2936);
   xor (n2938, n2924, n2937);
   not (n2939, n311);
   xnor (n294, n40, n39);
   not (n2940, n2899);
   or (n2941, n2939, n2940);
   and (n2942, n2846, n298);
   not (n2943, n2846);
   and (n2944, n2943, n38);
   nor (n2945, n2942, n2944);
   or (n2946, n2945, n296);
   nand (n2947, n2941, n2946);
   and (n2948, n2938, n2947);
   and (n2949, n2924, n2937);
   nand (n295, n293, n294);
   nor (n2950, n2948, n2949);
   and (n2951, n2934, n2849);
   and (n2952, n2845, n2762);
   nor (n2953, n2952, n2881);
   and (n2954, n2953, n2861);
   nor (n2955, n2951, n2954);
   nand (n2956, n2833, n40);
   nand (n2957, n2832, n276);
   and (n2958, n2956, n2957);
   and (n2959, n2958, n362);
   buf (n296, n295);
   nor (n2960, n2959, n277);
   xnor (n2961, n2955, n2960);
   or (n2962, n2950, n2961);
   or (n2963, n2955, n2960);
   nand (n2964, n2962, n2963);
   and (n2965, n2917, n2964);
   and (n2966, n2895, n2916);
   nor (n2967, n2965, n2966);
   not (n2968, n2967);
   or (n2969, n2887, n2968);
   not (n297, n296);
   or (n2970, n2967, n2886);
   nand (n2971, n2969, n2970);
   not (n2972, n2971);
   xnor (n2973, n2917, n2964);
   not (n2974, n2973);
   xnor (n2975, n2855, n40);
   not (n2976, n2975);
   and (n2977, n2976, n362);
   and (n2978, n2958, n274);
   nor (n2979, n2977, n2978);
   not (n298, n38);
   not (n2980, n2762);
   not (n2981, n2907);
   or (n2982, n2980, n2981);
   nand (n2983, n2982, n2909);
   not (n2984, n2983);
   not (n2985, n253);
   and (n2986, n2984, n2985);
   and (n2987, n3, n9);
   not (n2988, n3);
   and (n2989, n2988, n25);
   not (n299, n54);
   nor (n2990, n2987, n2989);
   buf (n2991, n2990);
   and (n2992, n2991, n2762);
   nor (n2993, n2992, n2924);
   and (n2994, n2993, n2848);
   nor (n2995, n2986, n2994);
   not (n2996, n2995);
   not (n2997, n353);
   and (n2998, n2996, n2997);
   and (n2999, n2995, n353);
   buf (n3, g2);
   buf (n30, g29);
   and (n300, n298, n299);
   nor (n3000, n2998, n2999);
   or (n3001, n2979, n3000);
   or (n3002, n2995, n352);
   nand (n3003, n3001, n3002);
   xor (n3004, n3003, n2960);
   xor (n3005, n2924, n2937);
   xor (n3006, n3005, n2947);
   and (n3007, n3004, n3006);
   and (n3008, n3003, n2960);
   nor (n3009, n3007, n3008);
   and (n301, n38, n54);
   xnor (n3010, n2950, n2961);
   xor (n3011, n2902, n2913);
   xor (n3012, n3010, n3011);
   and (n3013, n3009, n3012);
   and (n3014, n3010, n3011);
   nor (n3015, n3013, n3014);
   not (n3016, n3015);
   or (n3017, n2974, n3016);
   or (n3018, n2973, n3015);
   nand (n3019, n3017, n3018);
   nor (n302, n300, n301);
   not (n3020, n3019);
   xnor (n3021, n3009, n3012);
   not (n3022, n3021);
   xnor (n3023, n3004, n3006);
   xnor (n3024, n2932, n38);
   not (n3025, n3024);
   not (n3026, n297);
   or (n3027, n3025, n3026);
   or (n3028, n2945, n326);
   nand (n3029, n3027, n3028);
   and (n303, n297, n302);
   and (n3030, n3, n10);
   not (n3031, n3);
   and (n3032, n3031, n26);
   nor (n3033, n3030, n3032);
   buf (n3034, n3033);
   not (n3035, n3034);
   and (n3036, n36, n3035);
   xor (n3037, n3029, n3036);
   not (n3038, n40);
   and (n3039, n3, n6);
   not (n304, n263);
   not (n3040, n3);
   and (n3041, n3040, n22);
   nor (n3042, n3039, n3041);
   not (n3043, n3042);
   not (n3044, n3043);
   not (n3045, n3044);
   or (n3046, n3038, n3045);
   or (n3047, n2845, n40);
   nand (n3048, n3046, n3047);
   not (n3049, n3048);
   not (n305, n39);
   or (n3050, n266, n3049);
   or (n3051, n2975, n275);
   nand (n3052, n3050, n3051);
   and (n3053, n3037, n3052);
   and (n3054, n3029, n3036);
   nor (n3055, n3053, n3054);
   xnor (n3056, n3023, n3055);
   xor (n3057, n3000, n2979);
   not (n3058, n2831);
   xor (n3059, n42, n3058);
   not (n306, n305);
   and (n3060, n3059, n738);
   nor (n3061, n3060, n432);
   and (n3062, n3, n11);
   not (n3063, n3);
   and (n3064, n3063, n27);
   nor (n3065, n3062, n3064);
   buf (n3066, n3065);
   not (n3067, n3066);
   nand (n3068, n3067, n36);
   xor (n3069, n3061, n3068);
   or (n307, n304, n306);
   not (n3070, n3033);
   not (n3071, n3070);
   not (n3072, n3071);
   not (n3073, n37);
   and (n3074, n3072, n3073);
   and (n3075, n3071, n37);
   nor (n3076, n3074, n3075);
   and (n3077, n2848, n3076);
   and (n3078, n2993, n2861);
   nor (n3079, n3077, n3078);
   nand (n308, n39, n40);
   and (n3080, n3069, n3079);
   and (n3081, n3061, n3068);
   nor (n3082, n3080, n3081);
   xor (n3083, n3057, n3082);
   xor (n3084, n3037, n3052);
   and (n3085, n3083, n3084);
   and (n3086, n3057, n3082);
   nor (n3087, n3085, n3086);
   or (n3088, n3056, n3087);
   or (n3089, n3023, n3055);
   nand (n309, n307, n308);
   nand (n3090, n3088, n3089);
   not (n3091, n3090);
   or (n3092, n3022, n3091);
   xor (n3093, n3057, n3082);
   xor (n3094, n3093, n3084);
   not (n3095, n296);
   not (n3096, n38);
   not (n3097, n2907);
   or (n3098, n3096, n3097);
   or (n3099, n2907, n38);
   buf (n31, g30);
   not (n310, n309);
   nand (n3100, n3098, n3099);
   not (n3101, n3100);
   not (n3102, n3101);
   and (n3103, n3095, n3102);
   and (n3104, n3024, n311);
   nor (n3105, n3103, n3104);
   xor (n3106, n3105, n3052);
   not (n3107, n3106);
   not (n3108, n465);
   and (n3109, n3, n7);
   buf (n311, n310);
   not (n3110, n3);
   and (n3111, n3110, n23);
   or (n3112, n3109, n3111);
   not (n3113, n3112);
   and (n3114, n40, n3113);
   not (n3115, n40);
   and (n3116, n3115, n3112);
   or (n3117, n3114, n3116);
   not (n3118, n3117);
   or (n3119, n3108, n3118);
   not (n312, n53);
   nand (n3120, n3048, n274);
   nand (n3121, n3119, n3120);
   not (n3122, n3121);
   and (n3123, n3, n12);
   not (n3124, n3);
   and (n3125, n3124, n28);
   nor (n3126, n3123, n3125);
   buf (n3127, n3126);
   not (n3128, n3127);
   nand (n3129, n3128, n36);
   and (n313, n298, n312);
   not (n3130, n3129);
   and (n3131, n3122, n3130);
   and (n3132, n3121, n3129);
   nor (n3133, n3131, n3132);
   not (n3134, n2848);
   not (n3135, n3134);
   not (n3136, n2762);
   not (n3137, n3066);
   or (n3138, n3136, n3137);
   nand (n3139, n3138, n3068);
   and (n314, n38, n53);
   not (n3140, n3139);
   and (n3141, n3135, n3140);
   xor (n3142, n36, n3035);
   not (n3143, n3142);
   nor (n3144, n3143, n253);
   nor (n3145, n3141, n3144);
   or (n3146, n3133, n3145);
   not (n3147, n3121);
   or (n3148, n3147, n3129);
   nand (n3149, n3146, n3148);
   nor (n315, n313, n314);
   not (n3150, n3149);
   or (n3151, n3107, n3150);
   or (n3152, n3105, n3052);
   nand (n3153, n3151, n3152);
   xor (n3154, n3094, n3153);
   xor (n3155, n3061, n3068);
   xor (n3156, n3155, n3079);
   not (n3157, n38);
   not (n3158, n2991);
   or (n3159, n3157, n3158);
   and (n316, n311, n315);
   or (n3160, n2991, n38);
   nand (n3161, n3159, n3160);
   not (n3162, n3161);
   not (n3163, n376);
   or (n3164, n3162, n3163);
   nand (n3165, n3100, n311);
   nand (n3166, n3164, n3165);
   nand (n3167, n801, n44);
   and (n3168, n3166, n3167);
   not (n3169, n3166);
   nor (n317, n303, n316);
   not (n3170, n3167);
   and (n3171, n3169, n3170);
   nor (n3172, n3168, n3171);
   not (n3173, n515);
   not (n3174, n3059);
   or (n3175, n3173, n3174);
   not (n3176, n2855);
   and (n3177, n42, n3176);
   not (n3178, n42);
   and (n3179, n3178, n2855);
   or (n318, n292, n317);
   or (n3180, n3177, n3179);
   not (n3181, n3180);
   or (n3182, n737, n3181);
   nand (n3183, n3175, n3182);
   and (n3184, n3172, n3183);
   and (n3185, n3166, n3167);
   nor (n3186, n3184, n3185);
   xor (n3187, n3156, n3186);
   xnor (n3188, n3149, n3106);
   and (n3189, n3187, n3188);
   not (n319, n286);
   and (n3190, n3156, n3186);
   nor (n3191, n3189, n3190);
   and (n3192, n3154, n3191);
   and (n3193, n3094, n3153);
   nor (n3194, n3192, n3193);
   not (n3195, n3194);
   xor (n3196, n3056, n3087);
   nand (n3197, n3195, n3196);
   not (n3198, n3197);
   xnor (n3199, n3154, n3191);
   buf (n32, g31);
   or (n320, n319, n288);
   not (n3200, n3199);
   xor (n3201, n3156, n3186);
   xor (n3202, n3201, n3188);
   not (n3203, n3033);
   not (n3204, n3203);
   not (n3205, n38);
   and (n3206, n3204, n3205);
   not (n3207, n3204);
   and (n3208, n3207, n38);
   nor (n3209, n3206, n3208);
   nand (n321, n318, n320);
   not (n3210, n3209);
   or (n3211, n296, n3210);
   not (n3212, n3161);
   or (n3213, n3212, n326);
   nand (n3214, n3211, n3213);
   not (n3215, n3214);
   xor (n3216, n44, n3058);
   not (n3217, n3216);
   not (n3218, n44);
   not (n3219, n803);
   xor (n322, n280, n321);
   or (n3220, n3218, n3219);
   not (n3221, n44);
   nand (n3222, n3221, n45, n46);
   nand (n3223, n3220, n3222);
   buf (n3224, n3223);
   not (n3225, n3224);
   or (n3226, n3217, n3225);
   nand (n3227, n805, n44);
   nand (n3228, n3226, n3227);
   not (n3229, n3228);
   not (n323, n315);
   not (n3230, n3139);
   not (n3231, n253);
   and (n3232, n3230, n3231);
   and (n3233, n3, n12);
   not (n3234, n3);
   and (n3235, n3234, n28);
   nor (n3236, n3233, n3235);
   not (n3237, n3236);
   buf (n3238, n3237);
   not (n3239, n3238);
   not (n324, n297);
   not (n3240, n3239);
   not (n3241, n37);
   and (n3242, n3240, n3241);
   and (n3243, n3127, n37);
   nor (n3244, n3242, n3243);
   and (n3245, n3244, n2848);
   nor (n3246, n3232, n3245);
   not (n3247, n3246);
   or (n3248, n3229, n3247);
   or (n3249, n3228, n3246);
   or (n325, n323, n324);
   nand (n3250, n3248, n3249);
   not (n3251, n3250);
   or (n3252, n3215, n3251);
   not (n3253, n3246);
   nand (n3254, n3253, n3228);
   nand (n3255, n3252, n3254);
   not (n3256, n3255);
   not (n3257, n430);
   not (n3258, n3180);
   or (n3259, n3257, n3258);
   not (n326, n311);
   not (n3260, n42);
   not (n3261, n2845);
   or (n3262, n3260, n3261);
   or (n3263, n2845, n42);
   nand (n3264, n3262, n3263);
   nand (n3265, n3264, n867);
   nand (n3266, n3259, n3265);
   not (n3267, n3266);
   not (n3268, n3267);
   and (n3269, n3256, n3268);
   and (n327, n38, n267);
   and (n3270, n3255, n3267);
   nor (n3271, n3269, n3270);
   not (n3272, n3271);
   xor (n3273, n3133, n3145);
   and (n3274, n3272, n3273);
   and (n3275, n3255, n3266);
   nor (n3276, n3274, n3275);
   xor (n3277, n3202, n3276);
   not (n3278, n3273);
   not (n3279, n3278);
   not (n328, n38);
   not (n3280, n3272);
   or (n3281, n3279, n3280);
   nand (n3282, n3271, n3273);
   nand (n3283, n3281, n3282);
   xor (n3284, n3172, n3183);
   and (n3285, n3, n13);
   not (n3286, n3);
   and (n3287, n3286, n29);
   or (n3288, n3285, n3287);
   buf (n3289, n3288);
   and (n329, n328, n52);
   and (n3290, n36, n3289);
   not (n3291, n3290);
   and (n3292, n3267, n3291);
   and (n3293, n3266, n3290);
   nor (n3294, n3292, n3293);
   xor (n3295, n2907, n40);
   not (n3296, n3295);
   and (n3297, n3296, n362);
   and (n3298, n3117, n274);
   nor (n3299, n3297, n3298);
   buf (n33, g32);
   nor (n330, n327, n329);
   or (n3300, n3294, n3299);
   or (n3301, n3266, n3291);
   nand (n3302, n3300, n3301);
   xor (n3303, n3284, n3302);
   and (n3304, n3283, n3303);
   and (n3305, n3284, n3302);
   nor (n3306, n3304, n3305);
   and (n3307, n3277, n3306);
   and (n3308, n3202, n3276);
   nor (n3309, n3307, n3308);
   or (n331, n326, n330);
   nand (n3310, n3200, n3309);
   not (n3311, n3310);
   not (n3312, n3);
   nand (n3313, n3312, n35);
   not (n3314, n35);
   or (n3315, n3314, n19);
   nand (n3316, n3315, n3);
   nand (n3317, n3313, n3316);
   buf (n3318, n3317);
   buf (n3319, n3318);
   nand (n332, n325, n331);
   nand (n3320, n3319, n401);
   nand (n3321, n3320, n1267);
   not (n3322, n3321);
   not (n3323, n51);
   and (n3324, n3, n4);
   not (n3325, n3);
   and (n3326, n3325, n20);
   nor (n3327, n3324, n3326);
   not (n3328, n3327);
   or (n3329, n3328, n50);
   not (n333, n282);
   nand (n3330, n3328, n50);
   nand (n3331, n3329, n3330);
   not (n3332, n3331);
   or (n3333, n3323, n3332);
   not (n3334, n51);
   and (n3335, n2855, n3334);
   nor (n3336, n3335, n1274);
   nand (n3337, n3333, n3336);
   not (n3338, n3337);
   or (n3339, n3322, n3338);
   xor (n334, n332, n333);
   not (n3340, n3321);
   not (n3341, n3337);
   nand (n3342, n3340, n3341);
   nand (n3343, n3339, n3342);
   not (n3344, n311);
   not (n3345, n38);
   and (n3346, n3, n16);
   not (n3347, n3);
   and (n3348, n3347, n32);
   nor (n3349, n3346, n3348);
   not (n335, n41);
   not (n3350, n3349);
   not (n3351, n3350);
   not (n3352, n3351);
   or (n3353, n3345, n3352);
   not (n3354, n3350);
   or (n3355, n3354, n38);
   nand (n3356, n3353, n3355);
   not (n3357, n3356);
   or (n3358, n3344, n3357);
   and (n3359, n3, n17);
   or (n336, n335, n273);
   not (n3360, n3);
   and (n3361, n3360, n33);
   nor (n3362, n3359, n3361);
   buf (n3363, n3362);
   xor (n3364, n38, n3363);
   not (n3365, n3364);
   nand (n3366, n3365, n495);
   nand (n3367, n3358, n3366);
   not (n3368, n3367);
   xor (n3369, n3343, n3368);
   nand (n337, n336, n40);
   not (n3370, n1075);
   not (n3371, n2907);
   xor (n3372, n48, n3371);
   not (n3373, n3372);
   or (n3374, n3370, n3373);
   and (n3375, n48, n2868);
   not (n3376, n48);
   and (n3377, n3, n7);
   not (n3378, n3);
   and (n3379, n3378, n23);
   and (n338, n334, n337);
   nor (n3380, n3377, n3379);
   and (n3381, n3376, n3380);
   nor (n3382, n3375, n3381);
   nand (n3383, n3382, n1944);
   nand (n3384, n3374, n3383);
   not (n3385, n3384);
   not (n3386, n2845);
   and (n3387, n3386, n3334);
   and (n3388, n3, n5);
   not (n3389, n3);
   not (n339, n334);
   and (n3390, n3389, n21);
   nor (n3391, n3388, n3390);
   and (n3392, n1005, n3391);
   nor (n3393, n3387, n3392);
   and (n3394, n1574, n2855);
   nor (n3395, n3394, n1274);
   nand (n3396, n3393, n3395);
   and (n3397, n3396, n3320);
   not (n3398, n3396);
   not (n3399, n3320);
   buf (n34, g33);
   not (n340, n337);
   and (n3400, n3398, n3399);
   nor (n3401, n3397, n3400);
   not (n3402, n3401);
   or (n3403, n3385, n3402);
   not (n3404, n3396);
   nand (n3405, n3404, n3399);
   nand (n3406, n3403, n3405);
   not (n3407, n3406);
   and (n3408, n3369, n3407);
   and (n3409, n3343, n3368);
   and (n341, n339, n340);
   or (n3410, n3408, n3409);
   not (n3411, n3410);
   not (n3412, n3411);
   not (n3413, n274);
   not (n3414, n276);
   and (n3415, n3, n14);
   not (n3416, n3);
   and (n3417, n3416, n30);
   nor (n3418, n3415, n3417);
   buf (n3419, n3418);
   nor (n342, n338, n341);
   not (n3420, n3419);
   not (n3421, n3420);
   or (n3422, n3414, n3421);
   nand (n3423, n3419, n40);
   nand (n3424, n3422, n3423);
   not (n3425, n3424);
   or (n3426, n3413, n3425);
   and (n3427, n3, n15);
   not (n3428, n3);
   and (n3429, n3428, n31);
   xor (n343, n322, n342);
   nor (n3430, n3427, n3429);
   buf (n3431, n3430);
   and (n3432, n40, n3431);
   not (n3433, n40);
   not (n3434, n3431);
   and (n3435, n3433, n3434);
   or (n3436, n3432, n3435);
   nand (n3437, n3436, n362);
   nand (n3438, n3426, n3437);
   not (n3439, n430);
   xnor (n344, n292, n317);
   not (n3440, n3237);
   and (n3441, n42, n3440);
   not (n3442, n42);
   and (n3443, n3442, n3238);
   or (n3444, n3441, n3443);
   not (n3445, n3444);
   or (n3446, n3439, n3445);
   not (n3447, n42);
   and (n3448, n3, n13);
   not (n3449, n3);
   xnor (n345, n344, n279);
   and (n3450, n3449, n29);
   nor (n3451, n3448, n3450);
   not (n3452, n3451);
   or (n3453, n3447, n3452);
   and (n3454, n3, n13);
   not (n3455, n3);
   and (n3456, n3455, n29);
   nor (n3457, n3454, n3456);
   or (n3458, n3457, n42);
   nand (n3459, n3453, n3458);
   or (n346, n36, n57);
   nand (n3460, n3459, n867);
   nand (n3461, n3446, n3460);
   xor (n3462, n3438, n3461);
   not (n3463, n3462);
   and (n3464, n2991, n46);
   not (n3465, n2991);
   and (n3466, n3465, n504);
   nor (n3467, n3464, n3466);
   not (n3468, n533);
   nand (n3469, n3468, n532);
   nand (n347, n346, n288);
   not (n3470, n3469);
   buf (n3471, n3470);
   not (n3472, n3471);
   or (n3473, n3467, n3472);
   and (n3474, n2908, n504);
   not (n3475, n2908);
   and (n3476, n3475, n46);
   nor (n3477, n3474, n3476);
   or (n3478, n3477, n1019);
   nand (n3479, n3473, n3478);
   or (n348, n247, n347);
   not (n3480, n3479);
   or (n3481, n3463, n3480);
   nand (n3482, n3438, n3461);
   nand (n3483, n3481, n3482);
   not (n3484, n3483);
   not (n3485, n3484);
   buf (n3486, n3342);
   not (n3487, n3486);
   not (n3488, n252);
   not (n3489, n18);
   or (n349, n253, n283);
   and (n3490, n3489, n3);
   nor (n3491, n3, n34);
   nor (n3492, n3490, n3491);
   buf (n3493, n3492);
   nand (n3494, n3493, n36);
   not (n3495, n3493);
   nand (n3496, n3495, n2762);
   and (n3497, n3494, n3496);
   not (n3498, n3497);
   or (n3499, n3488, n3498);
   buf (n35, g34);
   nand (n350, n348, n349);
   not (n3500, n3317);
   buf (n3501, n3500);
   not (n3502, n3501);
   nor (n3503, n3502, n36);
   not (n3504, n3503);
   nand (n3505, n3319, n36);
   nand (n3506, n3504, n3505, n2848);
   nand (n3507, n3499, n3506);
   not (n3508, n3507);
   not (n3509, n3224);
   nand (n351, n43, n44);
   not (n3510, n3065);
   not (n3511, n3510);
   not (n3512, n44);
   and (n3513, n3511, n3512);
   and (n3514, n3510, n44);
   nor (n3515, n3513, n3514);
   not (n3516, n3515);
   or (n3517, n3509, n3516);
   and (n3518, n3, n10);
   not (n3519, n3);
   and (n352, n351, n42);
   and (n3520, n3519, n26);
   nor (n3521, n3518, n3520);
   not (n3522, n3521);
   not (n3523, n3522);
   not (n3524, n412);
   or (n3525, n3523, n3524);
   nand (n3526, n3521, n44);
   nand (n3527, n3525, n3526);
   nand (n3528, n805, n3527);
   nand (n3529, n3517, n3528);
   not (n353, n352);
   not (n3530, n3382);
   not (n3531, n1779);
   or (n3532, n3530, n3531);
   not (n3533, n48);
   not (n3534, n3533);
   not (n3535, n3043);
   or (n3536, n3534, n3535);
   nand (n3537, n3044, n48);
   nand (n3538, n3536, n3537);
   nand (n3539, n3538, n614);
   and (n354, n350, n353);
   nand (n3540, n3532, n3539);
   xor (n3541, n3529, n3540);
   not (n3542, n3541);
   or (n3543, n3508, n3542);
   nand (n3544, n3529, n3540);
   nand (n3545, n3543, n3544);
   not (n3546, n3545);
   or (n3547, n3487, n3546);
   or (n3548, n3545, n3486);
   nand (n3549, n3547, n3548);
   not (n355, n350);
   not (n3550, n3549);
   or (n3551, n3485, n3550);
   or (n3552, n3549, n3484);
   nand (n3553, n3551, n3552);
   not (n3554, n3553);
   or (n3555, n3412, n3554);
   xor (n3556, n3529, n3540);
   xor (n3557, n3507, n3556);
   not (n3558, n3557);
   not (n3559, n3467);
   and (n356, n355, n352);
   not (n3560, n543);
   and (n3561, n3559, n3560);
   not (n3562, n3070);
   not (n3563, n3562);
   not (n3564, n47);
   and (n3565, n3563, n3564);
   and (n3566, n3204, n47);
   nor (n3567, n3565, n3566);
   and (n3568, n3471, n3567);
   nor (n3569, n3561, n3568);
   nor (n357, n354, n356);
   not (n3570, n3569);
   not (n3571, n3570);
   not (n3572, n421);
   not (n3573, n42);
   not (n3574, n3419);
   or (n3575, n3573, n3574);
   or (n3576, n3419, n42);
   nand (n3577, n3575, n3576);
   not (n3578, n3577);
   or (n3579, n3572, n3578);
   and (n358, n276, n312);
   nand (n3580, n3459, n513);
   nand (n3581, n3579, n3580);
   not (n3582, n3581);
   and (n3583, n3515, n805);
   not (n3584, n44);
   not (n3585, n3126);
   or (n3586, n3584, n3585);
   or (n3587, n3440, n44);
   nand (n3588, n3586, n3587);
   not (n3589, n3588);
   and (n359, n40, n53);
   not (n3590, n3224);
   nor (n3591, n3589, n3590);
   nor (n3592, n3583, n3591);
   not (n3593, n3592);
   or (n3594, n3582, n3593);
   or (n3595, n3581, n3592);
   nand (n3596, n3594, n3595);
   not (n3597, n3596);
   or (n3598, n3571, n3597);
   and (n3599, n3515, n805);
   buf (n36, g35);
   nor (n360, n358, n359);
   nor (n3600, n3599, n3591);
   not (n3601, n3600);
   nand (n3602, n3601, n3581);
   nand (n3603, n3598, n3602);
   not (n3604, n3603);
   not (n3605, n3604);
   not (n3606, n3479);
   not (n3607, n3462);
   not (n3608, n3607);
   or (n3609, n3606, n3608);
   not (n361, n360);
   not (n3610, n3479);
   nand (n3611, n3610, n3462);
   nand (n3612, n3609, n3611);
   not (n3613, n3612);
   or (n3614, n3605, n3613);
   or (n3615, n3612, n3604);
   nand (n3616, n3614, n3615);
   not (n3617, n3616);
   or (n3618, n3558, n3617);
   not (n3619, n3604);
   not (n362, n266);
   nand (n3620, n3619, n3612);
   nand (n3621, n3618, n3620);
   not (n3622, n3621);
   not (n3623, n3553);
   not (n3624, n3410);
   and (n3625, n3623, n3624);
   and (n3626, n3553, n3410);
   nor (n3627, n3625, n3626);
   or (n3628, n3622, n3627);
   nand (n3629, n3555, n3628);
   not (n363, n362);
   not (n3630, n3629);
   not (n3631, n857);
   not (n3632, n3424);
   or (n3633, n3631, n3632);
   not (n3634, n40);
   not (n3635, n3457);
   or (n3636, n3634, n3635);
   or (n3637, n3457, n40);
   nand (n3638, n3636, n3637);
   nand (n3639, n3638, n274);
   or (n364, n361, n363);
   nand (n3640, n3633, n3639);
   not (n3641, n3640);
   and (n3642, n3, n8);
   not (n3643, n3);
   and (n3644, n3643, n24);
   nor (n3645, n3642, n3644);
   not (n3646, n3645);
   and (n3647, n47, n3646);
   not (n3648, n47);
   and (n3649, n3648, n3645);
   or (n365, n275, n271);
   or (n3650, n3647, n3649);
   and (n3651, n3471, n3650);
   and (n3652, n46, n3112);
   not (n3653, n46);
   and (n3654, n3653, n3380);
   nor (n3655, n3652, n3654);
   and (n3656, n3655, n542);
   nor (n3657, n3651, n3656);
   not (n3658, n3657);
   not (n3659, n376);
   nand (n366, n364, n365);
   not (n3660, n3356);
   or (n3661, n3659, n3660);
   not (n3662, n298);
   not (n3663, n3434);
   or (n3664, n3662, n3663);
   buf (n3665, n3431);
   not (n3666, n3665);
   or (n3667, n3666, n298);
   nand (n3668, n3664, n3667);
   nand (n3669, n3668, n311);
   and (n367, n357, n366);
   nand (n3670, n3661, n3669);
   not (n3671, n3670);
   or (n3672, n3658, n3671);
   or (n3673, n3657, n3670);
   nand (n3674, n3672, n3673);
   not (n3675, n3674);
   or (n3676, n3641, n3675);
   not (n3677, n3657);
   nand (n3678, n3677, n3670);
   nand (n3679, n3676, n3678);
   and (n368, n350, n353);
   not (n3680, n3679);
   not (n3681, n3505);
   not (n3682, n50);
   not (n3683, n2831);
   or (n3684, n3682, n3683);
   nand (n3685, n3684, n1480);
   not (n3686, n3685);
   and (n3687, n3681, n3686);
   and (n3688, n3505, n3685);
   nor (n3689, n3687, n3688);
   nor (n369, n367, n368);
   not (n3690, n3689);
   not (n3691, n3538);
   not (n3692, n1778);
   buf (n3693, n3692);
   not (n3694, n3693);
   or (n3695, n3691, n3694);
   not (n3696, n3533);
   not (n3697, n3391);
   not (n3698, n3697);
   or (n3699, n3696, n3698);
   buf (n37, g36);
   or (n370, n345, n369);
   or (n3700, n3697, n3533);
   nand (n3701, n3699, n3700);
   nand (n3702, n3701, n1039);
   nand (n3703, n3695, n3702);
   nand (n3704, n3690, n3703);
   not (n3705, n3505);
   nand (n3706, n3705, n3685);
   and (n3707, n3704, n3706);
   not (n3708, n3707);
   and (n3709, n3680, n3708);
   or (n371, n344, n279);
   and (n3710, n3679, n3707);
   nor (n3711, n3709, n3710);
   not (n3712, n421);
   not (n3713, n3444);
   or (n3714, n3712, n3713);
   not (n3715, n3510);
   not (n3716, n42);
   and (n3717, n3715, n3716);
   and (n3718, n3067, n42);
   nor (n3719, n3717, n3718);
   nand (n372, n370, n371);
   nand (n3720, n3719, n430);
   nand (n3721, n3714, n3720);
   not (n3722, n3721);
   not (n3723, n2923);
   not (n3724, n412);
   and (n3725, n3723, n3724);
   and (n3726, n2923, n412);
   nor (n3727, n3725, n3726);
   not (n3728, n3727);
   not (n3729, n556);
   xor (n373, n343, n372);
   and (n3730, n3728, n3729);
   and (n3731, n3224, n3527);
   nor (n3732, n3730, n3731);
   not (n3733, n3732);
   and (n3734, n3722, n3733);
   and (n3735, n3721, n3732);
   nor (n3736, n3734, n3735);
   not (n3737, n3363);
   nand (n3738, n3737, n36);
   not (n3739, n3737);
   not (n374, n373);
   nand (n3740, n3739, n2762);
   nand (n3741, n3738, n3740);
   not (n3742, n3741);
   not (n3743, n253);
   and (n3744, n3742, n3743);
   and (n3745, n2848, n3497);
   nor (n3746, n3744, n3745);
   or (n3747, n3736, n3746);
   not (n3748, n3721);
   or (n3749, n3748, n3732);
   xor (n375, n345, n369);
   nand (n3750, n3747, n3749);
   xor (n3751, n3711, n3750);
   not (n3752, n3483);
   not (n3753, n3549);
   or (n3754, n3752, n3753);
   not (n3755, n3486);
   nand (n3756, n3755, n3545);
   nand (n3757, n3754, n3756);
   not (n3758, n401);
   not (n3759, n16);
   not (n376, n295);
   and (n3760, n3, n3759);
   not (n3761, n3);
   not (n3762, n32);
   and (n3763, n3761, n3762);
   nor (n3764, n3760, n3763);
   buf (n3765, n3764);
   nor (n3766, n3765, n36);
   not (n3767, n3766);
   buf (n3768, n3765);
   nand (n3769, n3768, n36);
   not (n377, n55);
   nand (n3770, n3767, n3769);
   not (n3771, n3770);
   not (n3772, n3771);
   or (n3773, n3758, n3772);
   nand (n3774, n3738, n3740, n2848);
   nand (n3775, n3773, n3774);
   xor (n3776, n50, n3494);
   xor (n3777, n3775, n3776);
   and (n3778, n3719, n867);
   not (n3779, n42);
   and (n378, n298, n377);
   not (n3780, n3034);
   or (n3781, n3779, n3780);
   or (n3782, n3204, n42);
   nand (n3783, n3781, n3782);
   and (n3784, n3783, n430);
   nor (n3785, n3778, n3784);
   not (n3786, n3785);
   not (n3787, n3043);
   not (n3788, n504);
   and (n3789, n3787, n3788);
   and (n379, n38, n55);
   not (n3790, n2845);
   and (n3791, n3790, n504);
   nor (n3792, n3789, n3791);
   not (n3793, n3792);
   not (n3794, n1019);
   and (n3795, n3793, n3794);
   and (n3796, n3655, n3470);
   nor (n3797, n3795, n3796);
   not (n3798, n3797);
   not (n3799, n3798);
   buf (n38, g37);
   nor (n380, n378, n379);
   or (n3800, n3786, n3799);
   not (n3801, n3785);
   nand (n3802, n3801, n3797);
   nand (n3803, n3800, n3802);
   nor (n3804, n3058, n48);
   not (n3805, n3804);
   nand (n3806, n3058, n48);
   nand (n3807, n3805, n3806);
   not (n3808, n3807);
   not (n3809, n1038);
   and (n381, n376, n380);
   and (n3810, n3808, n3809);
   and (n3811, n3693, n3701);
   nor (n3812, n3810, n3811);
   and (n3813, n3803, n3812);
   not (n3814, n3803);
   not (n3815, n3812);
   and (n3816, n3814, n3815);
   nor (n3817, n3813, n3816);
   and (n3818, n3777, n3817);
   not (n3819, n3777);
   buf (n382, n310);
   not (n3820, n3817);
   and (n3821, n3819, n3820);
   or (n3822, n3818, n3821);
   xor (n3823, n3757, n3822);
   xor (n3824, n3751, n3823);
   not (n3825, n263);
   not (n3826, n3127);
   not (n3827, n3826);
   or (n3828, n3825, n3827);
   nand (n3829, n3127, n40);
   and (n383, n382, n302);
   nand (n3830, n3828, n3829);
   nand (n3831, n274, n3830);
   nand (n3832, n3638, n362);
   and (n3833, n3831, n3832);
   not (n3834, n311);
   not (n3835, n298);
   not (n3836, n3419);
   not (n3837, n3836);
   or (n3838, n3835, n3837);
   not (n3839, n3419);
   nor (n384, n381, n383);
   not (n3840, n3839);
   nand (n3841, n38, n3840);
   nand (n3842, n3838, n3841);
   not (n3843, n3842);
   or (n3844, n3834, n3843);
   nand (n3845, n376, n3668);
   nand (n3846, n3844, n3845);
   xor (n3847, n3833, n3846);
   xor (n3848, n2907, n44);
   nor (n3849, n3848, n556);
   nand (n385, n36, n58);
   nor (n3850, n3727, n3590);
   or (n3851, n3849, n3850);
   xor (n3852, n3847, n3851);
   xor (n3853, n3746, n3736);
   not (n3854, n3853);
   xor (n3855, n3689, n3703);
   not (n3856, n3855);
   not (n3857, n3674);
   not (n3858, n3640);
   not (n3859, n3858);
   xnor (n386, n384, n385);
   and (n3860, n3857, n3859);
   and (n3861, n3674, n3858);
   nor (n3862, n3860, n3861);
   not (n3863, n3862);
   not (n3864, n3863);
   or (n3865, n3856, n3864);
   not (n3866, n3855);
   nand (n3867, n3866, n3862);
   nand (n3868, n3865, n3867);
   not (n3869, n3868);
   and (n387, n40, n54);
   or (n3870, n3854, n3869);
   not (n3871, n3855);
   nand (n3872, n3871, n3863);
   nand (n3873, n3870, n3872);
   and (n3874, n3852, n3873);
   not (n3875, n3852);
   not (n3876, n3873);
   and (n3877, n3875, n3876);
   nor (n3878, n3874, n3877);
   xnor (n3879, n3824, n3878);
   nor (n388, n40, n54);
   not (n3880, n3879);
   or (n3881, n3630, n3880);
   not (n3882, n3751);
   xor (n3883, n3882, n3878);
   nand (n3884, n3823, n3883);
   nand (n3885, n3881, n3884);
   not (n3886, n3885);
   not (n3887, n3886);
   not (n3888, n3471);
   not (n3889, n3044);
   nor (n389, n387, n388);
   xor (n3890, n3564, n3889);
   not (n3891, n3890);
   or (n3892, n3888, n3891);
   not (n3893, n3697);
   not (n3894, n504);
   and (n3895, n3893, n3894);
   and (n3896, n2855, n504);
   nor (n3897, n3895, n3896);
   not (n3898, n3897);
   nand (n3899, n3898, n815);
   buf (n39, g38);
   and (n390, n362, n389);
   nand (n3900, n3892, n3899);
   not (n3901, n3738);
   and (n3902, n3900, n3901);
   not (n3903, n3900);
   and (n3904, n3903, n3738);
   nor (n3905, n3902, n3904);
   not (n3906, n3783);
   or (n3907, n3906, n737);
   and (n3908, n2923, n423);
   and (n3909, n2991, n42);
   and (n391, n274, n360);
   nor (n3910, n3908, n3909);
   or (n3911, n3910, n429);
   nand (n3912, n3907, n3911);
   xor (n3913, n3905, n3912);
   not (n3914, n3913);
   not (n3915, n3693);
   not (n3916, n610);
   not (n3917, n2831);
   or (n3918, n3916, n3917);
   nand (n3919, n3058, n49);
   nor (n392, n390, n391);
   nand (n3920, n3918, n3919);
   not (n3921, n3920);
   or (n3922, n3915, n3921);
   nand (n3923, n3922, n615);
   not (n3924, n3923);
   xor (n3925, n3924, n3851);
   not (n3926, n3770);
   not (n3927, n247);
   and (n3928, n3926, n3927);
   and (n3929, n3665, n2762);
   or (n393, n386, n392);
   nor (n3930, n3665, n2762);
   nor (n3931, n3929, n3930);
   and (n3932, n3931, n2861);
   nor (n3933, n3928, n3932);
   xnor (n3934, n3925, n3933);
   not (n3935, n3934);
   not (n3936, n3935);
   or (n3937, n3914, n3936);
   not (n3938, n3913);
   nand (n3939, n3938, n3934);
   or (n394, n384, n385);
   nand (n3940, n3937, n3939);
   not (n3941, n3750);
   not (n3942, n3711);
   not (n3943, n3942);
   or (n3944, n3941, n3943);
   not (n3945, n3707);
   nand (n3946, n3945, n3679);
   nand (n3947, n3944, n3946);
   xor (n3948, n3940, n3947);
   not (n3949, n3882);
   nand (n395, n393, n394);
   not (n3950, n3878);
   or (n3951, n3949, n3950);
   not (n3952, n3876);
   nand (n3953, n3952, n3852);
   nand (n3954, n3951, n3953);
   xor (n3955, n3948, n3954);
   not (n3956, n3955);
   not (n3957, n3848);
   and (n3958, n3957, n3224);
   and (n3959, n44, n3112);
   xor (n396, n375, n395);
   not (n3960, n44);
   and (n3961, n3960, n3113);
   nor (n3962, n3959, n3961);
   and (n3963, n3962, n805);
   nor (n3964, n3958, n3963);
   not (n3965, n3964);
   not (n3966, n3965);
   not (n3967, n376);
   not (n3968, n3842);
   or (n3969, n3967, n3968);
   or (n397, n36, n58);
   not (n3970, n38);
   not (n3971, n3457);
   or (n3972, n3970, n3971);
   or (n3973, n3457, n38);
   nand (n3974, n3972, n3973);
   nand (n3975, n3974, n382);
   nand (n3976, n3969, n3975);
   not (n3977, n3976);
   and (n3978, n362, n3830);
   not (n3979, n3510);
   nand (n398, n397, n385);
   not (n3980, n40);
   and (n3981, n3979, n3980);
   and (n3982, n3067, n40);
   nor (n3983, n3981, n3982);
   and (n3984, n3983, n274);
   nor (n3985, n3978, n3984);
   not (n3986, n3985);
   or (n3987, n3977, n3986);
   or (n3988, n3985, n3976);
   nand (n3989, n3987, n3988);
   or (n399, n247, n398);
   not (n3990, n3989);
   not (n3991, n3990);
   or (n3992, n3966, n3991);
   nand (n3993, n3989, n3964);
   nand (n3994, n3992, n3993);
   not (n3995, n3833);
   not (n3996, n3846);
   and (n3997, n3995, n3996);
   and (n3998, n3833, n3846);
   nor (n3999, n3997, n3998);
   buf (n4, g3);
   buf (n40, g39);
   buf (n400, n243);
   not (n4000, n3999);
   not (n4001, n3851);
   and (n4002, n4000, n4001);
   not (n4003, n3833);
   and (n4004, n3846, n4003);
   nor (n4005, n4002, n4004);
   xor (n4006, n3994, n4005);
   not (n4007, n3776);
   nor (n4008, n4007, n3775);
   and (n4009, n50, n3494);
   not (n401, n400);
   nor (n4010, n4008, n4009);
   not (n4011, n3815);
   not (n4012, n3803);
   or (n4013, n4011, n4012);
   not (n4014, n3785);
   nand (n4015, n4014, n3798);
   nand (n4016, n4013, n4015);
   xor (n4017, n4010, n4016);
   xnor (n4018, n4006, n4017);
   not (n4019, n3822);
   not (n402, n401);
   not (n4020, n3757);
   or (n4021, n4019, n4020);
   nand (n4022, n3777, n3820);
   nand (n4023, n4021, n4022);
   and (n4024, n4018, n4023);
   not (n4025, n4018);
   not (n4026, n4023);
   and (n4027, n4025, n4026);
   or (n4028, n4024, n4027);
   not (n4029, n4028);
   or (n403, n402, n347);
   and (n4030, n3956, n4029);
   and (n4031, n3955, n4028);
   nor (n4032, n4030, n4031);
   not (n4033, n4032);
   not (n4034, n4033);
   or (n4035, n3887, n4034);
   nand (n4036, n4032, n3885);
   nand (n4037, n4035, n4036);
   and (n4038, n3790, n50);
   and (n4039, n3044, n1005);
   nand (n404, n399, n403);
   nor (n4040, n4038, n4039);
   or (n4041, n4040, n3334);
   and (n4042, n2868, n3334);
   nor (n4043, n4042, n1274);
   nand (n4044, n4041, n4043);
   not (n4045, n4044);
   not (n4046, n3500);
   buf (n4047, n4046);
   nand (n4048, n4047, n311);
   nand (n4049, n4048, n1571);
   nand (n405, n36, n59);
   not (n4050, n4049);
   nand (n4051, n4045, n4050);
   not (n4052, n4051);
   not (n4053, n326);
   not (n4054, n3364);
   and (n4055, n4053, n4054);
   not (n4056, n38);
   and (n4057, n3, n3489);
   not (n4058, n3);
   not (n4059, n34);
   and (n406, n404, n405);
   and (n4060, n4058, n4059);
   nor (n4061, n4057, n4060);
   not (n4062, n4061);
   not (n4063, n4062);
   or (n4064, n4056, n4063);
   or (n4065, n3495, n38);
   nand (n4066, n4064, n4065);
   and (n4067, n4066, n376);
   nor (n4068, n4055, n4067);
   not (n4069, n4068);
   not (n407, n404);
   not (n4070, n3436);
   not (n4071, n274);
   or (n4072, n4070, n4071);
   not (n4073, n40);
   not (n4074, n3765);
   or (n4075, n4073, n4074);
   not (n4076, n3350);
   nand (n4077, n4076, n276);
   nand (n4078, n4075, n4077);
   not (n4079, n4078);
   not (n408, n405);
   nand (n4080, n4079, n857);
   nand (n4081, n4072, n4080);
   not (n4082, n4081);
   or (n4083, n4069, n4082);
   or (n4084, n4081, n4068);
   nand (n4085, n4083, n4084);
   nand (n4086, n4052, n4085);
   not (n4087, n4068);
   nand (n4088, n4087, n4081);
   and (n4089, n4086, n4088);
   and (n409, n407, n408);
   xor (n4090, n3368, n3343);
   xnor (n4091, n4090, n3406);
   xor (n4092, n4089, n4091);
   not (n4093, n310);
   not (n4094, n4066);
   or (n4095, n4093, n4094);
   not (n4096, n276);
   not (n4097, n4046);
   or (n4098, n4096, n4097);
   or (n4099, n4046, n263);
   buf (n41, g40);
   nor (n410, n406, n409);
   nand (n4100, n4098, n4099);
   or (n4101, n4100, n296);
   nand (n4102, n4095, n4101);
   not (n4103, n4102);
   not (n4104, n4078);
   not (n4105, n275);
   and (n4106, n4104, n4105);
   and (n4107, n3, n17);
   not (n4108, n3);
   and (n4109, n4108, n33);
   not (n411, n410);
   nor (n4110, n4107, n4109);
   not (n4111, n4110);
   and (n4112, n40, n4111);
   not (n4113, n40);
   and (n4114, n4113, n4110);
   or (n4115, n4112, n4114);
   nor (n4116, n4115, n266);
   nor (n4117, n4106, n4116);
   not (n4118, n4117);
   or (n4119, n4103, n4118);
   not (n412, n44);
   or (n4120, n4117, n4102);
   nand (n4121, n4119, n4120);
   not (n4122, n4121);
   not (n4123, n1019);
   and (n4124, n46, n3203);
   not (n4125, n46);
   and (n4126, n4125, n3204);
   or (n4127, n4124, n4126);
   not (n4128, n4127);
   and (n4129, n4123, n4128);
   not (n413, n412);
   and (n4130, n504, n3066);
   not (n4131, n504);
   and (n4132, n4131, n3510);
   nor (n4133, n4130, n4132);
   and (n4134, n3471, n4133);
   nor (n4135, n4129, n4134);
   not (n4136, n4135);
   not (n4137, n4136);
   or (n4138, n4122, n4137);
   not (n4139, n4117);
   not (n414, n42);
   nand (n4140, n4139, n4102);
   nand (n4141, n4138, n4140);
   not (n4142, n4141);
   xnor (n4143, n3401, n3384);
   not (n4144, n4143);
   not (n4145, n1944);
   not (n4146, n3372);
   or (n4147, n4145, n4146);
   and (n4148, n48, n2923);
   not (n4149, n48);
   nor (n415, n414, n43);
   and (n4150, n4149, n2991);
   nor (n4151, n4148, n4150);
   nand (n4152, n712, n4151);
   nand (n4153, n4147, n4152);
   not (n4154, n4153);
   not (n4155, n3224);
   not (n4156, n44);
   not (n4157, n3451);
   or (n4158, n4156, n4157);
   or (n4159, n3457, n44);
   not (n416, n415);
   nand (n4160, n4158, n4159);
   not (n4161, n4160);
   or (n4162, n4155, n4161);
   nand (n4163, n3588, n805);
   nand (n4164, n4162, n4163);
   not (n4165, n4164);
   not (n4166, n430);
   not (n4167, n3577);
   or (n4168, n4166, n4167);
   xnor (n4169, n42, n3431);
   or (n417, n413, n416);
   nand (n4170, n421, n4169);
   nand (n4171, n4168, n4170);
   not (n4172, n4171);
   not (n4173, n4172);
   or (n4174, n4165, n4173);
   or (n4175, n4172, n4164);
   nand (n4176, n4174, n4175);
   not (n4177, n4176);
   or (n4178, n4154, n4177);
   not (n4179, n4172);
   not (n418, n42);
   nand (n4180, n4179, n4164);
   nand (n4181, n4178, n4180);
   not (n4182, n4181);
   or (n4183, n4144, n4182);
   or (n4184, n4181, n4143);
   nand (n4185, n4183, n4184);
   nand (n4186, n4142, n4185);
   not (n4187, n4181);
   nand (n4188, n4187, n4143);
   nand (n4189, n4186, n4188);
   nand (n419, n418, n43, n44);
   not (n4190, n4189);
   and (n4191, n4092, n4190);
   not (n4192, n4092);
   and (n4193, n4192, n4189);
   nor (n4194, n4191, n4193);
   not (n4195, n4194);
   xor (n4196, n3557, n3604);
   xor (n4197, n4196, n3612);
   not (n4198, n4197);
   not (n4199, n4198);
   buf (n42, g41);
   nand (n420, n417, n419);
   xnor (n4200, n3596, n3569);
   not (n4201, n4200);
   xor (n4202, n4085, n4051);
   not (n4203, n4202);
   or (n4204, n4201, n4203);
   or (n4205, n4202, n4200);
   nand (n4206, n4204, n4205);
   not (n4207, n4206);
   nand (n4208, n4049, n4044);
   and (n4209, n4051, n4208);
   buf (n421, n420);
   not (n4210, n44);
   not (n4211, n3419);
   or (n4212, n4210, n4211);
   not (n4213, n3836);
   or (n4214, n4213, n44);
   nand (n4215, n4212, n4214);
   and (n4216, n4215, n3224);
   and (n4217, n4160, n805);
   nor (n4218, n4216, n4217);
   xor (n4219, n4048, n4218);
   buf (n422, n421);
   not (n4220, n3693);
   not (n4221, n4220);
   not (n4222, n610);
   not (n4223, n3035);
   or (n4224, n4222, n4223);
   nand (n4225, n3562, n49);
   nand (n4226, n4224, n4225);
   not (n4227, n4226);
   and (n4228, n4221, n4227);
   and (n4229, n4151, n1039);
   not (n423, n42);
   nor (n4230, n4228, n4229);
   and (n4231, n4219, n4230);
   and (n4232, n4048, n4218);
   nor (n4233, n4231, n4232);
   xor (n4234, n4209, n4233);
   not (n4235, n857);
   xor (n4236, n3493, n40);
   not (n4237, n4236);
   or (n4238, n4235, n4237);
   not (n4239, n4115);
   and (n424, n423, n267);
   nand (n4240, n4239, n274);
   nand (n4241, n4238, n4240);
   not (n4242, n4241);
   and (n4243, n1574, n2868);
   and (n4244, n2908, n3334);
   nor (n4245, n4243, n4244);
   and (n4246, n2932, n1005);
   nor (n4247, n4246, n1274);
   and (n4248, n4245, n4247);
   not (n4249, n738);
   and (n425, n42, n52);
   not (n4250, n3354);
   not (n4251, n423);
   and (n4252, n4250, n4251);
   and (n4253, n3351, n423);
   nor (n4254, n4252, n4253);
   not (n4255, n4254);
   or (n4256, n4249, n4255);
   nand (n4257, n4169, n430);
   nand (n4258, n4256, n4257);
   xor (n4259, n4248, n4258);
   nor (n426, n424, n425);
   not (n4260, n4259);
   or (n4261, n4242, n4260);
   nand (n4262, n4258, n4248);
   nand (n4263, n4261, n4262);
   and (n4264, n4234, n4263);
   and (n4265, n4209, n4233);
   nor (n4266, n4264, n4265);
   not (n4267, n4266);
   or (n4268, n4207, n4267);
   not (n4269, n4200);
   and (n427, n422, n426);
   nand (n4270, n4269, n4202);
   nand (n4271, n4268, n4270);
   not (n4272, n4271);
   or (n4273, n4199, n4272);
   not (n4274, n4271);
   nand (n4275, n4274, n4197);
   nand (n4276, n4273, n4275);
   not (n4277, n4276);
   or (n4278, n4195, n4277);
   nand (n4279, n4274, n4198);
   xor (n428, n43, n44);
   nand (n4280, n4278, n4279);
   not (n4281, n3622);
   not (n4282, n3627);
   not (n4283, n4282);
   or (n4284, n4281, n4283);
   nand (n4285, n3627, n3621);
   nand (n4286, n4284, n4285);
   and (n4287, n3868, n3853);
   not (n4288, n3868);
   not (n4289, n3853);
   not (n429, n428);
   and (n4290, n4288, n4289);
   or (n4291, n4287, n4290);
   not (n4292, n4291);
   and (n4293, n4189, n4092);
   and (n4294, n4089, n4091);
   nor (n4295, n4293, n4294);
   not (n4296, n4295);
   or (n4297, n4292, n4296);
   or (n4298, n4291, n4295);
   nand (n4299, n4297, n4298);
   buf (n43, g42);
   not (n430, n429);
   xor (n4300, n4286, n4299);
   xor (n4301, n4280, n4300);
   and (n4302, n4280, n4300);
   nor (n4303, n4301, n4302);
   xor (n4304, n3879, n3629);
   not (n4305, n4286);
   not (n4306, n4299);
   or (n4307, n4305, n4306);
   not (n4308, n4291);
   nand (n4309, n4308, n4295);
   not (n431, n430);
   nand (n4310, n4307, n4309);
   nor (n4311, n4304, n4310);
   nor (n4312, n4303, n4311);
   nand (n4313, n4037, n4312);
   not (n4314, n4141);
   not (n4315, n4185);
   or (n4316, n4314, n4315);
   buf (n4317, n4141);
   or (n4318, n4317, n4185);
   nand (n4319, n4316, n4318);
   nor (n432, n431, n423);
   not (n4320, n4319);
   not (n4321, n1956);
   not (n4322, n2991);
   or (n4323, n4321, n4322);
   not (n4324, n50);
   not (n4325, n3646);
   or (n4326, n4324, n4325);
   or (n4327, n2908, n50);
   nand (n4328, n4326, n4327);
   or (n4329, n4328, n3334);
   nor (n433, n427, n432);
   nand (n4330, n4323, n4329);
   not (n4331, n4330);
   not (n4332, n4331);
   not (n4333, n430);
   not (n4334, n4254);
   or (n4335, n4333, n4334);
   xor (n4336, n42, n4111);
   nand (n4337, n4336, n421);
   nand (n4338, n4335, n4337);
   not (n4339, n4338);
   not (n434, n433);
   or (n4340, n4332, n4339);
   or (n4341, n4338, n4331);
   nand (n4342, n4340, n4341);
   not (n4343, n4342);
   not (n4344, n805);
   not (n4345, n4215);
   or (n4346, n4344, n4345);
   not (n4347, n3431);
   and (n4348, n44, n4347);
   not (n4349, n44);
   and (n435, n411, n434);
   and (n4350, n4349, n3431);
   or (n4351, n4348, n4350);
   not (n4352, n4351);
   nand (n4353, n4352, n3224);
   nand (n4354, n4346, n4353);
   not (n4355, n4354);
   or (n4356, n4343, n4355);
   not (n4357, n4331);
   nand (n4358, n4357, n4338);
   nand (n4359, n4356, n4358);
   and (n436, n404, n408);
   not (n4360, n4359);
   not (n4361, n614);
   and (n4362, n48, n3521);
   not (n4363, n48);
   and (n4364, n4363, n3203);
   or (n4365, n4362, n4364);
   not (n4366, n4365);
   or (n4367, n4361, n4366);
   and (n4368, n48, n3065);
   not (n4369, n48);
   nor (n437, n435, n436);
   and (n4370, n3, n11);
   not (n4371, n3);
   and (n4372, n4371, n27);
   nor (n4373, n4370, n4372);
   not (n4374, n4373);
   and (n4375, n4369, n4374);
   or (n4376, n4368, n4375);
   nand (n4377, n711, n4376);
   nand (n4378, n4367, n4377);
   nand (n4379, n4046, n274);
   not (n438, n392);
   and (n4380, n4378, n4379, n340);
   and (n4381, n3440, n47);
   nor (n4382, n3127, n47);
   nor (n4383, n4381, n4382);
   and (n4384, n4383, n3471);
   and (n4385, n4133, n815);
   nor (n4386, n4384, n4385);
   not (n4387, n4386);
   and (n4388, n4380, n4387);
   not (n4389, n4380);
   and (n439, n386, n438);
   and (n4390, n4389, n4386);
   nor (n4391, n4388, n4390);
   not (n4392, n4391);
   or (n4393, n4360, n4392);
   nand (n4394, n4380, n4387);
   nand (n4395, n4393, n4394);
   not (n4396, n4395);
   not (n4397, n4153);
   not (n4398, n4397);
   not (n4399, n4176);
   buf (n44, g43);
   not (n440, n386);
   or (n4400, n4398, n4399);
   or (n4401, n4176, n4397);
   nand (n4402, n4400, n4401);
   not (n4403, n4402);
   not (n4404, n4121);
   not (n4405, n4135);
   and (n4406, n4404, n4405);
   and (n4407, n4121, n4135);
   nor (n4408, n4406, n4407);
   not (n4409, n4408);
   and (n441, n440, n392);
   or (n4410, n4403, n4409);
   or (n4411, n4408, n4402);
   nand (n4412, n4410, n4411);
   not (n4413, n4412);
   or (n4414, n4396, n4413);
   not (n4415, n4408);
   nand (n4416, n4415, n4402);
   nand (n4417, n4414, n4416);
   not (n4418, n4417);
   or (n4419, n4320, n4418);
   nor (n442, n439, n441);
   or (n4420, n4319, n4417);
   nand (n4421, n4419, n4420);
   not (n4422, n4421);
   not (n4423, n4266);
   not (n4424, n4423);
   buf (n4425, n4206);
   not (n4426, n4425);
   or (n4427, n4424, n4426);
   or (n4428, n4423, n4425);
   nand (n4429, n4427, n4428);
   xor (n443, n437, n442);
   not (n4430, n4429);
   not (n4431, n4430);
   or (n4432, n4422, n4431);
   not (n4433, n4319);
   nand (n4434, n4433, n4417);
   nand (n4435, n4432, n4434);
   not (n4436, n4435);
   and (n4437, n4276, n4194);
   not (n4438, n4276);
   not (n4439, n4194);
   xnor (n444, n357, n366);
   and (n4440, n4438, n4439);
   or (n4441, n4437, n4440);
   not (n4442, n4441);
   or (n4443, n4436, n4442);
   or (n4444, n4441, n4435);
   nand (n4445, n4443, n4444);
   xnor (n4446, n4412, n4395);
   not (n4447, n4446);
   not (n4448, n4447);
   not (n4449, n4230);
   and (n445, n443, n444);
   and (n4450, n4219, n4449);
   not (n4451, n4219);
   and (n4452, n4451, n4230);
   nor (n4453, n4450, n4452);
   not (n4454, n3471);
   xnor (n4455, n504, n3288);
   not (n4456, n4455);
   or (n4457, n4454, n4456);
   not (n4458, n46);
   not (n4459, n3127);
   and (n446, n437, n442);
   or (n4460, n4458, n4459);
   or (n4461, n3239, n46);
   nand (n4462, n4460, n4461);
   nand (n4463, n815, n4462);
   nand (n4464, n4457, n4463);
   not (n4465, n857);
   not (n4466, n4100);
   or (n4467, n4465, n4466);
   nand (n4468, n4236, n274);
   nand (n4469, n4467, n4468);
   nor (n447, n445, n446);
   xor (n4470, n4464, n4469);
   not (n4471, n4378);
   nand (n4472, n4379, n340);
   nand (n4473, n4471, n4472);
   not (n4474, n4473);
   nor (n4475, n4474, n4380);
   and (n4476, n4470, n4475);
   and (n4477, n4464, n4469);
   or (n4478, n4476, n4477);
   xor (n4479, n4453, n4478);
   and (n448, n396, n447);
   not (n4480, n4241);
   and (n4481, n4259, n4480);
   not (n4482, n4259);
   and (n4483, n4482, n4241);
   nor (n4484, n4481, n4483);
   not (n4485, n4484);
   and (n4486, n4479, n4485);
   and (n4487, n4453, n4478);
   nor (n4488, n4486, n4487);
   not (n4489, n4488);
   and (n449, n375, n395);
   xor (n4490, n4234, n4263);
   not (n4491, n4490);
   or (n4492, n4489, n4491);
   or (n4493, n4488, n4490);
   nand (n4494, n4492, n4493);
   not (n4495, n4494);
   or (n4496, n4448, n4495);
   not (n4497, n4488);
   nand (n4498, n4497, n4490);
   nand (n4499, n4496, n4498);
   buf (n45, g44);
   nor (n450, n448, n449);
   not (n4500, n4499);
   not (n4501, n4421);
   not (n4502, n4429);
   and (n4503, n4501, n4502);
   and (n4504, n4421, n4429);
   nor (n4505, n4503, n4504);
   nor (n4506, n4500, n4505);
   nand (n4507, n4445, n4506);
   not (n4508, n4507);
   and (n4509, n3318, n804);
   not (n451, n450);
   not (n4510, n4509);
   nand (n4511, n4510, n3170);
   not (n4512, n4511);
   not (n4513, n51);
   and (n4514, n50, n3440);
   not (n4515, n50);
   not (n4516, n3126);
   and (n4517, n4515, n4516);
   nor (n4518, n4514, n4517);
   not (n4519, n4518);
   not (n452, n451);
   or (n4520, n4513, n4519);
   and (n4521, n3289, n3334);
   nor (n4522, n4521, n1274);
   nand (n4523, n4520, n4522);
   not (n4524, n4523);
   or (n4525, n4512, n4524);
   not (n4526, n4511);
   not (n4527, n4523);
   nand (n4528, n4526, n4527);
   nand (n4529, n4525, n4528);
   or (n453, n374, n452);
   and (n4530, n3420, n3334);
   and (n4531, n3451, n1005);
   nor (n4532, n4530, n4531);
   and (n4533, n3288, n1829);
   nor (n4534, n4533, n1274);
   nand (n4535, n4532, n4534);
   not (n4536, n4535);
   not (n4537, n4510);
   and (n4538, n4536, n4537);
   and (n4539, n4535, n4509);
   xnor (n454, n396, n447);
   not (n4540, n4535);
   and (n4541, n4540, n4510);
   nor (n4542, n4539, n4541);
   not (n4543, n4542);
   not (n4544, n1075);
   not (n4545, n610);
   not (n4546, n3351);
   or (n4547, n4545, n4546);
   or (n4548, n3354, n610);
   nand (n4549, n4547, n4548);
   not (n455, n454);
   not (n4550, n4549);
   or (n4551, n4544, n4550);
   not (n4552, n48);
   not (n4553, n3431);
   or (n4554, n4552, n4553);
   not (n4555, n3431);
   not (n4556, n4555);
   or (n4557, n4556, n48);
   nand (n4558, n4554, n4557);
   nand (n4559, n4558, n1039);
   xor (n456, n437, n442);
   nand (n4560, n4551, n4559);
   and (n4561, n4543, n4560);
   nor (n4562, n4538, n4561);
   xor (n4563, n4529, n4562);
   not (n4564, n4563);
   not (n4565, n4564);
   not (n4566, n1944);
   not (n4567, n48);
   not (n4568, n3840);
   or (n4569, n4567, n4568);
   xor (n457, n456, n444);
   buf (n4570, n3419);
   or (n4571, n4570, n48);
   nand (n4572, n4569, n4571);
   not (n4573, n4572);
   or (n4574, n4566, n4573);
   not (n4575, n4558);
   or (n4576, n4575, n4220);
   nand (n4577, n4574, n4576);
   not (n4578, n4577);
   not (n4579, n3224);
   or (n458, n36, n59);
   not (n4580, n45);
   not (n4581, n4580);
   not (n4582, n3318);
   not (n4583, n4582);
   or (n4584, n4581, n4583);
   not (n4585, n4046);
   or (n4586, n4585, n504);
   nand (n4587, n4584, n4586);
   not (n4588, n4587);
   or (n4589, n4579, n4588);
   nand (n459, n458, n405);
   not (n4590, n412);
   not (n4591, n4061);
   or (n4592, n4590, n4591);
   or (n4593, n4061, n412);
   nand (n4594, n4592, n4593);
   nand (n4595, n4594, n805);
   nand (n4596, n4589, n4595);
   not (n4597, n815);
   not (n4598, n3765);
   not (n4599, n46);
   buf (n46, g45);
   or (n460, n247, n459);
   and (n4600, n4598, n4599);
   and (n4601, n3765, n46);
   nor (n4602, n4600, n4601);
   not (n4603, n4602);
   or (n4604, n4597, n4603);
   not (n4605, n4111);
   not (n4606, n504);
   or (n4607, n4605, n4606);
   nand (n4608, n4110, n46);
   nand (n4609, n4607, n4608);
   or (n461, n253, n398);
   nand (n4610, n4609, n3470);
   nand (n4611, n4604, n4610);
   and (n4612, n4596, n4611);
   not (n4613, n4596);
   not (n4614, n4611);
   and (n4615, n4613, n4614);
   nor (n4616, n4612, n4615);
   not (n4617, n4616);
   not (n4618, n4617);
   or (n4619, n4578, n4618);
   nand (n462, n460, n461);
   not (n4620, n4577);
   nand (n4621, n4620, n4616);
   nand (n4622, n4619, n4621);
   not (n4623, n4622);
   and (n4624, n4565, n4623);
   and (n4625, n4529, n4562);
   nor (n4626, n4624, n4625);
   not (n4627, n4626);
   not (n4628, n4627);
   not (n4629, n3471);
   not (n463, n462);
   not (n4630, n4602);
   or (n4631, n4629, n4630);
   and (n4632, n46, n3665);
   not (n4633, n46);
   and (n4634, n4633, n3434);
   or (n4635, n4632, n4634);
   nand (n4636, n4635, n1151);
   nand (n4637, n4631, n4636);
   not (n4638, n1075);
   and (n4639, n49, n4213);
   nand (n464, n36, n60);
   not (n4640, n49);
   and (n4641, n4640, n3836);
   nor (n4642, n4639, n4641);
   not (n4643, n4642);
   or (n4644, n4638, n4643);
   not (n4645, n1038);
   not (n4646, n48);
   not (n4647, n3451);
   or (n4648, n4646, n4647);
   or (n4649, n3457, n48);
   not (n465, n266);
   nand (n4650, n4648, n4649);
   nand (n4651, n4645, n4650);
   nand (n4652, n4644, n4651);
   xor (n4653, n4637, n4652);
   not (n4654, n4528);
   xor (n4655, n4653, n4654);
   not (n4656, n4655);
   not (n4657, n805);
   not (n4658, n412);
   not (n4659, n3737);
   and (n466, n40, n55);
   or (n4660, n4658, n4659);
   nand (n4661, n3363, n44);
   nand (n4662, n4660, n4661);
   not (n4663, n4662);
   or (n4664, n4657, n4663);
   nand (n4665, n4594, n3224);
   nand (n4666, n4664, n4665);
   not (n4667, n4582);
   nand (n4668, n4667, n1259);
   not (n4669, n4668);
   nor (n467, n40, n55);
   not (n4670, n4669);
   not (n4671, n4670);
   not (n4672, n3510);
   or (n4673, n4672, n1480);
   not (n4674, n1005);
   not (n4675, n3065);
   or (n4676, n4674, n4675);
   not (n4677, n1274);
   nand (n4678, n4676, n4677);
   not (n4679, n4678);
   nor (n468, n466, n467);
   nand (n4680, n3237, n3334);
   nand (n4681, n4673, n4679, n4680);
   not (n4682, n4681);
   not (n4683, n4682);
   or (n4684, n4671, n4683);
   nand (n4685, n4681, n4669);
   nand (n4686, n4684, n4685);
   xor (n4687, n4666, n4686);
   not (n4688, n4687);
   not (n4689, n4577);
   and (n469, n465, n468);
   not (n4690, n4616);
   or (n4691, n4689, n4690);
   nand (n4692, n4611, n4596);
   nand (n4693, n4691, n4692);
   not (n4694, n4693);
   not (n4695, n4694);
   or (n4696, n4688, n4695);
   not (n4697, n4687);
   nand (n4698, n4697, n4693);
   nand (n4699, n4696, n4698);
   buf (n47, g46);
   and (n470, n274, n389);
   not (n4700, n4699);
   or (n4701, n4656, n4700);
   or (n4702, n4699, n4655);
   nand (n4703, n4701, n4702);
   not (n4704, n4703);
   not (n4705, n4704);
   or (n4706, n4628, n4705);
   nand (n4707, n4703, n4626);
   nand (n4708, n4706, n4707);
   not (n4709, n4708);
   nor (n471, n469, n470);
   not (n4710, n4111);
   not (n4711, n3533);
   or (n4712, n4710, n4711);
   nand (n4713, n3363, n48);
   nand (n4714, n4712, n4713);
   and (n4715, n4714, n1944);
   not (n4716, n1779);
   not (n4717, n3493);
   not (n4718, n3533);
   and (n4719, n4717, n4718);
   xor (n472, n464, n471);
   and (n4720, n3493, n3533);
   nor (n4721, n4719, n4720);
   nor (n4722, n4716, n4721);
   nor (n4723, n4715, n4722);
   not (n4724, n4723);
   not (n4725, n4724);
   nand (n4726, n3318, n814);
   not (n4727, n4726);
   not (n4728, n4727);
   not (n4729, n4728);
   not (n473, n472);
   not (n4730, n3334);
   not (n4731, n3765);
   or (n4732, n4730, n4731);
   nand (n4733, n4556, n1005);
   nand (n4734, n4732, n4733);
   not (n4735, n1270);
   not (n4736, n4347);
   or (n4737, n4735, n4736);
   nand (n4738, n4737, n4677);
   nor (n4739, n4734, n4738);
   or (n474, n463, n473);
   not (n4740, n4739);
   or (n4741, n4729, n4740);
   or (n4742, n4728, n4739);
   nand (n4743, n4741, n4742);
   not (n4744, n4743);
   or (n4745, n4725, n4744);
   not (n4746, n4728);
   nand (n4747, n4746, n4739);
   nand (n4748, n4745, n4747);
   not (n4749, n4748);
   or (n475, n471, n464);
   not (n4750, n51);
   not (n4751, n50);
   and (n4752, n3, n14);
   not (n4753, n3);
   and (n4754, n4753, n30);
   nor (n4755, n4752, n4754);
   not (n4756, n4755);
   not (n4757, n4756);
   or (n4758, n4751, n4757);
   or (n4759, n3839, n50);
   nand (n476, n474, n475);
   nand (n4760, n4758, n4759);
   not (n4761, n4760);
   or (n4762, n4750, n4761);
   not (n4763, n3334);
   not (n4764, n4555);
   or (n4765, n4763, n4764);
   nand (n4766, n4765, n4677);
   not (n4767, n4766);
   nand (n4768, n4762, n4767);
   nand (n4769, n4726, n2369);
   and (n477, n38, n56);
   nor (n4770, n4768, n4769);
   not (n4771, n4770);
   nand (n4772, n4768, n4769);
   nand (n4773, n4771, n4772);
   not (n4774, n4773);
   not (n4775, n3470);
   xor (n4776, n3500, n48);
   not (n4777, n4776);
   or (n4778, n4775, n4777);
   not (n4779, n504);
   not (n478, n38);
   not (n4780, n3493);
   or (n4781, n4779, n4780);
   or (n4782, n3493, n504);
   nand (n4783, n4781, n4782);
   nand (n4784, n542, n4783);
   nand (n4785, n4778, n4784);
   not (n4786, n1039);
   not (n4787, n3765);
   not (n4788, n48);
   and (n4789, n4787, n4788);
   not (n479, n56);
   and (n4790, n3765, n48);
   nor (n4791, n4789, n4790);
   not (n4792, n4791);
   or (n4793, n4786, n4792);
   nand (n4794, n4714, n3693);
   nand (n4795, n4793, n4794);
   xor (n4796, n4785, n4795);
   not (n4797, n4796);
   or (n4798, n4774, n4797);
   or (n4799, n4796, n4773);
   buf (n48, g47);
   and (n480, n478, n479);
   nand (n4800, n4798, n4799);
   not (n4801, n4800);
   or (n4802, n4749, n4801);
   not (n4803, n4723);
   not (n4804, n4743);
   or (n4805, n4803, n4804);
   or (n4806, n4723, n4743);
   nand (n4807, n4805, n4806);
   not (n4808, n616);
   nor (n4809, n3501, n3692);
   nor (n481, n477, n480);
   nor (n4810, n4808, n4809);
   not (n4811, n1574);
   not (n4812, n3351);
   or (n4813, n4811, n4812);
   not (n4814, n3);
   nand (n4815, n4814, n3762);
   nand (n4816, n3759, n3);
   and (n4817, n1832, n4815, n4816);
   and (n4818, n3363, n1473);
   nor (n4819, n4817, n4818);
   not (n482, n481);
   nand (n4820, n4813, n4819);
   nand (n4821, n4810, n4820);
   buf (n4822, n4821);
   not (n4823, n4822);
   nand (n4824, n4807, n4823);
   nand (n4825, n4802, n4824);
   not (n4826, n4825);
   not (n4827, n4773);
   and (n4828, n4827, n4796);
   and (n4829, n4785, n4795);
   not (n483, n297);
   nor (n4830, n4828, n4829);
   not (n4831, n4830);
   not (n4832, n542);
   not (n4833, n4609);
   or (n4834, n4832, n4833);
   nand (n4835, n4783, n3470);
   nand (n4836, n4834, n4835);
   xor (n4837, n4770, n4836);
   not (n4838, n4837);
   not (n4839, n4560);
   or (n484, n482, n483);
   not (n4840, n4542);
   and (n4841, n4839, n4840);
   and (n4842, n4542, n4560);
   nor (n4843, n4841, n4842);
   not (n4844, n4843);
   or (n4845, n4838, n4844);
   or (n4846, n4843, n4837);
   nand (n4847, n4845, n4846);
   buf (n4848, n4847);
   nand (n4849, n4831, n4848);
   nand (n485, n311, n380);
   nand (n4850, n4826, n4849);
   xnor (n4851, n4622, n4563);
   not (n4852, n4843);
   nand (n4853, n4852, n4837);
   nand (n4854, n4770, n4836);
   and (n4855, n4853, n4854);
   nor (n4856, n4851, n4855);
   nor (n4857, n4810, n4820);
   not (n4858, n4857);
   nand (n4859, n4858, n4821);
   nand (n486, n484, n485);
   not (n4860, n4859);
   not (n4861, n4860);
   not (n4862, n3693);
   not (n4863, n4776);
   not (n4864, n4863);
   or (n4865, n4862, n4864);
   or (n4866, n4721, n1038);
   nand (n4867, n4865, n4866);
   not (n4868, n4867);
   or (n4869, n4861, n4868);
   and (n487, n486, n392);
   not (n4870, n4867);
   not (n4871, n4859);
   or (n4872, n4870, n4871);
   or (n4873, n4859, n4867);
   nand (n4874, n4872, n4873);
   nand (n4875, n3737, n51);
   or (n4876, n3501, n1480);
   nand (n4877, n3495, n50);
   nand (n4878, n4876, n4877);
   and (n4879, n4878, n1944);
   not (n488, n486);
   nor (n4880, n4047, n4877);
   nor (n4881, n4879, n4880);
   and (n4882, n4875, n4881);
   not (n4883, n4875);
   nand (n4884, n4047, n1944, n1005);
   and (n4885, n4883, n4884);
   nor (n4886, n4882, n4885);
   nand (n4887, n4874, n4886);
   nand (n4888, n4869, n4887);
   not (n4889, n4822);
   and (n489, n488, n438);
   not (n4890, n4807);
   or (n4891, n4889, n4890);
   or (n4892, n4822, n4807);
   nand (n4893, n4891, n4892);
   nand (n4894, n4888, n4893);
   not (n4895, n4894);
   nor (n4896, n4850, n4856, n4895);
   not (n4897, n4800);
   not (n4898, n4748);
   nand (n4899, n4897, n4898);
   buf (n49, g48);
   nor (n490, n487, n489);
   not (n4900, n4899);
   not (n4901, n4830);
   not (n4902, n4847);
   or (n4903, n4901, n4902);
   or (n4904, n4830, n4847);
   nand (n4905, n4903, n4904);
   not (n4906, n4905);
   or (n4907, n4900, n4906);
   nand (n4908, n4907, n4849);
   or (n4909, n4908, n4856);
   and (n491, n476, n490);
   nand (n4910, n4851, n4855);
   nand (n4911, n4909, n4910);
   nor (n4912, n4896, n4911);
   not (n4913, n4912);
   or (n4914, n4709, n4913);
   not (n4915, n4654);
   not (n4916, n4653);
   or (n4917, n4915, n4916);
   nand (n4918, n4637, n4652);
   nand (n4919, n4917, n4918);
   and (n492, n486, n392);
   not (n4920, n805);
   not (n4921, n3354);
   not (n4922, n412);
   and (n4923, n4921, n4922);
   buf (n4924, n4076);
   and (n4925, n4924, n412);
   nor (n4926, n4923, n4925);
   not (n4927, n4926);
   or (n4928, n4920, n4927);
   nand (n4929, n4662, n3224);
   nor (n493, n491, n492);
   nand (n4930, n4928, n4929);
   not (n4931, n4930);
   not (n4932, n4931);
   not (n4933, n3522);
   not (n4934, n1005);
   and (n4935, n4933, n4934);
   and (n4936, n3070, n1005);
   nor (n4937, n4935, n4936);
   and (n4938, n4937, n51);
   not (n4939, n3334);
   xor (n494, n457, n493);
   not (n4940, n3510);
   or (n4941, n4939, n4940);
   nand (n4942, n4941, n4677);
   nor (n4943, n4938, n4942);
   not (n4944, n43);
   and (n4945, n4944, n3318);
   not (n4946, n4944);
   and (n4947, n4946, n3500);
   or (n4948, n4945, n4947);
   nor (n4949, n4948, n736);
   not (n495, n296);
   not (n4950, n423);
   not (n4951, n4061);
   or (n4952, n4950, n4951);
   or (n4953, n4061, n423);
   nand (n4954, n4952, n4953);
   and (n4955, n4954, n513);
   or (n4956, n4949, n4955);
   and (n4957, n4943, n4956);
   not (n4958, n4943);
   nor (n4959, n4949, n4955);
   and (n496, n38, n57);
   and (n4960, n4958, n4959);
   nor (n4961, n4957, n4960);
   not (n4962, n4961);
   or (n4963, n4932, n4962);
   or (n4964, n4931, n4961);
   nand (n4965, n4963, n4964);
   xor (n4966, n4919, n4965);
   nand (n4967, n4635, n3471);
   not (n4968, n46);
   not (n4969, n4755);
   not (n497, n38);
   or (n4970, n4968, n4969);
   or (n4971, n3419, n46);
   nand (n4972, n4970, n4971);
   nand (n4973, n4972, n1151);
   and (n4974, n4967, n4973);
   not (n4975, n4974);
   nand (n4976, n4668, n352);
   not (n4977, n4976);
   not (n4978, n614);
   not (n4979, n3533);
   not (n498, n57);
   not (n4980, n3237);
   or (n4981, n4979, n4980);
   or (n4982, n3533, n3237);
   nand (n4983, n4981, n4982);
   not (n4984, n4983);
   or (n4985, n4978, n4984);
   nand (n4986, n4650, n1075);
   nand (n4987, n4985, n4986);
   not (n4988, n4987);
   not (n4989, n4988);
   and (n499, n497, n498);
   or (n4990, n4977, n4989);
   not (n4991, n4976);
   nand (n4992, n4991, n4987);
   nand (n4993, n4990, n4992);
   not (n4994, n4993);
   not (n4995, n4994);
   or (n4996, n4975, n4995);
   not (n4997, n4993);
   or (n4998, n4997, n4974);
   nand (n4999, n4996, n4998);
   buf (n5, g4);
   buf (n50, g49);
   nor (n500, n496, n499);
   not (n5000, n4666);
   not (n5001, n4686);
   or (n5002, n5000, n5001);
   not (n5003, n4670);
   nand (n5004, n5003, n4682);
   nand (n5005, n5002, n5004);
   not (n5006, n5005);
   and (n5007, n4999, n5006);
   not (n5008, n4999);
   and (n5009, n5008, n5005);
   and (n501, n495, n500);
   nor (n5010, n5007, n5009);
   nor (n5011, n4966, n5010);
   not (n5012, n5011);
   nand (n5013, n5010, n4966);
   nand (n5014, n5012, n5013);
   not (n5015, n4655);
   nand (n5016, n5015, n4699);
   not (n5017, n4687);
   nand (n5018, n5017, n4694);
   nand (n5019, n5016, n5018);
   and (n502, n311, n481);
   not (n5020, n5019);
   and (n5021, n5014, n5020);
   not (n5022, n4703);
   and (n5023, n5022, n4626);
   nor (n5024, n5021, n5023);
   nand (n5025, n4914, n5024);
   not (n5026, n4966);
   not (n5027, n5010);
   not (n5028, n5027);
   or (n5029, n5026, n5028);
   nor (n503, n501, n502);
   nand (n5030, n4919, n4965);
   nand (n5031, n5029, n5030);
   buf (n5032, n4992);
   not (n5033, n1779);
   not (n5034, n4983);
   or (n5035, n5033, n5034);
   nand (n5036, n4376, n614);
   nand (n5037, n5035, n5036);
   not (n5038, n5037);
   not (n5039, n4379);
   not (n504, n46);
   and (n5040, n5038, n5039);
   and (n5041, n5037, n4379);
   nor (n5042, n5040, n5041);
   not (n5043, n5042);
   not (n5044, n4351);
   not (n5045, n556);
   and (n5046, n5044, n5045);
   and (n5047, n4926, n3224);
   nor (n5048, n5046, n5047);
   not (n5049, n5048);
   and (n505, n504, n45);
   and (n5050, n5043, n5049);
   not (n5051, n5042);
   not (n5052, n5051);
   and (n5053, n5052, n5048);
   nor (n5054, n5050, n5053);
   xor (n5055, n5032, n5054);
   not (n5056, n4930);
   not (n5057, n4961);
   or (n5058, n5056, n5057);
   not (n5059, n4959);
   nor (n506, n505, n412);
   nand (n5060, n5059, n4943);
   nand (n5061, n5058, n5060);
   xnor (n5062, n5055, n5061);
   not (n5063, n513);
   not (n5064, n4336);
   or (n5065, n5063, n5064);
   nand (n5066, n1746, n4954);
   nand (n5067, n5065, n5066);
   not (n5068, n3470);
   not (n5069, n4972);
   xor (n507, n503, n506);
   or (n5070, n5068, n5069);
   nand (n5071, n4455, n815);
   nand (n5072, n5070, n5071);
   xor (n5073, n5067, n5072);
   not (n5074, n1956);
   not (n5075, n3071);
   or (n5076, n5074, n5075);
   and (n5077, n1477, n2923);
   and (n5078, n2991, n1574);
   nor (n5079, n5077, n5078);
   and (n508, n423, n312);
   nand (n5080, n5076, n5079);
   xor (n5081, n5073, n5080);
   not (n5082, n5005);
   not (n5083, n4999);
   or (n5084, n5082, n5083);
   not (n5085, n4974);
   nand (n5086, n5085, n4997);
   nand (n5087, n5084, n5086);
   xor (n5088, n5081, n5087);
   xor (n5089, n5062, n5088);
   and (n509, n42, n53);
   xor (n5090, n5031, n5089);
   not (n5091, n5014);
   not (n5092, n5019);
   and (n5093, n5091, n5092);
   and (n5094, n5014, n5019);
   nor (n5095, n5093, n5094);
   nand (n5096, n5020, n5014);
   nand (n5097, n5095, n5096);
   nand (n5098, n5025, n5090, n5097);
   not (n5099, n5098);
   buf (n51, g50);
   nor (n510, n508, n509);
   xor (n5100, n4464, n4469);
   xor (n5101, n5100, n4475);
   not (n5102, n5054);
   nand (n5103, n5102, n5032);
   not (n5104, n5103);
   not (n5105, n5061);
   or (n5106, n5104, n5105);
   not (n5107, n5032);
   nand (n5108, n5107, n5054);
   nand (n5109, n5106, n5108);
   and (n511, n422, n510);
   xor (n5110, n5101, n5109);
   xor (n5111, n4331, n4354);
   xnor (n5112, n5111, n4338);
   not (n5113, n5112);
   not (n5114, n5113);
   not (n5115, n5080);
   not (n5116, n5073);
   or (n5117, n5115, n5116);
   nand (n5118, n5067, n5072);
   nand (n5119, n5117, n5118);
   not (n512, n428);
   not (n5120, n5119);
   not (n5121, n5048);
   not (n5122, n5051);
   or (n5123, n5121, n5122);
   not (n5124, n5037);
   nand (n5125, n5124, n4379);
   nand (n5126, n5123, n5125);
   not (n5127, n5126);
   nand (n5128, n5120, n5127);
   nand (n5129, n5119, n5126);
   not (n513, n512);
   nand (n5130, n5128, n5129);
   not (n5131, n5130);
   and (n5132, n5114, n5131);
   buf (n5133, n5130);
   and (n5134, n5133, n5113);
   nor (n5135, n5132, n5134);
   xnor (n5136, n5110, n5135);
   not (n5137, n5062);
   not (n5138, n5088);
   or (n5139, n5137, n5138);
   not (n514, n513);
   nand (n5140, n5087, n5081);
   nand (n5141, n5139, n5140);
   nand (n5142, n5136, n5141);
   nand (n5143, n5089, n5031);
   nand (n5144, n5142, n5143);
   xnor (n5145, n4359, n4391);
   not (n5146, n5145);
   not (n5147, n5112);
   not (n5148, n5130);
   or (n5149, n5147, n5148);
   not (n515, n514);
   nand (n5150, n5127, n5119);
   nand (n5151, n5149, n5150);
   not (n5152, n5151);
   or (n5153, n5146, n5152);
   or (n5154, n5145, n5151);
   nand (n5155, n5153, n5154);
   not (n5156, n5155);
   xor (n5157, n4479, n4484);
   not (n5158, n5157);
   and (n5159, n5156, n5158);
   and (n516, n515, n426);
   and (n5160, n5155, n5157);
   nor (n5161, n5159, n5160);
   not (n5162, n5135);
   and (n5163, n5162, n5110);
   and (n5164, n5101, n5109);
   nor (n5165, n5163, n5164);
   nor (n5166, n5161, n5165);
   nor (n5167, n5144, n5166);
   not (n5168, n5167);
   or (n5169, n5099, n5168);
   nor (n517, n511, n516);
   not (n5170, n5166);
   nor (n5171, n5136, n5141);
   and (n5172, n5170, n5171);
   not (n5173, n5161);
   not (n5174, n5165);
   nor (n5175, n5173, n5174);
   nor (n5176, n5172, n5175);
   nand (n5177, n5169, n5176);
   not (n5178, n5157);
   not (n5179, n5178);
   and (n518, n507, n517);
   not (n5180, n5155);
   or (n5181, n5179, n5180);
   not (n5182, n5145);
   nand (n5183, n5182, n5151);
   nand (n5184, n5181, n5183);
   not (n5185, n4446);
   not (n5186, n4494);
   or (n5187, n5185, n5186);
   or (n5188, n4494, n4446);
   nand (n5189, n5187, n5188);
   and (n519, n503, n506);
   xnor (n5190, n5184, n5189);
   nor (n5191, n5177, n5190);
   not (n5192, n4505);
   not (n5193, n4499);
   and (n5194, n5192, n5193);
   and (n5195, n4505, n4499);
   nor (n5196, n5194, n5195);
   not (n5197, n5196);
   nand (n5198, n5191, n5197);
   not (n5199, n5198);
   buf (n52, g51);
   nor (n520, n518, n519);
   or (n5200, n4508, n5199);
   buf (n5201, n4445);
   nand (n5202, n5200, n5201);
   nor (n5203, n4313, n5202);
   not (n5204, n5203);
   nand (n5205, n5184, n5189);
   nor (n5206, n5196, n5205);
   buf (n5207, n5206);
   and (n5208, n5201, n5207);
   not (n5209, n4302);
   xor (n521, n433, n410);
   not (n5210, n4441);
   nand (n5211, n5210, n4435);
   nand (n5212, n5209, n5211);
   nor (n5213, n5208, n5212);
   nand (n5214, n4312, n4037);
   nor (n5215, n5213, n5214);
   not (n5216, n4304);
   not (n5217, n4310);
   nor (n5218, n5216, n5217);
   not (n5219, n5218);
   xor (n522, n520, n521);
   not (n5220, n4037);
   or (n5221, n5219, n5220);
   nand (n5222, n4033, n3885);
   nand (n5223, n5221, n5222);
   nor (n5224, n5215, n5223);
   nand (n5225, n5204, n5224);
   not (n5226, n4028);
   and (n5227, n5226, n3955);
   and (n5228, n3948, n3954);
   nor (n5229, n5227, n5228);
   xor (n523, n476, n490);
   not (n5230, n376);
   not (n5231, n3974);
   or (n5232, n5230, n5231);
   not (n5233, n38);
   not (n5234, n3239);
   or (n5235, n5233, n5234);
   or (n5236, n3239, n38);
   nand (n5237, n5235, n5236);
   nand (n5238, n5237, n310);
   nand (n5239, n5232, n5238);
   and (n524, n522, n523);
   xor (n5240, n3923, n5239);
   not (n5241, n2848);
   not (n5242, n3931);
   or (n5243, n5241, n5242);
   nand (n5244, n3840, n2762);
   not (n5245, n5244);
   not (n5246, n3420);
   nor (n5247, n5246, n2762);
   nor (n5248, n5245, n5247);
   nand (n5249, n2861, n5248);
   and (n525, n520, n521);
   nand (n5250, n5243, n5249);
   xor (n5251, n5240, n5250);
   not (n5252, n3851);
   nand (n5253, n3933, n3923);
   not (n5254, n5253);
   or (n5255, n5252, n5254);
   not (n5256, n3933);
   nand (n5257, n5256, n3924);
   nand (n5258, n5255, n5257);
   not (n5259, n274);
   nor (n526, n524, n525);
   not (n5260, n40);
   not (n5261, n3070);
   not (n5262, n5261);
   or (n5263, n5260, n5262);
   or (n5264, n3204, n40);
   nand (n5265, n5263, n5264);
   not (n5266, n5265);
   or (n5267, n5259, n5266);
   nand (n5268, n362, n3983);
   nand (n5269, n5267, n5268);
   and (n527, n494, n526);
   buf (n5270, n3769);
   xor (n5271, n5269, n5270);
   and (n5272, n3386, n412);
   not (n5273, n3386);
   and (n5274, n5273, n44);
   nor (n5275, n5272, n5274);
   not (n5276, n5275);
   not (n5277, n556);
   and (n5278, n5276, n5277);
   and (n5279, n3962, n3224);
   and (n528, n457, n493);
   nor (n5280, n5278, n5279);
   xnor (n5281, n5271, n5280);
   not (n5282, n5281);
   xor (n5283, n5258, n5282);
   xnor (n5284, n5251, n5283);
   not (n5285, n5284);
   not (n5286, n4023);
   not (n5287, n4018);
   or (n5288, n5286, n5287);
   not (n5289, n4005);
   nor (n529, n527, n528);
   xor (n5290, n3994, n4017);
   nand (n5291, n5289, n5290);
   nand (n5292, n5288, n5291);
   not (n5293, n5292);
   or (n5294, n5285, n5293);
   or (n5295, n5284, n5292);
   nand (n5296, n5294, n5295);
   or (n5297, n3990, n3964);
   not (n5298, n3976);
   or (n5299, n5298, n3985);
   buf (n53, g52);
   nand (n530, n455, n529);
   nand (n5300, n5297, n5299);
   not (n5301, n5300);
   not (n5302, n421);
   or (n5303, n3910, n5302);
   and (n5304, n2907, n42);
   not (n5305, n2907);
   and (n5306, n5305, n423);
   nor (n5307, n5304, n5306);
   or (n5308, n5307, n514);
   nand (n5309, n5303, n5308);
   not (n531, n530);
   not (n5310, n3897);
   not (n5311, n3469);
   and (n5312, n5310, n5311);
   not (n5313, n504);
   not (n5314, n2831);
   or (n5315, n5313, n5314);
   not (n5316, n3327);
   nand (n5317, n5316, n46);
   nand (n5318, n5315, n5317);
   nor (n5319, n5318, n627);
   xor (n532, n46, n47);
   nor (n5320, n5312, n5319);
   and (n5321, n5320, n616);
   not (n5322, n5320);
   and (n5323, n5322, n619);
   nor (n5324, n5321, n5323);
   xor (n5325, n5309, n5324);
   not (n5326, n3912);
   not (n5327, n3905);
   or (n5328, n5326, n5327);
   nand (n5329, n3900, n3901);
   xor (n533, n47, n48);
   nand (n5330, n5328, n5329);
   xor (n5331, n5325, n5330);
   not (n5332, n5331);
   not (n5333, n5332);
   or (n5334, n5301, n5333);
   not (n5335, n5300);
   nand (n5336, n5335, n5331);
   nand (n5337, n5334, n5336);
   not (n5338, n3994);
   not (n5339, n4017);
   nand (n534, n532, n533);
   or (n5340, n5338, n5339);
   nand (n5341, n4010, n4016);
   nand (n5342, n5340, n5341);
   xor (n5343, n5337, n5342);
   not (n5344, n3940);
   not (n5345, n3947);
   or (n5346, n5344, n5345);
   not (n5347, n3935);
   nand (n5348, n5347, n3913);
   nand (n5349, n5346, n5348);
   not (n535, n534);
   xor (n5350, n5343, n5349);
   not (n5351, n5350);
   and (n5352, n5296, n5351);
   not (n5353, n5296);
   and (n5354, n5353, n5350);
   nor (n5355, n5352, n5354);
   xor (n5356, n5229, n5355);
   nand (n5357, n5225, n5356);
   or (n5358, n5275, n3590);
   not (n5359, n2855);
   and (n536, n504, n267);
   not (n5360, n412);
   and (n5361, n5359, n5360);
   and (n5362, n2855, n412);
   nor (n5363, n5361, n5362);
   or (n5364, n5363, n556);
   nand (n5365, n5358, n5364);
   not (n5366, n5365);
   not (n5367, n465);
   not (n5368, n5265);
   or (n5369, n5367, n5368);
   and (n537, n46, n52);
   and (n5370, n40, n2991);
   not (n5371, n40);
   and (n5372, n5371, n2923);
   or (n5373, n5370, n5372);
   nand (n5374, n5373, n274);
   nand (n5375, n5369, n5374);
   not (n5376, n376);
   not (n5377, n5237);
   or (n5378, n5376, n5377);
   and (n5379, n38, n3066);
   nor (n538, n536, n537);
   not (n5380, n38);
   and (n5381, n5380, n3067);
   or (n5382, n5379, n5381);
   nand (n5383, n5382, n310);
   nand (n5384, n5378, n5383);
   xor (n5385, n5375, n5384);
   not (n5386, n5385);
   or (n5387, n5366, n5386);
   nand (n5388, n5384, n5375);
   nand (n5389, n5387, n5388);
   and (n539, n535, n538);
   not (n5390, n5389);
   not (n5391, n5247);
   not (n5392, n5318);
   nand (n5393, n5392, n3471);
   and (n5394, n5393, n816);
   not (n5395, n5394);
   and (n5396, n5391, n5395);
   not (n5397, n5391);
   and (n5398, n5397, n5394);
   nor (n5399, n5396, n5398);
   buf (n54, g53);
   not (n540, n533);
   or (n5400, n5390, n5399);
   or (n5401, n5394, n5391);
   nand (n5402, n5400, n5401);
   xor (n5403, n3294, n3299);
   xor (n5404, n5402, n5403);
   not (n5405, n805);
   not (n5406, n3216);
   or (n5407, n5405, n5406);
   not (n5408, n5363);
   nand (n5409, n5408, n3224);
   not (n541, n540);
   nand (n5410, n5407, n5409);
   xnor (n5411, n5410, n2369);
   not (n5412, n5373);
   not (n5413, n465);
   or (n5414, n5412, n5413);
   or (n5415, n3295, n275);
   nand (n5416, n5414, n5415);
   xor (n5417, n5411, n5416);
   not (n5418, n5417);
   not (n5419, n401);
   buf (n542, n541);
   xor (n5420, n36, n3289);
   not (n5421, n5420);
   or (n5422, n5419, n5421);
   not (n5423, n4213);
   not (n5424, n37);
   and (n5425, n5423, n5424);
   and (n5426, n4570, n37);
   nor (n5427, n5425, n5426);
   nand (n5428, n5427, n2848);
   nand (n5429, n5422, n5428);
   not (n543, n542);
   xor (n5430, n3930, n5429);
   not (n5431, n737);
   not (n5432, n5307);
   and (n5433, n5431, n5432);
   not (n5434, n2868);
   not (n5435, n42);
   and (n5436, n5434, n5435);
   and (n5437, n3112, n42);
   nor (n5438, n5436, n5437);
   and (n5439, n5438, n515);
   and (n544, n543, n46);
   nor (n5440, n5433, n5439);
   not (n5441, n5440);
   and (n5442, n5430, n5441);
   and (n5443, n3930, n5429);
   nor (n5444, n5442, n5443);
   not (n5445, n5444);
   not (n5446, n5445);
   or (n5447, n5418, n5446);
   and (n5448, n5438, n421);
   and (n5449, n3264, n1259);
   nor (n545, n539, n544);
   nor (n5450, n5448, n5449);
   not (n5451, n5450);
   not (n5452, n297);
   not (n5453, n5382);
   or (n5454, n5452, n5453);
   nand (n5455, n3209, n311);
   nand (n5456, n5454, n5455);
   not (n5457, n5456);
   and (n5458, n5451, n5457);
   and (n5459, n5456, n5450);
   and (n546, n44, n54);
   nor (n5460, n5458, n5459);
   not (n5461, n3127);
   not (n5462, n2762);
   or (n5463, n5461, n5462);
   nand (n5464, n5463, n3129);
   not (n5465, n5464);
   not (n5466, n253);
   and (n5467, n5465, n5466);
   and (n5468, n5420, n2848);
   nor (n5469, n5467, n5468);
   not (n547, n44);
   xnor (n5470, n5460, n5469);
   not (n5471, n5470);
   not (n5472, n5444);
   not (n5473, n5417);
   or (n5474, n5472, n5473);
   or (n5475, n5444, n5417);
   nand (n5476, n5474, n5475);
   nand (n5477, n5471, n5476);
   nand (n5478, n5447, n5477);
   not (n5479, n5478);
   and (n548, n547, n299);
   xor (n5480, n5404, n5479);
   not (n5481, n5480);
   not (n5482, n5481);
   not (n5483, n5365);
   and (n5484, n5385, n5483);
   not (n5485, n5385);
   and (n5486, n5485, n5365);
   nor (n5487, n5484, n5486);
   not (n5488, n5487);
   and (n5489, n5240, n5250);
   nor (n549, n546, n548);
   and (n5490, n3923, n5239);
   nor (n5491, n5489, n5490);
   not (n5492, n5491);
   not (n5493, n5440);
   not (n5494, n5430);
   or (n5495, n5493, n5494);
   or (n5496, n5430, n5440);
   nand (n5497, n5495, n5496);
   not (n5498, n5497);
   or (n5499, n5492, n5498);
   buf (n55, g54);
   not (n550, n549);
   or (n5500, n5497, n5491);
   nand (n5501, n5499, n5500);
   nand (n5502, n5488, n5501);
   not (n5503, n5491);
   nand (n5504, n5503, n5497);
   and (n5505, n5502, n5504);
   not (n5506, n5505);
   not (n5507, n5506);
   not (n5508, n5399);
   not (n5509, n5389);
   not (n551, n46);
   or (n5510, n5508, n5509);
   or (n5511, n5389, n5399);
   nand (n5512, n5510, n5511);
   not (n5513, n5512);
   or (n5514, n5271, n5280);
   not (n5515, n5269);
   or (n5516, n5515, n5270);
   nand (n5517, n5514, n5516);
   not (n5518, n5517);
   not (n5519, n5309);
   not (n552, n45);
   not (n5520, n5324);
   or (n5521, n5519, n5520);
   not (n5522, n5320);
   nand (n5523, n5522, n619);
   nand (n5524, n5521, n5523);
   and (n5525, n5394, n5524);
   not (n5526, n5394);
   not (n5527, n5524);
   and (n5528, n5526, n5527);
   nor (n5529, n5525, n5528);
   or (n553, n551, n552);
   not (n5530, n5529);
   or (n5531, n5518, n5530);
   not (n5532, n5527);
   nand (n5533, n5532, n5394);
   nand (n5534, n5531, n5533);
   not (n5535, n5534);
   not (n5536, n5535);
   or (n5537, n5513, n5536);
   not (n5538, n5512);
   nand (n5539, n5538, n5534);
   or (n554, n45, n46);
   nand (n5540, n5537, n5539);
   not (n5541, n5540);
   or (n5542, n5507, n5541);
   nand (n5543, n5534, n5512);
   nand (n5544, n5542, n5543);
   not (n5545, n5544);
   or (n5546, n5460, n5469);
   not (n5547, n5456);
   or (n5548, n5547, n5450);
   nand (n5549, n5546, n5548);
   nand (n555, n553, n554);
   not (n5550, n5549);
   not (n5551, n5410);
   not (n5552, n5551);
   not (n5553, n2369);
   and (n5554, n5552, n5553);
   and (n5555, n5411, n5416);
   nor (n5556, n5554, n5555);
   not (n5557, n5556);
   or (n5558, n5550, n5557);
   or (n5559, n5556, n5549);
   buf (n556, n555);
   nand (n5560, n5558, n5559);
   xor (n5561, n3250, n3214);
   not (n5562, n5561);
   and (n5563, n5560, n5562);
   not (n5564, n5560);
   and (n5565, n5564, n5561);
   nor (n5566, n5563, n5565);
   and (n5567, n5545, n5566);
   not (n5568, n5545);
   not (n5569, n5566);
   not (n557, n556);
   and (n5570, n5568, n5569);
   nor (n5571, n5567, n5570);
   not (n5572, n5571);
   or (n5573, n5482, n5572);
   or (n5574, n5545, n5566);
   nand (n5575, n5573, n5574);
   not (n5576, n3303);
   and (n5577, n3283, n5576);
   not (n5578, n3283);
   and (n5579, n5578, n3303);
   or (n558, n550, n557);
   nor (n5580, n5577, n5579);
   and (n5581, n5560, n5561);
   not (n5582, n5556);
   and (n5583, n5582, n5549);
   nor (n5584, n5581, n5583);
   not (n5585, n5584);
   and (n5586, n5580, n5585);
   not (n5587, n5580);
   and (n5588, n5587, n5584);
   nor (n5589, n5586, n5588);
   not (n559, n45);
   and (n5590, n5478, n5404);
   and (n5591, n5402, n5403);
   nor (n5592, n5590, n5591);
   and (n5593, n5589, n5592);
   not (n5594, n5589);
   not (n5595, n5592);
   and (n5596, n5594, n5595);
   nor (n5597, n5593, n5596);
   xor (n5598, n5575, n5597);
   not (n5599, n5480);
   buf (n56, g55);
   nor (n560, n44, n46);
   not (n5600, n5571);
   or (n5601, n5599, n5600);
   or (n5602, n5480, n5571);
   nand (n5603, n5601, n5602);
   not (n5604, n5476);
   not (n5605, n5470);
   and (n5606, n5604, n5605);
   and (n5607, n5476, n5470);
   nor (n5608, n5606, n5607);
   not (n5609, n5608);
   not (n561, n560);
   not (n5610, n5609);
   not (n5611, n5505);
   not (n5612, n5540);
   or (n5613, n5611, n5612);
   or (n5614, n5540, n5505);
   nand (n5615, n5613, n5614);
   not (n5616, n5615);
   not (n5617, n5616);
   or (n5618, n5610, n5617);
   nand (n5619, n5615, n5608);
   or (n562, n559, n561);
   nand (n5620, n5618, n5619);
   not (n5621, n5620);
   not (n5622, n5300);
   not (n5623, n5331);
   or (n5624, n5622, n5623);
   not (n5625, n3912);
   not (n5626, n3905);
   or (n5627, n5625, n5626);
   nand (n5628, n5627, n5329);
   nand (n5629, n5325, n5628);
   not (n563, n45);
   nand (n5630, n5624, n5629);
   not (n5631, n5630);
   not (n5632, n5631);
   xnor (n5633, n5517, n5529);
   not (n5634, n5633);
   and (n5635, n5632, n5634);
   not (n5636, n5501);
   not (n5637, n5487);
   and (n5638, n5636, n5637);
   and (n5639, n5487, n5501);
   nand (n564, n563, n44, n46);
   nor (n5640, n5638, n5639);
   not (n5641, n5640);
   xnor (n5642, n5633, n5630);
   and (n5643, n5641, n5642);
   nor (n5644, n5635, n5643);
   or (n5645, n5621, n5644);
   not (n5646, n5609);
   or (n5647, n5616, n5646);
   nand (n5648, n5645, n5647);
   xor (n5649, n5603, n5648);
   nand (n565, n562, n564);
   nand (n5650, n5598, n5649);
   not (n5651, n5650);
   not (n5652, n5644);
   not (n5653, n5620);
   or (n5654, n5652, n5653);
   or (n5655, n5644, n5620);
   nand (n5656, n5654, n5655);
   not (n5657, n5656);
   not (n5658, n5642);
   not (n5659, n5640);
   buf (n566, n565);
   and (n5660, n5658, n5659);
   and (n5661, n5642, n5640);
   nor (n5662, n5660, n5661);
   not (n5663, n5662);
   not (n5664, n5663);
   not (n5665, n5258);
   not (n5666, n5665);
   not (n5667, n5281);
   and (n5668, n5666, n5667);
   and (n5669, n5283, n5251);
   and (n567, n44, n55);
   nor (n5670, n5668, n5669);
   not (n5671, n5670);
   not (n5672, n5349);
   not (n5673, n5343);
   or (n5674, n5672, n5673);
   nand (n5675, n5342, n5337);
   nand (n5676, n5674, n5675);
   not (n5677, n5676);
   or (n5678, n5671, n5677);
   or (n5679, n5676, n5670);
   not (n568, n44);
   nand (n5680, n5678, n5679);
   not (n5681, n5680);
   or (n5682, n5664, n5681);
   not (n5683, n5670);
   nand (n5684, n5683, n5676);
   nand (n5685, n5682, n5684);
   not (n5686, n5685);
   not (n5687, n5686);
   or (n5688, n5657, n5687);
   not (n5689, n5685);
   and (n569, n568, n377);
   or (n5690, n5689, n5656);
   nand (n5691, n5688, n5690);
   buf (n5692, n5691);
   not (n5693, n5350);
   not (n5694, n5296);
   or (n5695, n5693, n5694);
   not (n5696, n5284);
   nand (n5697, n5696, n5292);
   nand (n5698, n5695, n5697);
   not (n5699, n5662);
   buf (n57, g56);
   nor (n570, n567, n569);
   not (n5700, n5680);
   or (n5701, n5699, n5700);
   or (n5702, n5680, n5662);
   nand (n5703, n5701, n5702);
   xor (n5704, n5698, n5703);
   nand (n5705, n5651, n5692, n5704);
   or (n5706, n5357, n5705);
   and (n5707, n5698, n5703);
   not (n5708, n5707);
   not (n5709, n5691);
   nand (n571, n566, n570);
   or (n5710, n5708, n5709);
   not (n5711, n5689);
   nand (n5712, n5711, n5656);
   nand (n5713, n5710, n5712);
   not (n5714, n5713);
   not (n5715, n5714);
   nor (n5716, n5229, n5355);
   nand (n5717, n5691, n5704, n5716);
   not (n5718, n5717);
   or (n5719, n5715, n5718);
   nand (n572, n558, n571);
   nand (n5720, n5719, n5651);
   and (n5721, n5603, n5648);
   nand (n5722, n5598, n5721);
   and (n5723, n5720, n5722);
   nand (n5724, n5706, n5723);
   and (n5725, n5575, n5597);
   or (n5726, n5724, n5725);
   xor (n5727, n3202, n3276);
   xor (n5728, n5727, n3306);
   not (n5729, n5728);
   nand (n573, n36, n64);
   or (n5730, n5592, n5589);
   or (n5731, n5580, n5584);
   nand (n5732, n5730, n5731);
   not (n5733, n5732);
   or (n5734, n5729, n5733);
   or (n5735, n5732, n5728);
   nand (n5736, n5734, n5735);
   nand (n5737, n5726, n5736);
   not (n5738, n5728);
   nand (n5739, n5738, n5732);
   xnor (n574, n572, n573);
   nand (n5740, n5737, n5739);
   not (n5741, n3199);
   not (n5742, n3309);
   or (n5743, n5741, n5742);
   or (n5744, n3199, n3309);
   nand (n5745, n5743, n5744);
   nand (n5746, n5740, n5745);
   not (n5747, n5746);
   or (n5748, n3311, n5747);
   not (n5749, n3196);
   not (n575, n574);
   not (n5750, n3194);
   or (n5751, n5749, n5750);
   or (n5752, n3196, n3194);
   nand (n5753, n5751, n5752);
   buf (n5754, n5753);
   nand (n5755, n5748, n5754);
   not (n5756, n5755);
   or (n5757, n3198, n5756);
   xor (n5758, n3021, n3090);
   nand (n5759, n5757, n5758);
   and (n576, n40, n59);
   nand (n5760, n3092, n5759);
   not (n5761, n5760);
   or (n5762, n3020, n5761);
   not (n5763, n2973);
   nand (n5764, n5763, n3015);
   nand (n5765, n5762, n5764);
   not (n5766, n5765);
   or (n5767, n2972, n5766);
   or (n5768, n2971, n5765);
   nand (n5769, n5767, n5768);
   not (n577, n40);
   nand (n5770, n5769, n2);
   nand (n5771, n2827, n5770);
   not (n5772, n2);
   not (n5773, n2971);
   not (n5774, n5765);
   or (n5775, n5773, n5774);
   not (n5776, n2967);
   nand (n5777, n5776, n2886);
   nand (n5778, n5775, n5777);
   or (n5779, n2833, n37);
   not (n578, n59);
   nand (n5780, n2833, n37);
   nand (n5781, n5779, n5780);
   and (n5782, n5781, n2849);
   nand (n5783, n2861, n36);
   not (n5784, n5783);
   nor (n5785, n5782, n5784);
   nand (n5786, n2855, n36);
   nand (n5787, n5785, n5786);
   not (n5788, n5787);
   nor (n5789, n5785, n5786);
   and (n579, n577, n578);
   nor (n5790, n5788, n5789);
   not (n5791, n5790);
   and (n5792, n2880, n2884);
   and (n5793, n2881, n2799);
   nor (n5794, n5792, n5793);
   not (n5795, n5794);
   and (n5796, n5791, n5795);
   and (n5797, n5790, n5794);
   nor (n5798, n5796, n5797);
   not (n5799, n5798);
   buf (n58, g57);
   nor (n580, n576, n579);
   and (n5800, n2873, n2885);
   nor (n5801, n5800, n2872);
   not (n5802, n5801);
   or (n5803, n5799, n5802);
   or (n5804, n5801, n5798);
   nand (n5805, n5803, n5804);
   not (n5806, n5805);
   and (n5807, n5778, n5806);
   not (n5808, n5778);
   and (n5809, n5808, n5805);
   and (n581, n465, n580);
   nor (n5810, n5807, n5809);
   not (n5811, n5810);
   or (n5812, n5772, n5811);
   not (n5813, n2805);
   nand (n5814, n5813, n2809);
   nand (n5815, n2824, n5814);
   or (n5816, n2791, n2804);
   nand (n5817, n5816, n2790);
   and (n5818, n2797, n2803);
   and (n5819, n2799, n2798);
   and (n582, n40, n58);
   nor (n5820, n5818, n5819);
   not (n5821, n5820);
   or (n5822, n247, n2795);
   nand (n5823, n5822, n5783);
   not (n5824, n5823);
   nand (n5825, n36, n53);
   nor (n5826, n5824, n5825);
   not (n5827, n5825);
   nor (n5828, n5827, n5823);
   nor (n5829, n5826, n5828);
   nor (n583, n40, n58);
   not (n5830, n5829);
   and (n5831, n5821, n5830);
   and (n5832, n5820, n5829);
   nor (n5833, n5831, n5832);
   xor (n5834, n5817, n5833);
   or (n5835, n5815, n5834);
   not (n5836, n5814);
   not (n5837, n2824);
   or (n5838, n5836, n5837);
   nand (n5839, n5838, n5834);
   nor (n584, n582, n583);
   nand (n5840, n5835, n5839);
   nand (n5841, n5840, n237);
   nand (n5842, n5812, n5841);
   not (n5843, n5842);
   and (n5844, n5771, n5843);
   not (n5845, n237);
   and (n5846, n2747, n2753, n530);
   not (n5847, n5846);
   nand (n5848, n5847, n2755);
   not (n5849, n5848);
   and (n585, n274, n584);
   or (n5850, n5845, n5849);
   nand (n5851, n5755, n3197);
   or (n5852, n5851, n5758);
   nand (n5853, n5852, n5759);
   nand (n5854, n5853, n2);
   nand (n5855, n5850, n5854);
   not (n5856, n5855);
   not (n5857, n5856);
   not (n5858, n5857);
   not (n5859, n237);
   nor (n586, n581, n585);
   or (n5860, n2756, n2786);
   nand (n5861, n5860, n2821);
   not (n5862, n5861);
   or (n5863, n5859, n5862);
   xnor (n5864, n5760, n3019);
   nand (n5865, n5864, n2);
   nand (n5866, n5863, n5865);
   not (n5867, n5866);
   or (n5868, n5858, n5867);
   not (n5869, n5855);
   not (n587, n586);
   nand (n5870, n5746, n3310);
   or (n5871, n5870, n5754);
   nand (n5872, n5871, n5755);
   not (n5873, n5872);
   not (n5874, n2);
   or (n5875, n5873, n5874);
   or (n5876, n2745, n2746);
   nand (n5877, n5876, n2747);
   nand (n5878, n5877, n237);
   nand (n5879, n5875, n5878);
   not (n588, n587);
   not (n5880, n5879);
   nand (n5881, n5869, n5880);
   nand (n5882, n5868, n5881);
   not (n5883, n5882);
   not (n5884, n5771);
   or (n5885, n5883, n5884);
   not (n5886, n5881);
   buf (n5887, n5866);
   not (n5888, n5887);
   nand (n5889, n5886, n5888);
   or (n589, n575, n588);
   nand (n5890, n5885, n5889);
   not (n5891, n237);
   not (n5892, n2730);
   nor (n5893, n2715, n5892);
   not (n5894, n2740);
   and (n5895, n5893, n5894);
   not (n5896, n5893);
   and (n5897, n5896, n2740);
   nor (n5898, n5895, n5897);
   not (n5899, n5898);
   buf (n59, g58);
   not (n590, n572);
   or (n5900, n5891, n5899);
   or (n5901, n5724, n5725);
   nand (n5902, n5901, n5736);
   not (n5903, n5902);
   not (n5904, n5739);
   or (n5905, n5903, n5904, n5745);
   nand (n5906, n5905, n5746);
   nand (n5907, n5906, n2);
   nand (n5908, n5900, n5907);
   not (n5909, n5908);
   or (n591, n590, n573);
   not (n5910, n5909);
   not (n5911, n237);
   not (n5912, n2721);
   nand (n5913, n5912, n2658);
   nand (n5914, n5913, n2692);
   buf (n5915, n2728);
   not (n5916, n5915);
   and (n5917, n5914, n5916);
   not (n5918, n5914);
   and (n5919, n5918, n5915);
   nand (n592, n589, n591);
   nor (n5920, n5917, n5919);
   not (n5921, n5920);
   or (n5922, n5911, n5921);
   buf (n5923, n5724);
   or (n5924, n5923, n5725, n5736);
   nand (n5925, n5924, n5902);
   nand (n5926, n5925, n2);
   nand (n5927, n5922, n5926);
   not (n5928, n5927);
   not (n5929, n237);
   xor (n593, n545, n592);
   not (n5930, n2721);
   not (n5931, n2658);
   not (n5932, n5931);
   or (n5933, n5930, n5932);
   nand (n5934, n5933, n5913);
   not (n5935, n5934);
   or (n5936, n5929, n5935);
   nor (n5937, n5598, n5721);
   not (n5938, n5937);
   buf (n5939, n5712);
   not (n594, n57);
   not (n5940, n5939);
   not (n5941, n5707);
   not (n5942, n5941);
   not (n5943, n5716);
   not (n5944, n5943);
   nand (n5945, n5225, n5356);
   not (n5946, n5945);
   or (n5947, n5944, n5946);
   nand (n5948, n5947, n5704);
   not (n5949, n5948);
   not (n595, n42);
   or (n5950, n5942, n5949);
   nand (n5951, n5950, n5692);
   not (n5952, n5951);
   or (n5953, n5940, n5952);
   buf (n5954, n5649);
   nand (n5955, n5953, n5954);
   not (n5956, n5955);
   or (n5957, n5938, n5956);
   not (n5958, n5923);
   nand (n5959, n5957, n5958);
   or (n596, n594, n595);
   nand (n5960, n5959, n2);
   nand (n5961, n5936, n5960);
   not (n5962, n5961);
   and (n5963, n5928, n5962);
   not (n5964, n5963);
   or (n5965, n5910, n5964);
   not (n5966, n5909);
   not (n5967, n5928);
   nand (n5968, n5966, n5967, n5879);
   nand (n5969, n5965, n5968);
   or (n597, n42, n57);
   not (n5970, n2);
   and (n5971, n5216, n4310);
   not (n5972, n5216);
   and (n5973, n5972, n5217);
   nor (n5974, n5971, n5973);
   not (n5975, n4301);
   not (n5976, n5198);
   and (n5977, n5976, n5201);
   not (n5978, n4445);
   not (n5979, n5206);
   nand (n598, n596, n597);
   or (n5980, n5978, n5979);
   nand (n5981, n5980, n4507);
   nor (n5982, n5977, n5981);
   nand (n5983, n5982, n5211);
   not (n5984, n5983);
   or (n5985, n5975, n5984);
   nand (n5986, n5985, n5209);
   xor (n5987, n5974, n5986);
   not (n5988, n5987);
   or (n5989, n5970, n5988);
   not (n599, n598);
   not (n5990, n2634);
   nor (n5991, n5990, n1721);
   not (n5992, n5991);
   buf (n5993, n2629);
   not (n5994, n5993);
   not (n5995, n5994);
   nand (n5996, n2582, n2611);
   not (n5997, n5996);
   or (n5998, n5995, n5997);
   nand (n5999, n5998, n2620);
   buf (n6, g5);
   buf (n60, g59);
   not (n600, n599);
   nand (n6000, n5999, n2632);
   not (n6001, n6000);
   or (n6002, n5992, n6001);
   nand (n6003, n1721, n2623, n2635);
   nand (n6004, n6002, n6003);
   nand (n6005, n6004, n237);
   nand (n6006, n5989, n6005);
   not (n6007, n85);
   nand (n6008, n6006, n6007);
   not (n6009, n84);
   not (n601, n421);
   not (n6010, n4037);
   not (n6011, n5218);
   nand (n6012, n5213, n5202, n6011);
   not (n6013, n4312);
   nand (n6014, n6013, n6011);
   nand (n6015, n6012, n6014);
   not (n6016, n6015);
   xor (n6017, n6010, n6016);
   not (n6018, n6017);
   not (n6019, n2);
   or (n602, n600, n601);
   or (n6020, n6018, n6019);
   not (n6021, n2637);
   not (n6022, n2642);
   or (n6023, n6021, n6022);
   or (n6024, n2637, n2642);
   nand (n6025, n6023, n6024);
   nand (n6026, n6025, n237);
   nand (n6027, n6020, n6026);
   xor (n6028, n6009, n6027);
   xor (n6029, n6008, n6028);
   and (n603, n42, n56);
   not (n6030, n2);
   not (n6031, n4301);
   not (n6032, n5983);
   or (n6033, n6031, n6032);
   or (n6034, n4301, n5983);
   nand (n6035, n6033, n6034);
   not (n6036, n6035);
   or (n6037, n6030, n6036);
   or (n6038, n5999, n2632);
   nand (n6039, n6038, n6000);
   nor (n604, n42, n56);
   nand (n6040, n6039, n237);
   nand (n6041, n6037, n6040);
   not (n6042, n6041);
   not (n6043, n86);
   and (n6044, n6042, n6043);
   and (n6045, n6041, n86);
   nor (n6046, n6044, n6045);
   not (n6047, n5982);
   not (n6048, n5191);
   nand (n6049, n6048, n5205);
   nor (n605, n603, n604);
   not (n6050, n6049);
   buf (n6051, n5197);
   not (n6052, n6051);
   or (n6053, n6050, n6052);
   nor (n6054, n5201, n4506);
   nand (n6055, n6053, n6054);
   not (n6056, n6055);
   or (n6057, n6047, n6056);
   nand (n6058, n6057, n2);
   not (n6059, n6058);
   nand (n606, n513, n605);
   not (n6060, n5994);
   not (n6061, n5996);
   or (n6062, n6060, n6061);
   or (n6063, n5996, n5994);
   nand (n6064, n6062, n6063);
   nand (n6065, n6064, n237);
   not (n6066, n6065);
   or (n6067, n6059, n6066);
   not (n6068, n87);
   nand (n6069, n6067, n6068);
   nand (n607, n602, n606);
   buf (n6070, n6069);
   nor (n6071, n6046, n6070);
   not (n6072, n6071);
   not (n6073, n86);
   and (n6074, n6041, n6073);
   not (n6075, n6074);
   and (n6076, n6072, n6075);
   and (n6077, n6006, n85);
   not (n6078, n6006);
   and (n6079, n6078, n6007);
   not (n608, n607);
   nor (n6080, n6077, n6079);
   nor (n6081, n6076, n6080);
   nor (n6082, n6029, n6081);
   not (n6083, n6082);
   not (n6084, n90);
   not (n6085, n2181);
   nor (n6086, n6085, n2050);
   not (n6087, n6086);
   buf (n6088, n2176);
   not (n6089, n6088);
   not (n609, n48);
   buf (n6090, n2298);
   not (n6091, n6090);
   not (n6092, n2527);
   or (n6093, n6091, n6092);
   buf (n6094, n2174);
   not (n6095, n6094);
   nand (n6096, n6093, n6095);
   not (n6097, n6096);
   or (n6098, n6089, n6097);
   buf (n6099, n2117);
   buf (n61, g60);
   not (n610, n49);
   nand (n6100, n6098, n6099);
   not (n6101, n6100);
   or (n6102, n6087, n6101);
   nand (n6103, n2299, n2527);
   nand (n6104, n6103, n2182, n2050);
   nand (n6105, n6102, n6104);
   not (n6106, n6105);
   not (n6107, n237);
   or (n6108, n6106, n6107);
   xor (n6109, n5136, n5141);
   not (n611, n610);
   not (n6110, n6109);
   not (n6111, n5095);
   not (n6112, n6111);
   nand (n6113, n4708, n4912);
   nand (n6114, n4626, n5022);
   nand (n6115, n6113, n6114);
   not (n6116, n6115);
   or (n6117, n6112, n6116);
   nand (n6118, n6117, n5096);
   buf (n6119, n5090);
   or (n612, n609, n611);
   nand (n6120, n6118, n6119);
   nand (n6121, n6120, n5143);
   not (n6122, n6121);
   or (n6123, n6110, n6122);
   nand (n6124, n6123, n5142);
   xor (n6125, n5174, n5173);
   not (n6126, n6125);
   and (n6127, n6124, n6126);
   not (n6128, n6124);
   and (n6129, n6128, n6125);
   xor (n613, n49, n50);
   nor (n6130, n6127, n6129);
   nand (n6131, n6130, n2);
   nand (n6132, n6108, n6131);
   xor (n6133, n6084, n6132);
   not (n6134, n91);
   not (n6135, n2);
   not (n6136, n6109);
   and (n6137, n6121, n6136);
   not (n6138, n6121);
   and (n6139, n6138, n6109);
   buf (n614, n613);
   nor (n6140, n6137, n6139);
   not (n6141, n6140);
   or (n6142, n6135, n6141);
   nand (n6143, n6096, n6088);
   or (n6144, n6143, n6099);
   nand (n6145, n6144, n6100);
   nand (n6146, n6145, n237);
   nand (n6147, n6142, n6146);
   and (n6148, n6134, n6147);
   or (n6149, n6133, n6148);
   nand (n615, n614, n48);
   not (n6150, n6149);
   not (n6151, n94);
   not (n6152, n237);
   or (n6153, n2347, n2522);
   nand (n6154, n6153, n2523);
   not (n6155, n6154);
   or (n6156, n6152, n6155);
   or (n6157, n4708, n4912);
   nand (n6158, n6157, n6113);
   nand (n6159, n6158, n2);
   nand (n616, n612, n615);
   nand (n6160, n6156, n6159);
   and (n6161, n6151, n6160);
   xor (n6162, n93, n6161);
   not (n6163, n6111);
   not (n6164, n6115);
   or (n6165, n6163, n6164);
   or (n6166, n6115, n6111);
   nand (n6167, n6165, n6166);
   not (n6168, n6167);
   not (n6169, n2);
   not (n617, n616);
   or (n6170, n6168, n6169);
   nand (n6171, n2523, n2345);
   or (n6172, n6171, n2526);
   nand (n6173, n6172, n2527);
   nand (n6174, n6173, n237);
   nand (n6175, n6170, n6174);
   xnor (n6176, n6162, n6175);
   not (n6177, n6176);
   and (n6178, n4851, n4855);
   not (n6179, n4851);
   and (n618, n608, n617);
   not (n6180, n4855);
   and (n6181, n6179, n6180);
   or (n6182, n6178, n6181);
   not (n6183, n6182);
   not (n6184, n4825);
   not (n6185, n6184);
   not (n6186, n4894);
   or (n6187, n6185, n6186);
   nand (n6188, n6187, n4899);
   not (n6189, n4905);
   not (n619, n616);
   nor (n6190, n6188, n6189);
   not (n6191, n4849);
   nor (n6192, n6190, n6191);
   not (n6193, n6192);
   or (n6194, n6183, n6193);
   or (n6195, n6192, n6182);
   nand (n6196, n6194, n6195);
   nand (n6197, n6196, n2);
   nand (n6198, n2516, n2518);
   not (n6199, n2352);
   buf (n62, g61);
   not (n620, n619);
   not (n6200, n2390);
   and (n6201, n6199, n6200);
   and (n6202, n2352, n2390);
   nor (n6203, n6201, n6202);
   and (n6204, n6198, n6203);
   not (n6205, n6198);
   not (n6206, n6203);
   and (n6207, n6205, n6206);
   nor (n6208, n6204, n6207);
   nand (n6209, n6208, n237);
   and (n621, n607, n620);
   nand (n6210, n6197, n6209);
   not (n6211, n6210);
   not (n6212, n6211);
   xor (n6213, n6151, n6160);
   not (n6214, n6213);
   or (n6215, n6212, n6214);
   or (n6216, n6213, n6211);
   nand (n6217, n6215, n6216);
   not (n6218, n6217);
   xor (n6219, n95, n6210);
   nor (n622, n618, n621);
   not (n6220, n237);
   xor (n6221, n2423, n2439);
   xor (n6222, n6221, n2495);
   not (n6223, n6222);
   or (n6224, n6220, n6223);
   nand (n6225, n4894, n4824);
   and (n6226, n4800, n4748);
   not (n6227, n4800);
   and (n6228, n6227, n4898);
   nor (n6229, n6226, n6228);
   and (n623, n504, n312);
   or (n6230, n6225, n6229);
   nand (n6231, n6225, n6229);
   nand (n6232, n6230, n6231, n2);
   nand (n6233, n6224, n6232);
   xor (n6234, n97, n6233);
   not (n6235, n4894);
   nor (n6236, n4893, n4888);
   nor (n6237, n6236, n237);
   not (n6238, n6237);
   or (n6239, n6235, n6238);
   and (n624, n46, n53);
   xor (n6240, n2490, n2477);
   nand (n6241, n6240, n237);
   nand (n6242, n6239, n6241);
   not (n6243, n6242);
   not (n6244, n98);
   not (n6245, n6244);
   and (n6246, n6243, n6245);
   and (n6247, n6242, n6244);
   nor (n6248, n6246, n6247);
   or (n6249, n4874, n4886);
   nor (n625, n623, n624);
   nand (n6250, n6249, n4887);
   and (n6251, n6250, n2);
   not (n6252, n2476);
   nand (n6253, n6252, n2474);
   xnor (n6254, n6253, n2458);
   and (n6255, n6254, n237);
   nor (n6256, n6251, n6255);
   nand (n6257, n99, n6256);
   or (n6258, n6248, n6257);
   not (n6259, n6244);
   and (n626, n535, n625);
   nand (n6260, n6259, n6242);
   nand (n6261, n6258, n6260);
   and (n6262, n6234, n6261);
   and (n6263, n97, n6233);
   or (n6264, n6262, n6263);
   nand (n6265, n6188, n6189);
   nand (n6266, n2, n6265);
   or (n6267, n6266, n6190);
   not (n6268, n2498);
   not (n6269, n6268);
   not (n627, n541);
   not (n6270, n2515);
   and (n6271, n6269, n6270);
   and (n6272, n6268, n2515);
   nor (n6273, n6271, n6272);
   or (n6274, n6273, n2);
   nand (n6275, n6267, n6274);
   xor (n6276, n96, n6275);
   and (n6277, n6264, n6276);
   and (n6278, n96, n6275);
   nor (n6279, n6277, n6278);
   and (n628, n627, n538);
   nand (n6280, n6219, n6279);
   not (n6281, n95);
   nand (n6282, n6211, n6281);
   and (n6283, n6280, n6282);
   not (n6284, n6283);
   or (n6285, n6218, n6284);
   not (n6286, n6213);
   nand (n6287, n6286, n6211);
   nand (n6288, n6285, n6287);
   not (n6289, n6288);
   nor (n629, n626, n628);
   or (n6290, n6177, n6289);
   not (n6291, n6161);
   not (n6292, n93);
   xnor (n6293, n6175, n6292);
   nand (n6294, n6291, n6293);
   nand (n6295, n6290, n6294);
   not (n6296, n6295);
   and (n6297, n6175, n6292);
   xor (n6298, n92, n6297);
   not (n6299, n6119);
   buf (n63, g62);
   or (n630, n622, n629);
   not (n6300, n6118);
   or (n6301, n6299, n6300);
   or (n6302, n6118, n6119);
   nand (n6303, n6301, n6302);
   nand (n6304, n6303, n2);
   nand (n6305, n2527, n6090, n6094);
   not (n6306, n6305);
   not (n6307, n6096);
   or (n6308, n6306, n6307);
   nand (n6309, n6308, n237);
   not (n631, n607);
   nand (n6310, n6304, n6309);
   xnor (n6311, n6298, n6310);
   not (n6312, n6311);
   or (n6313, n6296, n6312);
   nand (n6314, n6304, n6309);
   nor (n6315, n6314, n92);
   not (n6316, n6315);
   nand (n6317, n6314, n92);
   not (n6318, n6297);
   nand (n6319, n6316, n6317, n6318);
   or (n632, n631, n620);
   nand (n6320, n6313, n6319);
   not (n6321, n6320);
   xor (n6322, n6134, n6147);
   not (n6323, n6322);
   not (n6324, n92);
   nand (n6325, n6314, n6324);
   not (n6326, n6325);
   and (n6327, n6323, n6326);
   and (n6328, n6322, n6325);
   nor (n6329, n6327, n6328);
   nand (n633, n630, n632);
   or (n6330, n6321, n6329);
   not (n6331, n6322);
   nand (n6332, n6331, n6325);
   nand (n6333, n6330, n6332);
   not (n6334, n6333);
   not (n6335, n6334);
   or (n6336, n6150, n6335);
   and (n6337, n6084, n6132);
   not (n6338, n237);
   not (n6339, n6104);
   and (n634, n593, n633);
   buf (n6340, n2242);
   not (n6341, n6340);
   xor (n6342, n2189, n2579);
   nor (n6343, n6339, n6341, n6342);
   not (n6344, n6343);
   not (n6345, n6340);
   not (n6346, n6104);
   or (n6347, n6345, n6346);
   nand (n6348, n6347, n6342);
   nand (n6349, n6344, n6348);
   and (n635, n545, n592);
   not (n6350, n6349);
   or (n6351, n6338, n6350);
   not (n6352, n5191);
   nand (n6353, n5177, n5190);
   nand (n6354, n6352, n6353);
   nand (n6355, n2, n6354);
   nand (n6356, n6351, n6355);
   not (n6357, n89);
   nor (n6358, n6356, n6357);
   not (n6359, n6358);
   nor (n636, n634, n635);
   not (n6360, n89);
   nand (n6361, n6360, n6356);
   nand (n6362, n6359, n6361);
   and (n6363, n6337, n6362);
   not (n6364, n6337);
   not (n6365, n6362);
   and (n6366, n6364, n6365);
   nor (n6367, n6363, n6366);
   and (n6368, n6148, n6133);
   nor (n6369, n6367, n6368);
   and (n637, n362, n584);
   nand (n6370, n6336, n6369);
   not (n6371, n6084);
   not (n6372, n6132);
   or (n6373, n6371, n6372);
   nand (n6374, n6373, n6362);
   not (n6375, n6361);
   not (n6376, n6375);
   not (n6377, n2);
   not (n6378, n6051);
   xor (n6379, n6378, n6049);
   and (n638, n276, n498);
   not (n6380, n6379);
   or (n6381, n6377, n6380);
   nand (n6382, n6348, n2578, n2240);
   not (n6383, n6382);
   not (n6384, n2582);
   or (n6385, n6383, n6384);
   nand (n6386, n6385, n237);
   nand (n6387, n6381, n6386);
   not (n6388, n88);
   nor (n6389, n6387, n6388);
   and (n639, n40, n57);
   not (n6390, n6389);
   nand (n6391, n6387, n6388);
   nand (n6392, n6390, n6391);
   nand (n6393, n6376, n6392);
   and (n6394, n6374, n6393);
   nand (n6395, n6370, n6394);
   buf (n6396, n6393);
   xor (n6397, n6392, n6375);
   and (n6398, n6396, n6397);
   nand (n6399, n6065, n6058, n87);
   buf (n64, g63);
   nor (n640, n638, n639);
   nand (n6400, n6069, n6399);
   not (n6401, n6400);
   not (n6402, n6391);
   not (n6403, n6402);
   and (n6404, n6401, n6403);
   and (n6405, n6400, n6402);
   nor (n6406, n6404, n6405);
   nor (n6407, n6398, n6406);
   and (n6408, n6395, n6407);
   not (n6409, n6400);
   and (n641, n274, n640);
   nor (n6410, n6409, n6402);
   nor (n6411, n6408, n6410);
   not (n6412, n6074);
   and (n6413, n6080, n6412);
   not (n6414, n6070);
   not (n6415, n6046);
   nor (n6416, n6414, n6415);
   nor (n6417, n6413, n6416);
   nand (n6418, n6411, n6417);
   not (n6419, n6418);
   nor (n642, n637, n641);
   or (n6420, n6083, n6419);
   not (n6421, n6007);
   not (n6422, n6006);
   or (n6423, n6421, n6422);
   not (n6424, n6028);
   nand (n6425, n6423, n6424);
   nand (n6426, n6420, n6425);
   not (n6427, n2);
   buf (n6428, n5945);
   nand (n6429, n6428, n5943);
   not (n643, n642);
   or (n6430, n6429, n5704);
   nand (n6431, n6430, n5948);
   not (n6432, n6431);
   or (n6433, n6427, n6432);
   not (n6434, n2642);
   not (n6435, n2637);
   or (n6436, n6434, n6435);
   nand (n6437, n6436, n1565);
   buf (n6438, n2644);
   nand (n6439, n6437, n6438);
   not (n644, n643);
   buf (n6440, n6439);
   nand (n6441, n6440, n2648, n1429);
   not (n6442, n6441);
   not (n6443, n6439);
   not (n6444, n1429);
   or (n6445, n6443, n6444);
   not (n6446, n2648);
   nand (n6447, n6445, n6446);
   not (n6448, n6447);
   or (n6449, n6442, n6448);
   and (n645, n38, n60);
   nand (n6450, n6449, n237);
   nand (n6451, n6433, n6450);
   not (n6452, n6451);
   not (n6453, n6452);
   not (n6454, n2);
   not (n6455, n5224);
   or (n6456, n6455, n5203, n5356);
   nand (n6457, n6456, n6428);
   not (n6458, n6457);
   or (n6459, n6454, n6458);
   not (n646, n38);
   not (n6460, n6438);
   not (n6461, n6460);
   not (n6462, n6437);
   not (n6463, n6462);
   or (n6464, n6461, n6463);
   nand (n6465, n6464, n6440);
   nand (n6466, n6465, n237);
   nand (n6467, n6459, n6466);
   not (n6468, n6467);
   not (n6469, n6468);
   not (n647, n60);
   nand (n6470, n6453, n6469);
   and (n6471, n6009, n6027);
   not (n6472, n6471);
   nand (n6473, n6468, n6472);
   nand (n6474, n6470, n6473);
   nand (n6475, n6426, n6474);
   or (n6476, n2655, n2656);
   nand (n6477, n6476, n2657);
   and (n6478, n237, n6477);
   not (n6479, n237);
   and (n648, n646, n647);
   nand (n6480, n5951, n5939);
   or (n6481, n6480, n5954);
   nand (n6482, n6481, n5955);
   and (n6483, n6479, n6482);
   nor (n6484, n6478, n6483);
   not (n6485, n6484);
   not (n6486, n6485);
   not (n6487, n6486);
   not (n6488, n6487);
   not (n6489, n6452);
   nor (n649, n645, n648);
   not (n6490, n6489);
   not (n6491, n5692);
   not (n6492, n6491);
   and (n6493, n5948, n5941);
   not (n6494, n6493);
   or (n6495, n6492, n6494);
   nand (n6496, n6495, n5951);
   not (n6497, n6496);
   not (n6498, n2);
   or (n6499, n6497, n6498);
   buf (n65, g64);
   not (n650, n649);
   not (n6500, n1373);
   nor (n6501, n6500, n2651);
   not (n6502, n6501);
   not (n6503, n6447);
   or (n6504, n6502, n6503);
   nand (n6505, n6504, n2654);
   nand (n6506, n6505, n237);
   nand (n6507, n6499, n6506);
   not (n6508, n6507);
   nand (n6509, n6490, n6508);
   not (n651, n296);
   not (n6510, n6509);
   and (n6511, n6488, n6510);
   not (n6512, n5962);
   nor (n6513, n6511, n6512);
   nor (n6514, n6475, n6513);
   and (n6515, n5969, n6514);
   nand (n6516, n5890, n6515);
   nor (n6517, n5844, n6516);
   not (n6518, n5843);
   and (n6519, n5820, n5828);
   not (n652, n651);
   not (n6520, n5820);
   and (n6521, n6520, n5826);
   nor (n6522, n6519, n6521);
   nor (n6523, n2762, n242);
   and (n6524, n6523, n52);
   and (n6525, n1267, n267);
   nor (n6526, n6524, n6525);
   xor (n6527, n6522, n6526);
   not (n6528, n5833);
   not (n6529, n5817);
   or (n653, n650, n652);
   or (n6530, n6528, n6529);
   nand (n6531, n6530, n5839);
   xnor (n6532, n6527, n6531);
   and (n6533, n237, n6532);
   not (n6534, n237);
   not (n6535, n5787);
   not (n6536, n5794);
   or (n6537, n6535, n6536);
   or (n6538, n5794, n5789);
   nand (n6539, n6537, n6538);
   and (n654, n38, n59);
   not (n6540, n6539);
   and (n6541, n2833, n6523);
   not (n6542, n2833);
   and (n6543, n6542, n1267);
   nor (n6544, n6541, n6543);
   not (n6545, n6544);
   and (n6546, n6540, n6545);
   and (n6547, n6539, n6544);
   nor (n6548, n6546, n6547);
   not (n6549, n6548);
   not (n655, n38);
   not (n6550, n5805);
   not (n6551, n5778);
   or (n6552, n6550, n6551);
   not (n6553, n5801);
   nand (n6554, n6553, n5798);
   nand (n6555, n6552, n6554);
   not (n6556, n6555);
   or (n6557, n6549, n6556);
   or (n6558, n6555, n6548);
   nand (n6559, n6557, n6558);
   and (n656, n655, n578);
   and (n6560, n6534, n6559);
   nor (n6561, n6533, n6560);
   nand (n6562, n6518, n6561);
   nand (n6563, n6517, n6562);
   and (n6564, n237, n6532);
   not (n6565, n237);
   and (n6566, n6565, n6559);
   nor (n6567, n6564, n6566);
   buf (n6568, n5842);
   not (n6569, n1);
   nor (n657, n654, n656);
   nor (n6570, n6508, n6569, n6472, n6470);
   nand (n6571, n6512, n6487, n6570);
   nor (n6572, n5968, n6571);
   nand (n6573, n6568, n5890, n6572);
   nor (n6574, n6567, n6573);
   nand (n6575, n6563, n6574);
   not (n6576, n6575);
   not (n6577, n70);
   nor (n6578, n6577, n6007);
   not (n6579, n71);
   nand (n658, n310, n657);
   nor (n6580, n6007, n6579);
   nand (n6581, n68, n69);
   not (n6582, n6581);
   not (n6583, n6582);
   nand (n6584, n87, n88);
   nor (n6585, n6583, n6584);
   and (n6586, n68, n88);
   and (n6587, n69, n87);
   nor (n6588, n6586, n6587);
   nor (n6589, n6585, n6588);
   nand (n659, n653, n658);
   and (n6590, n6580, n6589);
   or (n6591, n6590, n6585);
   xor (n6592, n6578, n6591);
   nor (n6593, n6579, n6009);
   nand (n6594, n86, n87);
   nor (n6595, n6583, n6594);
   and (n6596, n68, n87);
   and (n6597, n69, n86);
   nor (n6598, n6596, n6597);
   nor (n6599, n6595, n6598);
   buf (n66, g65);
   not (n660, n659);
   xor (n6600, n6593, n6599);
   xor (n6601, n6592, n6600);
   nand (n6602, n70, n86);
   nand (n6603, n72, n84);
   and (n6604, n6602, n6603);
   nand (n6605, n70, n84);
   nand (n6606, n72, n86);
   nor (n6607, n6605, n6606);
   nor (n6608, n6604, n6607);
   not (n6609, n73);
   and (n661, n566, n549);
   nor (n6610, n6609, n6009);
   not (n6611, n6578);
   nand (n6612, n72, n87);
   nor (n6613, n6611, n6612);
   and (n6614, n70, n87);
   and (n6615, n72, n85);
   nor (n6616, n6614, n6615);
   nor (n6617, n6613, n6616);
   and (n6618, n6610, n6617);
   or (n6619, n6618, n6613);
   not (n662, n44);
   and (n6620, n6608, n6619);
   or (n6621, n6620, n6607);
   or (n6622, n6601, n6621);
   nand (n6623, n6601, n6621);
   nand (n6624, n6622, n6623);
   nor (n6625, n6579, n6073);
   nand (n6626, n88, n89);
   nor (n6627, n6583, n6626);
   and (n6628, n68, n89);
   and (n6629, n69, n88);
   not (n663, n53);
   nor (n6630, n6628, n6629);
   nor (n6631, n6627, n6630);
   and (n6632, n6625, n6631);
   or (n6633, n6632, n6627);
   xor (n6634, n6580, n6589);
   xor (n6635, n6633, n6634);
   xor (n6636, n6608, n6619);
   and (n6637, n6635, n6636);
   and (n6638, n6633, n6634);
   nor (n6639, n6637, n6638);
   and (n664, n662, n663);
   or (n6640, n6624, n6639);
   nand (n6641, n6640, n6623);
   xor (n6642, n6578, n6591);
   and (n6643, n6642, n6600);
   and (n6644, n6578, n6591);
   nor (n6645, n6643, n6644);
   nand (n6646, n85, n86);
   nor (n6647, n6583, n6646);
   and (n6648, n68, n86);
   and (n6649, n69, n85);
   and (n665, n44, n53);
   nor (n6650, n6648, n6649);
   nor (n6651, n6647, n6650);
   and (n6652, n6651, n6605);
   nor (n6653, n6651, n6605);
   nor (n6654, n6652, n6653);
   not (n6655, n6654);
   and (n6656, n6593, n6599);
   nor (n6657, n6656, n6595);
   not (n6658, n6657);
   or (n6659, n6655, n6658);
   nor (n666, n664, n665);
   or (n6660, n6657, n6654);
   nand (n6661, n6659, n6660);
   xor (n6662, n6645, n6661);
   or (n6663, n6641, n6662);
   not (n6664, n6663);
   and (n6665, n75, n85);
   and (n6666, n76, n84);
   nor (n6667, n6665, n6666);
   not (n6668, n6667);
   nand (n6669, n75, n76);
   and (n667, n556, n666);
   not (n6670, n6669);
   nand (n6671, n84, n85);
   not (n6672, n6671);
   nand (n6673, n6670, n6672);
   nand (n6674, n6668, n6673);
   nand (n6675, n72, n88);
   or (n6676, n6674, n6675);
   nand (n6677, n6676, n6673);
   and (n6678, n68, n92);
   and (n6679, n69, n91);
   nor (n668, n661, n667);
   nor (n6680, n6678, n6679);
   not (n6681, n6680);
   nand (n6682, n6582, n91, n92);
   nand (n6683, n6681, n6682);
   nand (n6684, n71, n89);
   nor (n6685, n6683, n6684);
   not (n6686, n6685);
   nand (n6687, n6686, n6682);
   xor (n6688, n6677, n6687);
   nor (n6689, n6388, n6579);
   not (n669, n668);
   nand (n6690, n90, n91);
   nor (n6691, n6583, n6690);
   and (n6692, n68, n91);
   and (n6693, n69, n90);
   nor (n6694, n6692, n6693);
   nor (n6695, n6691, n6694);
   xor (n6696, n6689, n6695);
   and (n6697, n6688, n6696);
   and (n6698, n6677, n6687);
   nor (n6699, n6697, n6698);
   buf (n67, g66);
   or (n670, n660, n669);
   nand (n6700, n74, n84);
   not (n6701, n6700);
   and (n6702, n6689, n6695);
   or (n6703, n6702, n6691);
   xor (n6704, n6701, n6703);
   nand (n6705, n75, n84);
   or (n6706, n6612, n6705);
   xnor (n6707, n6612, n6705);
   nand (n6708, n70, n89);
   nor (n6709, n6707, n6708);
   not (n671, n668);
   not (n6710, n6709);
   nand (n6711, n6706, n6710);
   xnor (n6712, n6704, n6711);
   xnor (n6713, n6699, n6712);
   nand (n6714, n70, n90);
   nand (n6715, n73, n87);
   or (n6716, n6714, n6715);
   xnor (n6717, n6715, n6714);
   nand (n6718, n74, n86);
   nor (n6719, n6717, n6718);
   not (n672, n659);
   not (n6720, n6719);
   nand (n6721, n6716, n6720);
   nand (n6722, n74, n85);
   nand (n6723, n73, n86);
   and (n6724, n6722, n6723);
   nand (n6725, n73, n74);
   nor (n6726, n6725, n6646);
   nor (n6727, n6724, n6726);
   xor (n6728, n6721, n6727);
   and (n6729, n6707, n6708);
   nand (n673, n671, n672);
   nor (n6730, n6729, n6709);
   and (n6731, n6728, n6730);
   xor (n6732, n6728, n6730);
   nor (n6733, n6609, n6388);
   and (n6734, n77, n91);
   not (n6735, n6734);
   nor (n6736, n6735, n6605);
   and (n6737, n70, n91);
   and (n6738, n77, n84);
   nor (n6739, n6737, n6738);
   nand (n674, n670, n673);
   nor (n6740, n6736, n6739);
   and (n6741, n6733, n6740);
   or (n6742, n6741, n6736);
   and (n6743, n75, n86);
   and (n6744, n76, n85);
   nor (n6745, n6743, n6744);
   not (n6746, n6745);
   not (n6747, n6646);
   nand (n6748, n6747, n6670);
   nand (n6749, n6746, n6748);
   not (n675, n674);
   nand (n6750, n72, n89);
   or (n6751, n6749, n6750);
   nand (n6752, n6751, n6748);
   nand (n6753, n6582, n92, n93);
   not (n6754, n6753);
   and (n6755, n68, n93);
   and (n6756, n69, n92);
   nor (n6757, n6755, n6756);
   nor (n6758, n6754, n6757);
   nor (n6759, n6084, n6579);
   or (n676, n644, n675);
   nand (n6760, n6758, n6759);
   nand (n6761, n6760, n6753);
   xor (n6762, n6752, n6761);
   and (n6763, n6742, n6762);
   and (n6764, n6752, n6761);
   or (n6765, n6763, n6764);
   and (n6766, n6732, n6765);
   nor (n6767, n6731, n6766);
   xor (n6768, n6713, n6767);
   nor (n6769, n6579, n6068);
   or (n677, n672, n668);
   nand (n6770, n89, n90);
   nor (n6771, n6583, n6770);
   and (n6772, n68, n90);
   and (n6773, n69, n89);
   nor (n6774, n6772, n6773);
   nor (n6775, n6771, n6774);
   xor (n6776, n6769, n6775);
   nor (n6777, n6609, n6007);
   nand (n6778, n70, n88);
   and (n6779, n6606, n6778);
   nand (n678, n676, n677);
   nor (n6780, n6675, n6602);
   nor (n6781, n6779, n6780);
   xor (n6782, n6777, n6781);
   xnor (n6783, n6776, n6782);
   and (n6784, n6721, n6727);
   nor (n6785, n6784, n6726);
   xor (n6786, n6783, n6785);
   xor (n6787, n6768, n6786);
   nor (n6788, n6581, n6151, n6292);
   and (n6789, n68, n94);
   nand (n679, n36, n62);
   and (n6790, n69, n93);
   nor (n6791, n6789, n6790);
   or (n6792, n6788, n6791);
   nand (n6793, n71, n91);
   nor (n6794, n6792, n6793);
   nor (n6795, n6794, n6788);
   nand (n6796, n74, n87);
   nor (n6797, n6795, n6796);
   not (n6798, n6797);
   and (n6799, n6795, n6796);
   buf (n68, g67);
   xnor (n680, n679, n545);
   nor (n6800, n6799, n6797);
   not (n6801, n72);
   nor (n6802, n6801, n6084);
   nor (n6803, n6669, n6594);
   and (n6804, n75, n87);
   and (n6805, n76, n86);
   nor (n6806, n6804, n6805);
   nor (n6807, n6803, n6806);
   and (n6808, n6802, n6807);
   or (n6809, n6808, n6803);
   xor (n681, n678, n680);
   nand (n6810, n6800, n6809);
   nand (n6811, n6798, n6810);
   xor (n6812, n6749, n6750);
   not (n6813, n6812);
   or (n6814, n6758, n6759);
   nand (n6815, n6814, n6760);
   nor (n6816, n6324, n6577);
   nand (n6817, n77, n78);
   nor (n6818, n6817, n6671);
   and (n6819, n77, n85);
   xor (n682, n636, n681);
   and (n6820, n78, n84);
   nor (n6821, n6819, n6820);
   nor (n6822, n6818, n6821);
   and (n6823, n6816, n6822);
   nor (n6824, n6823, n6818);
   and (n6825, n6815, n6824);
   nor (n6826, n6815, n6824);
   nor (n6827, n6825, n6826);
   not (n6828, n6827);
   or (n6829, n6813, n6828);
   not (n683, n642);
   not (n6830, n6826);
   nand (n6831, n6829, n6830);
   xor (n6832, n6811, n6831);
   xor (n6833, n6742, n6762);
   and (n6834, n6832, n6833);
   and (n6835, n6811, n6831);
   nor (n6836, n6834, n6835);
   xnor (n6837, n6688, n6696);
   and (n6838, n6683, n6684);
   nor (n6839, n6838, n6685);
   not (n684, n674);
   and (n6840, n6717, n6718);
   nor (n6841, n6840, n6719);
   xor (n6842, n6839, n6841);
   xor (n6843, n6674, n6675);
   and (n6844, n6842, n6843);
   and (n6845, n6839, n6841);
   nor (n6846, n6844, n6845);
   xor (n6847, n6837, n6846);
   and (n6848, n6836, n6847);
   and (n6849, n6846, n6837);
   or (n685, n683, n684);
   nor (n6850, n6848, n6849);
   and (n6851, n6787, n6850);
   and (n6852, n6768, n6786);
   nor (n6853, n6851, n6852);
   not (n6854, n6853);
   and (n6855, n6704, n6711);
   and (n6856, n6701, n6703);
   nor (n6857, n6855, n6856);
   xor (n6858, n6610, n6617);
   not (n6859, n6858);
   or (n686, n674, n642);
   xnor (n6860, n6857, n6859);
   and (n6861, n6777, n6781);
   or (n6862, n6861, n6780);
   and (n6863, n6769, n6775);
   or (n6864, n6863, n6771);
   xor (n6865, n6862, n6864);
   xor (n6866, n6625, n6631);
   xnor (n6867, n6865, n6866);
   xor (n6868, n6860, n6867);
   not (n6869, n6782);
   nand (n687, n685, n686);
   not (n6870, n6776);
   or (n6871, n6869, n6870);
   or (n6872, n6783, n6785);
   nand (n6873, n6871, n6872);
   xor (n6874, n6868, n6873);
   or (n6875, n6767, n6713);
   or (n6876, n6699, n6712);
   nand (n6877, n6875, n6876);
   xor (n6878, n6874, n6877);
   not (n6879, n6878);
   not (n688, n687);
   and (n6880, n6854, n6879);
   and (n6881, n6853, n6878);
   nor (n6882, n6880, n6881);
   xnor (n6883, n6624, n6639);
   or (n6884, n6860, n6867);
   or (n6885, n6857, n6859);
   nand (n6886, n6884, n6885);
   xor (n6887, n6633, n6634);
   xor (n6888, n6887, n6636);
   and (n6889, n6865, n6866);
   not (n689, n688);
   and (n6890, n6862, n6864);
   nor (n6891, n6889, n6890);
   not (n6892, n6891);
   and (n6893, n6888, n6892);
   not (n6894, n6888);
   and (n6895, n6894, n6891);
   nor (n6896, n6893, n6895);
   and (n6897, n6886, n6896);
   and (n6898, n6888, n6892);
   nor (n6899, n6897, n6898);
   buf (n69, g68);
   and (n690, n38, n61);
   xnor (n6900, n6883, n6899);
   not (n6901, n6900);
   xor (n6902, n6886, n6896);
   not (n6903, n6902);
   and (n6904, n6874, n6877);
   and (n6905, n6868, n6873);
   nor (n6906, n6904, n6905);
   not (n6907, n6906);
   or (n6908, n6903, n6907);
   or (n6909, n6906, n6902);
   not (n691, n38);
   nand (n6910, n6908, n6909);
   nand (n6911, n6901, n6910);
   nor (n6912, n6882, n6911);
   not (n6913, n6912);
   xor (n6914, n6768, n6786);
   xor (n6915, n6914, n6850);
   not (n6916, n6915);
   nor (n6917, n6725, n6626);
   and (n6918, n73, n89);
   and (n6919, n74, n88);
   not (n692, n61);
   nor (n6920, n6918, n6919);
   nor (n6921, n6917, n6920);
   nand (n6922, n73, n79);
   not (n6923, n6922);
   nand (n6924, n6923, n84, n90);
   not (n6925, n6924);
   and (n6926, n73, n90);
   and (n6927, n79, n84);
   nor (n6928, n6926, n6927);
   nor (n6929, n6925, n6928);
   and (n693, n691, n692);
   not (n6930, n74);
   nor (n6931, n6930, n6357);
   nand (n6932, n6929, n6931);
   nand (n6933, n6932, n6924);
   and (n6934, n6921, n6933);
   or (n6935, n6934, n6917);
   xor (n6936, n6733, n6740);
   nor (n6937, n6817, n6646);
   and (n6938, n77, n86);
   and (n6939, n78, n85);
   nor (n694, n690, n693);
   nor (n6940, n6938, n6939);
   nor (n6941, n6937, n6940);
   nor (n6942, n6292, n6577);
   nand (n6943, n6941, n6942);
   not (n6944, n6943);
   or (n6945, n6944, n6937);
   nand (n6946, n75, n88);
   nand (n6947, n76, n87);
   and (n6948, n6946, n6947);
   nor (n6949, n6669, n6584);
   not (n695, n694);
   nor (n6950, n6948, n6949);
   and (n6951, n72, n91);
   and (n6952, n6950, n6951);
   or (n6953, n6952, n6949);
   nand (n6954, n71, n92);
   not (n6955, n6954);
   nand (n6956, n6582, n94, n95);
   not (n6957, n6956);
   and (n6958, n68, n95);
   and (n6959, n69, n94);
   not (n696, n495);
   nor (n6960, n6958, n6959);
   nor (n6961, n6957, n6960);
   nand (n6962, n6955, n6961);
   nand (n6963, n6962, n6956);
   xor (n6964, n6953, n6963);
   and (n6965, n6945, n6964);
   and (n6966, n6953, n6963);
   or (n6967, n6965, n6966);
   xor (n6968, n6936, n6967);
   and (n6969, n6935, n6968);
   or (n697, n695, n696);
   and (n6970, n6936, n6967);
   nor (n6971, n6969, n6970);
   xnor (n6972, n6842, n6843);
   or (n6973, n6971, n6972);
   nand (n6974, n6971, n6972);
   nand (n6975, n6973, n6974);
   not (n6976, n6975);
   or (n6977, n6800, n6809);
   nand (n6978, n6977, n6810);
   xor (n6979, n6802, n6807);
   nand (n698, n311, n649);
   xor (n6980, n6816, n6822);
   xor (n6981, n6979, n6980);
   and (n6982, n6792, n6793);
   nor (n6983, n6982, n6794);
   and (n6984, n6981, n6983);
   and (n6985, n6979, n6980);
   nor (n6986, n6984, n6985);
   xor (n6987, n6978, n6986);
   xnor (n6988, n6827, n6812);
   and (n6989, n6987, n6988);
   nand (n699, n697, n698);
   and (n6990, n6978, n6986);
   nor (n6991, n6989, n6990);
   not (n6992, n6991);
   and (n6993, n6976, n6992);
   not (n6994, n6974);
   nor (n6995, n6993, n6994);
   xnor (n6996, n6836, n6847);
   xor (n6997, n6732, n6765);
   xor (n6998, n6996, n6997);
   and (n6999, n6995, n6998);
   buf (n7, g6);
   buf (n70, g69);
   and (n700, n48, n52);
   and (n7000, n6996, n6997);
   nor (n7001, n6999, n7000);
   not (n7002, n7001);
   or (n7003, n6916, n7002);
   or (n7004, n7001, n6915);
   nand (n7005, n7003, n7004);
   not (n7006, n7005);
   xnor (n7007, n6995, n6998);
   not (n7008, n7007);
   xor (n7009, n6975, n6991);
   not (n701, n48);
   xnor (n7010, n6832, n6833);
   xor (n7011, n7009, n7010);
   xor (n7012, n6945, n6964);
   xor (n7013, n6921, n6933);
   xor (n7014, n7012, n7013);
   nand (n7015, n72, n92);
   not (n7016, n7015);
   not (n7017, n7016);
   nand (n7018, n76, n88);
   nand (n7019, n75, n89);
   and (n702, n701, n267);
   and (n7020, n7018, n7019);
   nor (n7021, n6669, n6626);
   nor (n7022, n7020, n7021);
   not (n7023, n7022);
   or (n7024, n7017, n7023);
   not (n7025, n7021);
   nand (n7026, n7024, n7025);
   and (n7027, n73, n91);
   and (n7028, n79, n85);
   nor (n7029, n7027, n7028);
   nor (n703, n700, n702);
   not (n7030, n7029);
   nand (n7031, n6923, n85, n91);
   nand (n7032, n7030, n7031);
   nand (n7033, n80, n84);
   nor (n7034, n7032, n7033);
   not (n7035, n7034);
   nand (n7036, n7035, n7031);
   nand (n7037, n95, n96);
   nor (n7038, n6581, n7037);
   not (n7039, n7038);
   not (n704, n703);
   nand (n7040, n71, n93);
   not (n7041, n7040);
   and (n7042, n68, n96);
   and (n7043, n69, n95);
   nor (n7044, n7042, n7043);
   nor (n7045, n7038, n7044);
   nand (n7046, n7041, n7045);
   nand (n7047, n7039, n7046);
   xor (n7048, n7036, n7047);
   and (n7049, n7026, n7048);
   nand (n705, n48, n49);
   and (n7050, n7036, n7047);
   nor (n7051, n7049, n7050);
   not (n7052, n7051);
   and (n7053, n7014, n7052);
   and (n7054, n7012, n7013);
   or (n7055, n7053, n7054);
   xor (n7056, n6935, n6968);
   xnor (n7057, n7055, n7056);
   xnor (n7058, n6987, n6988);
   or (n7059, n7057, n7058);
   not (n706, n705);
   or (n7060, n7055, n7056);
   nand (n7061, n7059, n7060);
   and (n7062, n7011, n7061);
   and (n7063, n7009, n7010);
   nor (n7064, n7062, n7063);
   not (n7065, n7064);
   or (n7066, n7008, n7065);
   or (n7067, n7064, n7007);
   nand (n7068, n7066, n7067);
   not (n7069, n7068);
   and (n707, n50, n49);
   xor (n7070, n7057, n7058);
   xor (n7071, n6981, n6983);
   or (n7072, n6941, n6942);
   nand (n7073, n7072, n6943);
   and (n7074, n70, n94);
   nor (n7075, n6817, n6594);
   and (n7076, n77, n87);
   and (n7077, n78, n86);
   nor (n7078, n7076, n7077);
   nor (n7079, n7075, n7078);
   not (n708, n50);
   and (n7080, n7074, n7079);
   nor (n7081, n7080, n7075);
   xor (n7082, n7073, n7081);
   or (n7083, n6929, n6931);
   nand (n7084, n7083, n6932);
   and (n7085, n7082, n7084);
   and (n7086, n7073, n7081);
   nor (n7087, n7085, n7086);
   xor (n7088, n7071, n7087);
   not (n7089, n6961);
   and (n709, n708, n48);
   nand (n7090, n7089, n6954);
   and (n7091, n6962, n7090);
   not (n7092, n6950);
   not (n7093, n6951);
   and (n7094, n7092, n7093);
   nor (n7095, n7094, n6952);
   and (n7096, n7091, n7095);
   xor (n7097, n7091, n7095);
   and (n7098, n80, n85);
   nor (n7099, n6324, n6073, n6922);
   buf (n71, g70);
   nor (n710, n707, n709);
   and (n7100, n73, n92);
   and (n7101, n79, n86);
   nor (n7102, n7100, n7101);
   nor (n7103, n7099, n7102);
   and (n7104, n7098, n7103);
   or (n7105, n7104, n7099);
   nor (n7106, n6930, n6084);
   and (n7107, n70, n95);
   nand (n7108, n77, n88);
   nand (n7109, n78, n87);
   nor (n711, n706, n710);
   and (n7110, n7108, n7109);
   nor (n7111, n6817, n6584);
   nor (n7112, n7110, n7111);
   and (n7113, n7107, n7112);
   or (n7114, n7113, n7111);
   xor (n7115, n7106, n7114);
   and (n7116, n7105, n7115);
   and (n7117, n7106, n7114);
   or (n7118, n7116, n7117);
   and (n7119, n7097, n7118);
   buf (n712, n711);
   nor (n7120, n7096, n7119);
   not (n7121, n7120);
   and (n7122, n7088, n7121);
   and (n7123, n7071, n7087);
   nor (n7124, n7122, n7123);
   xnor (n7125, n7070, n7124);
   xor (n7126, n7012, n7013);
   not (n7127, n7051);
   xor (n7128, n7126, n7127);
   not (n7129, n7045);
   not (n713, n712);
   nand (n7130, n7129, n7040);
   and (n7131, n7046, n7130);
   xor (n7132, n7074, n7079);
   xor (n7133, n7131, n7132);
   not (n7134, n7015);
   not (n7135, n7022);
   or (n7136, n7134, n7135);
   or (n7137, n7022, n7015);
   nand (n7138, n7136, n7137);
   and (n7139, n7133, n7138);
   or (n714, n704, n713);
   and (n7140, n7131, n7132);
   nor (n7141, n7139, n7140);
   xor (n7142, n7026, n7048);
   and (n7143, n7141, n7142);
   not (n7144, n7141);
   not (n7145, n7142);
   and (n7146, n7144, n7145);
   nor (n7147, n7143, n7146);
   nand (n7148, n96, n97);
   nor (n7149, n6581, n7148);
   nand (n715, n714, n615);
   not (n7150, n7149);
   nand (n7151, n71, n94);
   not (n7152, n7151);
   and (n7153, n68, n97);
   and (n7154, n69, n96);
   nor (n7155, n7153, n7154);
   nor (n7156, n7149, n7155);
   nand (n7157, n7152, n7156);
   nand (n7158, n7150, n7157);
   and (n7159, n75, n90);
   xor (n716, n699, n715);
   and (n7160, n76, n89);
   nor (n7161, n7159, n7160);
   not (n7162, n7161);
   not (n7163, n6770);
   nand (n7164, n7163, n6670);
   nand (n7165, n7162, n7164);
   nand (n7166, n72, n93);
   nor (n7167, n7165, n7166);
   not (n7168, n7167);
   nand (n7169, n7168, n7164);
   or (n717, n36, n63);
   xor (n7170, n7158, n7169);
   and (n7171, n7032, n7033);
   nor (n7172, n7171, n7034);
   and (n7173, n7170, n7172);
   and (n7174, n7158, n7169);
   nor (n7175, n7173, n7174);
   or (n7176, n7147, n7175);
   or (n7177, n7141, n7145);
   nand (n7178, n7176, n7177);
   xor (n7179, n7128, n7178);
   nand (n718, n36, n63);
   and (n7180, n7088, n7121);
   not (n7181, n7088);
   and (n7182, n7181, n7120);
   nor (n7183, n7180, n7182);
   and (n7184, n7179, n7183);
   and (n7185, n7128, n7178);
   nor (n7186, n7184, n7185);
   or (n7187, n7125, n7186);
   or (n7188, n7070, n7124);
   nand (n7189, n7187, n7188);
   nand (n719, n717, n718);
   not (n7190, n7189);
   xor (n7191, n7009, n7010);
   xor (n7192, n7191, n7061);
   not (n7193, n7192);
   or (n7194, n7190, n7193);
   or (n7195, n7192, n7189);
   nand (n7196, n7194, n7195);
   not (n7197, n7196);
   xor (n7198, n7125, n7186);
   not (n7199, n7198);
   buf (n72, g71);
   or (n720, n247, n719);
   nand (n7200, n70, n74);
   nand (n7201, n93, n97);
   nor (n7202, n7200, n7201);
   not (n7203, n7202);
   and (n7204, n70, n97);
   and (n7205, n74, n93);
   nor (n7206, n7204, n7205);
   nor (n7207, n7202, n7206);
   and (n7208, n82, n85);
   nand (n7209, n7207, n7208);
   or (n721, n36, n62);
   nand (n7210, n7203, n7209);
   nand (n7211, n68, n99);
   not (n7212, n7211);
   nand (n7213, n7212, n4);
   not (n7214, n7213);
   nand (n7215, n7210, n7214);
   not (n7216, n7215);
   or (n7217, n7210, n7214);
   nand (n7218, n7217, n7215);
   not (n7219, n6705);
   nand (n722, n721, n679);
   and (n7220, n83, n92);
   nand (n7221, n7219, n7220);
   not (n7222, n7221);
   and (n7223, n75, n92);
   and (n7224, n83, n84);
   nor (n7225, n7223, n7224);
   not (n7226, n7225);
   nand (n7227, n7226, n7221);
   nand (n7228, n71, n96);
   nor (n7229, n7227, n7228);
   or (n723, n402, n722);
   nor (n7230, n7222, n7229);
   nor (n7231, n7218, n7230);
   nor (n7232, n7216, n7231);
   not (n7233, n7232);
   not (n7234, n7233);
   and (n7235, n76, n90);
   nand (n7236, n6734, n7235);
   not (n7237, n77);
   not (n7238, n90);
   or (n7239, n7237, n7238);
   nand (n724, n720, n723);
   nand (n7240, n76, n91);
   nand (n7241, n7239, n7240);
   nand (n7242, n7236, n7241);
   nand (n7243, n69, n98);
   or (n7244, n7242, n7243);
   nand (n7245, n7244, n7236);
   nand (n7246, n78, n95);
   nor (n7247, n6750, n7246);
   not (n7248, n7247);
   and (n7249, n72, n95);
   and (n725, n716, n724);
   and (n7250, n78, n89);
   nor (n7251, n7249, n7250);
   nor (n7252, n7247, n7251);
   and (n7253, n79, n88);
   nand (n7254, n7252, n7253);
   nand (n7255, n7248, n7254);
   nand (n7256, n7245, n7255);
   not (n7257, n7256);
   or (n7258, n7245, n7255);
   nand (n7259, n7258, n7256);
   and (n726, n699, n715);
   and (n7260, n81, n86);
   nand (n7261, n80, n94);
   nor (n7262, n7261, n6715);
   and (n7263, n73, n94);
   and (n7264, n80, n87);
   nor (n7265, n7263, n7264);
   nor (n7266, n7262, n7265);
   and (n7267, n7260, n7266);
   nor (n7268, n7267, n7262);
   nor (n7269, n7259, n7268);
   nor (n727, n725, n726);
   nor (n7270, n7257, n7269);
   not (n7271, n7270);
   not (n7272, n7271);
   or (n7273, n7234, n7272);
   nand (n7274, n7270, n7232);
   nand (n7275, n7273, n7274);
   and (n7276, n73, n93);
   and (n7277, n79, n87);
   nor (n7278, n7276, n7277);
   not (n7279, n7278);
   not (n728, n727);
   nand (n7280, n6923, n87, n93);
   nand (n7281, n7279, n7280);
   nand (n7282, n80, n86);
   nor (n7283, n7281, n7282);
   not (n7284, n7283);
   nand (n7285, n7284, n7280);
   and (n7286, n70, n96);
   nor (n7287, n6817, n6626);
   and (n7288, n77, n89);
   and (n7289, n78, n88);
   and (n729, n689, n728);
   nor (n7290, n7288, n7289);
   nor (n7291, n7287, n7290);
   and (n7292, n7286, n7291);
   or (n7293, n7292, n7287);
   and (n7294, n72, n94);
   nor (n7295, n6669, n6690);
   and (n7296, n75, n91);
   nor (n7297, n7296, n7235);
   nor (n7298, n7295, n7297);
   and (n7299, n7294, n7298);
   buf (n73, g72);
   not (n730, n727);
   or (n7300, n7299, n7295);
   xor (n7301, n7293, n7300);
   xor (n7302, n7285, n7301);
   or (n7303, n7275, n7302);
   nand (n7304, n7303, n7274);
   not (n7305, n7304);
   nand (n7306, n81, n91);
   nor (n7307, n6700, n7306);
   and (n7308, n74, n91);
   and (n7309, n81, n84);
   not (n731, n730);
   nor (n7310, n7308, n7309);
   nor (n7311, n7307, n7310);
   and (n7312, n82, n84);
   nand (n7313, n81, n92);
   nor (n7314, n7313, n6722);
   and (n7315, n74, n92);
   and (n7316, n81, n85);
   nor (n7317, n7315, n7316);
   nor (n7318, n7314, n7317);
   and (n7319, n7312, n7318);
   not (n732, n688);
   or (n7320, n7319, n7314);
   xor (n7321, n7311, n7320);
   xor (n7322, n7107, n7112);
   xor (n7323, n7098, n7103);
   xor (n7324, n7322, n7323);
   and (n7325, n7321, n7324);
   and (n7326, n7322, n7323);
   nor (n7327, n7325, n7326);
   not (n7328, n7327);
   and (n7329, n7305, n7328);
   or (n733, n731, n732);
   xor (n7330, n7304, n7327);
   and (n7331, n7311, n7320);
   or (n7332, n7331, n7307);
   and (n7333, n7285, n7301);
   and (n7334, n7293, n7300);
   or (n7335, n7333, n7334);
   xor (n7336, n7332, n7335);
   xor (n7337, n7105, n7115);
   xor (n7338, n7336, n7337);
   and (n7339, n7330, n7338);
   nand (n734, n687, n727);
   nor (n7340, n7329, n7339);
   xnor (n7341, n7147, n7175);
   nand (n7342, n6582, n97, n98);
   not (n7343, n7342);
   and (n7344, n68, n98);
   and (n7345, n69, n97);
   nor (n7346, n7344, n7345);
   not (n7347, n7346);
   nand (n7348, n7347, n7342);
   nand (n7349, n71, n95);
   nand (n735, n733, n734);
   nor (n7350, n7348, n7349);
   nor (n7351, n7343, n7350);
   not (n7352, n7166);
   not (n7353, n7165);
   or (n7354, n7352, n7353);
   not (n7355, n7167);
   nand (n7356, n7354, n7355);
   xor (n7357, n7351, n7356);
   not (n7358, n7151);
   not (n7359, n7156);
   not (n736, n420);
   not (n7360, n7359);
   or (n7361, n7358, n7360);
   nand (n7362, n7361, n7157);
   and (n7363, n7357, n7362);
   and (n7364, n7351, n7356);
   nor (n7365, n7363, n7364);
   xor (n7366, n7158, n7169);
   xor (n7367, n7366, n7172);
   xor (n7368, n7365, n7367);
   xor (n7369, n7133, n7138);
   buf (n737, n736);
   and (n7370, n7368, n7369);
   and (n7371, n7365, n7367);
   nor (n7372, n7370, n7371);
   xor (n7373, n7341, n7372);
   and (n7374, n7340, n7373);
   and (n7375, n7341, n7372);
   nor (n7376, n7374, n7375);
   xor (n7377, n7179, n7183);
   xor (n7378, n7073, n7081);
   xor (n7379, n7378, n7084);
   not (n738, n737);
   not (n7380, n7379);
   not (n7381, n7380);
   xor (n7382, n7097, n7118);
   not (n7383, n7382);
   or (n7384, n7381, n7383);
   xor (n7385, n7332, n7335);
   and (n7386, n7385, n7337);
   and (n7387, n7332, n7335);
   nor (n7388, n7386, n7387);
   xnor (n7389, n7382, n7380);
   and (n739, n738, n605);
   or (n7390, n7388, n7389);
   nand (n7391, n7384, n7390);
   xnor (n7392, n7377, n7391);
   or (n7393, n7376, n7392);
   or (n7394, n7377, n7391);
   nand (n7395, n7393, n7394);
   not (n7396, n7395);
   or (n7397, n7199, n7396);
   or (n7398, n7395, n7198);
   nand (n7399, n7397, n7398);
   buf (n74, g73);
   and (n740, n423, n377);
   not (n7400, n7399);
   xor (n7401, n7392, n7376);
   not (n7402, n7401);
   xor (n7403, n7373, n7340);
   xnor (n7404, n7388, n7389);
   xor (n7405, n7403, n7404);
   and (n7406, n7275, n7302);
   not (n7407, n7275);
   not (n7408, n7302);
   and (n7409, n7407, n7408);
   and (n741, n42, n55);
   nor (n7410, n7406, n7409);
   xor (n7411, n7286, n7291);
   and (n7412, n7281, n7282);
   nor (n7413, n7412, n7283);
   and (n7414, n7411, n7413);
   xor (n7415, n7411, n7413);
   nand (n7416, n79, n80);
   nor (n7417, n6626, n7416);
   not (n7418, n7417);
   and (n7419, n79, n89);
   nor (n742, n740, n741);
   and (n7420, n80, n88);
   nor (n7421, n7419, n7420);
   nor (n7422, n7417, n7421);
   and (n7423, n74, n94);
   nand (n7424, n7422, n7423);
   nand (n7425, n7418, n7424);
   not (n7426, n7425);
   nand (n7427, n78, n98);
   nor (n7428, n7427, n6714);
   not (n7429, n7428);
   and (n743, n430, n742);
   and (n7430, n70, n98);
   and (n7431, n78, n90);
   nor (n7432, n7430, n7431);
   nor (n7433, n7428, n7432);
   and (n7434, n73, n95);
   nand (n7435, n7433, n7434);
   nand (n7436, n7429, n7435);
   nand (n7437, n76, n96);
   nor (n7438, n7015, n7437);
   not (n7439, n7438);
   nor (n744, n739, n743);
   and (n7440, n72, n96);
   and (n7441, n76, n92);
   nor (n7442, n7440, n7441);
   nor (n7443, n7438, n7442);
   nand (n7444, n7443, n6734);
   nand (n7445, n7439, n7444);
   or (n7446, n7436, n7445);
   nand (n7447, n7445, n7436);
   nand (n7448, n7446, n7447);
   nor (n7449, n7426, n7448);
   not (n745, n722);
   not (n7450, n7447);
   or (n7451, n7449, n7450);
   and (n7452, n7415, n7451);
   nor (n7453, n7414, n7452);
   xnor (n7454, n7410, n7453);
   and (n7455, n7259, n7268);
   nor (n7456, n7455, n7269);
   not (n7457, n4);
   not (n7458, n7457);
   not (n7459, n7211);
   not (n746, n745);
   or (n7460, n7458, n7459);
   nand (n7461, n7460, n7213);
   and (n7462, n69, n99);
   nand (n7463, n7462, n5);
   or (n7464, n7461, n7463);
   nand (n7465, n71, n75);
   nor (n7466, n7201, n7465);
   not (n7467, n7466);
   and (n7468, n71, n97);
   and (n7469, n75, n93);
   and (n747, n243, n244);
   nor (n7470, n7468, n7469);
   nor (n7471, n7466, n7470);
   and (n7472, n83, n85);
   nand (n7473, n7471, n7472);
   nand (n7474, n7467, n7473);
   not (n7475, n7463);
   not (n7476, n7475);
   not (n7477, n7461);
   or (n7478, n7476, n7477);
   or (n7479, n7461, n7475);
   not (n748, n747);
   nand (n7480, n7478, n7479);
   nand (n7481, n7474, n7480);
   nand (n7482, n7464, n7481);
   xor (n7483, n7456, n7482);
   and (n7484, n7218, n7230);
   nor (n7485, n7484, n7231);
   and (n7486, n7483, n7485);
   and (n7487, n7456, n7482);
   nor (n7488, n7486, n7487);
   or (n7489, n7454, n7488);
   or (n749, n746, n748);
   or (n7490, n7410, n7453);
   nand (n7491, n7489, n7490);
   xor (n7492, n7365, n7367);
   xor (n7493, n7492, n7369);
   xor (n7494, n7324, n7321);
   not (n7495, n7494);
   xor (n7496, n7294, n7298);
   and (n7497, n7348, n7349);
   nor (n7498, n7497, n7350);
   xor (n7499, n7496, n7498);
   buf (n75, g74);
   or (n750, n36, n61);
   xor (n7500, n7312, n7318);
   and (n7501, n7499, n7500);
   and (n7502, n7496, n7498);
   nor (n7503, n7501, n7502);
   xor (n7504, n7351, n7356);
   xor (n7505, n7504, n7362);
   xor (n7506, n7503, n7505);
   not (n7507, n7506);
   or (n7508, n7495, n7507);
   or (n7509, n7503, n7505);
   nand (n751, n36, n61);
   nand (n7510, n7508, n7509);
   xor (n7511, n7493, n7510);
   and (n7512, n7491, n7511);
   and (n7513, n7493, n7510);
   nor (n7514, n7512, n7513);
   and (n7515, n7405, n7514);
   and (n7516, n7403, n7404);
   nor (n7517, n7515, n7516);
   not (n7518, n7517);
   or (n7519, n7402, n7518);
   nand (n752, n750, n751);
   or (n7520, n7517, n7401);
   nand (n7521, n7519, n7520);
   not (n7522, n7521);
   xor (n7523, n7403, n7404);
   xor (n7524, n7523, n7514);
   not (n7525, n7524);
   xor (n7526, n7491, n7511);
   xnor (n7527, n7330, n7338);
   xnor (n7528, n7526, n7527);
   xor (n7529, n7454, n7488);
   not (n753, n752);
   xor (n7530, n7506, n7494);
   or (n7531, n7207, n7208);
   and (n7532, n7209, n7531);
   xor (n7533, n7260, n7266);
   xor (n7534, n7532, n7533);
   and (n7535, n7227, n7228);
   nor (n7536, n7535, n7229);
   and (n7537, n7534, n7536);
   and (n7538, n7532, n7533);
   nor (n7539, n7537, n7538);
   nand (n754, n753, n252);
   not (n7540, n7539);
   not (n7541, n6);
   nand (n7542, n70, n99);
   nor (n7543, n7541, n7542);
   not (n7544, n7543);
   not (n7545, n6594);
   nand (n7546, n7545, n81, n82);
   not (n7547, n87);
   not (n7548, n81);
   or (n7549, n7547, n7548);
   nand (n755, n749, n754);
   nand (n7550, n82, n86);
   nand (n7551, n7549, n7550);
   and (n7552, n7546, n7551);
   not (n7553, n7552);
   or (n7554, n7544, n7553);
   nand (n7555, n7554, n7546);
   not (n7556, n7555);
   or (n7557, n7252, n7253);
   and (n7558, n7254, n7557);
   nand (n7559, n7242, n7243);
   and (n756, n755, n718);
   and (n7560, n7559, n7244);
   xor (n7561, n7558, n7560);
   not (n7562, n7561);
   or (n7563, n7556, n7562);
   nand (n7564, n7560, n7558);
   nand (n7565, n7563, n7564);
   not (n7566, n7565);
   and (n7567, n7540, n7566);
   and (n7568, n7565, n7539);
   nor (n7569, n7567, n7568);
   not (n757, n755);
   xnor (n7570, n7499, n7500);
   or (n7571, n7569, n7570);
   not (n7572, n7565);
   or (n7573, n7572, n7539);
   nand (n7574, n7571, n7573);
   xor (n7575, n7530, n7574);
   and (n7576, n7529, n7575);
   and (n7577, n7530, n7574);
   nor (n7578, n7576, n7577);
   and (n7579, n7528, n7578);
   not (n758, n718);
   xnor (n7580, n7491, n7511);
   and (n7581, n7580, n7527);
   nor (n7582, n7579, n7581);
   not (n7583, n7582);
   or (n7584, n7525, n7583);
   or (n7585, n7582, n7524);
   nand (n7586, n7584, n7585);
   not (n7587, n7586);
   xor (n7588, n7578, n7528);
   not (n7589, n7588);
   and (n759, n757, n758);
   xor (n7590, n7569, n7570);
   xor (n7591, n7456, n7482);
   xor (n7592, n7591, n7485);
   xor (n7593, n7590, n7592);
   not (n7594, n7543);
   not (n7595, n6);
   nand (n7596, n7595, n7542);
   nand (n7597, n7594, n7596);
   nand (n7598, n83, n86);
   nor (n7599, n7597, n7598);
   buf (n76, g75);
   nor (n760, n756, n759);
   not (n7600, n7599);
   not (n7601, n7599);
   nand (n7602, n7597, n7598);
   nand (n7603, n7601, n7602);
   not (n7604, n7603);
   nand (n7605, n71, n99);
   not (n7606, n7605);
   nand (n7607, n7606, n7);
   not (n7608, n7607);
   nand (n7609, n7604, n7608);
   xor (n761, n744, n760);
   nand (n7610, n7600, n7609);
   not (n7611, n7610);
   xnor (n7612, n7552, n7543);
   or (n7613, n7611, n7612);
   nand (n7614, n93, n97);
   nand (n7615, n73, n77);
   nor (n7616, n7614, n7615);
   not (n7617, n7616);
   and (n7618, n73, n97);
   and (n7619, n77, n93);
   and (n762, n735, n761);
   nor (n7620, n7618, n7619);
   nor (n7621, n7616, n7620);
   and (n7622, n78, n92);
   nand (n7623, n7621, n7622);
   nand (n7624, n7617, n7623);
   nand (n7625, n91, n96);
   nand (n7626, n74, n79);
   nor (n7627, n7625, n7626);
   not (n7628, n7627);
   and (n7629, n74, n96);
   nor (n763, n729, n762);
   and (n7630, n79, n91);
   nor (n7631, n7629, n7630);
   nor (n7632, n7627, n7631);
   and (n7633, n80, n90);
   nand (n7634, n7632, n7633);
   nand (n7635, n7628, n7634);
   or (n7636, n7624, n7635);
   nand (n7637, n7635, n7624);
   nand (n7638, n7636, n7637);
   and (n7639, n83, n87);
   and (n764, n682, n763);
   nand (n7640, n82, n94);
   nor (n7641, n7640, n7018);
   and (n7642, n76, n94);
   and (n7643, n82, n88);
   nor (n7644, n7642, n7643);
   nor (n7645, n7641, n7644);
   and (n7646, n7639, n7645);
   nor (n7647, n7646, n7641);
   or (n7648, n7638, n7647);
   nand (n7649, n7648, n7637);
   and (n765, n636, n681);
   not (n7650, n7612);
   not (n7651, n7610);
   or (n7652, n7650, n7651);
   or (n7653, n7610, n7612);
   nand (n7654, n7652, n7653);
   nand (n7655, n7649, n7654);
   nand (n7656, n7613, n7655);
   xor (n7657, n7532, n7533);
   xor (n7658, n7657, n7536);
   xor (n7659, n7656, n7658);
   nor (n766, n764, n765);
   nand (n7660, n81, n94);
   nor (n7661, n7660, n6946);
   and (n7662, n75, n94);
   and (n7663, n81, n88);
   nor (n7664, n7662, n7663);
   nor (n7665, n7661, n7664);
   and (n7666, n82, n87);
   nor (n7667, n7665, n7666);
   not (n7668, n7667);
   nand (n7669, n7665, n7666);
   and (n767, n38, n58);
   nand (n7670, n7668, n7669);
   nand (n7671, n95, n98);
   nand (n7672, n72, n75);
   nor (n7673, n7671, n7672);
   and (n7674, n72, n98);
   and (n7675, n75, n95);
   nor (n7676, n7674, n7675);
   nor (n7677, n7673, n7676);
   and (n7678, n81, n89);
   nand (n7679, n7677, n7678);
   not (n768, n38);
   not (n7680, n7673);
   and (n7681, n7679, n7680);
   nor (n7682, n7670, n7681);
   not (n7683, n7682);
   and (n7684, n7670, n7681);
   nor (n7685, n7684, n7682);
   nand (n7686, n77, n92);
   not (n7687, n7686);
   nand (n7688, n72, n76);
   nor (n7689, n7201, n7688);
   not (n769, n58);
   and (n7690, n72, n97);
   and (n7691, n76, n93);
   nor (n7692, n7690, n7691);
   nor (n7693, n7689, n7692);
   nand (n7694, n7687, n7693);
   not (n7695, n7693);
   nand (n7696, n7695, n7686);
   and (n7697, n7694, n7696);
   nand (n7698, n7685, n7697);
   nand (n7699, n7683, n7698);
   buf (n77, g76);
   and (n770, n768, n769);
   not (n7700, n7699);
   or (n7701, n7462, n5);
   nand (n7702, n7701, n7463);
   not (n7703, n7702);
   nand (n7704, n73, n78);
   nor (n7705, n7704, n7625);
   not (n7706, n7705);
   nand (n7707, n79, n90);
   not (n7708, n7707);
   and (n7709, n73, n96);
   nor (n771, n767, n770);
   and (n7710, n78, n91);
   nor (n7711, n7709, n7710);
   nor (n7712, n7705, n7711);
   nand (n7713, n7708, n7712);
   nand (n7714, n7706, n7713);
   nor (n7715, n7703, n7714);
   not (n7716, n7715);
   not (n7717, n7702);
   nand (n7718, n7717, n7714);
   nand (n7719, n7716, n7718);
   not (n772, n771);
   not (n7720, n7689);
   and (n7721, n7694, n7720);
   nor (n7722, n7719, n7721);
   not (n7723, n7722);
   nand (n7724, n7719, n7721);
   nand (n7725, n7723, n7724);
   not (n7726, n7725);
   and (n7727, n7700, n7726);
   and (n7728, n7699, n7725);
   nor (n7729, n7727, n7728);
   not (n773, n651);
   nand (n7730, n95, n98);
   nand (n7731, n71, n74);
   nor (n7732, n7730, n7731);
   not (n7733, n7732);
   nand (n7734, n80, n89);
   not (n7735, n7734);
   and (n7736, n71, n98);
   and (n7737, n74, n95);
   nor (n7738, n7736, n7737);
   nor (n7739, n7732, n7738);
   or (n774, n772, n773);
   nand (n7740, n7735, n7739);
   nand (n7741, n7733, n7740);
   not (n7742, n7661);
   nand (n7743, n7742, n7669);
   xor (n7744, n7741, n7743);
   or (n7745, n7471, n7472);
   and (n7746, n7473, n7745);
   xor (n7747, n7744, n7746);
   not (n7748, n7747);
   or (n7749, n7729, n7748);
   nand (n775, n310, n500);
   not (n7750, n7699);
   or (n7751, n7750, n7725);
   nand (n7752, n7749, n7751);
   and (n7753, n7659, n7752);
   and (n7754, n7656, n7658);
   nor (n7755, n7753, n7754);
   not (n7756, n7755);
   and (n7757, n7593, n7756);
   and (n7758, n7590, n7592);
   or (n7759, n7757, n7758);
   nand (n776, n774, n775);
   not (n7760, n7759);
   not (n7761, n7718);
   nor (n7762, n7761, n7722);
   or (n7763, n7480, n7474);
   nand (n7764, n7763, n7481);
   nor (n7765, n7762, n7764);
   not (n7766, n7765);
   nand (n7767, n7762, n7764);
   nand (n7768, n7766, n7767);
   not (n7769, n7424);
   not (n777, n776);
   nor (n7770, n7422, n7423);
   nor (n7771, n7769, n7770);
   not (n7772, n6735);
   not (n7773, n7443);
   or (n7774, n7772, n7773);
   or (n7775, n7443, n6735);
   nand (n7776, n7774, n7775);
   xor (n7777, n7771, n7776);
   or (n7778, n7433, n7434);
   and (n7779, n7435, n7778);
   or (n778, n36, n60);
   and (n7780, n7777, n7779);
   and (n7781, n7771, n7776);
   nor (n7782, n7780, n7781);
   nor (n7783, n7768, n7782);
   or (n7784, n7783, n7765);
   xor (n7785, n7415, n7451);
   xor (n7786, n7784, n7785);
   not (n7787, n7448);
   nor (n7788, n7787, n7425);
   nor (n7789, n7449, n7788);
   nand (n779, n778, n464);
   not (n7790, n7789);
   xor (n7791, n7741, n7743);
   and (n7792, n7791, n7746);
   and (n7793, n7741, n7743);
   nor (n7794, n7792, n7793);
   not (n7795, n7794);
   and (n7796, n7790, n7795);
   and (n7797, n7789, n7794);
   nor (n7798, n7796, n7797);
   xor (n7799, n7561, n7555);
   buf (n78, g77);
   not (n780, n779);
   not (n7800, n7799);
   or (n7801, n7798, n7800);
   not (n7802, n7789);
   or (n7803, n7794, n7802);
   nand (n7804, n7801, n7803);
   and (n7805, n7786, n7804);
   and (n7806, n7784, n7785);
   nor (n7807, n7805, n7806);
   xnor (n7808, n7760, n7807);
   xnor (n7809, n7529, n7575);
   not (n781, n780);
   or (n7810, n7808, n7809);
   or (n7811, n7760, n7807);
   nand (n7812, n7810, n7811);
   not (n7813, n7812);
   or (n7814, n7589, n7813);
   or (n7815, n7588, n7812);
   nand (n7816, n7814, n7815);
   not (n7817, n7816);
   xor (n7818, n7808, n7809);
   not (n7819, n7818);
   not (n782, n747);
   xor (n7820, n7786, n7804);
   and (n7821, n7798, n7799);
   not (n7822, n7798);
   and (n7823, n7822, n7800);
   nor (n7824, n7821, n7823);
   xor (n7825, n7782, n7768);
   and (n7826, n7824, n7825);
   not (n7827, n7824);
   not (n7828, n7825);
   and (n7829, n7827, n7828);
   or (n783, n781, n782);
   or (n7830, n7826, n7829);
   not (n7831, n7830);
   xor (n7832, n7771, n7776);
   xor (n7833, n7832, n7779);
   not (n7834, n7739);
   nand (n7835, n7834, n7734);
   and (n7836, n7740, n7835);
   not (n7837, n7707);
   not (n7838, n7712);
   not (n7839, n7838);
   not (n784, n459);
   or (n7840, n7837, n7839);
   nand (n7841, n7840, n7713);
   not (n7842, n7841);
   and (n7843, n7836, n7842);
   not (n7844, n7836);
   and (n7845, n7844, n7841);
   nor (n7846, n7843, n7845);
   not (n7847, n7608);
   not (n7848, n7603);
   or (n7849, n7847, n7848);
   nand (n785, n784, n252);
   or (n7850, n7603, n7608);
   nand (n7851, n7849, n7850);
   and (n7852, n7846, n7851);
   and (n7853, n7842, n7836);
   nor (n7854, n7852, n7853);
   not (n7855, n7854);
   and (n7856, n7833, n7855);
   not (n7857, n7833);
   and (n7858, n7857, n7854);
   nor (n7859, n7856, n7858);
   nand (n786, n783, n785);
   not (n7860, n7654);
   not (n7861, n7649);
   and (n7862, n7860, n7861);
   not (n7863, n7655);
   nor (n7864, n7862, n7863);
   and (n7865, n7859, n7864);
   and (n7866, n7833, n7855);
   nor (n7867, n7865, n7866);
   or (n7868, n7831, n7867);
   or (n7869, n7824, n7828);
   not (n787, n786);
   nand (n7870, n7868, n7869);
   xor (n7871, n7820, n7870);
   xnor (n7872, n7590, n7592);
   xor (n7873, n7872, n7755);
   and (n7874, n7871, n7873);
   and (n7875, n7820, n7870);
   nor (n7876, n7874, n7875);
   not (n7877, n7876);
   or (n7878, n7819, n7877);
   or (n7879, n7818, n7876);
   not (n788, n787);
   nand (n7880, n7878, n7879);
   not (n7881, n7880);
   xor (n7882, n7786, n7804);
   xnor (n7883, n7882, n7870);
   xor (n7884, n7883, n7873);
   not (n7885, n7867);
   not (n7886, n7830);
   or (n7887, n7885, n7886);
   or (n7888, n7830, n7867);
   nand (n7889, n7887, n7888);
   or (n789, n777, n788);
   xor (n7890, n7659, n7752);
   xor (n7891, n7889, n7890);
   and (n7892, n7729, n7747);
   not (n7893, n7729);
   and (n7894, n7893, n7748);
   nor (n7895, n7892, n7894);
   not (n7896, n7);
   not (n7897, n7896);
   not (n7898, n7605);
   or (n7899, n7897, n7898);
   buf (n79, g78);
   or (n790, n776, n787);
   nand (n7900, n7899, n7607);
   and (n7901, n72, n99);
   nand (n7902, n7901, n8);
   or (n7903, n7900, n7902);
   nand (n7904, n74, n78);
   nor (n7905, n7614, n7904);
   not (n7906, n7905);
   nand (n7907, n79, n92);
   not (n7908, n7907);
   and (n7909, n74, n97);
   nand (n791, n789, n790);
   and (n7910, n78, n93);
   nor (n7911, n7909, n7910);
   nor (n7912, n7905, n7911);
   nand (n7913, n7908, n7912);
   nand (n7914, n7906, n7913);
   xor (n7915, n7900, n7902);
   nand (n7916, n7914, n7915);
   nand (n7917, n7903, n7916);
   or (n7918, n7632, n7633);
   and (n7919, n7634, n7918);
   and (n792, n44, n52);
   or (n7920, n7621, n7622);
   and (n7921, n7623, n7920);
   xor (n7922, n7919, n7921);
   or (n7923, n7677, n7678);
   and (n7924, n7679, n7923);
   and (n7925, n7922, n7924);
   and (n7926, n7919, n7921);
   nor (n7927, n7925, n7926);
   not (n7928, n7927);
   and (n7929, n7917, n7928);
   not (n793, n44);
   not (n7930, n7917);
   and (n7931, n7930, n7927);
   nor (n7932, n7929, n7931);
   nand (n7933, n73, n76);
   nor (n7934, n7671, n7933);
   not (n7935, n7934);
   and (n7936, n73, n98);
   and (n7937, n76, n95);
   nor (n7938, n7936, n7937);
   nor (n7939, n7934, n7938);
   and (n794, n793, n267);
   and (n7940, n82, n89);
   nand (n7941, n7939, n7940);
   nand (n7942, n7935, n7941);
   nand (n7943, n75, n80);
   nor (n7944, n7625, n7943);
   not (n7945, n7944);
   nand (n7946, n81, n90);
   not (n7947, n7946);
   and (n7948, n75, n96);
   and (n7949, n80, n91);
   nor (n795, n792, n794);
   nor (n7950, n7948, n7949);
   nor (n7951, n7944, n7950);
   nand (n7952, n7947, n7951);
   nand (n7953, n7945, n7952);
   or (n7954, n7942, n7953);
   nand (n7955, n7953, n7942);
   nand (n7956, n7954, n7955);
   xor (n7957, n7639, n7645);
   not (n7958, n7957);
   or (n7959, n7956, n7958);
   not (n796, n795);
   nand (n7960, n7959, n7955);
   and (n7961, n7932, n7960);
   and (n7962, n7928, n7917);
   nor (n7963, n7961, n7962);
   xnor (n7964, n7895, n7963);
   or (n7965, n7914, n7915);
   nand (n7966, n7965, n7916);
   not (n7967, n7966);
   not (n7968, n7967);
   not (n7969, n7437);
   not (n797, n565);
   not (n7970, n7306);
   or (n7971, n7969, n7970);
   nand (n7972, n91, n96, n76, n81);
   nand (n7973, n7971, n7972);
   not (n7974, n7973);
   nand (n7975, n82, n90);
   not (n7976, n7975);
   nand (n7977, n7974, n7976);
   nand (n7978, n7977, n7972);
   nand (n7979, n73, n99);
   not (n798, n797);
   nor (n7980, n7979, n2918);
   nand (n7981, n7978, n7980);
   not (n7982, n7981);
   nor (n7983, n7978, n7980);
   nor (n7984, n7982, n7983);
   nand (n7985, n74, n77);
   nor (n7986, n7730, n7985);
   not (n7987, n7986);
   and (n7988, n74, n98);
   and (n7989, n77, n95);
   not (n799, n798);
   nor (n7990, n7988, n7989);
   nor (n7991, n7986, n7990);
   and (n7992, n83, n89);
   nand (n7993, n7991, n7992);
   nand (n7994, n7987, n7993);
   nand (n7995, n7984, n7994);
   nand (n7996, n7995, n7981);
   nand (n7997, n83, n94);
   nor (n7998, n7108, n7997);
   and (n7999, n77, n94);
   buf (n8, g7);
   buf (n80, g79);
   or (n800, n796, n799);
   and (n8000, n83, n88);
   nor (n8001, n7999, n8000);
   nor (n8002, n7998, n8001);
   not (n8003, n8002);
   or (n8004, n7901, n8);
   nand (n8005, n8004, n7902);
   or (n8006, n8003, n8005);
   not (n8007, n7998);
   nand (n8008, n8006, n8007);
   nand (n8009, n7996, n8008);
   nand (n801, n45, n46);
   or (n8010, n7996, n8008);
   and (n8011, n8009, n8010);
   not (n8012, n8011);
   or (n8013, n7968, n8012);
   nand (n8014, n8013, n8009);
   not (n8015, n7697);
   not (n8016, n7685);
   not (n8017, n8016);
   or (n8018, n8015, n8017);
   or (n8019, n8016, n7697);
   not (n802, n801);
   nand (n8020, n8018, n8019);
   nand (n8021, n7638, n7647);
   and (n8022, n7648, n8021);
   xor (n8023, n8020, n8022);
   and (n8024, n8014, n8023);
   and (n8025, n8020, n8022);
   nor (n8026, n8024, n8025);
   or (n8027, n7964, n8026);
   or (n8028, n7895, n7963);
   nand (n8029, n8027, n8028);
   nor (n803, n45, n46);
   and (n8030, n7891, n8029);
   and (n8031, n7889, n7890);
   nor (n8032, n8030, n8031);
   xor (n8033, n7884, n8032);
   not (n8034, n8033);
   xor (n8035, n7864, n7859);
   not (n8036, n8035);
   xor (n8037, n7846, n7851);
   not (n8038, n8037);
   not (n8039, n8038);
   nor (n804, n802, n803);
   xnor (n8040, n7924, n7922);
   not (n8041, n8040);
   not (n8042, n7957);
   not (n8043, n7956);
   or (n8044, n8042, n8043);
   or (n8045, n7956, n7957);
   nand (n8046, n8044, n8045);
   not (n8047, n8046);
   not (n8048, n7946);
   not (n8049, n7951);
   buf (n805, n804);
   not (n8050, n8049);
   or (n8051, n8048, n8050);
   nand (n8052, n8051, n7952);
   not (n8053, n8052);
   nand (n8054, n75, n79);
   nor (n8055, n7614, n8054);
   not (n8056, n8055);
   nand (n8057, n80, n92);
   not (n8058, n8057);
   and (n8059, n75, n97);
   or (n806, n805, n412);
   and (n8060, n79, n93);
   nor (n8061, n8059, n8060);
   nor (n8062, n8055, n8061);
   nand (n8063, n8058, n8062);
   nand (n8064, n8056, n8063);
   not (n8065, n8064);
   or (n8066, n7939, n7940);
   nand (n8067, n8066, n7941);
   nand (n8068, n8065, n8067);
   not (n8069, n8067);
   nand (n807, n800, n806);
   nand (n8070, n8069, n8064);
   and (n8071, n8068, n8070);
   not (n8072, n8071);
   or (n8073, n8053, n8072);
   nand (n8074, n8073, n8068);
   not (n8075, n8074);
   or (n8076, n8047, n8075);
   or (n8077, n8074, n8046);
   nand (n8078, n8076, n8077);
   not (n8079, n8078);
   xor (n808, n791, n807);
   or (n8080, n8041, n8079);
   not (n8081, n8046);
   nand (n8082, n8081, n8074);
   nand (n8083, n8080, n8082);
   not (n8084, n8083);
   or (n8085, n8039, n8084);
   xor (n8086, n7932, n7960);
   not (n8087, n8086);
   not (n8088, n8037);
   not (n8089, n8083);
   not (n809, n795);
   or (n8090, n8088, n8089);
   or (n8091, n8083, n8037);
   nand (n8092, n8090, n8091);
   nand (n8093, n8087, n8092);
   nand (n8094, n8085, n8093);
   not (n8095, n8094);
   or (n8096, n8036, n8095);
   or (n8097, n8094, n8035);
   nand (n8098, n8096, n8097);
   xor (n8099, n8026, n7964);
   buf (n81, g80);
   not (n810, n556);
   and (n8100, n8098, n8099);
   not (n8101, n8094);
   and (n8102, n8101, n8035);
   nor (n8103, n8100, n8102);
   not (n8104, n8103);
   xor (n8105, n7889, n7890);
   xor (n8106, n8105, n8029);
   not (n8107, n8106);
   or (n8108, n8104, n8107);
   or (n8109, n8106, n8103);
   or (n811, n809, n810);
   nand (n8110, n8108, n8109);
   not (n8111, n8110);
   xnor (n8112, n8011, n7966);
   not (n8113, n8112);
   not (n8114, n7980);
   not (n8115, n9);
   nand (n8116, n8115, n7979);
   nand (n8117, n8114, n8116);
   nand (n8118, n78, n94);
   nor (n8119, n8117, n8118);
   nand (n812, n566, n666);
   not (n8120, n8119);
   nand (n8121, n74, n99);
   not (n8122, n8121);
   nand (n8123, n8122, n10);
   not (n8124, n8123);
   not (n8125, n8119);
   nand (n8126, n8117, n8118);
   nand (n8127, n8125, n8126);
   not (n8128, n8127);
   nand (n8129, n8124, n8128);
   nand (n813, n811, n812);
   nand (n8130, n8120, n8129);
   not (n8131, n8130);
   not (n8132, n7907);
   not (n8133, n7912);
   not (n8134, n8133);
   or (n8135, n8132, n8134);
   nand (n8136, n8135, n7913);
   not (n8137, n8136);
   and (n8138, n8131, n8137);
   and (n8139, n8130, n8136);
   buf (n814, n533);
   nor (n8140, n8138, n8139);
   not (n8141, n8140);
   not (n8142, n8005);
   not (n8143, n8002);
   or (n8144, n8142, n8143);
   or (n8145, n8002, n8005);
   nand (n8146, n8144, n8145);
   and (n8147, n8141, n8146);
   not (n8148, n8136);
   and (n8149, n8130, n8148);
   buf (n815, n814);
   nor (n8150, n8147, n8149);
   not (n8151, n8150);
   or (n8152, n7984, n7994);
   nand (n8153, n8152, n7995);
   not (n8154, n8153);
   not (n8155, n8154);
   nand (n8156, n76, n80);
   nor (n8157, n7614, n8156);
   not (n8158, n8157);
   not (n8159, n7313);
   nand (n816, n815, n46);
   and (n8160, n76, n97);
   and (n8161, n80, n93);
   nor (n8162, n8160, n8161);
   nor (n8163, n8157, n8162);
   nand (n8164, n8159, n8163);
   nand (n8165, n8158, n8164);
   not (n8166, n8165);
   nand (n8167, n75, n78);
   nor (n8168, n7730, n8167);
   not (n8169, n8168);
   xor (n817, n813, n816);
   nand (n8170, n79, n94);
   not (n8171, n8170);
   nand (n8172, n75, n98);
   and (n8173, n7246, n8172);
   nor (n8174, n8173, n8168);
   nand (n8175, n8171, n8174);
   nand (n8176, n8169, n8175);
   not (n8177, n8176);
   or (n8178, n8166, n8177);
   xor (n8179, n8176, n8165);
   and (n818, n465, n640);
   nand (n8180, n77, n82);
   nor (n8181, n7625, n8180);
   not (n8182, n8181);
   nand (n8183, n83, n90);
   not (n8184, n8183);
   not (n8185, n91);
   not (n8186, n82);
   or (n8187, n8185, n8186);
   nand (n8188, n77, n96);
   nand (n8189, n8187, n8188);
   and (n819, n276, n479);
   not (n8190, n8189);
   nor (n8191, n8190, n8181);
   nand (n8192, n8184, n8191);
   nand (n8193, n8182, n8192);
   nand (n8194, n8179, n8193);
   nand (n8195, n8178, n8194);
   not (n8196, n8195);
   not (n8197, n8057);
   not (n8198, n8062);
   not (n8199, n8198);
   buf (n82, g81);
   and (n820, n40, n56);
   or (n8200, n8197, n8199);
   nand (n8201, n8200, n8063);
   not (n8202, n8201);
   or (n8203, n7991, n7992);
   nand (n8204, n8203, n7993);
   not (n8205, n8204);
   nand (n8206, n7973, n7975);
   and (n8207, n8206, n7977);
   not (n8208, n8207);
   or (n8209, n8205, n8208);
   nor (n821, n819, n820);
   or (n8210, n8207, n8204);
   nand (n8211, n8209, n8210);
   nand (n8212, n8202, n8211);
   not (n8213, n8204);
   nand (n8214, n8213, n8207);
   and (n8215, n8212, n8214);
   not (n8216, n8215);
   or (n8217, n8196, n8216);
   or (n8218, n8195, n8215);
   nand (n8219, n8217, n8218);
   and (n822, n274, n821);
   not (n8220, n8219);
   or (n8221, n8155, n8220);
   not (n8222, n8215);
   nand (n8223, n8222, n8195);
   nand (n8224, n8221, n8223);
   not (n8225, n8224);
   or (n8226, n8151, n8225);
   or (n8227, n8224, n8150);
   nand (n8228, n8226, n8227);
   not (n8229, n8228);
   nor (n823, n818, n822);
   or (n8230, n8113, n8229);
   not (n8231, n8150);
   nand (n8232, n8231, n8224);
   nand (n8233, n8230, n8232);
   not (n8234, n8233);
   not (n8235, n8023);
   xor (n8236, n8014, n8235);
   not (n8237, n8236);
   and (n8238, n8234, n8237);
   and (n8239, n8233, n8236);
   not (n824, n823);
   nor (n8240, n8238, n8239);
   not (n8241, n8086);
   not (n8242, n8092);
   or (n8243, n8241, n8242);
   or (n8244, n8092, n8086);
   nand (n8245, n8243, n8244);
   or (n8246, n8240, n8245);
   not (n8247, n8233);
   or (n8248, n8247, n8236);
   nand (n8249, n8246, n8248);
   and (n825, n817, n824);
   not (n8250, n8249);
   xnor (n8251, n8098, n8099);
   not (n8252, n8251);
   or (n8253, n8250, n8252);
   or (n8254, n8251, n8249);
   nand (n8255, n8253, n8254);
   not (n8256, n8255);
   xor (n8257, n8240, n8245);
   not (n8258, n8257);
   and (n8259, n8228, n8112);
   and (n826, n813, n816);
   not (n8260, n8228);
   not (n8261, n8112);
   and (n8262, n8260, n8261);
   nor (n8263, n8259, n8262);
   xnor (n8264, n8078, n8040);
   not (n8265, n8071);
   not (n8266, n8052);
   not (n8267, n8266);
   and (n8268, n8265, n8267);
   and (n8269, n8071, n8266);
   or (n827, n825, n826);
   nor (n8270, n8268, n8269);
   not (n8271, n8270);
   not (n8272, n8146);
   not (n8273, n8272);
   not (n8274, n8141);
   or (n8275, n8273, n8274);
   nand (n8276, n8140, n8146);
   nand (n8277, n8275, n8276);
   not (n8278, n8277);
   or (n8279, n8271, n8278);
   xor (n828, n808, n827);
   or (n8280, n8193, n8179);
   nand (n8281, n8280, n8194);
   not (n8282, n8281);
   not (n8283, n8123);
   not (n8284, n8128);
   or (n8285, n8283, n8284);
   not (n8286, n8123);
   nand (n8287, n8286, n8127);
   nand (n8288, n8285, n8287);
   not (n8289, n10);
   and (n829, n651, n657);
   not (n8290, n8289);
   not (n8291, n8121);
   or (n8292, n8290, n8291);
   nand (n8293, n8292, n8123);
   nand (n8294, n75, n99);
   not (n8295, n8294);
   nand (n8296, n8295, n11);
   or (n8297, n8293, n8296);
   nand (n8298, n78, n83);
   nor (n8299, n7625, n8298);
   buf (n83, g82);
   and (n830, n311, n771);
   not (n8300, n8299);
   nand (n8301, n76, n98);
   not (n8302, n8301);
   and (n8303, n78, n96);
   and (n8304, n83, n91);
   nor (n8305, n8303, n8304);
   nor (n8306, n8299, n8305);
   nand (n8307, n8302, n8306);
   nand (n8308, n8300, n8307);
   not (n8309, n8296);
   nor (n831, n829, n830);
   not (n8310, n8309);
   not (n8311, n8293);
   or (n8312, n8310, n8311);
   or (n8313, n8293, n8309);
   nand (n8314, n8312, n8313);
   nand (n8315, n8308, n8314);
   nand (n8316, n8297, n8315);
   xor (n8317, n8288, n8316);
   and (n8318, n8282, n8317);
   and (n8319, n8316, n8288);
   or (n832, n247, n752);
   nor (n8320, n8318, n8319);
   not (n8321, n8320);
   and (n8322, n8277, n8270);
   not (n8323, n8277);
   not (n8324, n8270);
   and (n8325, n8323, n8324);
   nor (n8326, n8322, n8325);
   nand (n8327, n8321, n8326);
   nand (n8328, n8279, n8327);
   xor (n8329, n8264, n8328);
   or (n833, n253, n779);
   and (n8330, n8263, n8329);
   and (n8331, n8328, n8264);
   nor (n8332, n8330, n8331);
   not (n8333, n8332);
   or (n8334, n8258, n8333);
   or (n8335, n8257, n8332);
   nand (n8336, n8334, n8335);
   not (n8337, n8336);
   not (n8338, n8163);
   not (n8339, n7313);
   nand (n834, n832, n833);
   and (n8340, n8338, n8339);
   and (n8341, n8163, n7313);
   nor (n8342, n8340, n8341);
   nand (n8343, n77, n81);
   nor (n8344, n7201, n8343);
   not (n8345, n8344);
   and (n8346, n77, n97);
   and (n8347, n81, n93);
   nor (n8348, n8346, n8347);
   not (n8349, n8348);
   and (n835, n831, n834);
   nand (n8350, n8345, n8349, n82, n92);
   not (n8351, n8344);
   and (n8352, n8350, n8351);
   xor (n8353, n8342, n8352);
   not (n8354, n8174);
   not (n8355, n8170);
   and (n8356, n8354, n8355);
   and (n8357, n8174, n8170);
   nor (n8358, n8356, n8357);
   and (n8359, n8353, n8358);
   not (n836, n831);
   and (n8360, n8342, n8352);
   nor (n8361, n8359, n8360);
   not (n8362, n8211);
   not (n8363, n8201);
   and (n8364, n8362, n8363);
   and (n8365, n8211, n8201);
   nor (n8366, n8364, n8365);
   and (n8367, n8361, n8366);
   not (n8368, n8361);
   not (n8369, n8366);
   not (n837, n834);
   and (n8370, n8368, n8369);
   or (n8371, n8367, n8370);
   nand (n8372, n79, n95);
   and (n8373, n7261, n8372);
   nand (n8374, n80, n95);
   nor (n8375, n8374, n8170);
   nor (n8376, n8373, n8375);
   not (n8377, n11);
   nand (n8378, n8377, n8294);
   nand (n8379, n8296, n8378);
   and (n838, n836, n837);
   not (n8380, n8379);
   and (n8381, n8376, n8380);
   nor (n8382, n8381, n8375);
   not (n8383, n8183);
   not (n8384, n8191);
   not (n8385, n8384);
   or (n8386, n8383, n8385);
   nand (n8387, n8386, n8192);
   not (n8388, n8387);
   and (n8389, n8382, n8388);
   nor (n839, n835, n838);
   not (n8390, n8382);
   and (n8391, n8390, n8387);
   nor (n8392, n8389, n8391);
   or (n8393, n8314, n8308);
   nand (n8394, n8393, n8315);
   or (n8395, n8392, n8394);
   or (n8396, n8382, n8387);
   nand (n8397, n8395, n8396);
   and (n8398, n8371, n8397);
   and (n8399, n8361, n8369);
   buf (n84, g83);
   and (n840, n422, n742);
   nor (n8400, n8398, n8399);
   and (n8401, n8219, n8153);
   not (n8402, n8219);
   and (n8403, n8402, n8154);
   nor (n8404, n8401, n8403);
   not (n8405, n8404);
   and (n8406, n8400, n8405);
   not (n8407, n8400);
   and (n8408, n8407, n8404);
   nor (n8409, n8406, n8408);
   and (n841, n423, n299);
   not (n8410, n8326);
   not (n8411, n8320);
   and (n8412, n8410, n8411);
   and (n8413, n8326, n8320);
   nor (n8414, n8412, n8413);
   or (n8415, n8409, n8414);
   not (n8416, n8405);
   or (n8417, n8400, n8416);
   nand (n8418, n8415, n8417);
   not (n8419, n8418);
   and (n842, n42, n54);
   xnor (n8420, n8263, n8329);
   not (n8421, n8420);
   or (n8422, n8419, n8421);
   or (n8423, n8420, n8418);
   nand (n8424, n8422, n8423);
   not (n8425, n8424);
   xor (n8426, n8317, n8281);
   not (n8427, n8426);
   nand (n8428, n79, n98);
   nor (n8429, n8188, n8428);
   nor (n843, n841, n842);
   not (n8430, n8429);
   not (n8431, n8374);
   and (n8432, n77, n98);
   and (n8433, n79, n96);
   nor (n8434, n8432, n8433);
   nor (n8435, n8429, n8434);
   nand (n8436, n8431, n8435);
   nand (n8437, n8430, n8436);
   not (n8438, n8437);
   nand (n8439, n76, n99);
   and (n844, n430, n843);
   not (n8440, n8439);
   nand (n8441, n8440, n12);
   not (n8442, n8441);
   and (n8443, n8438, n8442);
   and (n8444, n8437, n8441);
   nor (n8445, n8443, n8444);
   not (n8446, n97);
   not (n8447, n78);
   or (n8448, n8446, n8447);
   nand (n8449, n82, n93);
   nor (n845, n840, n844);
   nand (n8450, n8448, n8449);
   nand (n8451, n8450, n83, n92);
   not (n8452, n7614);
   nand (n8453, n8452, n78, n82);
   nand (n8454, n8451, n8453);
   not (n8455, n8454);
   or (n8456, n8445, n8455);
   not (n8457, n8437);
   or (n8458, n8457, n8441);
   nand (n8459, n8456, n8458);
   or (n846, n839, n845);
   not (n8460, n8459);
   xor (n8461, n8342, n8352);
   xor (n8462, n8461, n8358);
   not (n8463, n8462);
   or (n8464, n8460, n8463);
   or (n8465, n8462, n8459);
   nand (n8466, n8464, n8465);
   not (n8467, n8466);
   not (n8468, n82);
   not (n8469, n92);
   or (n847, n831, n837);
   or (n8470, n8468, n8469);
   or (n8471, n8344, n8348);
   nand (n8472, n8470, n8471);
   and (n8473, n8350, n8472);
   not (n8474, n8301);
   not (n8475, n8306);
   not (n8476, n8475);
   or (n8477, n8474, n8476);
   nand (n8478, n8477, n8307);
   not (n8479, n8478);
   nand (n848, n846, n847);
   and (n8480, n8473, n8479);
   not (n8481, n8473);
   and (n8482, n8481, n8478);
   nor (n8483, n8480, n8482);
   not (n8484, n12);
   nand (n8485, n8484, n8439);
   nand (n8486, n8441, n8485);
   xor (n8487, n8486, n7660);
   nand (n8488, n77, n99);
   not (n8489, n8488);
   xor (n849, n828, n848);
   nand (n8490, n8489, n13);
   and (n8491, n8487, n8490);
   and (n8492, n8486, n7660);
   nor (n8493, n8491, n8492);
   and (n8494, n8483, n8493);
   and (n8495, n8479, n8473);
   nor (n8496, n8494, n8495);
   not (n8497, n8496);
   not (n8498, n8497);
   or (n8499, n8467, n8498);
   buf (n85, g84);
   xor (n850, n766, n849);
   not (n8500, n8462);
   nand (n8501, n8500, n8459);
   nand (n8502, n8499, n8501);
   not (n8503, n8502);
   or (n8504, n8427, n8503);
   or (n8505, n8502, n8426);
   nand (n8506, n8504, n8505);
   xor (n8507, n8371, n8397);
   and (n8508, n8506, n8507);
   not (n8509, n8426);
   not (n851, n678);
   and (n8510, n8502, n8509);
   nor (n8511, n8508, n8510);
   not (n8512, n8511);
   xor (n8513, n8414, n8409);
   not (n8514, n8513);
   or (n8515, n8512, n8514);
   or (n8516, n8513, n8511);
   nand (n8517, n8515, n8516);
   not (n8518, n8517);
   xor (n8519, n8506, n8507);
   not (n852, n680);
   not (n8520, n8519);
   nand (n8521, n78, n81);
   nor (n8522, n7671, n8521);
   not (n8523, n8522);
   not (n8524, n95);
   not (n8525, n81);
   or (n8526, n8524, n8525);
   nand (n8527, n8526, n7427);
   not (n8528, n8527);
   nor (n8529, n8528, n8522);
   and (n853, n851, n852);
   not (n8530, n7640);
   nand (n8531, n8529, n8530);
   nand (n8532, n8523, n8531);
   nand (n8533, n79, n83);
   nor (n8534, n7201, n8533);
   not (n8535, n8534);
   nand (n8536, n80, n96);
   not (n8537, n8536);
   and (n8538, n79, n97);
   and (n8539, n83, n93);
   and (n854, n545, n679);
   nor (n8540, n8538, n8539);
   nor (n8541, n8534, n8540);
   nand (n8542, n8537, n8541);
   nand (n8543, n8535, n8542);
   nor (n8544, n8532, n8543);
   not (n8545, n8544);
   nand (n8546, n8532, n8543);
   nand (n8547, n8545, n8546);
   not (n8548, n8547);
   xnor (n8549, n8435, n8374);
   nor (n855, n853, n854);
   and (n8550, n8548, n8549);
   not (n8551, n8546);
   nor (n8552, n8550, n8551);
   not (n8553, n8552);
   not (n8554, n8379);
   not (n8555, n8376);
   or (n8556, n8554, n8555);
   or (n8557, n8376, n8379);
   nand (n8558, n8556, n8557);
   not (n8559, n8558);
   not (n856, n821);
   not (n8560, n8454);
   not (n8561, n8445);
   or (n8562, n8560, n8561);
   or (n8563, n8445, n8454);
   nand (n8564, n8562, n8563);
   not (n8565, n8564);
   not (n8566, n8565);
   or (n8567, n8559, n8566);
   not (n8568, n8558);
   nand (n8569, n8568, n8564);
   buf (n857, n265);
   nand (n8570, n8567, n8569);
   not (n8571, n8570);
   or (n8572, n8553, n8571);
   not (n8573, n8558);
   nand (n8574, n8573, n8565);
   nand (n8575, n8572, n8574);
   xor (n8576, n8392, n8394);
   xor (n8577, n8575, n8576);
   and (n8578, n8466, n8497);
   not (n8579, n8466);
   not (n858, n857);
   and (n8580, n8579, n8496);
   nor (n8581, n8578, n8580);
   or (n8582, n8577, n8581);
   not (n8583, n8575);
   or (n8584, n8583, n8576);
   nand (n8585, n8582, n8584);
   not (n8586, n8585);
   or (n8587, n8520, n8586);
   or (n8588, n8519, n8585);
   nand (n8589, n8587, n8588);
   or (n859, n856, n858);
   not (n8590, n8589);
   and (n8591, n8453, n8450);
   xor (n8592, n8591, n7220);
   and (n8593, n99, n78);
   and (n8594, n8593, n14);
   not (n8595, n8594);
   not (n8596, n13);
   not (n8597, n8596);
   not (n8598, n8488);
   or (n8599, n8597, n8598);
   buf (n86, g85);
   nand (n860, n274, n468);
   nand (n8600, n8599, n8490);
   not (n8601, n8600);
   not (n8602, n8601);
   or (n8603, n8595, n8602);
   nand (n8604, n80, n97);
   nand (n8605, n81, n96);
   nor (n8606, n8604, n8605);
   not (n8607, n8606);
   not (n8608, n8428);
   and (n8609, n8605, n8604);
   nand (n861, n859, n860);
   nor (n8610, n8609, n8606);
   nand (n8611, n8608, n8610);
   nand (n8612, n8607, n8611);
   not (n8613, n8594);
   not (n8614, n8600);
   or (n8615, n8613, n8614);
   or (n8616, n8600, n8594);
   nand (n8617, n8615, n8616);
   nand (n8618, n8612, n8617);
   nand (n8619, n8603, n8618);
   not (n862, n861);
   xor (n8620, n8592, n8619);
   xor (n8621, n8486, n7660);
   xor (n8622, n8621, n8490);
   not (n8623, n8622);
   and (n8624, n8620, n8623);
   and (n8625, n8592, n8619);
   nor (n8626, n8624, n8625);
   not (n8627, n8626);
   xor (n8628, n8483, n8493);
   not (n8629, n8628);
   not (n863, n751);
   or (n8630, n8627, n8629);
   not (n8631, n8626);
   not (n8632, n8631);
   or (n8633, n8632, n8628);
   nand (n8634, n8630, n8633);
   not (n8635, n8634);
   xor (n8636, n8570, n8552);
   or (n8637, n8635, n8636);
   not (n8638, n8628);
   or (n8639, n8632, n8638);
   and (n864, n862, n863);
   nand (n8640, n8637, n8639);
   buf (n8641, n8640);
   not (n8642, n8641);
   xor (n8643, n8577, n8581);
   not (n8644, n8643);
   or (n8645, n8642, n8644);
   or (n8646, n8643, n8641);
   nand (n8647, n8645, n8646);
   not (n8648, n8647);
   not (n8649, n8636);
   and (n865, n861, n751);
   not (n8650, n8634);
   or (n8651, n8649, n8650);
   or (n8652, n8634, n8636);
   nand (n8653, n8651, n8652);
   not (n8654, n8653);
   xnor (n8655, n8549, n8547);
   and (n8656, n83, n95);
   and (n8657, n8656, n8530);
   and (n8658, n82, n95);
   not (n8659, n7997);
   nor (n866, n864, n865);
   nor (n8660, n8658, n8659);
   nor (n8661, n8657, n8660);
   nand (n8662, n79, n99);
   not (n8663, n8662);
   nand (n8664, n8663, n15);
   not (n8665, n8664);
   and (n8666, n8661, n8665);
   nor (n8667, n8666, n8657);
   not (n8668, n8667);
   not (n8669, n8536);
   not (n867, n736);
   not (n8670, n8541);
   not (n8671, n8670);
   or (n8672, n8669, n8671);
   nand (n8673, n8672, n8542);
   and (n8674, n8529, n7640);
   not (n8675, n8529);
   and (n8676, n8675, n8530);
   or (n8677, n8674, n8676);
   xnor (n8678, n8673, n8677);
   not (n8679, n8678);
   and (n868, n867, n843);
   or (n8680, n8668, n8679);
   not (n8681, n8677);
   nand (n8682, n8681, n8673);
   nand (n8683, n8680, n8682);
   and (n8684, n8655, n8683);
   not (n8685, n8655);
   not (n8686, n8683);
   and (n8687, n8685, n8686);
   or (n8688, n8684, n8687);
   not (n8689, n8622);
   and (n869, n430, n510);
   not (n8690, n8620);
   or (n8691, n8689, n8690);
   or (n8692, n8620, n8622);
   nand (n8693, n8691, n8692);
   and (n8694, n8688, n8693);
   and (n8695, n8686, n8655);
   nor (n8696, n8694, n8695);
   not (n8697, n8696);
   or (n8698, n8654, n8697);
   or (n8699, n8653, n8696);
   buf (n87, g86);
   nor (n870, n868, n869);
   nand (n8700, n8698, n8699);
   not (n8701, n8700);
   not (n8702, n8693);
   and (n8703, n8688, n8702);
   not (n8704, n8688);
   and (n8705, n8704, n8693);
   nor (n8706, n8703, n8705);
   not (n8707, n8706);
   xnor (n8708, n8678, n8667);
   not (n8709, n8708);
   not (n871, n870);
   not (n8710, n8593);
   not (n8711, n14);
   and (n8712, n8710, n8711);
   nor (n8713, n8712, n8594);
   nand (n8714, n82, n97);
   not (n8715, n8714);
   nand (n8716, n81, n96);
   not (n8717, n8716);
   nand (n8718, n8715, n8717);
   not (n8719, n82);
   and (n872, n866, n871);
   not (n8720, n96);
   or (n8721, n8719, n8720);
   nand (n8722, n81, n97);
   nand (n8723, n8721, n8722);
   nand (n8724, n8718, n8723);
   nand (n8725, n80, n98);
   or (n8726, n8724, n8725);
   buf (n8727, n8718);
   nand (n8728, n8726, n8727);
   nor (n8729, n8713, n8728);
   not (n873, n866);
   not (n8730, n8729);
   nand (n8731, n8728, n8713);
   nand (n8732, n8730, n8731);
   not (n8733, n8732);
   not (n8734, n8428);
   not (n8735, n8610);
   or (n8736, n8734, n8735);
   or (n8737, n8610, n8428);
   nand (n8738, n8736, n8737);
   and (n8739, n8733, n8738);
   and (n874, n873, n870);
   not (n8740, n8731);
   nor (n8741, n8739, n8740);
   not (n8742, n8741);
   xor (n8743, n8612, n8617);
   not (n8744, n8743);
   and (n8745, n8742, n8744);
   and (n8746, n8741, n8743);
   nor (n8747, n8745, n8746);
   not (n8748, n8747);
   not (n8749, n8748);
   nor (n875, n872, n874);
   or (n8750, n8709, n8749);
   and (n8751, n8733, n8738);
   nor (n8752, n8751, n8740);
   not (n8753, n8743);
   or (n8754, n8752, n8753);
   nand (n8755, n8750, n8754);
   not (n8756, n8755);
   or (n8757, n8707, n8756);
   or (n8758, n8706, n8755);
   nand (n8759, n8757, n8758);
   xor (n876, n855, n875);
   not (n8760, n8759);
   not (n8761, n8747);
   not (n8762, n8708);
   and (n8763, n8761, n8762);
   and (n8764, n8747, n8708);
   nor (n8765, n8763, n8764);
   xnor (n8766, n8738, n8732);
   not (n8767, n8766);
   nand (n8768, n82, n97);
   nand (n8769, n83, n96);
   not (n877, n760);
   nor (n8770, n8768, n8769);
   not (n8771, n8770);
   nand (n8772, n8714, n8769);
   nand (n8773, n8771, n8772);
   nand (n8774, n81, n98);
   nor (n8775, n8773, n8774);
   buf (n8776, n8770);
   or (n8777, n8775, n8776);
   not (n8778, n8656);
   xor (n8779, n8662, n15);
   not (n878, n744);
   not (n8780, n8779);
   or (n8781, n8778, n8780);
   or (n8782, n8779, n8656);
   nand (n8783, n8781, n8782);
   nand (n8784, n8777, n8783);
   not (n8785, n8779);
   nand (n8786, n8785, n8656);
   and (n8787, n8784, n8786);
   and (n8788, n8661, n8664);
   not (n8789, n8661);
   and (n879, n877, n878);
   and (n8790, n8789, n8665);
   nor (n8791, n8788, n8790);
   and (n8792, n8787, n8791);
   not (n8793, n8787);
   not (n8794, n8791);
   and (n8795, n8793, n8794);
   nor (n8796, n8792, n8795);
   not (n8797, n8796);
   or (n8798, n8767, n8797);
   or (n8799, n8787, n8791);
   buf (n88, g87);
   and (n880, n755, n758);
   nand (n8800, n8798, n8799);
   not (n8801, n8800);
   and (n8802, n8765, n8801);
   not (n8803, n8765);
   and (n8804, n8803, n8800);
   nor (n8805, n8802, n8804);
   not (n8806, n8805);
   xor (n8807, n8796, n8766);
   not (n8808, n8783);
   nor (n8809, n8775, n8776);
   nor (n881, n879, n880);
   nand (n8810, n8808, n8809);
   and (n8811, n8784, n8810);
   not (n8812, n8726);
   and (n8813, n8724, n8725);
   nor (n8814, n8812, n8813);
   nand (n8815, n80, n99);
   nand (n8816, n8815, n3759);
   not (n8817, n8816);
   and (n8818, n8814, n8817);
   not (n8819, n8814);
   xor (n882, n813, n816);
   and (n8820, n8819, n8816);
   nor (n8821, n8818, n8820);
   or (n8822, n8811, n8821);
   or (n8823, n8814, n8816);
   nand (n8824, n8822, n8823);
   not (n8825, n8824);
   and (n8826, n8807, n8825);
   not (n8827, n8807);
   and (n8828, n8827, n8824);
   nor (n8829, n8826, n8828);
   not (n883, n823);
   not (n8830, n8829);
   not (n8831, n8821);
   and (n8832, n8811, n8831);
   not (n8833, n8811);
   and (n8834, n8833, n8821);
   nor (n8835, n8832, n8834);
   not (n8836, n8835);
   not (n8837, n16);
   not (n8838, n8815);
   not (n8839, n8838);
   xor (n884, n882, n883);
   or (n8840, n8837, n8839);
   nand (n8841, n8840, n8816);
   not (n8842, n8841);
   not (n8843, n8842);
   nand (n8844, n81, n99);
   not (n8845, n17);
   or (n8846, n8844, n8845);
   not (n8847, n8846);
   and (n8848, n8843, n8847);
   nand (n8849, n8773, n8774);
   not (n885, n884);
   not (n8850, n8849);
   nor (n8851, n8850, n8775);
   and (n8852, n8846, n8841);
   not (n8853, n8846);
   and (n8854, n8853, n8842);
   or (n8855, n8852, n8854);
   and (n8856, n8851, n8855);
   nor (n8857, n8848, n8856);
   not (n8858, n8857);
   and (n8859, n8836, n8858);
   xor (n886, n881, n885);
   and (n8860, n8835, n8857);
   nor (n8861, n8859, n8860);
   nand (n8862, n8844, n8845);
   and (n8863, n8846, n8862);
   nand (n8864, n83, n98);
   nor (n8865, n8864, n8768);
   and (n8866, n82, n98);
   and (n8867, n83, n97);
   nor (n8868, n8866, n8867);
   nor (n8869, n8865, n8868);
   xnor (n887, n839, n845);
   xnor (n8870, n8863, n8869);
   nand (n8871, n83, n19, n99);
   not (n8872, n8871);
   nand (n8873, n8872, n82);
   not (n8874, n99);
   not (n8875, n82);
   or (n8876, n8874, n8875);
   nand (n8877, n8876, n8871);
   and (n8878, n8873, n8877);
   and (n8879, n8864, n3489);
   and (n888, n886, n887);
   nor (n8880, n8864, n3489);
   nor (n8881, n8879, n8880);
   and (n8882, n8878, n8881);
   not (n8883, n8880);
   xor (n8884, n8873, n8883);
   nor (n8885, n8882, n8884);
   or (n8886, n8870, n8885);
   or (n8887, n8873, n8883);
   nand (n8888, n8886, n8887);
   not (n8889, n8888);
   and (n889, n881, n885);
   and (n8890, n8863, n8869);
   nor (n8891, n8890, n8865);
   buf (n8892, n8891);
   not (n8893, n8892);
   xor (n8894, n8851, n8855);
   not (n8895, n8894);
   or (n8896, n8893, n8895);
   or (n8897, n8892, n8894);
   nand (n8898, n8896, n8897);
   not (n8899, n8898);
   buf (n89, g88);
   nor (n890, n888, n889);
   or (n8900, n8889, n8899);
   not (n8901, n8892);
   nand (n8902, n8901, n8894);
   nand (n8903, n8900, n8902);
   or (n8904, n8861, n8903);
   not (n8905, n8835);
   nand (n8906, n8905, n8857);
   and (n8907, n8904, n8906);
   not (n8908, n8907);
   or (n8909, n8830, n8908);
   xor (n891, n876, n890);
   nand (n8910, n8807, n8825);
   nand (n8911, n8909, n8910);
   not (n8912, n8911);
   or (n8913, n8806, n8912);
   not (n8914, n8765);
   nand (n8915, n8914, n8800);
   nand (n8916, n8913, n8915);
   not (n8917, n8916);
   or (n8918, n8760, n8917);
   not (n8919, n8706);
   xor (n892, n850, n891);
   nand (n8920, n8919, n8755);
   nand (n8921, n8918, n8920);
   not (n8922, n8921);
   or (n8923, n8701, n8922);
   not (n8924, n8696);
   nand (n8925, n8924, n8653);
   nand (n8926, n8923, n8925);
   not (n8927, n8926);
   or (n8928, n8648, n8927);
   not (n8929, n8643);
   not (n893, n892);
   nand (n8930, n8929, n8641);
   nand (n8931, n8928, n8930);
   not (n8932, n8931);
   or (n8933, n8590, n8932);
   not (n8934, n8585);
   nand (n8935, n8934, n8519);
   nand (n8936, n8933, n8935);
   not (n8937, n8936);
   or (n8938, n8518, n8937);
   not (n8939, n8511);
   xor (n894, n636, n681);
   nand (n8940, n8939, n8513);
   nand (n8941, n8938, n8940);
   not (n8942, n8941);
   or (n8943, n8425, n8942);
   not (n8944, n8420);
   nand (n8945, n8944, n8418);
   nand (n8946, n8943, n8945);
   not (n8947, n8946);
   or (n8948, n8337, n8947);
   not (n8949, n8332);
   xor (n895, n894, n763);
   nand (n8950, n8949, n8257);
   nand (n8951, n8948, n8950);
   not (n8952, n8951);
   or (n8953, n8256, n8952);
   not (n8954, n8251);
   nand (n8955, n8954, n8249);
   nand (n8956, n8953, n8955);
   not (n8957, n8956);
   or (n8958, n8111, n8957);
   not (n8959, n8103);
   xor (n896, n881, n885);
   nand (n8960, n8959, n8106);
   nand (n8961, n8958, n8960);
   not (n8962, n8961);
   or (n8963, n8034, n8962);
   not (n8964, n8032);
   xor (n8965, n7820, n7870);
   xor (n8966, n8965, n7873);
   nand (n8967, n8964, n8966);
   nand (n8968, n8963, n8967);
   not (n8969, n8968);
   xor (n897, n896, n887);
   or (n8970, n7881, n8969);
   not (n8971, n7876);
   nand (n8972, n8971, n7818);
   nand (n8973, n8970, n8972);
   not (n8974, n8973);
   or (n8975, n7817, n8974);
   not (n8976, n7588);
   nand (n8977, n8976, n7812);
   nand (n8978, n8975, n8977);
   not (n8979, n8978);
   and (n898, n895, n897);
   or (n8980, n7587, n8979);
   not (n8981, n7524);
   nand (n8982, n8981, n7582);
   nand (n8983, n8980, n8982);
   not (n8984, n8983);
   or (n8985, n7522, n8984);
   not (n8986, n7401);
   nand (n8987, n8986, n7517);
   nand (n8988, n8985, n8987);
   not (n8989, n8988);
   not (n899, n895);
   or (n8990, n7400, n8989);
   not (n8991, n7395);
   nand (n8992, n8991, n7198);
   nand (n8993, n8990, n8992);
   not (n8994, n8993);
   or (n8995, n7197, n8994);
   not (n8996, n7192);
   nand (n8997, n8996, n7189);
   nand (n8998, n8995, n8997);
   not (n8999, n8998);
   buf (n9, g8);
   buf (n90, g89);
   not (n900, n897);
   or (n9000, n7069, n8999);
   not (n9001, n7007);
   nand (n9002, n9001, n7064);
   nand (n9003, n9000, n9002);
   not (n9004, n9003);
   or (n9005, n7006, n9004);
   not (n9006, n7001);
   nand (n9007, n9006, n6915);
   nand (n9008, n9005, n9007);
   not (n9009, n9008);
   and (n901, n899, n900);
   or (n9010, n6913, n9009);
   not (n9011, n6853);
   nand (n9012, n9011, n6878);
   or (n9013, n6911, n9012);
   not (n9014, n6906);
   nand (n9015, n9014, n6902);
   or (n9016, n9015, n6900);
   or (n9017, n6883, n6899);
   nand (n9018, n9013, n9016, n9017);
   not (n9019, n9018);
   nor (n902, n898, n901);
   nand (n9020, n9010, n9019);
   not (n9021, n9020);
   or (n9022, n6664, n9021);
   nand (n9023, n6641, n6662);
   nand (n9024, n9022, n9023);
   not (n9025, n6605);
   and (n9026, n6651, n9025);
   nor (n9027, n9026, n6647);
   and (n9028, n68, n85);
   and (n9029, n69, n84);
   xor (n903, n545, n592);
   nor (n9030, n9028, n9029);
   not (n9031, n9030);
   not (n9032, n6583);
   nand (n9033, n9032, n6672);
   nand (n9034, n9031, n9033);
   and (n9035, n9027, n9034);
   nor (n9036, n9027, n9034);
   nor (n9037, n9035, n9036);
   or (n9038, n6645, n6661);
   nand (n9039, n9038, n6660);
   xor (n904, n903, n633);
   xor (n9040, n9037, n9039);
   and (n9041, n9024, n9040);
   and (n9042, n9037, n9039);
   nor (n9043, n9041, n9042);
   not (n9044, n9043);
   not (n9045, n9036);
   nand (n9046, n68, n84);
   or (n9047, n9045, n9046);
   nand (n9048, n9047, n9033);
   or (n9049, n9044, n9048);
   nand (n905, n36, n65);
   and (n9050, n9045, n9046);
   nor (n9051, n9050, n1);
   nand (n9052, n9049, n9051);
   not (n9053, n9052);
   or (n9054, n6576, n9053);
   nand (n9055, n6569, n4814);
   nand (n9056, n1, n3);
   and (n9057, n9055, n9056, n2);
   or (n9058, n1, n3);
   or (n9059, n6569, n4814);
   not (n906, n429);
   nand (n9060, n9058, n9059);
   and (n9061, n237, n9060);
   nor (n9062, n9057, n9061);
   nand (n9063, n9054, n9062);
   not (n9064, n9063);
   nand (n9065, n5962, n5967);
   not (n9066, n9065);
   xor (n9067, n5928, n5962);
   not (n9068, n9067);
   or (n9069, n9066, n9068);
   not (n907, n598);
   nand (n9070, n6471, n6467);
   and (n9071, n6451, n9070);
   and (n9072, n6008, n6424);
   nor (n9073, n9071, n9072);
   not (n9074, n9073);
   nand (n9075, n6418, n6082);
   not (n9076, n9075);
   or (n9077, n9074, n9076);
   nand (n9078, n6452, n6473);
   nand (n9079, n9077, n9078);
   and (n908, n906, n907);
   not (n9080, n6452);
   not (n9081, n6508);
   and (n9082, n9080, n9081);
   and (n9083, n6508, n6452);
   nor (n9084, n9082, n9083);
   nor (n9085, n9079, n9084);
   not (n9086, n6508);
   not (n9087, n6485);
   or (n9088, n9086, n9087);
   nand (n9089, n6507, n6452);
   xor (n909, n42, n58);
   nand (n9090, n9088, n9089);
   nor (n9091, n9085, n9090);
   not (n9092, n6507);
   xnor (n9093, n6507, n6484);
   not (n9094, n9093);
   or (n9095, n9092, n9094);
   not (n9096, n5961);
   and (n9097, n237, n6477);
   not (n9098, n237);
   and (n9099, n9098, n6482);
   buf (n91, g90);
   and (n910, n421, n909);
   or (n9100, n9097, n9099);
   not (n9101, n9100);
   or (n9102, n9096, n9101);
   or (n9103, n9100, n5961);
   nand (n9104, n9102, n9103);
   nand (n9105, n9095, n9104);
   or (n9106, n9091, n9105);
   not (n9107, n5928);
   not (n9108, n5961);
   and (n9109, n9107, n9108);
   nor (n911, n908, n910);
   and (n9110, n5961, n6486);
   nor (n9111, n9109, n9110);
   nand (n9112, n9106, n9111);
   nand (n9113, n9069, n9112);
   xnor (n9114, n5927, n5908);
   buf (n9115, n9114);
   xnor (n9116, n9113, n9115);
   and (n9117, n9116, n1);
   buf (n9118, n8993);
   not (n9119, n9118);
   xor (n912, n905, n911);
   not (n9120, n7196);
   not (n9121, n9120);
   and (n9122, n9119, n9121);
   and (n9123, n9118, n9120);
   nor (n9124, n9122, n9123);
   nor (n9125, n9124, n1);
   nor (n9126, n9117, n9125);
   not (n9127, n9126);
   not (n9128, n1);
   and (n9129, n6329, n6321);
   buf (n913, n535);
   not (n9130, n6329);
   and (n9131, n9130, n6320);
   nor (n9132, n9129, n9131);
   not (n9133, n9132);
   or (n9134, n9128, n9133);
   xor (n9135, n8700, n8921);
   nand (n9136, n9135, n6569);
   nand (n9137, n9134, n9136);
   and (n9138, n9137, n16);
   not (n9139, n9137);
   and (n914, n46, n54);
   and (n9140, n9139, n3759);
   nor (n9141, n9138, n9140);
   not (n9142, n9141);
   not (n9143, n17);
   not (n9144, n18);
   not (n9145, n6569);
   xor (n9146, n8907, n8829);
   not (n9147, n9146);
   or (n9148, n9145, n9147);
   and (n9149, n6217, n6283);
   not (n915, n46);
   not (n9150, n6217);
   not (n9151, n6283);
   and (n9152, n9150, n9151);
   nor (n9153, n9149, n9152);
   nand (n9154, n9153, n1);
   nand (n9155, n9148, n9154);
   nand (n9156, n9155, n19);
   not (n9157, n9156);
   not (n9158, n9157);
   or (n9159, n9144, n9158);
   and (n916, n915, n299);
   not (n9160, n3489);
   not (n9161, n9156);
   or (n9162, n9160, n9161);
   buf (n9163, n6288);
   buf (n9164, n6176);
   and (n9165, n9163, n9164);
   not (n9166, n9163);
   not (n9167, n9164);
   and (n9168, n9166, n9167);
   nor (n9169, n9165, n9168);
   nor (n917, n914, n916);
   and (n9170, n1, n9169);
   not (n9171, n1);
   xor (n9172, n8911, n8805);
   and (n9173, n9171, n9172);
   or (n9174, n9170, n9173);
   nand (n9175, n9162, n9174);
   nand (n9176, n9159, n9175);
   not (n9177, n9176);
   or (n9178, n9143, n9177);
   xor (n9179, n6311, n6295);
   and (n918, n913, n917);
   and (n9180, n9179, n1);
   buf (n9181, n8759);
   xnor (n9182, n8916, n9181);
   nor (n9183, n9182, n1);
   nor (n9184, n9180, n9183);
   nand (n9185, n9178, n9184);
   or (n9186, n9176, n17);
   and (n9187, n9185, n9186);
   not (n9188, n9187);
   or (n9189, n9142, n9188);
   and (n919, n543, n625);
   nand (n9190, n16, n9137);
   nand (n9191, n9189, n9190);
   not (n9192, n9191);
   not (n9193, n6569);
   xor (n9194, n8926, n8647);
   not (n9195, n9194);
   or (n9196, n9193, n9195);
   xor (n9197, n6148, n6133);
   not (n9198, n6334);
   and (n9199, n9197, n9198);
   buf (n92, g91);
   nor (n920, n918, n919);
   not (n9200, n9197);
   and (n9201, n9200, n6334);
   nor (n9202, n9199, n9201);
   nand (n9203, n9202, n1);
   nand (n9204, n9196, n9203);
   and (n9205, n9204, n15);
   not (n9206, n9204);
   not (n9207, n15);
   and (n9208, n9206, n9207);
   nor (n9209, n9205, n9208);
   and (n921, n912, n920);
   not (n9210, n9209);
   or (n9211, n9192, n9210);
   nand (n9212, n15, n9204);
   nand (n9213, n9211, n9212);
   buf (n9214, n6374);
   nand (n9215, n6370, n9214);
   buf (n9216, n6397);
   not (n9217, n9216);
   and (n9218, n9215, n9217);
   not (n9219, n9215);
   and (n922, n905, n911);
   and (n9220, n9219, n9216);
   nor (n9221, n9218, n9220);
   nand (n9222, n1, n9221);
   xor (n9223, n8936, n8517);
   nand (n9224, n9223, n6569);
   nand (n9225, n9222, n9224);
   not (n9226, n6569);
   xor (n9227, n8589, n8931);
   not (n9228, n9227);
   or (n9229, n9226, n9228);
   nor (n923, n921, n922);
   not (n9230, n9197);
   not (n9231, n9198);
   or (n9232, n9230, n9231);
   nand (n9233, n9232, n6149);
   not (n9234, n6367);
   and (n9235, n9233, n9234);
   not (n9236, n9233);
   and (n9237, n9236, n6367);
   nor (n9238, n9235, n9237);
   nand (n9239, n1, n9238);
   not (n924, n923);
   nand (n9240, n9229, n9239);
   and (n9241, n9213, n9225, n9240);
   not (n9242, n9217);
   not (n9243, n9215);
   or (n9244, n9242, n9243);
   buf (n9245, n6396);
   nand (n9246, n9244, n9245);
   not (n9247, n6406);
   and (n9248, n9246, n9247);
   not (n9249, n9246);
   and (n925, n44, n56);
   and (n9250, n9249, n6406);
   nor (n9251, n9248, n9250);
   and (n9252, n9251, n1);
   xnor (n9253, n8941, n8424);
   nor (n9254, n9253, n1);
   nor (n9255, n9252, n9254);
   not (n9256, n6411);
   xnor (n9257, n6070, n6415);
   and (n9258, n9256, n9257);
   not (n9259, n9256);
   not (n926, n44);
   not (n9260, n9257);
   and (n9261, n9259, n9260);
   nor (n9262, n9258, n9261);
   and (n9263, n9262, n1);
   not (n9264, n8336);
   not (n9265, n8946);
   not (n9266, n9265);
   or (n9267, n9264, n9266);
   or (n9268, n9265, n8336);
   nand (n9269, n9267, n9268);
   and (n927, n926, n479);
   and (n9270, n9269, n6569);
   nor (n9271, n9263, n9270);
   nor (n9272, n9255, n9271);
   nand (n9273, n9241, n9272);
   not (n9274, n6569);
   xor (n9275, n8951, n8255);
   not (n9276, n9275);
   or (n9277, n9274, n9276);
   not (n9278, n9257);
   not (n9279, n9256);
   nor (n928, n925, n927);
   or (n9280, n9278, n9279);
   not (n9281, n6416);
   nand (n9282, n9280, n9281);
   and (n9283, n6080, n6074);
   not (n9284, n6080);
   and (n9285, n9284, n6412);
   nor (n9286, n9283, n9285);
   not (n9287, n9286);
   and (n9288, n9282, n9287);
   not (n9289, n9282);
   and (n929, n566, n928);
   and (n9290, n9289, n9286);
   nor (n9291, n9288, n9290);
   nand (n9292, n9291, n1);
   nand (n9293, n9277, n9292);
   not (n9294, n1);
   not (n9295, n6081);
   nand (n9296, n9295, n6418);
   xor (n9297, n9296, n6029);
   not (n9298, n9297);
   or (n9299, n9294, n9298);
   buf (n93, g92);
   and (n930, n556, n570);
   not (n9300, n8110);
   not (n9301, n8956);
   not (n9302, n9301);
   or (n9303, n9300, n9302);
   or (n9304, n9301, n8110);
   nand (n9305, n9303, n9304);
   nand (n9306, n9305, n6569);
   nand (n9307, n9299, n9306);
   nand (n9308, n9293, n9307);
   nor (n9309, n9273, n9308);
   nor (n931, n929, n930);
   nand (n9310, n6473, n9070);
   and (n9311, n6426, n9310);
   not (n9312, n6426);
   not (n9313, n9310);
   and (n9314, n9312, n9313);
   nor (n9315, n9311, n9314);
   not (n9316, n9315);
   not (n9317, n1);
   or (n9318, n9316, n9317);
   xor (n9319, n8961, n8033);
   not (n932, n931);
   nand (n9320, n9319, n6569);
   nand (n9321, n9318, n9320);
   nand (n9322, n9309, n9321);
   not (n9323, n1);
   and (n9324, n6469, n6472);
   or (n9325, n6426, n9324);
   or (n9326, n6469, n6472);
   nand (n9327, n9325, n9326);
   or (n9328, n6489, n6469);
   nand (n9329, n9328, n6470);
   not (n933, n932);
   xnor (n9330, n9327, n9329);
   not (n9331, n9330);
   or (n9332, n9323, n9331);
   xor (n9333, n8968, n7880);
   nand (n9334, n9333, n6569);
   nand (n9335, n9332, n9334);
   not (n9336, n1);
   xor (n9337, n9079, n9084);
   not (n9338, n9337);
   or (n9339, n9336, n9338);
   and (n934, n40, n60);
   not (n9340, n7816);
   not (n9341, n8973);
   not (n9342, n9341);
   or (n9343, n9340, n9342);
   or (n9344, n9341, n7816);
   nand (n9345, n9343, n9344);
   nand (n9346, n9345, n6569);
   nand (n9347, n9339, n9346);
   nand (n9348, n9335, n9347);
   nor (n9349, n9322, n9348);
   not (n935, n40);
   not (n9350, n1);
   nor (n9351, n6485, n6508);
   nor (n9352, n9351, n9091);
   xor (n9353, n9104, n9352);
   not (n9354, n9353);
   or (n9355, n9350, n9354);
   xor (n9356, n8983, n7521);
   nand (n9357, n9356, n6569);
   nand (n9358, n9355, n9357);
   buf (n9359, n8978);
   and (n936, n935, n647);
   xnor (n9360, n7586, n9359);
   and (n9361, n6569, n9360);
   not (n9362, n6569);
   buf (n9363, n9085);
   not (n9364, n9089);
   nor (n9365, n9363, n9364);
   not (n9366, n9365);
   buf (n9367, n9093);
   not (n9368, n9367);
   not (n9369, n9368);
   nor (n937, n934, n936);
   and (n9370, n9366, n9369);
   and (n9371, n9365, n9368);
   nor (n9372, n9370, n9371);
   and (n9373, n9362, n9372);
   nor (n9374, n9361, n9373);
   and (n9375, n9349, n9358, n9374);
   not (n9376, n1);
   not (n9377, n9352);
   not (n9378, n9104);
   or (n9379, n9377, n9378);
   not (n938, n937);
   nand (n9380, n6512, n6486);
   nand (n9381, n9379, n9380);
   xnor (n9382, n9381, n9067);
   not (n9383, n9382);
   or (n9384, n9376, n9383);
   xor (n9385, n8988, n7399);
   nand (n9386, n9385, n6569);
   nand (n9387, n9384, n9386);
   nand (n9388, n9127, n9375, n9387);
   not (n9389, n9388);
   not (n939, n265);
   not (n9390, n9115);
   not (n9391, n9113);
   not (n9392, n9391);
   or (n9393, n9390, n9392);
   nand (n9394, n5908, n5928);
   buf (n9395, n9394);
   nand (n9396, n9393, n9395);
   not (n9397, n5880);
   not (n9398, n9397);
   not (n9399, n5966);
   buf (n94, g93);
   or (n940, n938, n939);
   and (n9400, n9398, n9399);
   and (n9401, n5879, n5966);
   nor (n9402, n9400, n9401);
   not (n9403, n9402);
   and (n9404, n9396, n9403);
   not (n9405, n9396);
   and (n9406, n9405, n9402);
   nor (n9407, n9404, n9406);
   and (n9408, n1, n9407);
   not (n9409, n1);
   nand (n941, n274, n580);
   not (n9410, n8998);
   not (n9411, n7068);
   and (n9412, n9410, n9411);
   not (n9413, n9410);
   and (n9414, n9413, n7068);
   nor (n9415, n9412, n9414);
   and (n9416, n9409, n9415);
   nor (n9417, n9408, n9416);
   xor (n9418, n9003, n7005);
   and (n9419, n6569, n9418);
   nand (n942, n940, n941);
   not (n9420, n6569);
   not (n9421, n5909);
   not (n9422, n5872);
   not (n9423, n2);
   or (n9424, n9422, n9423);
   nand (n9425, n9424, n5878);
   not (n9426, n9425);
   or (n9427, n9421, n9426);
   nand (n9428, n9427, n9394);
   not (n9429, n9428);
   not (n943, n38);
   not (n9430, n9429);
   not (n9431, n9113);
   or (n9432, n9430, n9431);
   not (n9433, n9428);
   not (n9434, n9114);
   and (n9435, n9433, n9434);
   and (n9436, n5880, n5966);
   nor (n9437, n9435, n9436);
   nand (n9438, n9432, n9437);
   not (n9439, n5855);
   not (n944, n62);
   not (n9440, n5879);
   or (n9441, n9439, n9440);
   nand (n9442, n9441, n5881);
   not (n9443, n9442);
   and (n9444, n9438, n9443);
   not (n9445, n9438);
   and (n9446, n9445, n9442);
   nor (n9447, n9444, n9446);
   and (n9448, n9420, n9447);
   nor (n9449, n9419, n9448);
   and (n945, n943, n944);
   nor (n9450, n9417, n9449);
   nand (n9451, n9389, n9450);
   not (n9452, n9008);
   and (n9453, n9452, n6882);
   not (n9454, n9452);
   not (n9455, n6882);
   and (n9456, n9454, n9455);
   nor (n9457, n9453, n9456);
   and (n9458, n6569, n9457);
   not (n9459, n6569);
   and (n946, n38, n62);
   not (n9460, n9391);
   and (n9461, n5855, n5880);
   nor (n9462, n9461, n9428);
   and (n9463, n9460, n9462);
   or (n9464, n9437, n5857);
   not (n9465, n5855);
   nand (n9466, n9465, n9397);
   nand (n9467, n9464, n9466);
   nor (n9468, n9463, n9467);
   buf (n9469, n9468);
   nor (n947, n945, n946);
   and (n9470, n5866, n5856);
   not (n9471, n5866);
   and (n9472, n9471, n5857);
   nor (n9473, n9470, n9472);
   buf (n9474, n9473);
   xor (n9475, n9469, n9474);
   and (n9476, n9459, n9475);
   nor (n9477, n9458, n9476);
   nor (n9478, n9451, n9477);
   not (n9479, n9473);
   not (n948, n947);
   not (n9480, n9468);
   or (n9481, n9479, n9480);
   not (n9482, n5857);
   nand (n9483, n9482, n5887);
   nand (n9484, n9481, n9483);
   not (n9485, n5866);
   not (n9486, n5771);
   or (n9487, n9485, n9486);
   or (n9488, n5887, n5771);
   nand (n9489, n9487, n9488);
   not (n949, n376);
   xnor (n9490, n9484, n9489);
   or (n9491, n9490, n6569);
   not (n9492, n9455);
   not (n9493, n9008);
   or (n9494, n9492, n9493);
   nand (n9495, n9494, n9012);
   xnor (n9496, n9495, n6910);
   or (n9497, n9496, n1);
   nand (n9498, n9491, n9497);
   nand (n9499, n9478, n9498);
   buf (n95, g94);
   or (n950, n948, n949);
   not (n9500, n9499);
   not (n9501, n6910);
   not (n9502, n9495);
   or (n9503, n9501, n9502);
   nand (n9504, n9503, n9015);
   xnor (n9505, n9504, n6900);
   and (n9506, n6569, n9505);
   not (n9507, n6569);
   not (n9508, n5771);
   xor (n9509, n5842, n9508);
   nand (n951, n310, n694);
   not (n9510, n9489);
   not (n9511, n9484);
   or (n9512, n9510, n9511);
   nand (n9513, n5771, n5888);
   nand (n9514, n9512, n9513);
   and (n9515, n9509, n9514);
   not (n9516, n9509);
   not (n9517, n9514);
   and (n9518, n9516, n9517);
   nor (n9519, n9515, n9518);
   nand (n952, n950, n951);
   and (n9520, n9507, n9519);
   nor (n9521, n9506, n9520);
   not (n9522, n9521);
   nand (n9523, n9500, n9522);
   not (n9524, n9523);
   not (n9525, n6569);
   nor (n9526, n9048, n9050);
   not (n9527, n9526);
   not (n9528, n9043);
   or (n9529, n9527, n9528);
   xor (n953, n942, n952);
   or (n9530, n9043, n9526);
   nand (n9531, n9529, n9530);
   not (n9532, n9531);
   or (n9533, n9525, n9532);
   nand (n9534, n9533, n6575);
   buf (n9535, n9534);
   nand (n9536, n9524, n9535);
   nand (n9537, n9064, n9536);
   nand (n9538, n6663, n9023);
   xor (n9539, n9020, n9538);
   not (n954, n953);
   nor (n9540, n9539, n1);
   not (n9541, n9540);
   not (n9542, n9541);
   nand (n9543, n6568, n9508);
   and (n9544, n9517, n9543);
   nor (n9545, n6568, n9508);
   nor (n9546, n9544, n9545);
   nor (n9547, n6561, n6568);
   not (n9548, n9547);
   nand (n9549, n9548, n6562);
   or (n955, n933, n954);
   or (n9550, n9546, n9549, n6569);
   not (n9551, n9550);
   or (n9552, n9542, n9551);
   nand (n9553, n6567, n1);
   nor (n9554, n6563, n9553);
   not (n9555, n9554);
   xnor (n9556, n9024, n9040);
   nor (n9557, n9556, n1);
   not (n9558, n9557);
   nand (n9559, n9555, n9558, n6575);
   nand (n956, n942, n952);
   nand (n9560, n9552, n9559);
   not (n9561, n9560);
   or (n9562, n9044, n9048);
   nand (n9563, n9562, n9051);
   nand (n9564, n6575, n9563);
   not (n9565, n9062);
   nor (n9566, n9564, n9565);
   nand (n9567, n9524, n9561, n9566, n9535);
   not (n9568, n9063);
   nand (n9569, n9568, n9560);
   nand (n957, n955, n956);
   nor (n9570, n3645, n3380);
   not (n9571, n9570);
   not (n9572, n2845);
   or (n9573, n9571, n9572);
   nand (n9574, n3645, n3380);
   not (n9575, n9574);
   nand (n9576, n9575, n3043);
   nand (n9577, n9573, n9576);
   not (n9578, n9577);
   or (n9579, n9578, n2945);
   not (n958, n957);
   not (n9580, n9570);
   and (n9581, n9580, n9574);
   not (n9582, n9581);
   or (n9583, n9582, n2847);
   nand (n9584, n9579, n9583);
   not (n9585, n2833);
   nor (n9586, n9585, n335);
   xor (n9587, n9584, n9586);
   not (n9588, n2958);
   and (n9589, n3043, n3697);
   not (n959, n958);
   not (n9590, n9589);
   not (n9591, n2831);
   or (n9592, n9590, n9591);
   nand (n9593, n2845, n3176);
   or (n9594, n9593, n2832);
   nand (n9595, n9592, n9594);
   not (n9596, n9595);
   not (n9597, n9596);
   not (n9598, n9597);
   or (n9599, n9588, n9598);
   buf (n96, g95);
   or (n960, n924, n959);
   not (n9600, n9589);
   nand (n9601, n9600, n9593);
   not (n9602, n9601);
   not (n9603, n9602);
   and (n9604, n2834, n305);
   nor (n9605, n2834, n305);
   nor (n9606, n9604, n9605);
   not (n9607, n9606);
   or (n9608, n9603, n9607);
   nand (n9609, n9599, n9608);
   or (n961, n958, n923);
   and (n9610, n9587, n9609);
   and (n9611, n9584, n9586);
   nor (n9612, n9610, n9611);
   nand (n9613, n3034, n2991);
   not (n9614, n9613);
   not (n9615, n2907);
   and (n9616, n9614, n9615);
   nor (n9617, n3521, n2990);
   buf (n9618, n9617);
   and (n9619, n9618, n3475);
   nand (n962, n960, n961);
   nor (n9620, n9616, n9619);
   not (n9621, n9620);
   not (n9622, n2983);
   and (n9623, n9621, n9622);
   nor (n9624, n9618, n2907);
   and (n9625, n9624, n9613);
   nor (n9626, n9623, n9625);
   and (n9627, n9597, n9606);
   not (n9628, n9603);
   and (n9629, n9628, n2837);
   xor (n963, n629, n622);
   nor (n9630, n9627, n9629);
   xnor (n9631, n9626, n9630);
   xnor (n9632, n9612, n9631);
   not (n9633, n2847);
   and (n9634, n9577, n9633);
   and (n9635, n9581, n2953);
   nor (n9636, n9634, n9635);
   xor (n9637, n9636, n9624);
   xor (n9638, n9637, n2956);
   xor (n9639, n9632, n9638);
   nand (n964, n962, n963);
   not (n9640, n2930);
   and (n9641, n9621, n9640);
   not (n9642, n9617);
   nand (n9643, n9642, n9613);
   not (n9644, n9643);
   not (n9645, n9644);
   buf (n9646, n9645);
   not (n9647, n9646);
   and (n9648, n9647, n9622);
   nor (n9649, n9641, n9648);
   nand (n965, n957, n923);
   and (n9650, n3237, n4374);
   not (n9651, n9650);
   and (n9652, n9651, n3072);
   xnor (n9653, n9649, n9652);
   and (n9654, n2834, n335);
   nor (n9655, n9654, n9586);
   and (n9656, n9597, n9655);
   and (n9657, n9628, n2958);
   nor (n9658, n9656, n9657);
   or (n9659, n9653, n9658);
   and (n966, n964, n965);
   or (n9660, n9649, n9652);
   nand (n9661, n9659, n9660);
   xor (n9662, n9661, n9626);
   xor (n9663, n9587, n9609);
   and (n9664, n9662, n9663);
   and (n9665, n9661, n9626);
   nor (n9666, n9664, n9665);
   xor (n9667, n9639, n9666);
   not (n9668, n9667);
   xnor (n9669, n9662, n9663);
   not (n967, n966);
   and (n9670, n39, n2845);
   not (n9671, n39);
   and (n9672, n9671, n2846);
   nor (n9673, n9670, n9672);
   or (n9674, n9578, n9673);
   or (n9675, n9582, n2945);
   nand (n9676, n9674, n9675);
   and (n9677, n42, n3058);
   xor (n9678, n9676, n9677);
   not (n9679, n9621);
   and (n968, n904, n967);
   or (n9680, n9679, n3101);
   or (n9681, n9646, n2930);
   nand (n9682, n9680, n9681);
   and (n9683, n9678, n9682);
   and (n9684, n9676, n9677);
   nor (n9685, n9683, n9684);
   xnor (n9686, n9669, n9685);
   xor (n9687, n9653, n9658);
   and (n9688, n9597, n3059);
   and (n9689, n9628, n9655);
   not (n969, n904);
   nor (n9690, n9688, n9689);
   nand (n9691, n2833, n43);
   xor (n9692, n9690, n9691);
   nand (n9693, n3126, n4373);
   nor (n9694, n9693, n3521);
   not (n9695, n9694);
   nand (n9696, n9650, n3034);
   nand (n9697, n9695, n9696);
   and (n9698, n9697, n3142);
   and (n9699, n9652, n9693);
   buf (n97, g96);
   and (n970, n969, n966);
   nor (n9700, n9698, n9699);
   and (n9701, n9692, n9700);
   and (n9702, n9690, n9691);
   nor (n9703, n9701, n9702);
   xor (n9704, n9687, n9703);
   xor (n9705, n9678, n9682);
   and (n9706, n9704, n9705);
   and (n9707, n9687, n9703);
   nor (n9708, n9706, n9707);
   or (n9709, n9686, n9708);
   nor (n971, n968, n970);
   or (n9710, n9669, n9685);
   nand (n9711, n9709, n9710);
   not (n9712, n9711);
   or (n9713, n9668, n9712);
   or (n9714, n9711, n9667);
   nand (n9715, n9713, n9714);
   not (n9716, n9715);
   xor (n9717, n9686, n9708);
   not (n9718, n9717);
   xor (n9719, n9687, n9703);
   xor (n972, n735, n761);
   xor (n9720, n9719, n9705);
   xnor (n9721, n2928, n39);
   or (n9722, n9679, n9721);
   or (n9723, n9646, n3101);
   nand (n9724, n9722, n9723);
   not (n9725, n3059);
   not (n9726, n9628);
   or (n9727, n9725, n9726);
   or (n9728, n2833, n43);
   nand (n9729, n9728, n9691);
   and (n973, n971, n972);
   or (n9730, n9596, n9729);
   nand (n9731, n9727, n9730);
   xor (n9732, n9724, n9731);
   and (n9733, n44, n3058);
   and (n9734, n9732, n9733);
   and (n9735, n9724, n9731);
   nor (n9736, n9734, n9735);
   and (n9737, n9577, n3048);
   not (n9738, n9673);
   and (n9739, n9581, n9738);
   and (n974, n967, n904);
   nor (n9740, n9737, n9739);
   xnor (n9741, n9740, n9682);
   or (n9742, n9736, n9741);
   or (n9743, n9740, n9682);
   nand (n9744, n9742, n9743);
   xor (n9745, n9720, n9744);
   xnor (n9746, n9736, n9741);
   xor (n9747, n9690, n9691);
   xor (n9748, n9747, n9700);
   not (n9749, n9697);
   nor (n975, n973, n974);
   or (n9750, n9749, n3076);
   nand (n9751, n9693, n9651);
   not (n9752, n9751);
   not (n9753, n9752);
   not (n9754, n3142);
   or (n9755, n9753, n9754);
   nand (n9756, n9750, n9755);
   and (n9757, n3, n13);
   not (n9758, n3);
   and (n9759, n9758, n29);
   and (n976, n902, n975);
   or (n9760, n9757, n9759);
   and (n9761, n4756, n9760);
   not (n9762, n9761);
   and (n9763, n9762, n3238);
   or (n9764, n9756, n9763);
   nand (n9765, n9756, n9763);
   nand (n9766, n9764, n9765);
   and (n9767, n2846, n335);
   and (n9768, n2845, n41);
   nor (n9769, n9767, n9768);
   and (n977, n895, n897);
   or (n9770, n9578, n9769);
   or (n9771, n9582, n3049);
   nand (n9772, n9770, n9771);
   and (n9773, n9766, n9772);
   not (n9774, n9763);
   and (n9775, n9756, n9774);
   nor (n9776, n9773, n9775);
   xor (n9777, n9748, n9776);
   and (n9778, n9746, n9777);
   and (n9779, n9776, n9748);
   nor (n978, n976, n977);
   nor (n9780, n9778, n9779);
   and (n9781, n9745, n9780);
   and (n9782, n9720, n9744);
   nor (n9783, n9781, n9782);
   not (n9784, n9783);
   or (n9785, n9718, n9784);
   or (n9786, n9783, n9717);
   nand (n9787, n9785, n9786);
   not (n9788, n9787);
   xnor (n9789, n9745, n9780);
   not (n979, n978);
   not (n9790, n9789);
   xor (n9791, n9777, n9746);
   not (n9792, n3264);
   or (n9793, n9578, n9792);
   or (n9794, n9582, n9769);
   nand (n9795, n9793, n9794);
   not (n9796, n9795);
   and (n9797, n9597, n3216);
   not (n9798, n9729);
   and (n9799, n9798, n9602);
   buf (n98, g97);
   or (n980, n893, n979);
   nor (n9800, n9797, n9799);
   not (n9801, n9800);
   and (n9802, n9796, n9801);
   and (n9803, n9795, n9800);
   nor (n9804, n9802, n9803);
   not (n9805, n3127);
   not (n9806, n9761);
   or (n9807, n9805, n9806);
   nand (n9808, n3419, n3451);
   or (n9809, n9808, n3127);
   not (n981, n975);
   nand (n9810, n9807, n9809);
   buf (n9811, n9810);
   not (n9812, n5464);
   and (n9813, n9811, n9812);
   and (n9814, n9763, n9808);
   nor (n9815, n9813, n9814);
   or (n9816, n9804, n9815);
   not (n9817, n9795);
   or (n9818, n9817, n9800);
   nand (n9819, n9816, n9818);
   and (n982, n902, n981);
   or (n9820, n9749, n3210);
   or (n9821, n9753, n3076);
   nand (n9822, n9820, n9821);
   xor (n9823, n9819, n9822);
   xor (n9824, n9732, n9733);
   and (n9825, n9823, n9824);
   and (n9826, n9819, n9822);
   nor (n9827, n9825, n9826);
   xor (n9828, n9791, n9827);
   xor (n9829, n9823, n9824);
   not (n983, n902);
   xor (n9830, n9766, n9772);
   or (n9831, n9679, n3295);
   or (n9832, n9646, n9721);
   nand (n9833, n9831, n9832);
   nand (n9834, n3058, n45);
   not (n9835, n9834);
   xor (n9836, n9833, n9835);
   not (n9837, n9822);
   and (n9838, n9836, n9837);
   and (n9839, n9833, n9835);
   and (n984, n983, n975);
   nor (n9840, n9838, n9839);
   not (n9841, n9840);
   and (n9842, n9830, n9841);
   not (n9843, n9830);
   and (n9844, n9843, n9840);
   nor (n9845, n9842, n9844);
   and (n9846, n9829, n9845);
   and (n9847, n9830, n9841);
   nor (n9848, n9846, n9847);
   and (n9849, n9828, n9848);
   nor (n985, n982, n984);
   and (n9850, n9791, n9827);
   nor (n9851, n9849, n9850);
   not (n9852, n9851);
   or (n9853, n9790, n9852);
   or (n9854, n9851, n9789);
   nand (n9855, n9853, n9854);
   not (n9856, n9855);
   xor (n9857, n9791, n9827);
   xor (n9858, n9857, n9848);
   not (n9859, n9858);
   not (n986, n985);
   xnor (n9860, n9829, n9845);
   xnor (n9861, n2846, n43);
   or (n9862, n9578, n9861);
   or (n9863, n9582, n9792);
   nand (n9864, n9862, n9863);
   xnor (n9865, n3072, n39);
   or (n9866, n9749, n9865);
   or (n9867, n9753, n3210);
   nand (n9868, n9866, n9867);
   xor (n9869, n9864, n9868);
   not (n987, n963);
   or (n9870, n2833, n45);
   nand (n9871, n9870, n9834);
   or (n9872, n9596, n9871);
   not (n9873, n3216);
   or (n9874, n9603, n9873);
   nand (n9875, n9872, n9874);
   and (n9876, n9869, n9875);
   and (n9877, n9864, n9868);
   nor (n9878, n9876, n9877);
   not (n9879, n9878);
   not (n988, n962);
   not (n9880, n9811);
   or (n9881, n9880, n3244);
   not (n9882, n9761);
   nand (n9883, n9882, n9808);
   not (n9884, n9883);
   not (n9885, n9884);
   or (n9886, n9885, n5464);
   nand (n9887, n9881, n9886);
   not (n9888, n3836);
   nor (n9889, n3351, n3665);
   not (n989, n988);
   nor (n9890, n9888, n9889);
   not (n9891, n9890);
   xor (n9892, n9887, n9891);
   and (n9893, n2928, n335);
   and (n9894, n2925, n41);
   nor (n9895, n9893, n9894);
   or (n9896, n9679, n9895);
   or (n9897, n9646, n3295);
   nand (n9898, n9896, n9897);
   and (n9899, n9892, n9898);
   buf (n99, g98);
   or (n990, n987, n989);
   and (n9900, n9887, n9891);
   nor (n9901, n9899, n9900);
   not (n9902, n9901);
   and (n9903, n9879, n9902);
   xor (n9904, n9878, n9901);
   xor (n9905, n9804, n9815);
   and (n9906, n9904, n9905);
   nor (n9907, n9903, n9906);
   xor (n9908, n9860, n9907);
   xnor (n9909, n9869, n9875);
   not (n991, n963);
   not (n9910, n9697);
   not (n9911, n5265);
   or (n9912, n9910, n9911);
   or (n9913, n9753, n9865);
   nand (n9914, n9912, n9913);
   or (n9915, n9596, n5318);
   or (n9916, n9603, n9871);
   nand (n9917, n9915, n9916);
   xor (n9918, n9914, n9917);
   and (n9919, n3058, n47);
   nand (n992, n991, n962);
   and (n9920, n9918, n9919);
   and (n9921, n9914, n9917);
   nor (n9922, n9920, n9921);
   xor (n9923, n9909, n9922);
   xnor (n9924, n9892, n9898);
   and (n9925, n9923, n9924);
   and (n9926, n9909, n9922);
   nor (n9927, n9925, n9926);
   not (n9928, n9811);
   not (n9929, n5237);
   nand (n993, n990, n992);
   or (n9930, n9928, n9929);
   or (n9931, n9885, n3244);
   nand (n9932, n9930, n9931);
   or (n9933, n9679, n5307);
   or (n9934, n9645, n9895);
   nand (n9935, n9933, n9934);
   xor (n9936, n9932, n9935);
   or (n9937, n9578, n5275);
   or (n9938, n9582, n9861);
   nand (n9939, n9937, n9938);
   or (n994, n36, n65);
   and (n9940, n9936, n9939);
   and (n9941, n9932, n9935);
   nor (n9942, n9940, n9941);
   nand (n9943, n3431, n4756, n3349);
   not (n9944, n3431);
   nand (n9945, n3765, n4755, n9944);
   and (n9946, n9943, n9945);
   not (n9947, n9946);
   not (n9948, n9947);
   not (n9949, n9948);
   nand (n995, n994, n905);
   and (n9950, n9949, n5248);
   not (n9951, n3431);
   not (n9952, n3764);
   or (n9953, n9951, n9952);
   not (n9954, n3430);
   nand (n9955, n9954, n3349);
   nand (n9956, n9953, n9955);
   not (n9957, n9956);
   not (n9958, n9957);
   not (n9959, n4570);
   or (n996, n247, n995);
   and (n9960, n9958, n9959);
   nor (n9961, n9950, n9960);
   not (n9962, n9961);
   not (n9963, n9962);
   not (n9964, n5317);
   and (n9965, n9963, n9964);
   and (n9966, n9962, n5317);
   nor (n9967, n9965, n9966);
   or (n9968, n9942, n9967);
   or (n9969, n9961, n5317);
   or (n997, n36, n64);
   nand (n9970, n9968, n9969);
   and (n9971, n9836, n9837);
   not (n9972, n9836);
   and (n9973, n9972, n9822);
   nor (n9974, n9971, n9973);
   xnor (n9975, n9970, n9974);
   or (n9976, n9927, n9975);
   or (n9977, n9970, n9974);
   nand (n9978, n9976, n9977);
   and (n9979, n9908, n9978);
   nand (n998, n997, n573);
   and (n9980, n9860, n9907);
   nor (n9981, n9979, n9980);
   not (n9982, n9981);
   or (n9983, n9859, n9982);
   or (n9984, n9981, n9858);
   nand (n9985, n9983, n9984);
   not (n9986, n9985);
   xor (n9987, n9927, n9975);
   xnor (n9988, n9904, n9905);
   xor (n9989, n9987, n9988);
   or (n999, n253, n998);
   xor (n9990, n9942, n9967);
   and (n9991, n5261, n41);
   not (n9992, n5261);
   and (n9993, n9992, n335);
   nor (n9994, n9991, n9993);
   or (n9995, n9749, n9994);
   or (n9996, n9753, n9911);
   nand (n9997, n9995, n9996);
   not (n9998, n3806);
   xor (n9999, n9997, n9998);
endmodule
