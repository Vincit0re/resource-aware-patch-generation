module top ( g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 , g98 , g99 , g100 , g101 , g102 , g103 , g104 , g105 , g106 , g107 , g108 , g109 , g110 , g111 , g112 , g113 , g114 , g115 , g116 , g117 , g118 , g119 , g120 , g121 , g122 , g123 , g124 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g136 , g137 , g138 , g139 , g140 , g141 , g142 , g143 , g144 , g145 , g146 , g147 , g148 , g149 , g150 , g151 , g152 , g153 , g154 , g155 , g156 , g157 , g158 , g159 , g160 , g161 , g162 , g163 , g164 , g165 , g166 , g167 , g168 , g169 , g170 , g171 , g172 , g173 , g174 , g175 , g176 , g177 , g178 , g179 , g180 , g181 , g182 , g183 , g184 , g185 , g186 , g187 , g188 , g189 , g190 , g191 , g192 , g193 , g194 , g195 , g196 , g197 , g198 , g199 , g200 , g201 , g202 , g203 , g204 , g205 , g206 , g207 , g208 , g209 , g210 , g211 , g212 , g213 , g214 , g215 , g216 , g217 , g218 , g219 , g220 , g221 , g222 , g223 , g224 , g225 , g226 );
input g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 , g98 ;
output g99 , g100 , g101 , g102 , g103 , g104 , g105 , g106 , g107 , g108 , g109 , g110 , g111 , g112 , g113 , g114 , g115 , g116 , g117 , g118 , g119 , g120 , g121 , g122 , g123 , g124 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g136 , g137 , g138 , g139 , g140 , g141 , g142 , g143 , g144 , g145 , g146 , g147 , g148 , g149 , g150 , g151 , g152 , g153 , g154 , g155 , g156 , g157 , g158 , g159 , g160 , g161 , g162 , g163 , g164 , g165 , g166 , g167 , g168 , g169 , g170 , g171 , g172 , g173 , g174 , g175 , g176 , g177 , g178 , g179 , g180 , g181 , g182 , g183 , g184 , g185 , g186 , g187 , g188 , g189 , g190 , g191 , g192 , g193 , g194 , g195 , g196 , g197 , g198 , g199 , g200 , g201 , g202 , g203 , g204 , g205 , g206 , g207 , g208 , g209 , g210 , g211 , g212 , g213 , g214 , g215 , g216 , g217 , g218 , g219 , g220 , g221 , g222 , g223 , g224 , g225 , g226 ;

wire n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , 
     n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , 
     n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , 
     n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , 
     n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , 
     n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , 
     n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , 
     n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , 
     n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , 
     n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , 
     n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , 
     n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , 
     n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , 
     n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , 
     n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , 
     n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , 
     n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , 
     n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , 
     n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , 
     n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , 
     n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , 
     n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , 
     n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , 
     n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , 
     n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , 
     n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , 
     n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , 
     n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , 
     n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , 
     n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , 
     n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , 
     n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , 
     n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , 
     n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , 
     n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , 
     n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , 
     n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , 
     n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , 
     n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , 
     n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , 
     n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , 
     n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , 
     n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , 
     n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , 
     n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , 
     n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , 
     n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , 
     n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , 
     n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , 
     n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , 
     n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , 
     n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , 
     n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , 
     n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , 
     n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , 
     n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , 
     n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , 
     n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , 
     n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , 
     n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , 
     n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , 
     n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , 
     n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , 
     n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , 
     n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , 
     n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , 
     n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , 
     n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , 
     n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , 
     n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , 
     n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , 
     n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , 
     n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , 
     n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , 
     n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , 
     n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , 
     n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , 
     n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , 
     n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , 
     n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , 
     n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , 
     n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , 
     n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , 
     n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , 
     n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , 
     n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , 
     n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , 
     n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , 
     n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , 
     n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , 
     n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , 
     n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , 
     n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , 
     n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , 
     n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , 
     n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , 
     n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , 
     n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , 
     n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , 
     n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , 
     n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , 
     n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , 
     n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , 
     n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , 
     n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , 
     n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , 
     n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , 
     n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , 
     n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , 
     n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , 
     n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , 
     n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , 
     n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , 
     n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , 
     n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , 
     n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , 
     n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , 
     n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , 
     n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , 
     n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , 
     n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , 
     n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , 
     n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , 
     n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , 
     n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , 
     n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , 
     n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , 
     n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , 
     n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , 
     n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , 
     n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , 
     n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , 
     n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , 
     n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , 
     n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , 
     n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , 
     n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , 
     n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , 
     n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , 
     n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , 
     n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , 
     n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , 
     n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , 
     n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , 
     n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , 
     n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , 
     n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , 
     n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , 
     n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , 
     n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , 
     n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , 
     n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , 
     n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , 
     n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , 
     n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , 
     n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , 
     n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , 
     n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , 
     n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , 
     n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , 
     n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , 
     n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , 
     n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , 
     n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , 
     n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , 
     n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , 
     n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , 
     n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , 
     n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , 
     n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , 
     n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , 
     n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , 
     n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , 
     n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , 
     n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , 
     n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , 
     n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , 
     n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , 
     n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , 
     n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , 
     n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , 
     n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , 
     n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , 
     n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , 
     n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , 
     n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , 
     n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , 
     n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , 
     n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , 
     n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , 
     n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , 
     n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , 
     n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , 
     n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , 
     n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , 
     n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , 
     n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , 
     n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , 
     n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , 
     n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , 
     n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , 
     n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , 
     n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , 
     n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , 
     n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , 
     n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , 
     n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , 
     n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , 
     n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , 
     n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , 
     n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , 
     n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , 
     n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , 
     n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , 
     n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , 
     n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , 
     n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , 
     n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , 
     n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , 
     n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , 
     n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , 
     n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , 
     n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , 
     n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , 
     n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , 
     n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , 
     n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , 
     n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , 
     n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , 
     n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , 
     n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , 
     n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , 
     n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , 
     n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , 
     n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , 
     n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , 
     n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , 
     n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , 
     n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , 
     n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , 
     n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , 
     n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , 
     n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , 
     n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , 
     n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , 
     n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , 
     n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , 
     n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , 
     n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , 
     n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , 
     n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , 
     n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , 
     n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , 
     n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , 
     n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , 
     n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , 
     n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , 
     n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , 
     n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , 
     n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , 
     n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , 
     n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , 
     n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , 
     n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , 
     n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , 
     n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , 
     n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , 
     n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , 
     n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , 
     n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , 
     n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , 
     n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , 
     n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , 
     n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , 
     n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , 
     n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , 
     n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , 
     n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , 
     n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , 
     n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , 
     n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , 
     n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , 
     n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , 
     n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , 
     n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , 
     n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , 
     n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , 
     n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , 
     n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , 
     n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , 
     n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , 
     n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , 
     n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , 
     n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , 
     n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , 
     n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , 
     n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , 
     n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , 
     n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , 
     n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , 
     n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , 
     n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , 
     n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , 
     n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , 
     n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , 
     n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , 
     n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , 
     n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , 
     n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , 
     n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , 
     n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , 
     n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , 
     n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , 
     n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , 
     n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , 
     n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , 
     n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , 
     n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , 
     n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , 
     n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , 
     n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , 
     n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , 
     n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , 
     n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , 
     n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , 
     n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , 
     n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , 
     n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , 
     n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , 
     n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , 
     n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , 
     n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , 
     n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , 
     n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , 
     n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , 
     n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , 
     n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , 
     n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , 
     n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , 
     n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , 
     n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , 
     n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , 
     n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , 
     n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , 
     n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , 
     n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , 
     n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , 
     n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , 
     n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , 
     n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , 
     n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , 
     n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , 
     n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , 
     n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , 
     n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , 
     n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , 
     n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , 
     n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , 
     n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , 
     n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , 
     n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , 
     n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , 
     n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , 
     n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , 
     n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , 
     n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , 
     n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , 
     n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , 
     n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , 
     n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , 
     n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , 
     n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , 
     n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , 
     n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , 
     n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , 
     n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , 
     n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , 
     n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , 
     n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , 
     n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , 
     n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , 
     n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , 
     n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , 
     n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , 
     n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , 
     n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , 
     n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , 
     n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , 
     n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , 
     n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , 
     n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , 
     n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , 
     n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , 
     n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , 
     n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , 
     n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , 
     n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , 
     n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , 
     n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , 
     n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , 
     n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , 
     n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , 
     n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , 
     n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , 
     n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , 
     n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , 
     n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , 
     n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , 
     n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , 
     n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , 
     n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , 
     n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , 
     n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , 
     n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , 
     n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , 
     n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , 
     n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , 
     n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , 
     n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , 
     n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , 
     n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , 
     n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , 
     n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , 
     n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , 
     n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , 
     n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , 
     n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , 
     n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , 
     n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , 
     n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , 
     n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , 
     n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , 
     n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , 
     n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , 
     n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , 
     n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , 
     n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , 
     n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , 
     n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , 
     n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , 
     n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , 
     n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , 
     n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , 
     n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , 
     n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , 
     n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , 
     n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , 
     n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , 
     n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , 
     n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , 
     n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , 
     n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , 
     n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , 
     n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , 
     n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , 
     n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , 
     n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , 
     n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , 
     n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , 
     n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , 
     n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , 
     n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , 
     n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , 
     n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , 
     n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , 
     n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , 
     n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , 
     n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , 
     n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , 
     n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , 
     n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , 
     n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , 
     n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , 
     n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , 
     n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , 
     n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , 
     n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , 
     n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , 
     n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , 
     n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , 
     n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , 
     n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , 
     n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , 
     n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , 
     n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , 
     n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , 
     n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , 
     n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , 
     n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , 
     n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , 
     n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , 
     n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , 
     n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , 
     n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , 
     n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , 
     n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , 
     n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , 
     n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , 
     n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , 
     n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , 
     n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , 
     n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , 
     n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , 
     n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , 
     n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , 
     n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , 
     n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , 
     n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , 
     n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , 
     n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , 
     n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , 
     n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , 
     n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , 
     n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , 
     n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , 
     n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , 
     n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , 
     n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , 
     n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , 
     n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , 
     n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , 
     n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , 
     n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , 
     n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , 
     n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , 
     n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , 
     n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , 
     n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , 
     n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , 
     n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , 
     n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , 
     n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , 
     n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , 
     n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , 
     n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , 
     n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , 
     n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , 
     n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , 
     n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , 
     n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , 
     n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , 
     n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , 
     n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , 
     n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , 
     n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , 
     n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , 
     n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , 
     n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , 
     n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , 
     n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , 
     n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , 
     n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , 
     n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , 
     n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , 
     n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , 
     n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , 
     n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , 
     n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , 
     n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , 
     n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , 
     n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , 
     n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , 
     n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , 
     n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , 
     n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , 
     n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , 
     n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , 
     n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , 
     n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , 
     n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , 
     n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , 
     n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , 
     n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , 
     n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , 
     n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , 
     n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , 
     n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , 
     n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , 
     n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , 
     n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , 
     n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , 
     n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , 
     n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , 
     n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , 
     n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , 
     n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , 
     n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , 
     n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , 
     n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , 
     n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , 
     n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , 
     n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , 
     n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , 
     n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , 
     n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , 
     n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , 
     n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , 
     n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , 
     n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , 
     n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , 
     n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , 
     n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , 
     n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , 
     n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , 
     n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , 
     n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , 
     n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , 
     n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , 
     n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , 
     n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , 
     n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , 
     n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , 
     n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , 
     n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , 
     n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , 
     n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , 
     n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , 
     n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , 
     n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , 
     n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , 
     n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , 
     n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , 
     n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , 
     n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , 
     n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , 
     n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , 
     n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , 
     n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , 
     n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , 
     n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , 
     n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , 
     n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , 
     n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , 
     n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , 
     n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , 
     n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , 
     n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , 
     n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , 
     n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , 
     n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , 
     n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , 
     n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , 
     n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , 
     n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , 
     n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , 
     n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , 
     n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , 
     n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , 
     n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , 
     n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , 
     n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , 
     n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , 
     n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , 
     n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , 
     n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , 
     n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , 
     n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , 
     n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , 
     n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , 
     n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , 
     n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , 
     n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , 
     n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , 
     n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , 
     n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , 
     n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , 
     n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , 
     n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , 
     n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , 
     n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , 
     n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , 
     n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , 
     n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , 
     n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , 
     n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , 
     n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , 
     n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , 
     n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , 
     n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , 
     n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , 
     n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , 
     n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , 
     n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , 
     n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , 
     n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , 
     n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , 
     n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , 
     n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , 
     n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , 
     n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , 
     n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , 
     n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , 
     n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , 
     n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , 
     n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , 
     n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , 
     n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , 
     n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , 
     n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , 
     n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , 
     n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , 
     n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , 
     n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , 
     n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , 
     n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , 
     n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , 
     n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , 
     n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , 
     n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , 
     n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , 
     n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , 
     n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , 
     n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , 
     n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , 
     n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , 
     n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , 
     n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , 
     n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , 
     n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , 
     n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , 
     n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , 
     n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , 
     n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , 
     n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , 
     n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , 
     n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , 
     n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , 
     n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , 
     n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , 
     n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , 
     n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , 
     n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , 
     n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , 
     n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , 
     n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , 
     n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , 
     n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , 
     n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , 
     n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , 
     n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , 
     n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , 
     n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , 
     n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , 
     n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , 
     n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , 
     n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , 
     n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , 
     n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , 
     n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , 
     n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , 
     n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , 
     n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , 
     n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , 
     n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , 
     n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , 
     n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , 
     n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , 
     n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , 
     n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , 
     n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , 
     n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , 
     n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , 
     n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , 
     n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , 
     n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , 
     n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , 
     n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , 
     n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , 
     n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , 
     n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , 
     n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , 
     n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , 
     n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , 
     n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , 
     n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , 
     n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , 
     n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , 
     n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , 
     n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , 
     n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , 
     n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , 
     n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , 
     n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , 
     n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , 
     n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , 
     n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , 
     n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , 
     n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , 
     n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , 
     n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , 
     n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , 
     n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , 
     n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , 
     n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , 
     n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , 
     n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , 
     n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , 
     n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , 
     n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , 
     n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , 
     n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , 
     n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , 
     n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , 
     n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , 
     n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , 
     n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , 
     n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , 
     n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , 
     n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , 
     n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , 
     n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , 
     n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , 
     n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , 
     n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , 
     n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , 
     n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , 
     n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , 
     n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , 
     n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , 
     n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , 
     n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , 
     n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , 
     n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , 
     n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , 
     n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , 
     n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , 
     n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , 
     n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , 
     n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , 
     n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , 
     n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , 
     n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , 
     n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , 
     n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , 
     n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , 
     n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , 
     n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , 
     n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , 
     n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , 
     n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , 
     n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , 
     n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , 
     n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , 
     n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , 
     n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , 
     n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , 
     n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , 
     n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , 
     n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , 
     n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , 
     n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , 
     n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , 
     n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , 
     n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , 
     n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , 
     n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , 
     n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , 
     n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , 
     n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , 
     n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , 
     n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , 
     n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , 
     n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , 
     n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , 
     n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , 
     n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , 
     n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , 
     n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , 
     n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , 
     n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , 
     n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , 
     n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , 
     n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , 
     n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , 
     n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , 
     n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , 
     n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , 
     n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , 
     n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , 
     n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , 
     n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , 
     n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , 
     n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , 
     n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , 
     n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , 
     n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , 
     n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , 
     n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , 
     n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , 
     n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , 
     n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , 
     n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , 
     n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , 
     n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , 
     n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , 
     n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , 
     n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , 
     n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , 
     n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , 
     n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , 
     n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , 
     n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , 
     n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , 
     n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , 
     n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , 
     n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , 
     n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , 
     n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , 
     n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , 
     n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , 
     n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , 
     n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , 
     n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , 
     n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , 
     n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , 
     n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , 
     n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , 
     n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , 
     n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , 
     n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , 
     n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , 
     n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , 
     n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , 
     n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , 
     n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , 
     n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , 
     n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , 
     n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , 
     n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , 
     n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , 
     n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , 
     n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , 
     n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , 
     n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , 
     n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , 
     n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , 
     n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , 
     n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , 
     n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , 
     n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , 
     n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , 
     n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , 
     n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , 
     n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , 
     n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , 
     n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , 
     n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , 
     n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , 
     n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , 
     n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , 
     n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , 
     n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , 
     n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , 
     n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , 
     n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , 
     n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , 
     n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , 
     n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , 
     n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , 
     n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , 
     n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , 
     n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , 
     n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , 
     n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , 
     n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , 
     n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , 
     n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , 
     n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , 
     n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , 
     n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , 
     n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , 
     n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , 
     n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , 
     n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , 
     n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , 
     n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , 
     n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , 
     n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , 
     n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , 
     n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , 
     n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , 
     n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , 
     n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , 
     n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , 
     n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , 
     n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , 
     n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , 
     n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , 
     n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , 
     n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , 
     n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , 
     n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , 
     n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , 
     n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , 
     n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , 
     n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , 
     n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , 
     n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , 
     n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , 
     n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , 
     n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , 
     n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , 
     n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , 
     n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , 
     n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , 
     n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , 
     n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , 
     n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , 
     n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , 
     n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , 
     n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , 
     n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , 
     n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , 
     n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , 
     n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , 
     n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , 
     n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , 
     n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , 
     n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , 
     n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , 
     n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , 
     n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , 
     n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , 
     n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , 
     n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , 
     n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , 
     n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , 
     n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , 
     n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , 
     n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , 
     n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , 
     n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , 
     n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , 
     n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , 
     n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , 
     n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , 
     n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , 
     n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , 
     n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , 
     n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , 
     n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , 
     n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , 
     n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , 
     n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , 
     n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , 
     n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , 
     n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , 
     n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , 
     n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , 
     n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , 
     n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , 
     n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , 
     n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , 
     n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , 
     n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , 
     n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , 
     n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , 
     n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , 
     n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , 
     n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , 
     n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , 
     n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , 
     n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , 
     n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , 
     n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , 
     n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , 
     n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , 
     n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , 
     n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , 
     n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , 
     n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , 
     n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , 
     n10720 , n10721 , n10722 , n10723 , n10724 , n10725 ;
buf ( n1 , g0 );
buf ( n2 , g1 );
buf ( n3 , g2 );
buf ( n4 , g3 );
buf ( n5 , g4 );
buf ( n6 , g5 );
buf ( n7 , g6 );
buf ( n8 , g7 );
buf ( n9 , g8 );
buf ( n10 , g9 );
buf ( n11 , g10 );
buf ( n12 , g11 );
buf ( n13 , g12 );
buf ( n14 , g13 );
buf ( n15 , g14 );
buf ( n16 , g15 );
buf ( n17 , g16 );
buf ( n18 , g17 );
buf ( n19 , g18 );
buf ( n20 , g19 );
buf ( n21 , g20 );
buf ( n22 , g21 );
buf ( n23 , g22 );
buf ( n24 , g23 );
buf ( n25 , g24 );
buf ( n26 , g25 );
buf ( n27 , g26 );
buf ( n28 , g27 );
buf ( n29 , g28 );
buf ( n30 , g29 );
buf ( n31 , g30 );
buf ( n32 , g31 );
buf ( n33 , g32 );
buf ( n34 , g33 );
buf ( n35 , g34 );
buf ( n36 , g35 );
buf ( n37 , g36 );
buf ( n38 , g37 );
buf ( n39 , g38 );
buf ( n40 , g39 );
buf ( n41 , g40 );
buf ( n42 , g41 );
buf ( n43 , g42 );
buf ( n44 , g43 );
buf ( n45 , g44 );
buf ( n46 , g45 );
buf ( n47 , g46 );
buf ( n48 , g47 );
buf ( n49 , g48 );
buf ( n50 , g49 );
buf ( n51 , g50 );
buf ( n52 , g51 );
buf ( n53 , g52 );
buf ( n54 , g53 );
buf ( n55 , g54 );
buf ( n56 , g55 );
buf ( n57 , g56 );
buf ( n58 , g57 );
buf ( n59 , g58 );
buf ( n60 , g59 );
buf ( n61 , g60 );
buf ( n62 , g61 );
buf ( n63 , g62 );
buf ( n64 , g63 );
buf ( n65 , g64 );
buf ( n66 , g65 );
buf ( n67 , g66 );
buf ( n68 , g67 );
buf ( n69 , g68 );
buf ( n70 , g69 );
buf ( n71 , g70 );
buf ( n72 , g71 );
buf ( n73 , g72 );
buf ( n74 , g73 );
buf ( n75 , g74 );
buf ( n76 , g75 );
buf ( n77 , g76 );
buf ( n78 , g77 );
buf ( n79 , g78 );
buf ( n80 , g79 );
buf ( n81 , g80 );
buf ( n82 , g81 );
buf ( n83 , g82 );
buf ( n84 , g83 );
buf ( n85 , g84 );
buf ( n86 , g85 );
buf ( n87 , g86 );
buf ( n88 , g87 );
buf ( n89 , g88 );
buf ( n90 , g89 );
buf ( n91 , g90 );
buf ( n92 , g91 );
buf ( n93 , g92 );
buf ( n94 , g93 );
buf ( n95 , g94 );
buf ( n96 , g95 );
buf ( n97 , g96 );
buf ( n98 , g97 );
buf ( n99 , g98 );
buf ( g99 , n100 );
buf ( g100 , n101 );
buf ( g101 , n102 );
buf ( g102 , n103 );
buf ( g103 , n104 );
buf ( g104 , n105 );
buf ( g105 , n106 );
buf ( g106 , n107 );
buf ( g107 , n108 );
buf ( g108 , n109 );
buf ( g109 , n110 );
buf ( g110 , n111 );
buf ( g111 , n112 );
buf ( g112 , n113 );
buf ( g113 , n114 );
buf ( g114 , n115 );
buf ( g115 , n116 );
buf ( g116 , n117 );
buf ( g117 , n118 );
buf ( g118 , n119 );
buf ( g119 , n120 );
buf ( g120 , n121 );
buf ( g121 , n122 );
buf ( g122 , n123 );
buf ( g123 , n124 );
buf ( g124 , n125 );
buf ( g125 , n126 );
buf ( g126 , n127 );
buf ( g127 , n128 );
buf ( g128 , n129 );
buf ( g129 , n130 );
buf ( g130 , n131 );
buf ( g131 , n132 );
buf ( g132 , n133 );
buf ( g133 , n134 );
buf ( g134 , n135 );
buf ( g135 , n136 );
buf ( g136 , n137 );
buf ( g137 , n138 );
buf ( g138 , n139 );
buf ( g139 , n140 );
buf ( g140 , n141 );
buf ( g141 , n142 );
buf ( g142 , n143 );
buf ( g143 , n144 );
buf ( g144 , n145 );
buf ( g145 , n146 );
buf ( g146 , n147 );
buf ( g147 , n148 );
buf ( g148 , n149 );
buf ( g149 , n150 );
buf ( g150 , n151 );
buf ( g151 , n152 );
buf ( g152 , n153 );
buf ( g153 , n154 );
buf ( g154 , n155 );
buf ( g155 , n156 );
buf ( g156 , n157 );
buf ( g157 , n158 );
buf ( g158 , n159 );
buf ( g159 , n160 );
buf ( g160 , n161 );
buf ( g161 , n162 );
buf ( g162 , n163 );
buf ( g163 , n164 );
buf ( g164 , n165 );
buf ( g165 , n166 );
buf ( g166 , n167 );
buf ( g167 , n168 );
buf ( g168 , n169 );
buf ( g169 , n170 );
buf ( g170 , n171 );
buf ( g171 , n172 );
buf ( g172 , n173 );
buf ( g173 , n174 );
buf ( g174 , n175 );
buf ( g175 , n176 );
buf ( g176 , n177 );
buf ( g177 , n178 );
buf ( g178 , n179 );
buf ( g179 , n180 );
buf ( g180 , n181 );
buf ( g181 , n182 );
buf ( g182 , n183 );
buf ( g183 , n184 );
buf ( g184 , n185 );
buf ( g185 , n186 );
buf ( g186 , n187 );
buf ( g187 , n188 );
buf ( g188 , n189 );
buf ( g189 , n190 );
buf ( g190 , n191 );
buf ( g191 , n192 );
buf ( g192 , n193 );
buf ( g193 , n194 );
buf ( g194 , n195 );
buf ( g195 , n196 );
buf ( g196 , n197 );
buf ( g197 , n198 );
buf ( g198 , n199 );
buf ( g199 , n200 );
buf ( g200 , n201 );
buf ( g201 , n202 );
buf ( g202 , n203 );
buf ( g203 , n204 );
buf ( g204 , n205 );
buf ( g205 , n206 );
buf ( g206 , n207 );
buf ( g207 , n208 );
buf ( g208 , n209 );
buf ( g209 , n210 );
buf ( g210 , n211 );
buf ( g211 , n212 );
buf ( g212 , n213 );
buf ( g213 , n214 );
buf ( g214 , n215 );
buf ( g215 , n216 );
buf ( g216 , n217 );
buf ( g217 , n218 );
buf ( g218 , n219 );
buf ( g219 , n220 );
buf ( g220 , n221 );
buf ( g221 , n222 );
buf ( g222 , n223 );
buf ( g223 , n224 );
buf ( g224 , n225 );
buf ( g225 , n226 );
buf ( g226 , n227 );
buf ( n100 , 1'b0 );
buf ( n101 , 1'b0 );
buf ( n102 , 1'b0 );
buf ( n103 , 1'b0 );
buf ( n104 , 1'b0 );
buf ( n105 , 1'b0 );
buf ( n106 , 1'b0 );
buf ( n107 , 1'b0 );
buf ( n108 , 1'b0 );
buf ( n109 , 1'b0 );
buf ( n110 , 1'b0 );
buf ( n111 , 1'b0 );
buf ( n112 , 1'b0 );
buf ( n113 , 1'b0 );
buf ( n114 , 1'b0 );
buf ( n115 , 1'b0 );
buf ( n116 , 1'b0 );
buf ( n117 , 1'b0 );
buf ( n118 , 1'b0 );
buf ( n119 , 1'b0 );
buf ( n120 , 1'b0 );
buf ( n121 , 1'b0 );
buf ( n122 , 1'b0 );
buf ( n123 , 1'b0 );
buf ( n124 , 1'b0 );
buf ( n125 , 1'b0 );
buf ( n126 , 1'b0 );
buf ( n127 , 1'b0 );
buf ( n128 , 1'b0 );
buf ( n129 , 1'b0 );
buf ( n130 , 1'b0 );
buf ( n131 , n10424 );
buf ( n132 , n10416 );
buf ( n133 , n10427 );
buf ( n134 , n10358 );
buf ( n135 , n10447 );
buf ( n136 , n10445 );
buf ( n137 , n10531 );
buf ( n138 , n9989 );
buf ( n139 , n9995 );
buf ( n140 , n9684 );
buf ( n141 , n10539 );
buf ( n142 , n9267 );
buf ( n143 , n8903 );
buf ( n144 , n10579 );
buf ( n145 , n10584 );
buf ( n146 , n10567 );
buf ( n147 , n10568 );
buf ( n148 , n10619 );
buf ( n149 , n9024 );
buf ( n150 , n9035 );
buf ( n151 , n10631 );
buf ( n152 , n9007 );
buf ( n153 , n8998 );
buf ( n154 , n8988 );
buf ( n155 , n8984 );
buf ( n156 , n10701 );
buf ( n157 , n8976 );
buf ( n158 , n8965 );
buf ( n159 , n10720 );
buf ( n160 , n10707 );
buf ( n161 , n10709 );
buf ( n162 , n10711 );
buf ( n163 , n10713 );
buf ( n164 , 1'b0 );
buf ( n165 , 1'b0 );
buf ( n166 , 1'b0 );
buf ( n167 , 1'b0 );
buf ( n168 , 1'b0 );
buf ( n169 , 1'b0 );
buf ( n170 , 1'b0 );
buf ( n171 , 1'b0 );
buf ( n172 , 1'b0 );
buf ( n173 , 1'b0 );
buf ( n174 , 1'b0 );
buf ( n175 , 1'b0 );
buf ( n176 , 1'b0 );
buf ( n177 , 1'b0 );
buf ( n178 , 1'b0 );
buf ( n179 , 1'b0 );
buf ( n180 , 1'b0 );
buf ( n181 , 1'b0 );
buf ( n182 , 1'b0 );
buf ( n183 , 1'b0 );
buf ( n184 , 1'b0 );
buf ( n185 , 1'b0 );
buf ( n186 , 1'b0 );
buf ( n187 , 1'b0 );
buf ( n188 , 1'b0 );
buf ( n189 , 1'b0 );
buf ( n190 , 1'b0 );
buf ( n191 , 1'b0 );
buf ( n192 , 1'b0 );
buf ( n193 , 1'b0 );
buf ( n194 , 1'b0 );
buf ( n195 , 1'b0 );
buf ( n196 , 1'b0 );
buf ( n197 , 1'b0 );
buf ( n198 , n10530 );
buf ( n199 , n10426 );
buf ( n200 , n10725 );
buf ( n201 , n10719 );
buf ( n202 , n10434 );
buf ( n203 , n10443 );
buf ( n204 , n10453 );
buf ( n205 , n10462 );
buf ( n206 , n10472 );
buf ( n207 , n10483 );
buf ( n208 , n10493 );
buf ( n209 , n10505 );
buf ( n210 , n10543 );
buf ( n211 , n10557 );
buf ( n212 , n10564 );
buf ( n213 , n10582 );
buf ( n214 , n10590 );
buf ( n215 , n10600 );
buf ( n216 , n10613 );
buf ( n217 , n10625 );
buf ( n218 , n10638 );
buf ( n219 , n10646 );
buf ( n220 , n10656 );
buf ( n221 , n10668 );
buf ( n222 , n10674 );
buf ( n223 , n10680 );
buf ( n224 , n10685 );
buf ( n225 , n10693 );
buf ( n226 , n10700 );
buf ( n227 , n10705 );
and ( n295 , n3 , n4 );
not ( n296 , n3 );
and ( n297 , n296 , n20 );
nor ( n298 , n295 , n297 );
buf ( n299 , n298 );
not ( n300 , n299 );
buf ( n301 , n300 );
not ( n302 , n301 );
buf ( n303 , n302 );
not ( n304 , n38 );
and ( n305 , n303 , n304 );
nor ( n306 , n302 , n304 );
nor ( n307 , n305 , n306 );
not ( n308 , n307 );
and ( n309 , n3 , n6 );
not ( n310 , n3 );
and ( n311 , n310 , n22 );
nor ( n312 , n309 , n311 );
not ( n313 , n312 );
not ( n314 , n313 );
and ( n315 , n3 , n5 );
not ( n316 , n3 );
and ( n317 , n316 , n21 );
nor ( n318 , n315 , n317 );
nand ( n319 , n314 , n318 );
and ( n320 , n300 , n319 );
not ( n321 , n300 );
not ( n322 , n318 );
nand ( n323 , n313 , n322 );
and ( n324 , n321 , n323 );
or ( n325 , n320 , n324 );
not ( n326 , n325 );
not ( n327 , n326 );
not ( n328 , n327 );
not ( n329 , n328 );
or ( n330 , n308 , n329 );
nand ( n331 , n323 , n319 );
not ( n332 , n331 );
buf ( n333 , n332 );
not ( n334 , n333 );
not ( n335 , n303 );
or ( n336 , n335 , n37 );
not ( n337 , n37 );
nor ( n338 , n303 , n337 );
not ( n339 , n338 );
nand ( n340 , n336 , n339 );
or ( n341 , n334 , n340 );
nand ( n342 , n330 , n341 );
not ( n343 , n39 );
nor ( n344 , n303 , n343 );
xor ( n345 , n342 , n344 );
and ( n346 , n3 , n6 );
not ( n347 , n3 );
and ( n348 , n347 , n22 );
nor ( n349 , n346 , n348 );
not ( n350 , n349 );
not ( n351 , n350 );
not ( n352 , n351 );
and ( n353 , n3 , n8 );
not ( n354 , n3 );
and ( n355 , n354 , n24 );
nor ( n356 , n353 , n355 );
and ( n357 , n3 , n7 );
not ( n358 , n3 );
and ( n359 , n358 , n23 );
nor ( n360 , n357 , n359 );
nor ( n361 , n356 , n360 );
not ( n362 , n361 );
or ( n363 , n352 , n362 );
buf ( n364 , n356 );
nand ( n365 , n364 , n360 );
not ( n366 , n350 );
or ( n367 , n365 , n366 );
nand ( n368 , n363 , n367 );
not ( n369 , n368 );
buf ( n370 , n369 );
not ( n371 , n370 );
not ( n372 , n351 );
not ( n373 , n372 );
not ( n374 , n36 );
and ( n375 , n373 , n374 );
nor ( n376 , n373 , n374 );
nor ( n377 , n375 , n376 );
and ( n378 , n371 , n377 );
buf ( n379 , n349 );
not ( n380 , n379 );
not ( n381 , n380 );
or ( n382 , n361 , n381 );
not ( n383 , n382 );
and ( n384 , n383 , n365 );
nor ( n385 , n378 , n384 );
xor ( n386 , n345 , n385 );
not ( n387 , n361 );
nand ( n388 , n387 , n365 );
not ( n389 , n388 );
and ( n390 , n389 , n377 );
and ( n391 , n372 , n337 );
and ( n392 , n373 , n37 );
nor ( n393 , n391 , n392 );
nor ( n394 , n370 , n393 );
nor ( n395 , n390 , n394 );
not ( n396 , n10 );
and ( n397 , n396 , n3 );
nor ( n398 , n3 , n26 );
nor ( n399 , n397 , n398 );
not ( n400 , n25 );
or ( n401 , n400 , n3 );
nand ( n402 , n3 , n9 );
nand ( n403 , n401 , n402 );
and ( n404 , n399 , n403 );
and ( n405 , n3 , n8 );
not ( n406 , n3 );
and ( n407 , n406 , n24 );
nor ( n408 , n405 , n407 );
buf ( n409 , n408 );
nor ( n410 , n404 , n409 );
xor ( n411 , n395 , n410 );
nand ( n412 , n301 , n40 );
and ( n413 , n411 , n412 );
and ( n414 , n395 , n410 );
nor ( n415 , n413 , n414 );
xor ( n416 , n386 , n415 );
and ( n417 , n372 , n304 );
and ( n418 , n373 , n38 );
nor ( n419 , n417 , n418 );
or ( n420 , n370 , n419 );
not ( n421 , n389 );
or ( n422 , n421 , n393 );
nand ( n423 , n420 , n422 );
not ( n424 , n41 );
nor ( n425 , n302 , n424 );
xor ( n426 , n423 , n425 );
not ( n427 , n40 );
nand ( n428 , n302 , n427 );
and ( n429 , n412 , n428 );
not ( n430 , n429 );
not ( n431 , n328 );
or ( n432 , n430 , n431 );
and ( n433 , n303 , n343 );
nor ( n434 , n433 , n344 );
not ( n435 , n434 );
or ( n436 , n334 , n435 );
nand ( n437 , n432 , n436 );
and ( n438 , n426 , n437 );
and ( n439 , n423 , n425 );
nor ( n440 , n438 , n439 );
and ( n441 , n328 , n434 );
and ( n442 , n333 , n307 );
nor ( n443 , n441 , n442 );
not ( n444 , n403 );
and ( n445 , n3 , n10 );
not ( n446 , n3 );
and ( n447 , n446 , n26 );
nor ( n448 , n445 , n447 );
buf ( n449 , n448 );
nand ( n450 , n444 , n449 );
not ( n451 , n450 );
not ( n452 , n356 );
and ( n453 , n451 , n452 );
and ( n454 , n404 , n364 );
nor ( n455 , n453 , n454 );
not ( n456 , n455 );
and ( n457 , n409 , n374 );
not ( n458 , n409 );
and ( n459 , n458 , n36 );
nor ( n460 , n457 , n459 );
and ( n461 , n456 , n460 );
and ( n462 , n410 , n450 );
nor ( n463 , n461 , n462 );
xnor ( n464 , n443 , n463 );
or ( n465 , n440 , n464 );
or ( n466 , n443 , n463 );
nand ( n467 , n465 , n466 );
and ( n468 , n416 , n467 );
and ( n469 , n386 , n415 );
nor ( n470 , n468 , n469 );
not ( n471 , n470 );
or ( n472 , n327 , n340 );
and ( n473 , n335 , n374 );
and ( n474 , n303 , n36 );
nor ( n475 , n473 , n474 );
or ( n476 , n334 , n475 );
nand ( n477 , n472 , n476 );
or ( n478 , n477 , n383 );
nand ( n479 , n477 , n383 );
nand ( n480 , n478 , n479 );
xnor ( n481 , n480 , n306 );
xnor ( n482 , n481 , n385 );
and ( n483 , n345 , n385 );
and ( n484 , n342 , n344 );
nor ( n485 , n483 , n484 );
xor ( n486 , n482 , n485 );
not ( n487 , n486 );
and ( n488 , n471 , n487 );
and ( n489 , n470 , n486 );
nor ( n490 , n488 , n489 );
not ( n491 , n490 );
not ( n492 , n491 );
xnor ( n493 , n416 , n467 );
not ( n494 , n493 );
xnor ( n495 , n440 , n464 );
xor ( n496 , n395 , n410 );
xor ( n497 , n496 , n412 );
xor ( n498 , n495 , n497 );
not ( n499 , n404 );
nand ( n500 , n499 , n450 );
not ( n501 , n500 );
and ( n502 , n501 , n460 );
not ( n503 , n456 );
buf ( n504 , n409 );
not ( n505 , n504 );
not ( n506 , n37 );
and ( n507 , n505 , n506 );
and ( n508 , n504 , n37 );
nor ( n509 , n507 , n508 );
nor ( n510 , n503 , n509 );
nor ( n511 , n502 , n510 );
not ( n512 , n12 );
and ( n513 , n512 , n3 );
nor ( n514 , n3 , n28 );
nor ( n515 , n513 , n514 );
not ( n516 , n11 );
and ( n517 , n3 , n516 );
not ( n518 , n3 );
not ( n519 , n27 );
and ( n520 , n518 , n519 );
nor ( n521 , n517 , n520 );
nand ( n522 , n515 , n521 );
not ( n523 , n522 );
buf ( n524 , n449 );
nor ( n525 , n523 , n524 );
xnor ( n526 , n511 , n525 );
and ( n527 , n303 , n424 );
nor ( n528 , n527 , n425 );
and ( n529 , n328 , n528 );
and ( n530 , n333 , n429 );
nor ( n531 , n529 , n530 );
or ( n532 , n526 , n531 );
or ( n533 , n511 , n525 );
nand ( n534 , n532 , n533 );
xor ( n535 , n534 , n463 );
xor ( n536 , n426 , n437 );
and ( n537 , n535 , n536 );
and ( n538 , n534 , n463 );
nor ( n539 , n537 , n538 );
and ( n540 , n498 , n539 );
and ( n541 , n495 , n497 );
nor ( n542 , n540 , n541 );
not ( n543 , n542 );
or ( n544 , n494 , n543 );
or ( n545 , n542 , n493 );
nand ( n546 , n544 , n545 );
not ( n547 , n546 );
xor ( n548 , n495 , n497 );
xor ( n549 , n548 , n539 );
not ( n550 , n549 );
xnor ( n551 , n535 , n536 );
xnor ( n552 , n372 , n39 );
or ( n553 , n370 , n552 );
or ( n554 , n421 , n419 );
nand ( n555 , n553 , n554 );
and ( n556 , n42 , n300 );
xor ( n557 , n555 , n556 );
and ( n558 , n409 , n38 );
not ( n559 , n409 );
and ( n560 , n559 , n304 );
nor ( n561 , n558 , n560 );
or ( n562 , n503 , n561 );
not ( n563 , n501 );
or ( n564 , n563 , n509 );
nand ( n565 , n562 , n564 );
and ( n566 , n557 , n565 );
and ( n567 , n555 , n556 );
nor ( n568 , n566 , n567 );
xnor ( n569 , n551 , n568 );
xor ( n570 , n42 , n300 );
and ( n571 , n328 , n570 );
and ( n572 , n333 , n528 );
nor ( n573 , n571 , n572 );
nand ( n574 , n301 , n43 );
xor ( n575 , n573 , n574 );
not ( n576 , n524 );
not ( n577 , n523 );
or ( n578 , n576 , n577 );
and ( n579 , n3 , n12 );
not ( n580 , n3 );
and ( n581 , n580 , n28 );
nor ( n582 , n579 , n581 );
and ( n583 , n3 , n11 );
not ( n584 , n3 );
and ( n585 , n584 , n27 );
nor ( n586 , n583 , n585 );
buf ( n587 , n586 );
nand ( n588 , n582 , n587 );
not ( n589 , n588 );
buf ( n590 , n399 );
nand ( n591 , n589 , n590 );
nand ( n592 , n578 , n591 );
not ( n593 , n592 );
not ( n594 , n593 );
buf ( n595 , n590 );
xor ( n596 , n36 , n595 );
and ( n597 , n594 , n596 );
and ( n598 , n525 , n588 );
nor ( n599 , n597 , n598 );
and ( n600 , n575 , n599 );
and ( n601 , n573 , n574 );
nor ( n602 , n600 , n601 );
xor ( n603 , n526 , n531 );
xor ( n604 , n602 , n603 );
xor ( n605 , n557 , n565 );
and ( n606 , n604 , n605 );
and ( n607 , n602 , n603 );
nor ( n608 , n606 , n607 );
or ( n609 , n569 , n608 );
or ( n610 , n551 , n568 );
nand ( n611 , n609 , n610 );
not ( n612 , n611 );
or ( n613 , n550 , n612 );
or ( n614 , n611 , n549 );
nand ( n615 , n613 , n614 );
not ( n616 , n615 );
xor ( n617 , n569 , n608 );
not ( n618 , n617 );
xor ( n619 , n602 , n603 );
xor ( n620 , n619 , n605 );
or ( n621 , n301 , n43 );
nand ( n622 , n621 , n574 );
or ( n623 , n327 , n622 );
not ( n624 , n570 );
or ( n625 , n334 , n624 );
nand ( n626 , n623 , n625 );
xnor ( n627 , n505 , n39 );
or ( n628 , n503 , n627 );
or ( n629 , n563 , n561 );
nand ( n630 , n628 , n629 );
xor ( n631 , n626 , n630 );
and ( n632 , n44 , n300 );
and ( n633 , n631 , n632 );
and ( n634 , n626 , n630 );
nor ( n635 , n633 , n634 );
not ( n636 , n40 );
not ( n637 , n312 );
or ( n638 , n636 , n637 );
or ( n639 , n379 , n40 );
nand ( n640 , n638 , n639 );
not ( n641 , n640 );
or ( n642 , n370 , n641 );
or ( n643 , n421 , n552 );
nand ( n644 , n642 , n643 );
and ( n645 , n565 , n644 );
not ( n646 , n565 );
not ( n647 , n644 );
and ( n648 , n646 , n647 );
nor ( n649 , n645 , n648 );
or ( n650 , n635 , n649 );
or ( n651 , n647 , n565 );
nand ( n652 , n650 , n651 );
xor ( n653 , n620 , n652 );
xor ( n654 , n573 , n574 );
xor ( n655 , n654 , n599 );
not ( n656 , n596 );
and ( n657 , n588 , n522 );
not ( n658 , n657 );
or ( n659 , n656 , n658 );
and ( n660 , n37 , n524 );
not ( n661 , n37 );
and ( n662 , n661 , n595 );
nor ( n663 , n660 , n662 );
or ( n664 , n593 , n663 );
nand ( n665 , n659 , n664 );
not ( n666 , n515 );
not ( n667 , n666 );
not ( n668 , n13 );
and ( n669 , n3 , n668 );
not ( n670 , n3 );
not ( n671 , n29 );
and ( n672 , n670 , n671 );
nor ( n673 , n669 , n672 );
not ( n674 , n673 );
not ( n675 , n674 );
and ( n676 , n3 , n14 );
not ( n677 , n3 );
and ( n678 , n677 , n30 );
or ( n679 , n676 , n678 );
nand ( n680 , n675 , n679 );
nand ( n681 , n667 , n680 );
not ( n682 , n681 );
or ( n683 , n665 , n682 );
nand ( n684 , n665 , n682 );
nand ( n685 , n683 , n684 );
and ( n686 , n372 , n424 );
not ( n687 , n372 );
and ( n688 , n687 , n41 );
nor ( n689 , n686 , n688 );
or ( n690 , n370 , n689 );
or ( n691 , n421 , n641 );
nand ( n692 , n690 , n691 );
and ( n693 , n685 , n692 );
and ( n694 , n665 , n681 );
nor ( n695 , n693 , n694 );
xor ( n696 , n655 , n695 );
xnor ( n697 , n635 , n649 );
and ( n698 , n696 , n697 );
and ( n699 , n655 , n695 );
or ( n700 , n698 , n699 );
not ( n701 , n700 );
and ( n702 , n653 , n701 );
and ( n703 , n620 , n652 );
nor ( n704 , n702 , n703 );
not ( n705 , n704 );
or ( n706 , n618 , n705 );
or ( n707 , n704 , n617 );
nand ( n708 , n706 , n707 );
not ( n709 , n708 );
xor ( n710 , n44 , n300 );
not ( n711 , n710 );
or ( n712 , n325 , n711 );
or ( n713 , n334 , n622 );
nand ( n714 , n712 , n713 );
not ( n715 , n714 );
not ( n716 , n42 );
not ( n717 , n312 );
or ( n718 , n716 , n717 );
or ( n719 , n379 , n42 );
nand ( n720 , n718 , n719 );
not ( n721 , n720 );
or ( n722 , n370 , n721 );
or ( n723 , n421 , n689 );
nand ( n724 , n722 , n723 );
and ( n725 , n715 , n724 );
not ( n726 , n724 );
and ( n727 , n726 , n714 );
nor ( n728 , n725 , n727 );
not ( n729 , n666 );
nor ( n730 , n680 , n729 );
not ( n731 , n730 );
and ( n732 , n3 , n14 );
not ( n733 , n3 );
and ( n734 , n733 , n30 );
nor ( n735 , n732 , n734 );
and ( n736 , n3 , n13 );
not ( n737 , n3 );
and ( n738 , n737 , n29 );
nor ( n739 , n736 , n738 );
and ( n740 , n735 , n739 );
nand ( n741 , n740 , n729 );
nand ( n742 , n731 , n741 );
and ( n743 , n3 , n12 );
not ( n744 , n3 );
and ( n745 , n744 , n28 );
nor ( n746 , n743 , n745 );
buf ( n747 , n746 );
not ( n748 , n747 );
nand ( n749 , n748 , n36 );
not ( n750 , n749 );
not ( n751 , n746 );
not ( n752 , n751 );
and ( n753 , n752 , n374 );
nor ( n754 , n750 , n753 );
and ( n755 , n742 , n754 );
buf ( n756 , n739 );
nand ( n757 , n735 , n756 );
and ( n758 , n682 , n757 );
nor ( n759 , n755 , n758 );
or ( n760 , n728 , n759 );
or ( n761 , n726 , n715 );
nand ( n762 , n760 , n761 );
not ( n763 , n449 );
not ( n764 , n38 );
and ( n765 , n763 , n764 );
not ( n766 , n448 );
not ( n767 , n766 );
and ( n768 , n767 , n38 );
nor ( n769 , n765 , n768 );
or ( n770 , n593 , n769 );
not ( n771 , n657 );
or ( n772 , n771 , n663 );
nand ( n773 , n770 , n772 );
xor ( n774 , n762 , n773 );
xor ( n775 , n631 , n632 );
and ( n776 , n774 , n775 );
and ( n777 , n762 , n773 );
nor ( n778 , n776 , n777 );
xor ( n779 , n655 , n695 );
xor ( n780 , n779 , n697 );
and ( n781 , n778 , n780 );
xor ( n782 , n774 , n775 );
xor ( n783 , n685 , n692 );
not ( n784 , n409 );
not ( n785 , n40 );
and ( n786 , n784 , n785 );
and ( n787 , n409 , n40 );
nor ( n788 , n786 , n787 );
or ( n789 , n503 , n788 );
or ( n790 , n563 , n627 );
nand ( n791 , n789 , n790 );
nand ( n792 , n300 , n45 );
not ( n793 , n792 );
xor ( n794 , n791 , n793 );
not ( n795 , n773 );
and ( n796 , n794 , n795 );
and ( n797 , n791 , n793 );
nor ( n798 , n796 , n797 );
not ( n799 , n798 );
and ( n800 , n783 , n799 );
not ( n801 , n783 );
and ( n802 , n801 , n798 );
nor ( n803 , n800 , n802 );
and ( n804 , n782 , n803 );
and ( n805 , n783 , n799 );
nor ( n806 , n804 , n805 );
xor ( n807 , n655 , n695 );
xor ( n808 , n807 , n697 );
and ( n809 , n806 , n808 );
and ( n810 , n778 , n806 );
or ( n811 , n781 , n809 , n810 );
not ( n812 , n811 );
not ( n813 , n812 );
xnor ( n814 , n653 , n701 );
not ( n815 , n814 );
or ( n816 , n813 , n815 );
or ( n817 , n814 , n812 );
nand ( n818 , n816 , n817 );
not ( n819 , n818 );
xor ( n820 , n655 , n695 );
xor ( n821 , n820 , n697 );
xor ( n822 , n778 , n806 );
xor ( n823 , n821 , n822 );
not ( n824 , n823 );
not ( n825 , n43 );
and ( n826 , n372 , n825 );
not ( n827 , n372 );
and ( n828 , n827 , n43 );
nor ( n829 , n826 , n828 );
or ( n830 , n369 , n829 );
or ( n831 , n421 , n721 );
nand ( n832 , n830 , n831 );
and ( n833 , n595 , n343 );
and ( n834 , n524 , n39 );
nor ( n835 , n833 , n834 );
or ( n836 , n593 , n835 );
or ( n837 , n771 , n769 );
nand ( n838 , n836 , n837 );
xor ( n839 , n832 , n838 );
not ( n840 , n45 );
not ( n841 , n840 );
not ( n842 , n299 );
or ( n843 , n841 , n842 );
nand ( n844 , n843 , n792 );
or ( n845 , n327 , n844 );
or ( n846 , n334 , n711 );
nand ( n847 , n845 , n846 );
and ( n848 , n839 , n847 );
and ( n849 , n832 , n838 );
nor ( n850 , n848 , n849 );
not ( n851 , n754 );
not ( n852 , n740 );
nand ( n853 , n852 , n680 );
buf ( n854 , n853 );
not ( n855 , n854 );
not ( n856 , n855 );
or ( n857 , n851 , n856 );
not ( n858 , n757 );
not ( n859 , n747 );
and ( n860 , n858 , n859 );
not ( n861 , n751 );
not ( n862 , n861 );
nor ( n863 , n862 , n680 );
nor ( n864 , n860 , n863 );
not ( n865 , n37 );
not ( n866 , n747 );
or ( n867 , n865 , n866 );
or ( n868 , n747 , n37 );
nand ( n869 , n867 , n868 );
not ( n870 , n869 );
or ( n871 , n864 , n870 );
nand ( n872 , n857 , n871 );
not ( n873 , n15 );
and ( n874 , n3 , n873 );
not ( n875 , n3 );
not ( n876 , n31 );
and ( n877 , n875 , n876 );
nor ( n878 , n874 , n877 );
buf ( n879 , n878 );
not ( n880 , n16 );
and ( n881 , n880 , n3 );
nor ( n882 , n3 , n32 );
nor ( n883 , n881 , n882 );
nand ( n884 , n879 , n883 );
not ( n885 , n884 );
and ( n886 , n3 , n14 );
not ( n887 , n3 );
and ( n888 , n887 , n30 );
nor ( n889 , n886 , n888 );
buf ( n890 , n889 );
nor ( n891 , n885 , n890 );
or ( n892 , n872 , n891 );
nand ( n893 , n872 , n891 );
nand ( n894 , n892 , n893 );
and ( n895 , n505 , n424 );
and ( n896 , n409 , n41 );
nor ( n897 , n895 , n896 );
or ( n898 , n503 , n897 );
or ( n899 , n563 , n788 );
nand ( n900 , n898 , n899 );
and ( n901 , n894 , n900 );
not ( n902 , n891 );
and ( n903 , n872 , n902 );
nor ( n904 , n901 , n903 );
xor ( n905 , n850 , n904 );
xnor ( n906 , n728 , n759 );
and ( n907 , n905 , n906 );
and ( n908 , n850 , n904 );
nor ( n909 , n907 , n908 );
not ( n910 , n909 );
xor ( n911 , n782 , n803 );
not ( n912 , n911 );
or ( n913 , n910 , n912 );
xnor ( n914 , n911 , n909 );
xnor ( n915 , n839 , n847 );
not ( n916 , n46 );
not ( n917 , n916 );
not ( n918 , n299 );
or ( n919 , n917 , n918 );
nand ( n920 , n300 , n46 );
nand ( n921 , n919 , n920 );
not ( n922 , n921 );
not ( n923 , n922 );
not ( n924 , n326 );
or ( n925 , n923 , n924 );
not ( n926 , n844 );
nand ( n927 , n926 , n332 );
nand ( n928 , n925 , n927 );
not ( n929 , n449 );
and ( n930 , n40 , n929 );
not ( n931 , n40 );
and ( n932 , n931 , n767 );
nor ( n933 , n930 , n932 );
not ( n934 , n933 );
or ( n935 , n593 , n934 );
or ( n936 , n771 , n835 );
nand ( n937 , n935 , n936 );
xor ( n938 , n928 , n937 );
and ( n939 , n47 , n300 );
and ( n940 , n938 , n939 );
and ( n941 , n928 , n937 );
nor ( n942 , n940 , n941 );
xor ( n943 , n915 , n942 );
xnor ( n944 , n894 , n900 );
and ( n945 , n943 , n944 );
and ( n946 , n915 , n942 );
nor ( n947 , n945 , n946 );
not ( n948 , n304 );
not ( n949 , n729 );
or ( n950 , n948 , n949 );
nand ( n951 , n861 , n38 );
nand ( n952 , n950 , n951 );
not ( n953 , n952 );
or ( n954 , n864 , n953 );
or ( n955 , n854 , n870 );
nand ( n956 , n954 , n955 );
not ( n957 , n42 );
not ( n958 , n409 );
or ( n959 , n957 , n958 );
or ( n960 , n409 , n42 );
nand ( n961 , n959 , n960 );
not ( n962 , n961 );
or ( n963 , n503 , n962 );
or ( n964 , n563 , n897 );
nand ( n965 , n963 , n964 );
xor ( n966 , n956 , n965 );
not ( n967 , n366 );
not ( n968 , n44 );
and ( n969 , n967 , n968 );
and ( n970 , n351 , n44 );
nor ( n971 , n969 , n970 );
or ( n972 , n370 , n971 );
or ( n973 , n421 , n829 );
nand ( n974 , n972 , n973 );
and ( n975 , n966 , n974 );
and ( n976 , n956 , n965 );
nor ( n977 , n975 , n976 );
and ( n978 , n3 , n15 );
not ( n979 , n3 );
and ( n980 , n979 , n31 );
nor ( n981 , n978 , n980 );
and ( n982 , n3 , n16 );
not ( n983 , n3 );
and ( n984 , n983 , n32 );
nor ( n985 , n982 , n984 );
nand ( n986 , n981 , n985 );
not ( n987 , n986 );
and ( n988 , n3 , n14 );
not ( n989 , n3 );
and ( n990 , n989 , n30 );
nor ( n991 , n988 , n990 );
buf ( n992 , n991 );
not ( n993 , n992 );
and ( n994 , n987 , n993 );
and ( n995 , n885 , n890 );
nor ( n996 , n994 , n995 );
not ( n997 , n996 );
not ( n998 , n997 );
not ( n999 , n374 );
not ( n1000 , n889 );
or ( n1001 , n999 , n1000 );
or ( n1002 , n992 , n374 );
nand ( n1003 , n1001 , n1002 );
or ( n1004 , n998 , n1003 );
not ( n1005 , n986 );
or ( n1006 , n902 , n1005 );
nand ( n1007 , n1004 , n1006 );
not ( n1008 , n1007 );
not ( n1009 , n920 );
and ( n1010 , n1008 , n1009 );
and ( n1011 , n1007 , n920 );
nor ( n1012 , n1010 , n1011 );
or ( n1013 , n977 , n1012 );
not ( n1014 , n1007 );
or ( n1015 , n1014 , n920 );
nand ( n1016 , n1013 , n1015 );
and ( n1017 , n794 , n795 );
not ( n1018 , n794 );
and ( n1019 , n1018 , n773 );
nor ( n1020 , n1017 , n1019 );
xnor ( n1021 , n1016 , n1020 );
or ( n1022 , n947 , n1021 );
or ( n1023 , n1016 , n1020 );
nand ( n1024 , n1022 , n1023 );
or ( n1025 , n914 , n1024 );
nand ( n1026 , n913 , n1025 );
not ( n1027 , n1026 );
or ( n1028 , n824 , n1027 );
or ( n1029 , n1026 , n823 );
nand ( n1030 , n1028 , n1029 );
not ( n1031 , n1030 );
xnor ( n1032 , n914 , n1024 );
not ( n1033 , n1032 );
xor ( n1034 , n947 , n1021 );
xor ( n1035 , n850 , n904 );
xor ( n1036 , n1035 , n906 );
xor ( n1037 , n1034 , n1036 );
and ( n1038 , n372 , n840 );
and ( n1039 , n366 , n45 );
nor ( n1040 , n1038 , n1039 );
or ( n1041 , n369 , n1040 );
or ( n1042 , n388 , n971 );
nand ( n1043 , n1041 , n1042 );
and ( n1044 , n667 , n343 );
and ( n1045 , n747 , n39 );
nor ( n1046 , n1044 , n1045 );
or ( n1047 , n864 , n1046 );
or ( n1048 , n854 , n953 );
nand ( n1049 , n1047 , n1048 );
xor ( n1050 , n1043 , n1049 );
not ( n1051 , n1050 );
not ( n1052 , n1051 );
xor ( n1053 , n47 , n300 );
and ( n1054 , n326 , n1053 );
and ( n1055 , n333 , n922 );
nor ( n1056 , n1054 , n1055 );
not ( n1057 , n1056 );
and ( n1058 , n1052 , n1057 );
and ( n1059 , n1043 , n1049 );
nor ( n1060 , n1058 , n1059 );
xnor ( n1061 , n938 , n939 );
xnor ( n1062 , n1060 , n1061 );
not ( n1063 , n1062 );
xor ( n1064 , n966 , n974 );
not ( n1065 , n1064 );
and ( n1066 , n1063 , n1065 );
and ( n1067 , n1060 , n1061 );
nor ( n1068 , n1066 , n1067 );
xor ( n1069 , n977 , n1012 );
and ( n1070 , n524 , n424 );
not ( n1071 , n524 );
and ( n1072 , n1071 , n41 );
nor ( n1073 , n1070 , n1072 );
not ( n1074 , n1073 );
or ( n1075 , n593 , n1074 );
or ( n1076 , n771 , n934 );
nand ( n1077 , n1075 , n1076 );
and ( n1078 , n3 , n4 );
not ( n1079 , n3 );
and ( n1080 , n1079 , n20 );
nor ( n1081 , n1078 , n1080 );
not ( n1082 , n1081 );
nand ( n1083 , n1082 , n48 );
not ( n1084 , n1083 );
xor ( n1085 , n1077 , n1084 );
and ( n1086 , n505 , n825 );
and ( n1087 , n504 , n43 );
nor ( n1088 , n1086 , n1087 );
or ( n1089 , n503 , n1088 );
or ( n1090 , n563 , n962 );
nand ( n1091 , n1089 , n1090 );
and ( n1092 , n1085 , n1091 );
and ( n1093 , n1077 , n1084 );
nor ( n1094 , n1092 , n1093 );
not ( n1095 , n991 );
not ( n1096 , n1095 );
not ( n1097 , n1096 );
not ( n1098 , n37 );
and ( n1099 , n1097 , n1098 );
and ( n1100 , n992 , n37 );
nor ( n1101 , n1099 , n1100 );
or ( n1102 , n998 , n1101 );
and ( n1103 , n884 , n986 );
buf ( n1104 , n1103 );
not ( n1105 , n1104 );
or ( n1106 , n1105 , n1003 );
nand ( n1107 , n1102 , n1106 );
buf ( n1108 , n985 );
buf ( n1109 , n1108 );
nor ( n1110 , n1107 , n1109 );
and ( n1111 , n1110 , n1014 );
not ( n1112 , n1110 );
and ( n1113 , n1112 , n1007 );
nor ( n1114 , n1111 , n1113 );
or ( n1115 , n1094 , n1114 );
or ( n1116 , n1110 , n1007 );
nand ( n1117 , n1115 , n1116 );
xor ( n1118 , n1069 , n1117 );
and ( n1119 , n1068 , n1118 );
and ( n1120 , n1069 , n1117 );
nor ( n1121 , n1119 , n1120 );
and ( n1122 , n1037 , n1121 );
and ( n1123 , n1034 , n1036 );
nor ( n1124 , n1122 , n1123 );
not ( n1125 , n1124 );
or ( n1126 , n1033 , n1125 );
or ( n1127 , n1124 , n1032 );
nand ( n1128 , n1126 , n1127 );
not ( n1129 , n1128 );
xnor ( n1130 , n1068 , n1118 );
xor ( n1131 , n943 , n944 );
xnor ( n1132 , n1130 , n1131 );
xor ( n1133 , n1094 , n1114 );
not ( n1134 , n299 );
nand ( n1135 , n1134 , n49 );
not ( n1136 , n1135 );
not ( n1137 , n1136 );
not ( n1138 , n42 );
not ( n1139 , n449 );
or ( n1140 , n1138 , n1139 );
or ( n1141 , n767 , n42 );
nand ( n1142 , n1140 , n1141 );
not ( n1143 , n1142 );
not ( n1144 , n592 );
or ( n1145 , n1143 , n1144 );
nand ( n1146 , n657 , n1073 );
nand ( n1147 , n1145 , n1146 );
not ( n1148 , n1147 );
or ( n1149 , n1137 , n1148 );
not ( n1150 , n1135 );
not ( n1151 , n1147 );
or ( n1152 , n1150 , n1151 );
or ( n1153 , n1147 , n1135 );
nand ( n1154 , n1152 , n1153 );
not ( n1155 , n44 );
not ( n1156 , n409 );
or ( n1157 , n1155 , n1156 );
or ( n1158 , n409 , n44 );
nand ( n1159 , n1157 , n1158 );
not ( n1160 , n1159 );
or ( n1161 , n503 , n1160 );
or ( n1162 , n563 , n1088 );
nand ( n1163 , n1161 , n1162 );
nand ( n1164 , n1154 , n1163 );
nand ( n1165 , n1149 , n1164 );
not ( n1166 , n1165 );
not ( n1167 , n38 );
not ( n1168 , n889 );
or ( n1169 , n1167 , n1168 );
or ( n1170 , n992 , n38 );
nand ( n1171 , n1169 , n1170 );
not ( n1172 , n1171 );
or ( n1173 , n998 , n1172 );
buf ( n1174 , n1103 );
not ( n1175 , n1174 );
or ( n1176 , n1175 , n1101 );
nand ( n1177 , n1173 , n1176 );
not ( n1178 , n374 );
buf ( n1179 , n883 );
not ( n1180 , n1179 );
or ( n1181 , n1178 , n1180 );
and ( n1182 , n3 , n17 );
not ( n1183 , n3 );
and ( n1184 , n1183 , n33 );
nor ( n1185 , n1182 , n1184 );
not ( n1186 , n1185 );
and ( n1187 , n883 , n1186 );
not ( n1188 , n1187 );
nand ( n1189 , n1181 , n1188 );
nand ( n1190 , n1177 , n1189 );
not ( n1191 , n1190 );
and ( n1192 , n1166 , n1191 );
and ( n1193 , n1165 , n1190 );
nor ( n1194 , n1192 , n1193 );
not ( n1195 , n312 );
not ( n1196 , n46 );
and ( n1197 , n1195 , n1196 );
and ( n1198 , n351 , n46 );
nor ( n1199 , n1197 , n1198 );
not ( n1200 , n1199 );
not ( n1201 , n1200 );
not ( n1202 , n368 );
or ( n1203 , n1201 , n1202 );
or ( n1204 , n388 , n1040 );
nand ( n1205 , n1203 , n1204 );
not ( n1206 , n40 );
not ( n1207 , n861 );
or ( n1208 , n1206 , n1207 );
or ( n1209 , n747 , n40 );
nand ( n1210 , n1208 , n1209 );
not ( n1211 , n1210 );
not ( n1212 , n742 );
or ( n1213 , n1211 , n1212 );
not ( n1214 , n1046 );
nand ( n1215 , n1214 , n855 );
nand ( n1216 , n1213 , n1215 );
xor ( n1217 , n1205 , n1216 );
not ( n1218 , n48 );
nand ( n1219 , n1218 , n1081 );
nand ( n1220 , n1219 , n1083 );
not ( n1221 , n1220 );
buf ( n1222 , n1221 );
not ( n1223 , n1222 );
not ( n1224 , n326 );
or ( n1225 , n1223 , n1224 );
not ( n1226 , n1053 );
or ( n1227 , n334 , n1226 );
nand ( n1228 , n1225 , n1227 );
and ( n1229 , n1217 , n1228 );
and ( n1230 , n1205 , n1216 );
nor ( n1231 , n1229 , n1230 );
or ( n1232 , n1194 , n1231 );
not ( n1233 , n1165 );
or ( n1234 , n1233 , n1190 );
nand ( n1235 , n1232 , n1234 );
xor ( n1236 , n1133 , n1235 );
not ( n1237 , n1050 );
not ( n1238 , n1056 );
and ( n1239 , n1237 , n1238 );
and ( n1240 , n1050 , n1056 );
nor ( n1241 , n1239 , n1240 );
and ( n1242 , n1107 , n1109 );
nor ( n1243 , n1242 , n1110 );
xor ( n1244 , n1241 , n1243 );
xnor ( n1245 , n1085 , n1091 );
and ( n1246 , n1244 , n1245 );
and ( n1247 , n1241 , n1243 );
nor ( n1248 , n1246 , n1247 );
and ( n1249 , n1236 , n1248 );
and ( n1250 , n1235 , n1133 );
nor ( n1251 , n1249 , n1250 );
or ( n1252 , n1132 , n1251 );
or ( n1253 , n1130 , n1131 );
nand ( n1254 , n1252 , n1253 );
not ( n1255 , n1254 );
xor ( n1256 , n1034 , n1036 );
xor ( n1257 , n1256 , n1121 );
not ( n1258 , n1257 );
or ( n1259 , n1255 , n1258 );
or ( n1260 , n1257 , n1254 );
nand ( n1261 , n1259 , n1260 );
not ( n1262 , n1261 );
xor ( n1263 , n1132 , n1251 );
not ( n1264 , n1263 );
xnor ( n1265 , n1062 , n1064 );
not ( n1266 , n1265 );
xor ( n1267 , n1194 , n1231 );
or ( n1268 , n1177 , n1189 );
nand ( n1269 , n1268 , n1190 );
not ( n1270 , n1269 );
not ( n1271 , n524 );
not ( n1272 , n43 );
and ( n1273 , n1271 , n1272 );
and ( n1274 , n524 , n43 );
nor ( n1275 , n1273 , n1274 );
or ( n1276 , n593 , n1275 );
not ( n1277 , n1142 );
or ( n1278 , n771 , n1277 );
nand ( n1279 , n1276 , n1278 );
not ( n1280 , n1279 );
nand ( n1281 , n1082 , n50 );
not ( n1282 , n1281 );
xor ( n1283 , n890 , n39 );
not ( n1284 , n1283 );
not ( n1285 , n1284 );
not ( n1286 , n997 );
or ( n1287 , n1285 , n1286 );
nand ( n1288 , n1104 , n1171 );
nand ( n1289 , n1287 , n1288 );
not ( n1290 , n1289 );
or ( n1291 , n1282 , n1290 );
or ( n1292 , n1289 , n1281 );
nand ( n1293 , n1291 , n1292 );
not ( n1294 , n1293 );
or ( n1295 , n1280 , n1294 );
not ( n1296 , n1281 );
nand ( n1297 , n1296 , n1289 );
nand ( n1298 , n1295 , n1297 );
nand ( n1299 , n1270 , n1298 );
not ( n1300 , n1299 );
xnor ( n1301 , n1267 , n1300 );
xnor ( n1302 , n1217 , n1228 );
and ( n1303 , n409 , n840 );
not ( n1304 , n409 );
and ( n1305 , n1304 , n45 );
nor ( n1306 , n1303 , n1305 );
not ( n1307 , n1306 );
not ( n1308 , n456 );
or ( n1309 , n1307 , n1308 );
nand ( n1310 , n501 , n1159 );
nand ( n1311 , n1309 , n1310 );
not ( n1312 , n1311 );
and ( n1313 , n861 , n41 );
not ( n1314 , n861 );
and ( n1315 , n1314 , n424 );
nor ( n1316 , n1313 , n1315 );
not ( n1317 , n1316 );
and ( n1318 , n742 , n1317 );
not ( n1319 , n1210 );
nor ( n1320 , n1319 , n854 );
nor ( n1321 , n1318 , n1320 );
not ( n1322 , n1321 );
or ( n1323 , n1312 , n1322 );
or ( n1324 , n1311 , n1321 );
nand ( n1325 , n1323 , n1324 );
and ( n1326 , n47 , n351 );
not ( n1327 , n47 );
and ( n1328 , n1327 , n380 );
nor ( n1329 , n1326 , n1328 );
or ( n1330 , n369 , n1329 );
or ( n1331 , n421 , n1199 );
nand ( n1332 , n1330 , n1331 );
and ( n1333 , n1325 , n1332 );
not ( n1334 , n1321 );
and ( n1335 , n1334 , n1311 );
nor ( n1336 , n1333 , n1335 );
xnor ( n1337 , n1302 , n1336 );
xnor ( n1338 , n1154 , n1163 );
or ( n1339 , n1337 , n1338 );
or ( n1340 , n1302 , n1336 );
nand ( n1341 , n1339 , n1340 );
or ( n1342 , n1301 , n1341 );
or ( n1343 , n1267 , n1300 );
nand ( n1344 , n1342 , n1343 );
not ( n1345 , n1344 );
or ( n1346 , n1266 , n1345 );
or ( n1347 , n1344 , n1265 );
nand ( n1348 , n1346 , n1347 );
xor ( n1349 , n1236 , n1248 );
and ( n1350 , n1348 , n1349 );
not ( n1351 , n1344 );
and ( n1352 , n1351 , n1265 );
nor ( n1353 , n1350 , n1352 );
not ( n1354 , n1353 );
or ( n1355 , n1264 , n1354 );
or ( n1356 , n1353 , n1263 );
nand ( n1357 , n1355 , n1356 );
not ( n1358 , n1357 );
not ( n1359 , n1298 );
nand ( n1360 , n1359 , n1269 );
and ( n1361 , n1360 , n1299 );
not ( n1362 , n325 );
not ( n1363 , n49 );
not ( n1364 , n1363 );
not ( n1365 , n299 );
or ( n1366 , n1364 , n1365 );
nand ( n1367 , n1366 , n1135 );
not ( n1368 , n1367 );
and ( n1369 , n1362 , n1368 );
and ( n1370 , n332 , n1222 );
nor ( n1371 , n1369 , n1370 );
xor ( n1372 , n36 , n1179 );
and ( n1373 , n3 , n17 );
not ( n1374 , n3 );
and ( n1375 , n1374 , n33 );
nor ( n1376 , n1373 , n1375 );
buf ( n1377 , n1376 );
not ( n1378 , n1377 );
buf ( n1379 , n1378 );
and ( n1380 , n1372 , n1379 );
nand ( n1381 , n883 , n1185 );
not ( n1382 , n1381 );
and ( n1383 , n1382 , n337 );
nor ( n1384 , n1380 , n1383 );
xor ( n1385 , n1371 , n1384 );
not ( n1386 , n1385 );
and ( n1387 , n40 , n1095 );
not ( n1388 , n40 );
and ( n1389 , n1388 , n992 );
nor ( n1390 , n1387 , n1389 );
not ( n1391 , n1390 );
or ( n1392 , n998 , n1391 );
buf ( n1393 , n1103 );
not ( n1394 , n1393 );
or ( n1395 , n1394 , n1283 );
nand ( n1396 , n1392 , n1395 );
not ( n1397 , n1396 );
nand ( n1398 , n300 , n51 );
not ( n1399 , n1398 );
not ( n1400 , n1185 );
nand ( n1401 , n1109 , n1400 );
not ( n1402 , n1401 );
not ( n1403 , n506 );
and ( n1404 , n1402 , n1403 );
and ( n1405 , n1187 , n337 );
nor ( n1406 , n1404 , n1405 );
nand ( n1407 , n1382 , n304 );
nand ( n1408 , n1406 , n1407 );
nand ( n1409 , n1399 , n1408 );
not ( n1410 , n1408 );
nand ( n1411 , n1410 , n1398 );
and ( n1412 , n1409 , n1411 );
not ( n1413 , n1412 );
or ( n1414 , n1397 , n1413 );
nand ( n1415 , n1414 , n1409 );
not ( n1416 , n1415 );
or ( n1417 , n1386 , n1416 );
or ( n1418 , n1371 , n1384 );
nand ( n1419 , n1417 , n1418 );
xor ( n1420 , n1361 , n1419 );
xor ( n1421 , n1293 , n1279 );
not ( n1422 , n1421 );
xor ( n1423 , n1332 , n1325 );
not ( n1424 , n44 );
not ( n1425 , n449 );
or ( n1426 , n1424 , n1425 );
nand ( n1427 , n590 , n968 );
nand ( n1428 , n1426 , n1427 );
not ( n1429 , n1428 );
not ( n1430 , n592 );
or ( n1431 , n1429 , n1430 );
not ( n1432 , n1275 );
nand ( n1433 , n1432 , n657 );
nand ( n1434 , n1431 , n1433 );
and ( n1435 , n409 , n46 );
not ( n1436 , n409 );
and ( n1437 , n1436 , n916 );
nor ( n1438 , n1435 , n1437 );
not ( n1439 , n1438 );
not ( n1440 , n1439 );
not ( n1441 , n456 );
or ( n1442 , n1440 , n1441 );
nand ( n1443 , n501 , n1306 );
nand ( n1444 , n1442 , n1443 );
xor ( n1445 , n1434 , n1444 );
and ( n1446 , n42 , n751 );
not ( n1447 , n42 );
and ( n1448 , n1447 , n747 );
nor ( n1449 , n1446 , n1448 );
not ( n1450 , n1449 );
not ( n1451 , n742 );
or ( n1452 , n1450 , n1451 );
or ( n1453 , n854 , n1316 );
nand ( n1454 , n1452 , n1453 );
and ( n1455 , n1445 , n1454 );
and ( n1456 , n1434 , n1444 );
nor ( n1457 , n1455 , n1456 );
not ( n1458 , n1457 );
and ( n1459 , n1423 , n1458 );
not ( n1460 , n1423 );
and ( n1461 , n1460 , n1457 );
nor ( n1462 , n1459 , n1461 );
not ( n1463 , n1462 );
or ( n1464 , n1422 , n1463 );
nand ( n1465 , n1423 , n1458 );
nand ( n1466 , n1464 , n1465 );
and ( n1467 , n1420 , n1466 );
and ( n1468 , n1361 , n1419 );
nor ( n1469 , n1467 , n1468 );
xor ( n1470 , n1241 , n1243 );
xor ( n1471 , n1470 , n1245 );
xnor ( n1472 , n1469 , n1471 );
xor ( n1473 , n1301 , n1341 );
or ( n1474 , n1472 , n1473 );
or ( n1475 , n1469 , n1471 );
nand ( n1476 , n1474 , n1475 );
not ( n1477 , n1476 );
xnor ( n1478 , n1348 , n1349 );
not ( n1479 , n1478 );
or ( n1480 , n1477 , n1479 );
or ( n1481 , n1478 , n1476 );
nand ( n1482 , n1480 , n1481 );
not ( n1483 , n1482 );
xor ( n1484 , n1472 , n1473 );
not ( n1485 , n1484 );
xor ( n1486 , n1420 , n1466 );
xor ( n1487 , n1337 , n1338 );
xor ( n1488 , n1486 , n1487 );
xnor ( n1489 , n1415 , n1385 );
not ( n1490 , n50 );
not ( n1491 , n1490 );
not ( n1492 , n299 );
or ( n1493 , n1491 , n1492 );
nand ( n1494 , n1493 , n1281 );
or ( n1495 , n325 , n1494 );
or ( n1496 , n1367 , n331 );
nand ( n1497 , n1495 , n1496 );
not ( n1498 , n1497 );
and ( n1499 , n48 , n312 );
not ( n1500 , n48 );
and ( n1501 , n1500 , n350 );
or ( n1502 , n1499 , n1501 );
not ( n1503 , n1502 );
not ( n1504 , n368 );
or ( n1505 , n1503 , n1504 );
not ( n1506 , n1329 );
nand ( n1507 , n1506 , n389 );
nand ( n1508 , n1505 , n1507 );
not ( n1509 , n1508 );
not ( n1510 , n1509 );
or ( n1511 , n1498 , n1510 );
not ( n1512 , n1497 );
nand ( n1513 , n1512 , n1508 );
nand ( n1514 , n1511 , n1513 );
nand ( n1515 , n332 , n51 );
and ( n1516 , n323 , n301 );
and ( n1517 , n1515 , n1516 );
not ( n1518 , n38 );
not ( n1519 , n1108 );
or ( n1520 , n1518 , n1519 );
or ( n1521 , n1108 , n38 );
nand ( n1522 , n1520 , n1521 );
not ( n1523 , n1522 );
not ( n1524 , n1379 );
or ( n1525 , n1523 , n1524 );
or ( n1526 , n1381 , n39 );
nand ( n1527 , n1525 , n1526 );
and ( n1528 , n1517 , n1527 );
and ( n1529 , n1514 , n1528 );
and ( n1530 , n1508 , n1497 );
nor ( n1531 , n1529 , n1530 );
xor ( n1532 , n1489 , n1531 );
not ( n1533 , n1532 );
and ( n1534 , n524 , n45 );
not ( n1535 , n524 );
and ( n1536 , n1535 , n840 );
nor ( n1537 , n1534 , n1536 );
or ( n1538 , n593 , n1537 );
not ( n1539 , n1428 );
or ( n1540 , n771 , n1539 );
nand ( n1541 , n1538 , n1540 );
not ( n1542 , n1393 );
not ( n1543 , n1390 );
or ( n1544 , n1542 , n1543 );
not ( n1545 , n890 );
not ( n1546 , n41 );
and ( n1547 , n1545 , n1546 );
buf ( n1548 , n992 );
and ( n1549 , n1548 , n41 );
nor ( n1550 , n1547 , n1549 );
not ( n1551 , n1550 );
not ( n1552 , n996 );
nand ( n1553 , n1551 , n1552 );
nand ( n1554 , n1544 , n1553 );
xor ( n1555 , n1541 , n1554 );
not ( n1556 , n47 );
not ( n1557 , n409 );
or ( n1558 , n1556 , n1557 );
or ( n1559 , n409 , n47 );
nand ( n1560 , n1558 , n1559 );
not ( n1561 , n1560 );
or ( n1562 , n503 , n1561 );
or ( n1563 , n563 , n1438 );
nand ( n1564 , n1562 , n1563 );
and ( n1565 , n1555 , n1564 );
and ( n1566 , n1541 , n1554 );
nor ( n1567 , n1565 , n1566 );
not ( n1568 , n747 );
not ( n1569 , n43 );
and ( n1570 , n1568 , n1569 );
and ( n1571 , n752 , n43 );
nor ( n1572 , n1570 , n1571 );
not ( n1573 , n1572 );
not ( n1574 , n1573 );
not ( n1575 , n742 );
or ( n1576 , n1574 , n1575 );
nand ( n1577 , n855 , n1449 );
nand ( n1578 , n1576 , n1577 );
and ( n1579 , n366 , n49 );
not ( n1580 , n366 );
and ( n1581 , n1580 , n1363 );
nor ( n1582 , n1579 , n1581 );
not ( n1583 , n1582 );
not ( n1584 , n1583 );
not ( n1585 , n368 );
or ( n1586 , n1584 , n1585 );
nand ( n1587 , n389 , n1502 );
nand ( n1588 , n1586 , n1587 );
xor ( n1589 , n1578 , n1588 );
and ( n1590 , n381 , n51 );
nor ( n1591 , n379 , n51 );
nor ( n1592 , n1590 , n1591 );
and ( n1593 , n326 , n1592 );
not ( n1594 , n1494 );
and ( n1595 , n332 , n1594 );
nor ( n1596 , n1593 , n1595 );
not ( n1597 , n1596 );
and ( n1598 , n1589 , n1597 );
and ( n1599 , n1578 , n1588 );
or ( n1600 , n1598 , n1599 );
not ( n1601 , n1600 );
xor ( n1602 , n1567 , n1601 );
xnor ( n1603 , n1412 , n1396 );
and ( n1604 , n1602 , n1603 );
and ( n1605 , n1567 , n1601 );
nor ( n1606 , n1604 , n1605 );
not ( n1607 , n1606 );
or ( n1608 , n1533 , n1607 );
or ( n1609 , n1489 , n1531 );
nand ( n1610 , n1608 , n1609 );
and ( n1611 , n1488 , n1610 );
and ( n1612 , n1486 , n1487 );
nor ( n1613 , n1611 , n1612 );
not ( n1614 , n1613 );
or ( n1615 , n1485 , n1614 );
or ( n1616 , n1613 , n1484 );
nand ( n1617 , n1615 , n1616 );
not ( n1618 , n1617 );
not ( n1619 , n356 );
not ( n1620 , n1619 );
not ( n1621 , n48 );
not ( n1622 , n1621 );
or ( n1623 , n1620 , n1622 );
not ( n1624 , n48 );
or ( n1625 , n1624 , n1619 );
nand ( n1626 , n1623 , n1625 );
and ( n1627 , n456 , n1626 );
and ( n1628 , n501 , n1560 );
nor ( n1629 , n1627 , n1628 );
not ( n1630 , n388 );
not ( n1631 , n1582 );
and ( n1632 , n1630 , n1631 );
and ( n1633 , n50 , n350 );
not ( n1634 , n50 );
and ( n1635 , n1634 , n312 );
nor ( n1636 , n1633 , n1635 );
and ( n1637 , n368 , n1636 );
nor ( n1638 , n1632 , n1637 );
xor ( n1639 , n1629 , n1638 );
not ( n1640 , n427 );
not ( n1641 , n1382 );
or ( n1642 , n1640 , n1641 );
not ( n1643 , n1401 );
and ( n1644 , n39 , n1643 );
not ( n1645 , n39 );
and ( n1646 , n1645 , n1187 );
nor ( n1647 , n1644 , n1646 );
nand ( n1648 , n1642 , n1647 );
not ( n1649 , n1648 );
and ( n1650 , n1639 , n1649 );
and ( n1651 , n1629 , n1638 );
or ( n1652 , n1650 , n1651 );
not ( n1653 , n1652 );
not ( n1654 , n1653 );
not ( n1655 , n1517 );
not ( n1656 , n1527 );
and ( n1657 , n1655 , n1656 );
nor ( n1658 , n1657 , n1528 );
not ( n1659 , n1658 );
not ( n1660 , n1515 );
not ( n1661 , n42 );
not ( n1662 , n889 );
or ( n1663 , n1661 , n1662 );
or ( n1664 , n992 , n42 );
nand ( n1665 , n1663 , n1664 );
not ( n1666 , n1665 );
not ( n1667 , n1552 );
or ( n1668 , n1666 , n1667 );
not ( n1669 , n1550 );
nand ( n1670 , n1669 , n1393 );
nand ( n1671 , n1668 , n1670 );
not ( n1672 , n1671 );
or ( n1673 , n1660 , n1672 );
or ( n1674 , n1515 , n1671 );
nand ( n1675 , n1673 , n1674 );
not ( n1676 , n46 );
not ( n1677 , n449 );
or ( n1678 , n1676 , n1677 );
or ( n1679 , n449 , n46 );
nand ( n1680 , n1678 , n1679 );
not ( n1681 , n1680 );
or ( n1682 , n593 , n1681 );
or ( n1683 , n771 , n1537 );
nand ( n1684 , n1682 , n1683 );
nand ( n1685 , n1675 , n1684 );
not ( n1686 , n1515 );
nand ( n1687 , n1686 , n1671 );
and ( n1688 , n1685 , n1687 );
not ( n1689 , n1688 );
or ( n1690 , n1659 , n1689 );
or ( n1691 , n1658 , n1688 );
nand ( n1692 , n1690 , n1691 );
not ( n1693 , n1692 );
or ( n1694 , n1654 , n1693 );
not ( n1695 , n1688 );
nand ( n1696 , n1695 , n1658 );
nand ( n1697 , n1694 , n1696 );
and ( n1698 , n1514 , n1528 );
not ( n1699 , n1514 );
not ( n1700 , n1528 );
and ( n1701 , n1699 , n1700 );
nor ( n1702 , n1698 , n1701 );
xor ( n1703 , n1434 , n1444 );
xor ( n1704 , n1703 , n1454 );
xor ( n1705 , n1702 , n1704 );
not ( n1706 , n1705 );
or ( n1707 , n1697 , n1706 );
or ( n1708 , n1702 , n1704 );
nand ( n1709 , n1707 , n1708 );
xnor ( n1710 , n1462 , n1421 );
xor ( n1711 , n1709 , n1710 );
xnor ( n1712 , n1606 , n1532 );
and ( n1713 , n1711 , n1712 );
and ( n1714 , n1709 , n1710 );
nor ( n1715 , n1713 , n1714 );
not ( n1716 , n1715 );
xnor ( n1717 , n1488 , n1610 );
not ( n1718 , n1717 );
or ( n1719 , n1716 , n1718 );
or ( n1720 , n1717 , n1715 );
nand ( n1721 , n1719 , n1720 );
not ( n1722 , n1721 );
xor ( n1723 , n1709 , n1710 );
xor ( n1724 , n1723 , n1712 );
not ( n1725 , n1724 );
and ( n1726 , n1697 , n1706 );
not ( n1727 , n1697 );
and ( n1728 , n1727 , n1705 );
nor ( n1729 , n1726 , n1728 );
xor ( n1730 , n1567 , n1601 );
xor ( n1731 , n1730 , n1603 );
and ( n1732 , n1729 , n1731 );
not ( n1733 , n1729 );
not ( n1734 , n1731 );
and ( n1735 , n1733 , n1734 );
nor ( n1736 , n1732 , n1735 );
xor ( n1737 , n1541 , n1554 );
xor ( n1738 , n1737 , n1564 );
xor ( n1739 , n1578 , n1588 );
not ( n1740 , n1596 );
xor ( n1741 , n1739 , n1740 );
xor ( n1742 , n1738 , n1741 );
not ( n1743 , n47 );
not ( n1744 , n524 );
or ( n1745 , n1743 , n1744 );
or ( n1746 , n524 , n47 );
nand ( n1747 , n1745 , n1746 );
not ( n1748 , n1747 );
not ( n1749 , n592 );
or ( n1750 , n1748 , n1749 );
nand ( n1751 , n657 , n1680 );
nand ( n1752 , n1750 , n1751 );
and ( n1753 , n409 , n1363 );
not ( n1754 , n409 );
and ( n1755 , n1754 , n49 );
nor ( n1756 , n1753 , n1755 );
not ( n1757 , n1756 );
not ( n1758 , n456 );
or ( n1759 , n1757 , n1758 );
nand ( n1760 , n501 , n1626 );
nand ( n1761 , n1759 , n1760 );
xor ( n1762 , n1752 , n1761 );
not ( n1763 , n424 );
not ( n1764 , n1382 );
or ( n1765 , n1763 , n1764 );
not ( n1766 , n427 );
not ( n1767 , n1179 );
or ( n1768 , n1766 , n1767 );
nand ( n1769 , n1108 , n40 );
nand ( n1770 , n1768 , n1769 );
not ( n1771 , n1770 );
or ( n1772 , n1771 , n1524 );
nand ( n1773 , n1765 , n1772 );
and ( n1774 , n1762 , n1773 );
and ( n1775 , n1761 , n1752 );
nor ( n1776 , n1774 , n1775 );
not ( n1777 , n1393 );
not ( n1778 , n1665 );
or ( n1779 , n1777 , n1778 );
not ( n1780 , n1552 );
not ( n1781 , n1096 );
not ( n1782 , n43 );
and ( n1783 , n1781 , n1782 );
and ( n1784 , n992 , n43 );
nor ( n1785 , n1783 , n1784 );
or ( n1786 , n1780 , n1785 );
nand ( n1787 , n1779 , n1786 );
not ( n1788 , n51 );
nor ( n1789 , n388 , n1788 );
nor ( n1790 , n1789 , n382 );
nand ( n1791 , n1787 , n1790 );
xor ( n1792 , n747 , n44 );
or ( n1793 , n864 , n1792 );
or ( n1794 , n854 , n1572 );
nand ( n1795 , n1793 , n1794 );
and ( n1796 , n1791 , n1795 );
not ( n1797 , n1791 );
not ( n1798 , n1795 );
and ( n1799 , n1797 , n1798 );
nor ( n1800 , n1796 , n1799 );
or ( n1801 , n1776 , n1800 );
or ( n1802 , n1791 , n1798 );
nand ( n1803 , n1801 , n1802 );
and ( n1804 , n1742 , n1803 );
and ( n1805 , n1738 , n1741 );
nor ( n1806 , n1804 , n1805 );
and ( n1807 , n1736 , n1806 );
and ( n1808 , n1729 , n1731 );
nor ( n1809 , n1807 , n1808 );
not ( n1810 , n1809 );
or ( n1811 , n1725 , n1810 );
or ( n1812 , n1809 , n1724 );
nand ( n1813 , n1811 , n1812 );
not ( n1814 , n1813 );
not ( n1815 , n1675 );
not ( n1816 , n1684 );
not ( n1817 , n1816 );
and ( n1818 , n1815 , n1817 );
and ( n1819 , n1675 , n1816 );
nor ( n1820 , n1818 , n1819 );
not ( n1821 , n1820 );
not ( n1822 , n1821 );
xor ( n1823 , n1629 , n1638 );
not ( n1824 , n1648 );
xor ( n1825 , n1823 , n1824 );
not ( n1826 , n1825 );
not ( n1827 , n1826 );
and ( n1828 , n1822 , n1827 );
or ( n1829 , n1787 , n1790 );
nand ( n1830 , n1829 , n1791 );
not ( n1831 , n1830 );
and ( n1832 , n45 , n752 );
not ( n1833 , n45 );
and ( n1834 , n1833 , n667 );
nor ( n1835 , n1832 , n1834 );
or ( n1836 , n1835 , n864 );
or ( n1837 , n854 , n1792 );
nand ( n1838 , n1836 , n1837 );
not ( n1839 , n389 );
not ( n1840 , n1636 );
or ( n1841 , n1839 , n1840 );
or ( n1842 , n369 , n1592 );
nand ( n1843 , n1841 , n1842 );
xnor ( n1844 , n1838 , n1843 );
not ( n1845 , n1844 );
and ( n1846 , n1831 , n1845 );
and ( n1847 , n1838 , n1843 );
nor ( n1848 , n1846 , n1847 );
and ( n1849 , n1826 , n1820 );
not ( n1850 , n1826 );
and ( n1851 , n1850 , n1821 );
or ( n1852 , n1849 , n1851 );
and ( n1853 , n1848 , n1852 );
nor ( n1854 , n1828 , n1853 );
xor ( n1855 , n1692 , n1653 );
xor ( n1856 , n1854 , n1855 );
xor ( n1857 , n1742 , n1803 );
and ( n1858 , n1856 , n1857 );
and ( n1859 , n1854 , n1855 );
nor ( n1860 , n1858 , n1859 );
not ( n1861 , n1860 );
not ( n1862 , n1806 );
and ( n1863 , n1736 , n1862 );
not ( n1864 , n1736 );
and ( n1865 , n1864 , n1806 );
nor ( n1866 , n1863 , n1865 );
not ( n1867 , n1866 );
or ( n1868 , n1861 , n1867 );
or ( n1869 , n1866 , n1860 );
nand ( n1870 , n1868 , n1869 );
not ( n1871 , n1870 );
not ( n1872 , n889 );
not ( n1873 , n44 );
and ( n1874 , n1872 , n1873 );
and ( n1875 , n1096 , n44 );
nor ( n1876 , n1874 , n1875 );
not ( n1877 , n1876 );
not ( n1878 , n1877 );
not ( n1879 , n1552 );
or ( n1880 , n1878 , n1879 );
not ( n1881 , n1785 );
nand ( n1882 , n1881 , n1103 );
nand ( n1883 , n1880 , n1882 );
xor ( n1884 , n1789 , n1883 );
not ( n1885 , n48 );
not ( n1886 , n1885 );
not ( n1887 , n590 );
or ( n1888 , n1886 , n1887 );
or ( n1889 , n1885 , n590 );
nand ( n1890 , n1888 , n1889 );
not ( n1891 , n1890 );
or ( n1892 , n593 , n1891 );
not ( n1893 , n1747 );
or ( n1894 , n771 , n1893 );
nand ( n1895 , n1892 , n1894 );
and ( n1896 , n1884 , n1895 );
and ( n1897 , n1789 , n1883 );
nor ( n1898 , n1896 , n1897 );
not ( n1899 , n42 );
not ( n1900 , n1899 );
not ( n1901 , n1382 );
or ( n1902 , n1900 , n1901 );
and ( n1903 , n41 , n1643 );
not ( n1904 , n41 );
and ( n1905 , n1904 , n1187 );
nor ( n1906 , n1903 , n1905 );
nand ( n1907 , n1902 , n1906 );
not ( n1908 , n1756 );
not ( n1909 , n501 );
or ( n1910 , n1908 , n1909 );
not ( n1911 , n1619 );
not ( n1912 , n50 );
and ( n1913 , n1911 , n1912 );
not ( n1914 , n409 );
and ( n1915 , n1914 , n50 );
nor ( n1916 , n1913 , n1915 );
nand ( n1917 , n456 , n1916 );
nand ( n1918 , n1910 , n1917 );
xor ( n1919 , n1907 , n1918 );
not ( n1920 , n916 );
not ( n1921 , n729 );
or ( n1922 , n1920 , n1921 );
nand ( n1923 , n861 , n46 );
nand ( n1924 , n1922 , n1923 );
not ( n1925 , n1924 );
not ( n1926 , n742 );
or ( n1927 , n1925 , n1926 );
or ( n1928 , n854 , n1835 );
nand ( n1929 , n1927 , n1928 );
nand ( n1930 , n1919 , n1929 );
nand ( n1931 , n1918 , n1907 );
and ( n1932 , n1930 , n1931 );
xor ( n1933 , n1898 , n1932 );
xnor ( n1934 , n1762 , n1773 );
and ( n1935 , n1933 , n1934 );
and ( n1936 , n1898 , n1932 );
nor ( n1937 , n1935 , n1936 );
xor ( n1938 , n1776 , n1800 );
xnor ( n1939 , n1937 , n1938 );
xnor ( n1940 , n1852 , n1848 );
or ( n1941 , n1939 , n1940 );
or ( n1942 , n1937 , n1938 );
nand ( n1943 , n1941 , n1942 );
not ( n1944 , n1943 );
xor ( n1945 , n1854 , n1855 );
xor ( n1946 , n1945 , n1857 );
not ( n1947 , n1946 );
or ( n1948 , n1944 , n1947 );
or ( n1949 , n1946 , n1943 );
nand ( n1950 , n1948 , n1949 );
not ( n1951 , n1950 );
nand ( n1952 , n657 , n51 );
nand ( n1953 , n1952 , n525 );
not ( n1954 , n44 );
not ( n1955 , n1108 );
or ( n1956 , n1954 , n1955 );
or ( n1957 , n1108 , n44 );
nand ( n1958 , n1956 , n1957 );
and ( n1959 , n1958 , n1379 );
and ( n1960 , n1382 , n840 );
nor ( n1961 , n1959 , n1960 );
or ( n1962 , n1953 , n1961 );
not ( n1963 , n1962 );
not ( n1964 , n1963 );
and ( n1965 , n1548 , n840 );
not ( n1966 , n1548 );
and ( n1967 , n1966 , n45 );
nor ( n1968 , n1965 , n1967 );
not ( n1969 , n1968 );
not ( n1970 , n1174 );
or ( n1971 , n1969 , n1970 );
not ( n1972 , n46 );
not ( n1973 , n992 );
or ( n1974 , n1972 , n1973 );
or ( n1975 , n889 , n46 );
nand ( n1976 , n1974 , n1975 );
nand ( n1977 , n997 , n1976 );
nand ( n1978 , n1971 , n1977 );
not ( n1979 , n1885 );
not ( n1980 , n515 );
or ( n1981 , n1979 , n1980 );
or ( n1982 , n667 , n1621 );
nand ( n1983 , n1981 , n1982 );
not ( n1984 , n1983 );
or ( n1985 , n1984 , n864 );
and ( n1986 , n47 , n747 );
not ( n1987 , n47 );
and ( n1988 , n1987 , n667 );
nor ( n1989 , n1986 , n1988 );
or ( n1990 , n854 , n1989 );
nand ( n1991 , n1985 , n1990 );
and ( n1992 , n1978 , n1991 );
not ( n1993 , n1978 );
not ( n1994 , n1991 );
and ( n1995 , n1993 , n1994 );
nor ( n1996 , n1992 , n1995 );
not ( n1997 , n1996 );
or ( n1998 , n1964 , n1997 );
nand ( n1999 , n1978 , n1991 );
nand ( n2000 , n1998 , n1999 );
not ( n2001 , n449 );
not ( n2002 , n49 );
and ( n2003 , n2001 , n2002 );
and ( n2004 , n767 , n49 );
nor ( n2005 , n2003 , n2004 );
not ( n2006 , n2005 );
not ( n2007 , n2006 );
not ( n2008 , n592 );
or ( n2009 , n2007 , n2008 );
nand ( n2010 , n657 , n1890 );
nand ( n2011 , n2009 , n2010 );
not ( n2012 , n2011 );
nand ( n2013 , n524 , n51 );
nand ( n2014 , n590 , n1788 );
and ( n2015 , n2013 , n2014 );
and ( n2016 , n2015 , n456 );
not ( n2017 , n1916 );
nor ( n2018 , n2017 , n500 );
nor ( n2019 , n2016 , n2018 );
not ( n2020 , n2019 );
or ( n2021 , n2012 , n2020 );
or ( n2022 , n2011 , n2019 );
nand ( n2023 , n2021 , n2022 );
xnor ( n2024 , n42 , n1108 );
not ( n2025 , n2024 );
or ( n2026 , n2025 , n1524 );
or ( n2027 , n1381 , n43 );
nand ( n2028 , n2026 , n2027 );
xor ( n2029 , n2023 , n2028 );
xor ( n2030 , n2000 , n2029 );
not ( n2031 , n771 );
not ( n2032 , n2005 );
and ( n2033 , n2031 , n2032 );
and ( n2034 , n595 , n50 );
and ( n2035 , n524 , n1490 );
nor ( n2036 , n2034 , n2035 );
and ( n2037 , n592 , n2036 );
nor ( n2038 , n2033 , n2037 );
not ( n2039 , n2038 );
nand ( n2040 , n501 , n51 );
not ( n2041 , n2040 );
nand ( n2042 , n1643 , n43 );
nand ( n2043 , n1187 , n825 );
nand ( n2044 , n1382 , n968 );
and ( n2045 , n2042 , n2043 , n2044 );
xnor ( n2046 , n2041 , n2045 );
nand ( n2047 , n2039 , n2046 );
not ( n2048 , n2045 );
nand ( n2049 , n2048 , n2041 );
and ( n2050 , n2047 , n2049 );
not ( n2051 , n1968 );
not ( n2052 , n997 );
or ( n2053 , n2051 , n2052 );
nand ( n2054 , n1174 , n1877 );
nand ( n2055 , n2053 , n2054 );
and ( n2056 , n2040 , n410 );
nor ( n2057 , n2055 , n2056 );
not ( n2058 , n2057 );
nand ( n2059 , n2055 , n2056 );
nand ( n2060 , n2058 , n2059 );
or ( n2061 , n864 , n1989 );
not ( n2062 , n1924 );
or ( n2063 , n854 , n2062 );
nand ( n2064 , n2061 , n2063 );
nor ( n2065 , n2060 , n2064 );
not ( n2066 , n2065 );
nand ( n2067 , n2060 , n2064 );
nand ( n2068 , n2066 , n2067 );
xnor ( n2069 , n2050 , n2068 );
and ( n2070 , n2030 , n2069 );
and ( n2071 , n2000 , n2029 );
nor ( n2072 , n2070 , n2071 );
not ( n2073 , n2072 );
not ( n2074 , n2028 );
not ( n2075 , n2023 );
or ( n2076 , n2074 , n2075 );
not ( n2077 , n2019 );
nand ( n2078 , n2077 , n2011 );
nand ( n2079 , n2076 , n2078 );
not ( n2080 , n2079 );
xor ( n2081 , n2080 , n2059 );
xor ( n2082 , n1789 , n1883 );
xor ( n2083 , n2082 , n1895 );
not ( n2084 , n2083 );
xor ( n2085 , n2081 , n2084 );
not ( n2086 , n2068 );
not ( n2087 , n2050 );
not ( n2088 , n2087 );
or ( n2089 , n2086 , n2088 );
not ( n2090 , n2060 );
nand ( n2091 , n2090 , n2064 );
nand ( n2092 , n2089 , n2091 );
not ( n2093 , n2092 );
not ( n2094 , n1919 );
not ( n2095 , n2094 );
not ( n2096 , n1929 );
and ( n2097 , n2095 , n2096 );
and ( n2098 , n2094 , n1929 );
nor ( n2099 , n2097 , n2098 );
not ( n2100 , n2099 );
and ( n2101 , n2093 , n2100 );
and ( n2102 , n2092 , n2099 );
nor ( n2103 , n2101 , n2102 );
xor ( n2104 , n2085 , n2103 );
not ( n2105 , n2104 );
or ( n2106 , n2073 , n2105 );
or ( n2107 , n2104 , n2072 );
nand ( n2108 , n2106 , n2107 );
not ( n2109 , n2108 );
and ( n2110 , n747 , n49 );
not ( n2111 , n747 );
and ( n2112 , n2111 , n1363 );
nor ( n2113 , n2110 , n2112 );
or ( n2114 , n864 , n2113 );
or ( n2115 , n854 , n1984 );
nand ( n2116 , n2114 , n2115 );
not ( n2117 , n2116 );
not ( n2118 , n1976 );
not ( n2119 , n1393 );
or ( n2120 , n2118 , n2119 );
not ( n2121 , n47 );
and ( n2122 , n1548 , n2121 );
not ( n2123 , n1548 );
and ( n2124 , n2123 , n47 );
nor ( n2125 , n2122 , n2124 );
nand ( n2126 , n1552 , n2125 );
nand ( n2127 , n2120 , n2126 );
not ( n2128 , n593 );
not ( n2129 , n2015 );
and ( n2130 , n2128 , n2129 );
and ( n2131 , n657 , n2036 );
nor ( n2132 , n2130 , n2131 );
xnor ( n2133 , n2127 , n2132 );
not ( n2134 , n2133 );
or ( n2135 , n2117 , n2134 );
not ( n2136 , n2132 );
nand ( n2137 , n2136 , n2127 );
nand ( n2138 , n2135 , n2137 );
not ( n2139 , n2046 );
not ( n2140 , n2038 );
and ( n2141 , n2139 , n2140 );
and ( n2142 , n2046 , n2038 );
nor ( n2143 , n2141 , n2142 );
xor ( n2144 , n2138 , n2143 );
not ( n2145 , n1963 );
xor ( n2146 , n1996 , n2145 );
or ( n2147 , n2144 , n2146 );
not ( n2148 , n2138 );
or ( n2149 , n2148 , n2143 );
nand ( n2150 , n2147 , n2149 );
not ( n2151 , n2069 );
and ( n2152 , n2030 , n2151 );
not ( n2153 , n2030 );
and ( n2154 , n2153 , n2069 );
nor ( n2155 , n2152 , n2154 );
xnor ( n2156 , n2150 , n2155 );
not ( n2157 , n2156 );
and ( n2158 , n2144 , n2146 );
not ( n2159 , n2144 );
not ( n2160 , n2146 );
and ( n2161 , n2159 , n2160 );
nor ( n2162 , n2158 , n2161 );
xor ( n2163 , n2133 , n2116 );
not ( n2164 , n2163 );
not ( n2165 , n1952 );
and ( n2166 , n1187 , n840 );
nor ( n2167 , n1401 , n840 );
nor ( n2168 , n2166 , n2167 );
nand ( n2169 , n1382 , n916 );
nand ( n2170 , n2168 , n2169 );
xor ( n2171 , n2165 , n2170 );
not ( n2172 , n2125 );
not ( n2173 , n1393 );
or ( n2174 , n2172 , n2173 );
not ( n2175 , n48 );
not ( n2176 , n889 );
or ( n2177 , n2175 , n2176 );
or ( n2178 , n992 , n48 );
nand ( n2179 , n2177 , n2178 );
nand ( n2180 , n1552 , n2179 );
nand ( n2181 , n2174 , n2180 );
and ( n2182 , n2171 , n2181 );
and ( n2183 , n2165 , n2170 );
nor ( n2184 , n2182 , n2183 );
not ( n2185 , n1961 );
not ( n2186 , n1953 );
or ( n2187 , n2185 , n2186 );
nand ( n2188 , n2187 , n1962 );
xor ( n2189 , n2184 , n2188 );
not ( n2190 , n2189 );
or ( n2191 , n2164 , n2190 );
or ( n2192 , n2184 , n2188 );
nand ( n2193 , n2191 , n2192 );
and ( n2194 , n2162 , n2193 );
not ( n2195 , n2162 );
not ( n2196 , n2193 );
and ( n2197 , n2195 , n2196 );
nor ( n2198 , n2194 , n2197 );
not ( n2199 , n2198 );
xor ( n2200 , n2163 , n2189 );
xnor ( n2201 , n2171 , n2181 );
nor ( n2202 , n853 , n1788 );
nor ( n2203 , n2202 , n681 );
not ( n2204 , n46 );
not ( n2205 , n1108 );
or ( n2206 , n2204 , n2205 );
or ( n2207 , n1108 , n46 );
nand ( n2208 , n2206 , n2207 );
not ( n2209 , n2208 );
or ( n2210 , n2209 , n1524 );
or ( n2211 , n1381 , n47 );
nand ( n2212 , n2210 , n2211 );
nand ( n2213 , n2203 , n2212 );
not ( n2214 , n854 );
not ( n2215 , n2113 );
and ( n2216 , n2214 , n2215 );
and ( n2217 , n747 , n1490 );
not ( n2218 , n747 );
and ( n2219 , n2218 , n50 );
nor ( n2220 , n2217 , n2219 );
buf ( n2221 , n2220 );
and ( n2222 , n742 , n2221 );
nor ( n2223 , n2216 , n2222 );
xor ( n2224 , n2213 , n2223 );
and ( n2225 , n2201 , n2224 );
and ( n2226 , n2213 , n2223 );
nor ( n2227 , n2225 , n2226 );
and ( n2228 , n2200 , n2227 );
not ( n2229 , n2200 );
not ( n2230 , n2227 );
and ( n2231 , n2229 , n2230 );
nor ( n2232 , n2228 , n2231 );
not ( n2233 , n2232 );
or ( n2234 , n2203 , n2212 );
nand ( n2235 , n2234 , n2213 );
xor ( n2236 , n49 , n992 );
not ( n2237 , n2236 );
not ( n2238 , n2237 );
not ( n2239 , n997 );
or ( n2240 , n2238 , n2239 );
nand ( n2241 , n2179 , n1103 );
nand ( n2242 , n2240 , n2241 );
not ( n2243 , n51 );
nand ( n2244 , n2243 , n679 );
nand ( n2245 , n890 , n51 );
and ( n2246 , n2244 , n2245 );
and ( n2247 , n2246 , n742 );
not ( n2248 , n2221 );
nor ( n2249 , n2248 , n853 );
nor ( n2250 , n2247 , n2249 );
xnor ( n2251 , n2242 , n2250 );
and ( n2252 , n2235 , n2251 );
not ( n2253 , n2235 );
xor ( n2254 , n2242 , n2250 );
and ( n2255 , n2253 , n2254 );
or ( n2256 , n2252 , n2255 );
not ( n2257 , n2202 );
not ( n2258 , n996 );
not ( n2259 , n679 );
not ( n2260 , n50 );
and ( n2261 , n2259 , n2260 );
and ( n2262 , n679 , n50 );
nor ( n2263 , n2261 , n2262 );
not ( n2264 , n2263 );
not ( n2265 , n2264 );
and ( n2266 , n2258 , n2265 );
and ( n2267 , n1103 , n2237 );
nor ( n2268 , n2266 , n2267 );
not ( n2269 , n2268 );
or ( n2270 , n2257 , n2269 );
or ( n2271 , n2268 , n2202 );
nand ( n2272 , n2270 , n2271 );
not ( n2273 , n2272 );
and ( n2274 , n47 , n1643 );
not ( n2275 , n47 );
and ( n2276 , n2275 , n1187 );
nor ( n2277 , n2274 , n2276 );
nand ( n2278 , n1382 , n1621 );
and ( n2279 , n2277 , n2278 );
or ( n2280 , n2273 , n2279 );
not ( n2281 , n2268 );
nand ( n2282 , n2281 , n2202 );
nand ( n2283 , n2280 , n2282 );
and ( n2284 , n2256 , n2283 );
not ( n2285 , n2256 );
not ( n2286 , n2283 );
and ( n2287 , n2285 , n2286 );
nor ( n2288 , n2284 , n2287 );
not ( n2289 , n2288 );
not ( n2290 , n2279 );
not ( n2291 , n2290 );
not ( n2292 , n2273 );
or ( n2293 , n2291 , n2292 );
nand ( n2294 , n2272 , n2279 );
nand ( n2295 , n2293 , n2294 );
and ( n2296 , n1108 , n1621 );
not ( n2297 , n1108 );
and ( n2298 , n2297 , n48 );
nor ( n2299 , n2296 , n2298 );
not ( n2300 , n2299 );
or ( n2301 , n2300 , n1524 );
or ( n2302 , n1381 , n49 );
nand ( n2303 , n2301 , n2302 );
nand ( n2304 , n1103 , n51 );
and ( n2305 , n2304 , n891 );
and ( n2306 , n2303 , n2305 );
and ( n2307 , n2295 , n2306 );
not ( n2308 , n2295 );
not ( n2309 , n2306 );
and ( n2310 , n2308 , n2309 );
nor ( n2311 , n2307 , n2310 );
not ( n2312 , n2311 );
not ( n2313 , n2304 );
nor ( n2314 , n50 , n51 );
not ( n2315 , n2314 );
not ( n2316 , n1179 );
or ( n2317 , n2315 , n2316 );
or ( n2318 , n1381 , n51 );
nand ( n2319 , n2317 , n2318 );
nor ( n2320 , n2313 , n2319 );
not ( n2321 , n1363 );
not ( n2322 , n1179 );
or ( n2323 , n2321 , n2322 );
nand ( n2324 , n2323 , n1381 );
and ( n2325 , n1185 , n50 );
not ( n2326 , n2325 );
and ( n2327 , n2324 , n2326 );
and ( n2328 , n1643 , n49 );
nor ( n2329 , n2327 , n2328 );
nor ( n2330 , n2320 , n2329 );
not ( n2331 , n2330 );
not ( n2332 , n998 );
not ( n2333 , n2246 );
and ( n2334 , n2332 , n2333 );
not ( n2335 , n2264 );
and ( n2336 , n1104 , n2335 );
nor ( n2337 , n2334 , n2336 );
not ( n2338 , n2337 );
xor ( n2339 , n2303 , n2305 );
not ( n2340 , n2339 );
or ( n2341 , n2338 , n2340 );
or ( n2342 , n2337 , n2339 );
nand ( n2343 , n2341 , n2342 );
not ( n2344 , n2343 );
or ( n2345 , n2331 , n2344 );
not ( n2346 , n2337 );
nand ( n2347 , n2346 , n2339 );
nand ( n2348 , n2345 , n2347 );
not ( n2349 , n2348 );
or ( n2350 , n2312 , n2349 );
nand ( n2351 , n2295 , n2306 );
nand ( n2352 , n2350 , n2351 );
not ( n2353 , n2352 );
or ( n2354 , n2289 , n2353 );
nand ( n2355 , n2256 , n2283 );
nand ( n2356 , n2354 , n2355 );
not ( n2357 , n2356 );
xor ( n2358 , n2224 , n2201 );
not ( n2359 , n2358 );
or ( n2360 , n2254 , n2235 );
not ( n2361 , n2242 );
or ( n2362 , n2361 , n2250 );
nand ( n2363 , n2360 , n2362 );
not ( n2364 , n2363 );
and ( n2365 , n2359 , n2364 );
and ( n2366 , n2358 , n2363 );
nor ( n2367 , n2365 , n2366 );
not ( n2368 , n2367 );
and ( n2369 , n2357 , n2368 );
not ( n2370 , n2363 );
and ( n2371 , n2358 , n2370 );
nor ( n2372 , n2369 , n2371 );
not ( n2373 , n2372 );
or ( n2374 , n2233 , n2373 );
nand ( n2375 , n2200 , n2227 );
nand ( n2376 , n2374 , n2375 );
not ( n2377 , n2376 );
or ( n2378 , n2199 , n2377 );
nand ( n2379 , n2193 , n2162 );
nand ( n2380 , n2378 , n2379 );
not ( n2381 , n2380 );
or ( n2382 , n2157 , n2381 );
not ( n2383 , n2155 );
nand ( n2384 , n2383 , n2150 );
nand ( n2385 , n2382 , n2384 );
not ( n2386 , n2385 );
or ( n2387 , n2109 , n2386 );
not ( n2388 , n2072 );
nand ( n2389 , n2388 , n2104 );
nand ( n2390 , n2387 , n2389 );
or ( n2391 , n2103 , n2085 );
not ( n2392 , n2092 );
or ( n2393 , n2392 , n2099 );
nand ( n2394 , n2391 , n2393 );
not ( n2395 , n2394 );
xor ( n2396 , n1830 , n1844 );
xor ( n2397 , n2080 , n2059 );
and ( n2398 , n2397 , n2084 );
and ( n2399 , n2080 , n2059 );
nor ( n2400 , n2398 , n2399 );
xor ( n2401 , n2396 , n2400 );
xor ( n2402 , n1898 , n1932 );
xor ( n2403 , n2402 , n1934 );
not ( n2404 , n2403 );
xor ( n2405 , n2401 , n2404 );
not ( n2406 , n2405 );
nor ( n2407 , n2395 , n2406 );
or ( n2408 , n2390 , n2407 );
not ( n2409 , n2394 );
nand ( n2410 , n2409 , n2406 );
nand ( n2411 , n2408 , n2410 );
and ( n2412 , n1939 , n1940 );
not ( n2413 , n1939 );
not ( n2414 , n1940 );
and ( n2415 , n2413 , n2414 );
nor ( n2416 , n2412 , n2415 );
xor ( n2417 , n2396 , n2400 );
not ( n2418 , n2403 );
and ( n2419 , n2417 , n2418 );
and ( n2420 , n2396 , n2400 );
or ( n2421 , n2419 , n2420 );
not ( n2422 , n2421 );
xnor ( n2423 , n2416 , n2422 );
or ( n2424 , n2411 , n2423 );
or ( n2425 , n2416 , n2422 );
nand ( n2426 , n2424 , n2425 );
not ( n2427 , n2426 );
or ( n2428 , n1951 , n2427 );
not ( n2429 , n1943 );
nand ( n2430 , n2429 , n1946 );
nand ( n2431 , n2428 , n2430 );
not ( n2432 , n2431 );
or ( n2433 , n1871 , n2432 );
not ( n2434 , n1860 );
nand ( n2435 , n2434 , n1866 );
nand ( n2436 , n2433 , n2435 );
not ( n2437 , n2436 );
or ( n2438 , n1814 , n2437 );
not ( n2439 , n1724 );
nand ( n2440 , n2439 , n1809 );
nand ( n2441 , n2438 , n2440 );
not ( n2442 , n2441 );
or ( n2443 , n1722 , n2442 );
not ( n2444 , n1717 );
nand ( n2445 , n2444 , n1715 );
nand ( n2446 , n2443 , n2445 );
not ( n2447 , n2446 );
or ( n2448 , n1618 , n2447 );
not ( n2449 , n1613 );
nand ( n2450 , n2449 , n1484 );
nand ( n2451 , n2448 , n2450 );
not ( n2452 , n2451 );
or ( n2453 , n1483 , n2452 );
not ( n2454 , n1478 );
nand ( n2455 , n2454 , n1476 );
nand ( n2456 , n2453 , n2455 );
not ( n2457 , n2456 );
or ( n2458 , n1358 , n2457 );
not ( n2459 , n1353 );
nand ( n2460 , n2459 , n1263 );
nand ( n2461 , n2458 , n2460 );
not ( n2462 , n2461 );
or ( n2463 , n1262 , n2462 );
not ( n2464 , n1257 );
nand ( n2465 , n2464 , n1254 );
nand ( n2466 , n2463 , n2465 );
not ( n2467 , n2466 );
or ( n2468 , n1129 , n2467 );
not ( n2469 , n1032 );
nand ( n2470 , n2469 , n1124 );
nand ( n2471 , n2468 , n2470 );
not ( n2472 , n2471 );
or ( n2473 , n1031 , n2472 );
not ( n2474 , n823 );
nand ( n2475 , n2474 , n1026 );
nand ( n2476 , n2473 , n2475 );
not ( n2477 , n2476 );
or ( n2478 , n819 , n2477 );
not ( n2479 , n814 );
nand ( n2480 , n2479 , n812 );
nand ( n2481 , n2478 , n2480 );
not ( n2482 , n2481 );
or ( n2483 , n709 , n2482 );
not ( n2484 , n704 );
nand ( n2485 , n2484 , n617 );
nand ( n2486 , n2483 , n2485 );
not ( n2487 , n2486 );
or ( n2488 , n616 , n2487 );
not ( n2489 , n549 );
nand ( n2490 , n2489 , n611 );
nand ( n2491 , n2488 , n2490 );
not ( n2492 , n2491 );
or ( n2493 , n547 , n2492 );
not ( n2494 , n493 );
nand ( n2495 , n2494 , n542 );
nand ( n2496 , n2493 , n2495 );
not ( n2497 , n2496 );
or ( n2498 , n492 , n2497 );
not ( n2499 , n470 );
nand ( n2500 , n2499 , n486 );
nand ( n2501 , n2498 , n2500 );
not ( n2502 , n2501 );
or ( n2503 , n482 , n485 );
or ( n2504 , n481 , n385 );
nand ( n2505 , n2503 , n2504 );
not ( n2506 , n2505 );
and ( n2507 , n480 , n306 );
and ( n2508 , n477 , n382 );
nor ( n2509 , n2507 , n2508 );
not ( n2510 , n475 );
and ( n2511 , n328 , n2510 );
and ( n2512 , n1516 , n319 );
nor ( n2513 , n2511 , n2512 );
xnor ( n2514 , n2513 , n338 );
xnor ( n2515 , n2509 , n2514 );
not ( n2516 , n2515 );
and ( n2517 , n2506 , n2516 );
and ( n2518 , n2505 , n2515 );
nor ( n2519 , n2517 , n2518 );
not ( n2520 , n2519 );
and ( n2521 , n2502 , n2520 );
and ( n2522 , n2501 , n2519 );
nor ( n2523 , n2521 , n2522 );
and ( n2524 , n3 , n1 );
not ( n2525 , n3 );
not ( n2526 , n1 );
and ( n2527 , n2525 , n2526 );
nor ( n2528 , n2524 , n2527 );
xor ( n2529 , n2528 , n2 );
buf ( n2530 , n2529 );
buf ( n2531 , n2530 );
or ( n2532 , n2523 , n2531 );
nand ( n2533 , n41 , n42 );
not ( n2534 , n2533 );
not ( n2535 , n427 );
or ( n2536 , n2534 , n2535 );
or ( n2537 , n41 , n42 );
nand ( n2538 , n2537 , n40 );
nand ( n2539 , n2536 , n2538 );
buf ( n2540 , n2539 );
not ( n2541 , n2540 );
not ( n2542 , n2541 );
not ( n2543 , n1210 );
or ( n2544 , n2542 , n2543 );
not ( n2545 , n41 );
not ( n2546 , n42 );
and ( n2547 , n2545 , n2546 );
and ( n2548 , n41 , n42 );
nor ( n2549 , n2547 , n2548 );
buf ( n2550 , n2549 );
not ( n2551 , n2550 );
not ( n2552 , n521 );
not ( n2553 , n427 );
and ( n2554 , n2552 , n2553 );
buf ( n2555 , n521 );
and ( n2556 , n2555 , n427 );
nor ( n2557 , n2554 , n2556 );
or ( n2558 , n2551 , n2557 );
nand ( n2559 , n2544 , n2558 );
not ( n2560 , n2559 );
xnor ( n2561 , n39 , n38 );
xor ( n2562 , n39 , n40 );
nor ( n2563 , n2561 , n2562 );
buf ( n2564 , n2563 );
not ( n2565 , n2564 );
not ( n2566 , n1171 );
or ( n2567 , n2565 , n2566 );
not ( n2568 , n38 );
not ( n2569 , n756 );
or ( n2570 , n2568 , n2569 );
or ( n2571 , n756 , n38 );
nand ( n2572 , n2570 , n2571 );
buf ( n2573 , n2562 );
nand ( n2574 , n2572 , n2573 );
nand ( n2575 , n2567 , n2574 );
nor ( n2576 , n45 , n46 );
nand ( n2577 , n2576 , n44 );
not ( n2578 , n44 );
nand ( n2579 , n2578 , n45 , n46 );
nand ( n2580 , n2577 , n2579 );
buf ( n2581 , n2580 );
not ( n2582 , n2581 );
not ( n2583 , n1159 );
or ( n2584 , n2582 , n2583 );
xor ( n2585 , n45 , n46 );
not ( n2586 , n2585 );
not ( n2587 , n2586 );
not ( n2588 , n44 );
not ( n2589 , n360 );
or ( n2590 , n2588 , n2589 );
and ( n2591 , n3 , n7 );
not ( n2592 , n3 );
and ( n2593 , n2592 , n23 );
nor ( n2594 , n2591 , n2593 );
buf ( n2595 , n2594 );
or ( n2596 , n44 , n2595 );
nand ( n2597 , n2590 , n2596 );
nand ( n2598 , n2587 , n2597 );
nand ( n2599 , n2584 , n2598 );
xor ( n2600 , n2575 , n2599 );
not ( n2601 , n2600 );
not ( n2602 , n2601 );
or ( n2603 , n2560 , n2602 );
not ( n2604 , n2559 );
nand ( n2605 , n2604 , n2600 );
nand ( n2606 , n2603 , n2605 );
not ( n2607 , n1171 );
not ( n2608 , n2573 );
or ( n2609 , n2607 , n2608 );
xor ( n2610 , n38 , n878 );
nand ( n2611 , n2610 , n2564 );
nand ( n2612 , n2609 , n2611 );
not ( n2613 , n2612 );
not ( n2614 , n2613 );
not ( n2615 , n40 );
not ( n2616 , n756 );
or ( n2617 , n2615 , n2616 );
or ( n2618 , n756 , n40 );
nand ( n2619 , n2617 , n2618 );
not ( n2620 , n2619 );
not ( n2621 , n2620 );
not ( n2622 , n2540 );
and ( n2623 , n2621 , n2622 );
and ( n2624 , n1210 , n2550 );
nor ( n2625 , n2623 , n2624 );
not ( n2626 , n2625 );
not ( n2627 , n2626 );
or ( n2628 , n2614 , n2627 );
nand ( n2629 , n2612 , n2625 );
nand ( n2630 , n2628 , n2629 );
buf ( n2631 , n2585 );
buf ( n2632 , n2631 );
not ( n2633 , n2632 );
not ( n2634 , n2633 );
not ( n2635 , n1160 );
and ( n2636 , n2634 , n2635 );
and ( n2637 , n3 , n9 );
not ( n2638 , n3 );
and ( n2639 , n2638 , n25 );
or ( n2640 , n2637 , n2639 );
not ( n2641 , n2640 );
and ( n2642 , n2641 , n968 );
not ( n2643 , n3 );
nand ( n2644 , n2643 , n25 );
nand ( n2645 , n2644 , n402 );
buf ( n2646 , n2645 );
and ( n2647 , n2646 , n44 );
nor ( n2648 , n2642 , n2647 );
and ( n2649 , n2648 , n2581 );
nor ( n2650 , n2636 , n2649 );
buf ( n2651 , n2650 );
and ( n2652 , n2630 , n2651 );
and ( n2653 , n2612 , n2626 );
nor ( n2654 , n2652 , n2653 );
xor ( n2655 , n2606 , n2654 );
and ( n2656 , n3 , n18 );
not ( n2657 , n3 );
and ( n2658 , n2657 , n34 );
nor ( n2659 , n2656 , n2658 );
buf ( n2660 , n2659 );
nor ( n2661 , n2660 , n374 );
buf ( n2662 , n2661 );
not ( n2663 , n2662 );
not ( n2664 , n1490 );
and ( n2665 , n2663 , n2664 );
and ( n2666 , n1377 , n374 );
nor ( n2667 , n1377 , n374 );
nor ( n2668 , n2666 , n2667 );
not ( n2669 , n2668 );
not ( n2670 , n2669 );
not ( n2671 , n37 );
not ( n2672 , n38 );
nand ( n2673 , n2671 , n2672 );
nand ( n2674 , n37 , n38 );
nand ( n2675 , n2673 , n2674 );
xor ( n2676 , n36 , n37 );
nand ( n2677 , n2675 , n2676 );
buf ( n2678 , n2677 );
not ( n2679 , n2678 );
and ( n2680 , n2670 , n2679 );
xor ( n2681 , n37 , n38 );
buf ( n2682 , n2681 );
and ( n2683 , n2682 , n1372 );
nor ( n2684 , n2680 , n2683 );
and ( n2685 , n2662 , n1490 );
not ( n2686 , n2662 );
and ( n2687 , n2686 , n50 );
nor ( n2688 , n2685 , n2687 );
and ( n2689 , n2684 , n2688 );
nor ( n2690 , n2665 , n2689 );
not ( n2691 , n2690 );
not ( n2692 , n48 );
not ( n2693 , n47 );
nor ( n2694 , n2693 , n46 );
not ( n2695 , n2694 );
or ( n2696 , n2692 , n2695 );
nand ( n2697 , n2121 , n1624 , n46 );
nand ( n2698 , n2696 , n2697 );
buf ( n2699 , n2698 );
not ( n2700 , n2699 );
not ( n2701 , n2595 );
and ( n2702 , n2701 , n916 );
and ( n2703 , n2595 , n46 );
nor ( n2704 , n2702 , n2703 );
or ( n2705 , n2700 , n2704 );
and ( n2706 , n48 , n47 );
not ( n2707 , n48 );
and ( n2708 , n2707 , n2121 );
or ( n2709 , n2706 , n2708 );
or ( n2710 , n1199 , n2709 );
nand ( n2711 , n2705 , n2710 );
not ( n2712 , n2711 );
xor ( n2713 , n43 , n44 );
not ( n2714 , n2713 );
not ( n2715 , n2714 );
not ( n2716 , n2715 );
not ( n2717 , n1142 );
or ( n2718 , n2716 , n2717 );
nand ( n2719 , n968 , n825 , n42 );
nand ( n2720 , n1899 , n43 , n44 );
nand ( n2721 , n2719 , n2720 );
buf ( n2722 , n2721 );
xor ( n2723 , n42 , n2555 );
nand ( n2724 , n2722 , n2723 );
nand ( n2725 , n2718 , n2724 );
not ( n2726 , n2725 );
not ( n2727 , n49 );
not ( n2728 , n50 );
and ( n2729 , n2727 , n2728 );
and ( n2730 , n49 , n50 );
nor ( n2731 , n2729 , n2730 );
buf ( n2732 , n2731 );
buf ( n2733 , n2732 );
not ( n2734 , n2733 );
not ( n2735 , n2734 );
not ( n2736 , n1220 );
and ( n2737 , n2735 , n2736 );
not ( n2738 , n1363 );
not ( n2739 , n48 );
nor ( n2740 , n2739 , n50 );
not ( n2741 , n2740 );
or ( n2742 , n2738 , n2741 );
not ( n2743 , n48 );
nand ( n2744 , n2743 , n49 , n50 );
nand ( n2745 , n2742 , n2744 );
not ( n2746 , n2745 );
not ( n2747 , n2746 );
buf ( n2748 , n2747 );
and ( n2749 , n48 , n318 );
not ( n2750 , n48 );
and ( n2751 , n2750 , n322 );
or ( n2752 , n2749 , n2751 );
and ( n2753 , n2748 , n2752 );
nor ( n2754 , n2737 , n2753 );
not ( n2755 , n2754 );
or ( n2756 , n2726 , n2755 );
or ( n2757 , n2725 , n2754 );
nand ( n2758 , n2756 , n2757 );
not ( n2759 , n2758 );
or ( n2760 , n2712 , n2759 );
not ( n2761 , n2754 );
nand ( n2762 , n2761 , n2725 );
nand ( n2763 , n2760 , n2762 );
not ( n2764 , n2763 );
not ( n2765 , n2764 );
or ( n2766 , n2691 , n2765 );
not ( n2767 , n2690 );
nand ( n2768 , n2767 , n2763 );
nand ( n2769 , n2766 , n2768 );
xor ( n2770 , n2655 , n2769 );
xnor ( n2771 , n2684 , n2688 );
xor ( n2772 , n2758 , n2711 );
xor ( n2773 , n2771 , n2772 );
and ( n2774 , n2674 , n36 );
not ( n2775 , n2774 );
not ( n2776 , n2681 );
and ( n2777 , n3 , n19 );
not ( n2778 , n3 );
and ( n2779 , n2778 , n35 );
nor ( n2780 , n2777 , n2779 );
not ( n2781 , n2780 );
not ( n2782 , n2781 );
nor ( n2783 , n2776 , n2782 );
nor ( n2784 , n2775 , n2783 );
or ( n2785 , n1494 , n1788 );
and ( n2786 , n3 , n5 );
not ( n2787 , n3 );
and ( n2788 , n2787 , n21 );
nor ( n2789 , n2786 , n2788 );
not ( n2790 , n2789 );
not ( n2791 , n2790 );
not ( n2792 , n51 );
nand ( n2793 , n2792 , n50 );
not ( n2794 , n2793 );
buf ( n2795 , n2794 );
nand ( n2796 , n2791 , n2795 );
nand ( n2797 , n2785 , n2796 );
nand ( n2798 , n2784 , n2797 );
buf ( n2799 , n2798 );
not ( n2800 , n2581 );
not ( n2801 , n44 );
not ( n2802 , n587 );
or ( n2803 , n2801 , n2802 );
or ( n2804 , n587 , n44 );
nand ( n2805 , n2803 , n2804 );
not ( n2806 , n2805 );
or ( n2807 , n2800 , n2806 );
nand ( n2808 , n2587 , n1428 );
nand ( n2809 , n2807 , n2808 );
not ( n2810 , n2661 );
nand ( n2811 , n2660 , n374 );
nand ( n2812 , n2810 , n2811 );
not ( n2813 , n2675 );
not ( n2814 , n2813 );
or ( n2815 , n2812 , n2814 );
nand ( n2816 , n2781 , n36 );
nand ( n2817 , n2782 , n374 );
not ( n2818 , n2677 );
nand ( n2819 , n2816 , n2817 , n2818 );
nand ( n2820 , n2815 , n2819 );
xor ( n2821 , n2809 , n2820 );
not ( n2822 , n1502 );
xor ( n2823 , n49 , n50 );
buf ( n2824 , n2823 );
not ( n2825 , n2824 );
or ( n2826 , n2822 , n2825 );
and ( n2827 , n48 , n2595 );
not ( n2828 , n48 );
and ( n2829 , n2828 , n2701 );
or ( n2830 , n2827 , n2829 );
nand ( n2831 , n2748 , n2830 );
nand ( n2832 , n2826 , n2831 );
and ( n2833 , n2821 , n2832 );
and ( n2834 , n2809 , n2820 );
nor ( n2835 , n2833 , n2834 );
xor ( n2836 , n2799 , n2835 );
not ( n2837 , n42 );
not ( n2838 , n756 );
or ( n2839 , n2837 , n2838 );
or ( n2840 , n756 , n42 );
nand ( n2841 , n2839 , n2840 );
not ( n2842 , n2841 );
not ( n2843 , n2722 );
or ( n2844 , n2842 , n2843 );
not ( n2845 , n2714 );
nand ( n2846 , n2845 , n1449 );
nand ( n2847 , n2844 , n2846 );
not ( n2848 , n2847 );
not ( n2849 , n2540 );
not ( n2850 , n981 );
not ( n2851 , n40 );
or ( n2852 , n2850 , n2851 );
buf ( n2853 , n981 );
or ( n2854 , n2853 , n40 );
nand ( n2855 , n2852 , n2854 );
nand ( n2856 , n2849 , n2855 );
nand ( n2857 , n1390 , n2550 );
and ( n2858 , n2856 , n2857 );
not ( n2859 , n2858 );
or ( n2860 , n2848 , n2859 );
or ( n2861 , n2847 , n2858 );
nand ( n2862 , n2860 , n2861 );
and ( n2863 , n2640 , n46 );
not ( n2864 , n2640 );
and ( n2865 , n2864 , n916 );
nor ( n2866 , n2863 , n2865 );
not ( n2867 , n2866 );
not ( n2868 , n2698 );
not ( n2869 , n2868 );
buf ( n2870 , n2869 );
not ( n2871 , n2870 );
or ( n2872 , n2867 , n2871 );
or ( n2873 , n1438 , n2709 );
nand ( n2874 , n2872 , n2873 );
nand ( n2875 , n2862 , n2874 );
not ( n2876 , n2858 );
nand ( n2877 , n2876 , n2847 );
and ( n2878 , n2875 , n2877 );
and ( n2879 , n2836 , n2878 );
and ( n2880 , n2799 , n2835 );
nor ( n2881 , n2879 , n2880 );
and ( n2882 , n2773 , n2881 );
and ( n2883 , n2771 , n2772 );
nor ( n2884 , n2882 , n2883 );
buf ( n2885 , n2884 );
or ( n2886 , n2770 , n2885 );
not ( n2887 , n2606 );
not ( n2888 , n2769 );
or ( n2889 , n2887 , n2888 );
or ( n2890 , n2769 , n2606 );
nand ( n2891 , n2889 , n2890 );
buf ( n2892 , n2654 );
or ( n2893 , n2891 , n2892 );
nand ( n2894 , n2886 , n2893 );
not ( n2895 , n2682 );
and ( n2896 , n2853 , n374 );
nor ( n2897 , n2853 , n374 );
nor ( n2898 , n2896 , n2897 );
not ( n2899 , n2898 );
or ( n2900 , n2895 , n2899 );
not ( n2901 , n2677 );
nand ( n2902 , n1523 , n2901 );
nand ( n2903 , n2900 , n2902 );
not ( n2904 , n1221 );
buf ( n2905 , n2745 );
not ( n2906 , n2905 );
or ( n2907 , n2904 , n2906 );
nand ( n2908 , n2823 , n48 );
buf ( n2909 , n2908 );
nand ( n2910 , n2907 , n2909 );
and ( n2911 , n2903 , n2910 );
not ( n2912 , n2903 );
not ( n2913 , n2910 );
and ( n2914 , n2912 , n2913 );
nor ( n2915 , n2911 , n2914 );
not ( n2916 , n2915 );
not ( n2917 , n2916 );
not ( n2918 , n2651 );
not ( n2919 , n2918 );
or ( n2920 , n2917 , n2919 );
nand ( n2921 , n2903 , n2913 );
nand ( n2922 , n2920 , n2921 );
not ( n2923 , n2564 );
not ( n2924 , n2572 );
or ( n2925 , n2923 , n2924 );
not ( n2926 , n2573 );
not ( n2927 , n2926 );
nand ( n2928 , n952 , n2927 );
nand ( n2929 , n2925 , n2928 );
not ( n2930 , n2929 );
not ( n2931 , n2913 );
or ( n2932 , n2930 , n2931 );
or ( n2933 , n2929 , n2913 );
nand ( n2934 , n2932 , n2933 );
not ( n2935 , n2818 );
not ( n2936 , n2898 );
or ( n2937 , n2935 , n2936 );
or ( n2938 , n1003 , n2814 );
nand ( n2939 , n2937 , n2938 );
and ( n2940 , n2934 , n2939 );
not ( n2941 , n2934 );
not ( n2942 , n2939 );
and ( n2943 , n2941 , n2942 );
nor ( n2944 , n2940 , n2943 );
xor ( n2945 , n2922 , n2944 );
and ( n2946 , n36 , n1179 );
not ( n2947 , n2550 );
not ( n2948 , n933 );
or ( n2949 , n2947 , n2948 );
not ( n2950 , n2557 );
not ( n2951 , n2540 );
nand ( n2952 , n2950 , n2951 );
nand ( n2953 , n2949 , n2952 );
xor ( n2954 , n2946 , n2953 );
not ( n2955 , n2581 );
not ( n2956 , n2597 );
or ( n2957 , n2955 , n2956 );
or ( n2958 , n2633 , n971 );
nand ( n2959 , n2957 , n2958 );
xor ( n2960 , n2954 , n2959 );
xor ( n2961 , n2945 , n2960 );
and ( n2962 , n2894 , n2961 );
not ( n2963 , n2894 );
not ( n2964 , n2961 );
and ( n2965 , n2963 , n2964 );
nor ( n2966 , n2962 , n2965 );
not ( n2967 , n2651 );
not ( n2968 , n2916 );
or ( n2969 , n2967 , n2968 );
nand ( n2970 , n2915 , n2918 );
nand ( n2971 , n2969 , n2970 );
or ( n2972 , n1377 , n374 );
not ( n2973 , n1200 );
not ( n2974 , n2699 );
or ( n2975 , n2973 , n2974 );
and ( n2976 , n2790 , n46 );
not ( n2977 , n2790 );
and ( n2978 , n2977 , n916 );
nor ( n2979 , n2976 , n2978 );
xor ( n2980 , n47 , n48 );
not ( n2981 , n2980 );
not ( n2982 , n2981 );
nand ( n2983 , n2979 , n2982 );
nand ( n2984 , n2975 , n2983 );
xor ( n2985 , n2972 , n2984 );
not ( n2986 , n2722 );
not ( n2987 , n2986 );
and ( n2988 , n1275 , n2987 );
not ( n2989 , n2640 );
not ( n2990 , n42 );
and ( n2991 , n2989 , n2990 );
and ( n2992 , n2646 , n42 );
nor ( n2993 , n2991 , n2992 );
and ( n2994 , n2993 , n2715 );
nor ( n2995 , n2988 , n2994 );
xor ( n2996 , n2985 , n2995 );
xnor ( n2997 , n2971 , n2996 );
not ( n2998 , n1539 );
not ( n2999 , n2955 );
and ( n3000 , n2998 , n2999 );
and ( n3001 , n2648 , n2632 );
nor ( n3002 , n3000 , n3001 );
not ( n3003 , n3002 );
not ( n3004 , n2722 );
not ( n3005 , n1449 );
or ( n3006 , n3004 , n3005 );
buf ( n3007 , n2713 );
nand ( n3008 , n2723 , n3007 );
nand ( n3009 , n3006 , n3008 );
not ( n3010 , n3009 );
not ( n3011 , n2814 );
not ( n3012 , n3011 );
not ( n3013 , n2668 );
or ( n3014 , n3012 , n3013 );
not ( n3015 , n2661 );
nand ( n3016 , n3015 , n2901 , n2811 );
nand ( n3017 , n3014 , n3016 );
not ( n3018 , n3017 );
not ( n3019 , n3018 );
or ( n3020 , n3010 , n3019 );
not ( n3021 , n3009 );
not ( n3022 , n3011 );
not ( n3023 , n2668 );
or ( n3024 , n3022 , n3023 );
nand ( n3025 , n3024 , n3016 );
nand ( n3026 , n3021 , n3025 );
nand ( n3027 , n3020 , n3026 );
nand ( n3028 , n3003 , n3027 );
not ( n3029 , n3018 );
nand ( n3030 , n3029 , n3009 );
nand ( n3031 , n3028 , n3030 );
not ( n3032 , n3031 );
not ( n3033 , n2704 );
not ( n3034 , n2709 );
and ( n3035 , n3033 , n3034 );
not ( n3036 , n1626 );
not ( n3037 , n2868 );
and ( n3038 , n3036 , n3037 );
nor ( n3039 , n3035 , n3038 );
not ( n3040 , n3039 );
not ( n3041 , n1390 );
not ( n3042 , n2539 );
buf ( n3043 , n3042 );
not ( n3044 , n3043 );
or ( n3045 , n3041 , n3044 );
nand ( n3046 , n2619 , n2550 );
nand ( n3047 , n3045 , n3046 );
not ( n3048 , n1522 );
not ( n3049 , n2564 );
or ( n3050 , n3048 , n3049 );
nand ( n3051 , n2610 , n2573 );
nand ( n3052 , n3050 , n3051 );
xor ( n3053 , n3047 , n3052 );
nand ( n3054 , n3040 , n3053 );
nand ( n3055 , n3047 , n3052 );
and ( n3056 , n3054 , n3055 );
not ( n3057 , n50 );
not ( n3058 , n299 );
or ( n3059 , n3057 , n3058 );
nand ( n3060 , n50 , n51 );
not ( n3061 , n3060 );
not ( n3062 , n3061 );
nand ( n3063 , n3059 , n3062 );
not ( n3064 , n3063 );
not ( n3065 , n3064 );
not ( n3066 , n2816 );
and ( n3067 , n3065 , n3066 );
not ( n3068 , n3063 );
not ( n3069 , n2816 );
and ( n3070 , n3068 , n3069 );
and ( n3071 , n2816 , n3063 );
nor ( n3072 , n3070 , n3071 );
not ( n3073 , n3072 );
not ( n3074 , n1502 );
not ( n3075 , n2747 );
or ( n3076 , n3074 , n3075 );
nand ( n3077 , n2752 , n2824 );
nand ( n3078 , n3076 , n3077 );
and ( n3079 , n3073 , n3078 );
nor ( n3080 , n3067 , n3079 );
and ( n3081 , n3056 , n3080 );
not ( n3082 , n3056 );
not ( n3083 , n3080 );
and ( n3084 , n3082 , n3083 );
nor ( n3085 , n3081 , n3084 );
not ( n3086 , n3085 );
or ( n3087 , n3032 , n3086 );
not ( n3088 , n3056 );
nand ( n3089 , n3088 , n3083 );
nand ( n3090 , n3087 , n3089 );
or ( n3091 , n2997 , n3090 );
or ( n3092 , n2971 , n2996 );
nand ( n3093 , n3091 , n3092 );
not ( n3094 , n2767 );
not ( n3095 , n2764 );
or ( n3096 , n3094 , n3095 );
not ( n3097 , n2606 );
nand ( n3098 , n3097 , n2769 );
nand ( n3099 , n3096 , n3098 );
not ( n3100 , n2993 );
not ( n3101 , n2722 );
or ( n3102 , n3100 , n3101 );
nand ( n3103 , n961 , n2715 );
nand ( n3104 , n3102 , n3103 );
not ( n3105 , n48 );
not ( n3106 , n1363 );
or ( n3107 , n3105 , n3106 );
nand ( n3108 , n3107 , n2908 );
not ( n3109 , n3108 );
and ( n3110 , n3104 , n3109 );
not ( n3111 , n3104 );
and ( n3112 , n3111 , n3108 );
nor ( n3113 , n3110 , n3112 );
not ( n3114 , n2979 );
or ( n3115 , n2700 , n3114 );
or ( n3116 , n921 , n2709 );
nand ( n3117 , n3115 , n3116 );
xnor ( n3118 , n3113 , n3117 );
not ( n3119 , n3118 );
not ( n3120 , n2600 );
not ( n3121 , n2559 );
or ( n3122 , n3120 , n3121 );
nand ( n3123 , n2575 , n2599 );
nand ( n3124 , n3122 , n3123 );
not ( n3125 , n3124 );
not ( n3126 , n3125 );
not ( n3127 , n2995 );
not ( n3128 , n2667 );
not ( n3129 , n3128 );
not ( n3130 , n2984 );
or ( n3131 , n3129 , n3130 );
or ( n3132 , n2984 , n3128 );
nand ( n3133 , n3131 , n3132 );
not ( n3134 , n3133 );
or ( n3135 , n3127 , n3134 );
not ( n3136 , n2984 );
nand ( n3137 , n3136 , n3128 );
nand ( n3138 , n3135 , n3137 );
not ( n3139 , n3138 );
not ( n3140 , n3139 );
or ( n3141 , n3126 , n3140 );
nand ( n3142 , n3138 , n3124 );
nand ( n3143 , n3141 , n3142 );
not ( n3144 , n3143 );
or ( n3145 , n3119 , n3144 );
or ( n3146 , n3143 , n3118 );
nand ( n3147 , n3145 , n3146 );
xor ( n3148 , n3099 , n3147 );
xor ( n3149 , n3093 , n3148 );
xnor ( n3150 , n2966 , n3149 );
not ( n3151 , n3150 );
xnor ( n3152 , n2770 , n2885 );
not ( n3153 , n3152 );
not ( n3154 , n3153 );
xnor ( n3155 , n3090 , n2997 );
not ( n3156 , n3155 );
buf ( n3157 , n3002 );
not ( n3158 , n3157 );
buf ( n3159 , n3027 );
not ( n3160 , n3159 );
or ( n3161 , n3158 , n3160 );
or ( n3162 , n3159 , n3157 );
nand ( n3163 , n3161 , n3162 );
not ( n3164 , n3163 );
and ( n3165 , n3078 , n3072 );
not ( n3166 , n3078 );
and ( n3167 , n3166 , n3073 );
or ( n3168 , n3165 , n3167 );
not ( n3169 , n3168 );
and ( n3170 , n3164 , n3169 );
xor ( n3171 , n3002 , n3168 );
xnor ( n3172 , n3171 , n3159 );
not ( n3173 , n3053 );
not ( n3174 , n3039 );
and ( n3175 , n3173 , n3174 );
and ( n3176 , n3053 , n3039 );
nor ( n3177 , n3175 , n3176 );
and ( n3178 , n3172 , n3177 );
nor ( n3179 , n3170 , n3178 );
not ( n3180 , n3179 );
and ( n3181 , n2630 , n2918 );
not ( n3182 , n2630 );
and ( n3183 , n3182 , n2651 );
or ( n3184 , n3181 , n3183 );
xor ( n3185 , n3031 , n3184 );
xor ( n3186 , n3185 , n3085 );
not ( n3187 , n3186 );
or ( n3188 , n3180 , n3187 );
and ( n3189 , n2630 , n2918 );
not ( n3190 , n2630 );
and ( n3191 , n3190 , n2651 );
or ( n3192 , n3189 , n3191 );
xor ( n3193 , n3085 , n3031 );
nand ( n3194 , n3192 , n3193 );
nand ( n3195 , n3188 , n3194 );
not ( n3196 , n3195 );
not ( n3197 , n3196 );
or ( n3198 , n3156 , n3197 );
not ( n3199 , n3155 );
nand ( n3200 , n3199 , n3195 );
nand ( n3201 , n3198 , n3200 );
not ( n3202 , n3201 );
or ( n3203 , n3154 , n3202 );
nand ( n3204 , n3195 , n3155 );
nand ( n3205 , n3203 , n3204 );
not ( n3206 , n3205 );
not ( n3207 , n3206 );
or ( n3208 , n3151 , n3207 );
not ( n3209 , n752 );
not ( n3210 , n2795 );
not ( n3211 , n3210 );
not ( n3212 , n3211 );
or ( n3213 , n3209 , n3212 );
not ( n3214 , n50 );
nand ( n3215 , n3214 , n51 );
not ( n3216 , n3215 );
and ( n3217 , n2555 , n3216 );
not ( n3218 , n3062 );
and ( n3219 , n587 , n3218 );
nor ( n3220 , n3217 , n3219 );
nand ( n3221 , n3213 , n3220 );
not ( n3222 , n3221 );
nor ( n3223 , n2782 , n2714 );
not ( n3224 , n3223 );
and ( n3225 , n3 , n17 );
not ( n3226 , n3 );
and ( n3227 , n3226 , n33 );
or ( n3228 , n3225 , n3227 );
not ( n3229 , n3228 );
not ( n3230 , n44 );
and ( n3231 , n3229 , n3230 );
and ( n3232 , n1378 , n44 );
nor ( n3233 , n3231 , n3232 );
not ( n3234 , n3233 );
not ( n3235 , n2632 );
or ( n3236 , n3234 , n3235 );
xnor ( n3237 , n44 , n2660 );
nand ( n3238 , n3237 , n2581 );
nand ( n3239 , n3236 , n3238 );
not ( n3240 , n3239 );
not ( n3241 , n3240 );
or ( n3242 , n3224 , n3241 );
not ( n3243 , n3223 );
nand ( n3244 , n3243 , n3239 );
nand ( n3245 , n3242 , n3244 );
not ( n3246 , n3245 );
or ( n3247 , n3222 , n3246 );
nand ( n3248 , n3239 , n3223 );
nand ( n3249 , n3247 , n3248 );
not ( n3250 , n3249 );
not ( n3251 , n3250 );
not ( n3252 , n878 );
not ( n3253 , n916 );
and ( n3254 , n3252 , n3253 );
and ( n3255 , n878 , n916 );
nor ( n3256 , n3254 , n3255 );
or ( n3257 , n2700 , n3256 );
not ( n3258 , n1976 );
or ( n3259 , n3258 , n2709 );
nand ( n3260 , n3257 , n3259 );
not ( n3261 , n3260 );
not ( n3262 , n2905 );
not ( n3263 , n1624 );
not ( n3264 , n675 );
or ( n3265 , n3263 , n3264 );
or ( n3266 , n675 , n1624 );
nand ( n3267 , n3265 , n3266 );
not ( n3268 , n3267 );
or ( n3269 , n3262 , n3268 );
nand ( n3270 , n2824 , n1983 );
nand ( n3271 , n3269 , n3270 );
nand ( n3272 , n43 , n44 );
and ( n3273 , n3272 , n42 );
not ( n3274 , n3273 );
nor ( n3275 , n3223 , n3274 );
nor ( n3276 , n3271 , n3275 );
not ( n3277 , n3276 );
nand ( n3278 , n3271 , n3275 );
nand ( n3279 , n3277 , n3278 );
not ( n3280 , n3279 );
or ( n3281 , n3261 , n3280 );
or ( n3282 , n3260 , n3279 );
nand ( n3283 , n3281 , n3282 );
not ( n3284 , n3283 );
or ( n3285 , n3251 , n3284 );
or ( n3286 , n3250 , n3283 );
nand ( n3287 , n3285 , n3286 );
not ( n3288 , n3287 );
and ( n3289 , n2036 , n51 );
and ( n3290 , n3211 , n587 );
nor ( n3291 , n3289 , n3290 );
not ( n3292 , n3007 );
and ( n3293 , n3 , n18 );
not ( n3294 , n3 );
and ( n3295 , n3294 , n34 );
nor ( n3296 , n3293 , n3295 );
not ( n3297 , n3296 );
xor ( n3298 , n42 , n3297 );
not ( n3299 , n3298 );
or ( n3300 , n3292 , n3299 );
not ( n3301 , n43 );
not ( n3302 , n2781 );
or ( n3303 , n3301 , n3302 );
or ( n3304 , n2781 , n43 );
nand ( n3305 , n3303 , n3304 );
nand ( n3306 , n2722 , n3305 );
nand ( n3307 , n3300 , n3306 );
not ( n3308 , n3307 );
not ( n3309 , n2632 );
not ( n3310 , n1958 );
or ( n3311 , n3309 , n3310 );
nand ( n3312 , n3233 , n2581 );
nand ( n3313 , n3311 , n3312 );
not ( n3314 , n3313 );
not ( n3315 , n3314 );
or ( n3316 , n3308 , n3315 );
or ( n3317 , n3314 , n3307 );
nand ( n3318 , n3316 , n3317 );
xnor ( n3319 , n3291 , n3318 );
not ( n3320 , n3319 );
not ( n3321 , n3320 );
not ( n3322 , n51 );
not ( n3323 , n2220 );
or ( n3324 , n3322 , n3323 );
not ( n3325 , n2793 );
nand ( n3326 , n3325 , n756 );
nand ( n3327 , n3324 , n3326 );
nand ( n3328 , n840 , n44 );
not ( n3329 , n3328 );
nand ( n3330 , n3329 , n2782 );
nand ( n3331 , n2782 , n916 , n44 );
buf ( n3332 , n2577 );
nand ( n3333 , n3330 , n3331 , n3332 );
nand ( n3334 , n3327 , n3333 );
not ( n3335 , n3334 );
or ( n3336 , n2209 , n2700 );
or ( n3337 , n3256 , n2709 );
nand ( n3338 , n3336 , n3337 );
not ( n3339 , n3338 );
not ( n3340 , n3267 );
not ( n3341 , n2733 );
or ( n3342 , n3340 , n3341 );
nand ( n3343 , n2905 , n2236 );
nand ( n3344 , n3342 , n3343 );
not ( n3345 , n3344 );
not ( n3346 , n3345 );
or ( n3347 , n3339 , n3346 );
or ( n3348 , n3338 , n3345 );
nand ( n3349 , n3347 , n3348 );
and ( n3350 , n3335 , n3349 );
and ( n3351 , n3338 , n3344 );
nor ( n3352 , n3350 , n3351 );
not ( n3353 , n3352 );
not ( n3354 , n3353 );
or ( n3355 , n3321 , n3354 );
nand ( n3356 , n3319 , n3352 );
nand ( n3357 , n3355 , n3356 );
not ( n3358 , n3357 );
or ( n3359 , n3288 , n3358 );
or ( n3360 , n3357 , n3287 );
nand ( n3361 , n3359 , n3360 );
not ( n3362 , n3361 );
not ( n3363 , n2747 );
not ( n3364 , n3363 );
xor ( n3365 , n48 , n878 );
not ( n3366 , n3365 );
not ( n3367 , n3366 );
and ( n3368 , n3364 , n3367 );
and ( n3369 , n2179 , n2824 );
nor ( n3370 , n3368 , n3369 );
not ( n3371 , n3370 );
not ( n3372 , n3228 );
not ( n3373 , n46 );
and ( n3374 , n3372 , n3373 );
not ( n3375 , n1376 );
and ( n3376 , n3375 , n46 );
nor ( n3377 , n3374 , n3376 );
not ( n3378 , n3377 );
not ( n3379 , n3037 );
or ( n3380 , n3378 , n3379 );
buf ( n3381 , n2980 );
nand ( n3382 , n2208 , n3381 );
nand ( n3383 , n3380 , n3382 );
not ( n3384 , n3383 );
not ( n3385 , n2632 );
not ( n3386 , n3237 );
or ( n3387 , n3385 , n3386 );
and ( n3388 , n3 , n19 );
not ( n3389 , n3 );
and ( n3390 , n3389 , n35 );
nor ( n3391 , n3388 , n3390 );
and ( n3392 , n3391 , n45 );
not ( n3393 , n3391 );
and ( n3394 , n3393 , n840 );
nor ( n3395 , n3392 , n3394 );
nand ( n3396 , n2577 , n2579 );
nand ( n3397 , n3395 , n3396 );
nand ( n3398 , n3387 , n3397 );
not ( n3399 , n3398 );
not ( n3400 , n3399 );
or ( n3401 , n3384 , n3400 );
or ( n3402 , n3383 , n3399 );
nand ( n3403 , n3401 , n3402 );
nand ( n3404 , n3371 , n3403 );
nand ( n3405 , n3383 , n3398 );
and ( n3406 , n3404 , n3405 );
xnor ( n3407 , n3245 , n3221 );
not ( n3408 , n3407 );
and ( n3409 , n3406 , n3408 );
not ( n3410 , n3406 );
and ( n3411 , n3410 , n3407 );
nor ( n3412 , n3409 , n3411 );
and ( n3413 , n3349 , n3334 );
not ( n3414 , n3349 );
and ( n3415 , n3414 , n3335 );
nor ( n3416 , n3413 , n3415 );
or ( n3417 , n3412 , n3416 );
or ( n3418 , n3406 , n3407 );
nand ( n3419 , n3417 , n3418 );
nand ( n3420 , n3362 , n3419 );
not ( n3421 , n3420 );
xor ( n3422 , n3403 , n3370 );
not ( n3423 , n3422 );
not ( n3424 , n2905 );
not ( n3425 , n2299 );
or ( n3426 , n3424 , n3425 );
nand ( n3427 , n3365 , n2733 );
nand ( n3428 , n3426 , n3427 );
not ( n3429 , n3428 );
and ( n3430 , n50 , n51 );
not ( n3431 , n3430 );
not ( n3432 , n673 );
or ( n3433 , n3431 , n3432 );
not ( n3434 , n2314 );
nand ( n3435 , n3433 , n3434 );
not ( n3436 , n3435 );
nand ( n3437 , n1490 , n739 );
nand ( n3438 , n3436 , n2244 , n3437 );
not ( n3439 , n3438 );
not ( n3440 , n3391 );
nand ( n3441 , n3440 , n2585 );
not ( n3442 , n3441 );
or ( n3443 , n3439 , n3442 );
not ( n3444 , n3438 );
not ( n3445 , n3441 );
nand ( n3446 , n3444 , n3445 );
nand ( n3447 , n3443 , n3446 );
or ( n3448 , n3429 , n3447 );
nand ( n3449 , n3448 , n3446 );
not ( n3450 , n3449 );
nor ( n3451 , n3327 , n3333 );
not ( n3452 , n3451 );
nand ( n3453 , n3452 , n3334 );
not ( n3454 , n3453 );
and ( n3455 , n3450 , n3454 );
and ( n3456 , n3453 , n3449 );
nor ( n3457 , n3455 , n3456 );
not ( n3458 , n3457 );
or ( n3459 , n3423 , n3458 );
or ( n3460 , n3457 , n3422 );
nand ( n3461 , n3459 , n3460 );
and ( n3462 , n3447 , n3429 );
not ( n3463 , n3447 );
and ( n3464 , n3463 , n3428 );
nor ( n3465 , n3462 , n3464 );
not ( n3466 , n3465 );
not ( n3467 , n3466 );
not ( n3468 , n51 );
not ( n3469 , n2263 );
or ( n3470 , n3468 , n3469 );
not ( n3471 , n2793 );
nand ( n3472 , n2853 , n3471 );
nand ( n3473 , n3470 , n3472 );
nand ( n3474 , n2980 , n46 );
not ( n3475 , n3474 );
nand ( n3476 , n3475 , n2782 );
buf ( n3477 , n2697 );
nand ( n3478 , n3476 , n3477 );
nand ( n3479 , n3473 , n3478 );
not ( n3480 , n3479 );
not ( n3481 , n2869 );
not ( n3482 , n916 );
not ( n3483 , n3297 );
or ( n3484 , n3482 , n3483 );
or ( n3485 , n3297 , n916 );
nand ( n3486 , n3484 , n3485 );
not ( n3487 , n3486 );
or ( n3488 , n3481 , n3487 );
nand ( n3489 , n3377 , n3381 );
nand ( n3490 , n3488 , n3489 );
not ( n3491 , n3490 );
and ( n3492 , n3480 , n3491 );
and ( n3493 , n3479 , n3490 );
nor ( n3494 , n3492 , n3493 );
not ( n3495 , n3494 );
and ( n3496 , n3467 , n3495 );
not ( n3497 , n3479 );
and ( n3498 , n3497 , n3490 );
nor ( n3499 , n3496 , n3498 );
nor ( n3500 , n3461 , n3499 );
not ( n3501 , n3500 );
nand ( n3502 , n3461 , n3499 );
nand ( n3503 , n3501 , n3502 );
and ( n3504 , n2853 , n3218 );
not ( n3505 , n2853 );
and ( n3506 , n3505 , n3216 );
nor ( n3507 , n3504 , n3506 );
nand ( n3508 , n1109 , n3325 );
and ( n3509 , n3507 , n3508 );
not ( n3510 , n3509 );
and ( n3511 , n2781 , n3381 );
not ( n3512 , n3511 );
not ( n3513 , n2823 );
not ( n3514 , n3513 );
not ( n3515 , n48 );
not ( n3516 , n1185 );
not ( n3517 , n3516 );
or ( n3518 , n3515 , n3517 );
or ( n3519 , n1400 , n48 );
nand ( n3520 , n3518 , n3519 );
not ( n3521 , n3520 );
and ( n3522 , n3514 , n3521 );
not ( n3523 , n1624 );
not ( n3524 , n3297 );
or ( n3525 , n3523 , n3524 );
or ( n3526 , n3297 , n1621 );
nand ( n3527 , n3525 , n3526 );
and ( n3528 , n2905 , n3527 );
nor ( n3529 , n3522 , n3528 );
not ( n3530 , n3529 );
or ( n3531 , n3512 , n3530 );
or ( n3532 , n3529 , n3511 );
nand ( n3533 , n3531 , n3532 );
nand ( n3534 , n3510 , n3533 );
not ( n3535 , n3529 );
nand ( n3536 , n3535 , n3511 );
and ( n3537 , n3534 , n3536 );
not ( n3538 , n3537 );
not ( n3539 , n3391 );
not ( n3540 , n48 );
and ( n3541 , n3539 , n3540 );
not ( n3542 , n3440 );
and ( n3543 , n3542 , n48 );
nor ( n3544 , n3541 , n3543 );
not ( n3545 , n3544 );
not ( n3546 , n2869 );
or ( n3547 , n3545 , n3546 );
nand ( n3548 , n3486 , n2982 );
nand ( n3549 , n3547 , n3548 );
not ( n3550 , n3549 );
not ( n3551 , n2905 );
not ( n3552 , n3551 );
not ( n3553 , n3520 );
and ( n3554 , n3552 , n3553 );
and ( n3555 , n2299 , n2733 );
nor ( n3556 , n3554 , n3555 );
not ( n3557 , n3556 );
or ( n3558 , n3550 , n3557 );
or ( n3559 , n3549 , n3556 );
nand ( n3560 , n3558 , n3559 );
not ( n3561 , n3560 );
not ( n3562 , n3561 );
nor ( n3563 , n3473 , n3478 );
not ( n3564 , n3563 );
nand ( n3565 , n3564 , n3479 );
not ( n3566 , n3565 );
not ( n3567 , n3566 );
or ( n3568 , n3562 , n3567 );
nand ( n3569 , n3565 , n3560 );
nand ( n3570 , n3568 , n3569 );
not ( n3571 , n3570 );
or ( n3572 , n3538 , n3571 );
or ( n3573 , n3537 , n3570 );
nand ( n3574 , n3572 , n3573 );
and ( n3575 , n1788 , n2325 );
not ( n3576 , n1788 );
not ( n3577 , n1108 );
not ( n3578 , n1490 );
and ( n3579 , n3577 , n3578 );
and ( n3580 , n1108 , n1490 );
nor ( n3581 , n3579 , n3580 );
and ( n3582 , n3576 , n3581 );
nor ( n3583 , n3575 , n3582 );
nand ( n3584 , n2823 , n3440 );
nand ( n3585 , n3584 , n3108 );
nor ( n3586 , n3583 , n3585 );
not ( n3587 , n3586 );
xor ( n3588 , n3509 , n3533 );
xor ( n3589 , n3587 , n3588 );
not ( n3590 , n3527 );
not ( n3591 , n2733 );
or ( n3592 , n3590 , n3591 );
not ( n3593 , n2905 );
or ( n3594 , n3593 , n3544 );
nand ( n3595 , n3592 , n3594 );
not ( n3596 , n3584 );
not ( n3597 , n3596 );
not ( n3598 , n51 );
not ( n3599 , n2325 );
or ( n3600 , n3598 , n3599 );
nand ( n3601 , n1378 , n3216 );
nand ( n3602 , n3600 , n3601 );
not ( n3603 , n3602 );
or ( n3604 , n3597 , n3603 );
not ( n3605 , n3471 );
nand ( n3606 , n3605 , n2326 );
not ( n3607 , n2732 );
nand ( n3608 , n3607 , n2781 );
nand ( n3609 , n3606 , n3608 , n2660 );
nand ( n3610 , n3604 , n3609 );
xor ( n3611 , n3595 , n3610 );
and ( n3612 , n3583 , n3585 );
nor ( n3613 , n3612 , n3586 );
and ( n3614 , n3611 , n3613 );
and ( n3615 , n3595 , n3610 );
or ( n3616 , n3614 , n3615 );
not ( n3617 , n3616 );
and ( n3618 , n3589 , n3617 );
and ( n3619 , n3587 , n3588 );
or ( n3620 , n3618 , n3619 );
nand ( n3621 , n3574 , n3620 );
not ( n3622 , n3621 );
not ( n3623 , n3465 );
not ( n3624 , n3494 );
and ( n3625 , n3623 , n3624 );
and ( n3626 , n3494 , n3465 );
nor ( n3627 , n3625 , n3626 );
nand ( n3628 , n3566 , n3560 );
not ( n3629 , n3556 );
nand ( n3630 , n3629 , n3549 );
and ( n3631 , n3628 , n3630 );
nand ( n3632 , n3627 , n3631 );
not ( n3633 , n3570 );
nand ( n3634 , n3633 , n3537 );
and ( n3635 , n3632 , n3634 );
not ( n3636 , n3635 );
or ( n3637 , n3622 , n3636 );
not ( n3638 , n3631 );
not ( n3639 , n3627 );
nand ( n3640 , n3638 , n3639 );
nand ( n3641 , n3637 , n3640 );
nor ( n3642 , n3503 , n3641 );
not ( n3643 , n3502 );
nor ( n3644 , n3642 , n3643 );
not ( n3645 , n3457 );
not ( n3646 , n3422 );
not ( n3647 , n3646 );
and ( n3648 , n3645 , n3647 );
not ( n3649 , n3449 );
and ( n3650 , n3649 , n3453 );
nor ( n3651 , n3648 , n3650 );
and ( n3652 , n3412 , n3416 );
not ( n3653 , n3412 );
not ( n3654 , n3416 );
and ( n3655 , n3653 , n3654 );
nor ( n3656 , n3652 , n3655 );
not ( n3657 , n3656 );
and ( n3658 , n3651 , n3657 );
not ( n3659 , n3651 );
and ( n3660 , n3659 , n3656 );
nor ( n3661 , n3658 , n3660 );
nor ( n3662 , n3644 , n3661 );
not ( n3663 , n3662 );
or ( n3664 , n3421 , n3663 );
or ( n3665 , n3656 , n3651 );
not ( n3666 , n3665 );
not ( n3667 , n3419 );
not ( n3668 , n3667 );
not ( n3669 , n3361 );
not ( n3670 , n3669 );
or ( n3671 , n3668 , n3670 );
nand ( n3672 , n3361 , n3419 );
nand ( n3673 , n3671 , n3672 );
not ( n3674 , n3673 );
or ( n3675 , n3666 , n3674 );
nand ( n3676 , n3669 , n3419 );
nand ( n3677 , n3675 , n3676 );
nand ( n3678 , n3664 , n3677 );
not ( n3679 , n3287 );
and ( n3680 , n3357 , n3679 );
and ( n3681 , n3320 , n3352 );
nor ( n3682 , n3680 , n3681 );
not ( n3683 , n3682 );
not ( n3684 , n3283 );
not ( n3685 , n3249 );
or ( n3686 , n3684 , n3685 );
not ( n3687 , n3279 );
nand ( n3688 , n3687 , n3260 );
nand ( n3689 , n3686 , n3688 );
not ( n3690 , n3689 );
not ( n3691 , n2715 );
not ( n3692 , n3228 );
not ( n3693 , n42 );
and ( n3694 , n3692 , n3693 );
and ( n3695 , n3375 , n42 );
nor ( n3696 , n3694 , n3695 );
not ( n3697 , n3696 );
or ( n3698 , n3691 , n3697 );
nand ( n3699 , n3298 , n2722 );
nand ( n3700 , n3698 , n3699 );
not ( n3701 , n2640 );
not ( n3702 , n50 );
and ( n3703 , n3701 , n3702 );
nor ( n3704 , n3703 , n2314 );
not ( n3705 , n3060 );
nand ( n3706 , n2640 , n3705 );
and ( n3707 , n3704 , n2014 , n3706 );
xnor ( n3708 , n3700 , n3707 );
not ( n3709 , n1976 );
not ( n3710 , n3037 );
or ( n3711 , n3709 , n3710 );
not ( n3712 , n916 );
not ( n3713 , n675 );
or ( n3714 , n3712 , n3713 );
nand ( n3715 , n756 , n46 );
nand ( n3716 , n3714 , n3715 );
nand ( n3717 , n3716 , n3381 );
nand ( n3718 , n3711 , n3717 );
xor ( n3719 , n3708 , n3718 );
not ( n3720 , n3719 );
and ( n3721 , n3690 , n3720 );
and ( n3722 , n3689 , n3719 );
nor ( n3723 , n3721 , n3722 );
not ( n3724 , n2581 );
not ( n3725 , n1958 );
or ( n3726 , n3724 , n3725 );
not ( n3727 , n44 );
not ( n3728 , n2853 );
or ( n3729 , n3727 , n3728 );
or ( n3730 , n2853 , n44 );
nand ( n3731 , n3729 , n3730 );
nand ( n3732 , n3731 , n2587 );
nand ( n3733 , n3726 , n3732 );
xor ( n3734 , n3733 , n3278 );
nand ( n3735 , n2905 , n1983 );
xor ( n3736 , n48 , n521 );
nand ( n3737 , n2733 , n3736 );
nand ( n3738 , n3735 , n3737 );
not ( n3739 , n3738 );
not ( n3740 , n2533 );
nor ( n3741 , n41 , n42 );
nor ( n3742 , n3740 , n3741 );
nand ( n3743 , n2781 , n3742 );
buf ( n3744 , n3743 );
not ( n3745 , n3744 );
and ( n3746 , n3739 , n3745 );
and ( n3747 , n3738 , n3744 );
nor ( n3748 , n3746 , n3747 );
xnor ( n3749 , n3734 , n3748 );
not ( n3750 , n3307 );
not ( n3751 , n3313 );
or ( n3752 , n3750 , n3751 );
not ( n3753 , n3291 );
nand ( n3754 , n3753 , n3318 );
nand ( n3755 , n3752 , n3754 );
not ( n3756 , n3755 );
and ( n3757 , n3749 , n3756 );
not ( n3758 , n3749 );
and ( n3759 , n3758 , n3755 );
nor ( n3760 , n3757 , n3759 );
xor ( n3761 , n3723 , n3760 );
not ( n3762 , n3761 );
or ( n3763 , n3683 , n3762 );
or ( n3764 , n3761 , n3682 );
nand ( n3765 , n3763 , n3764 );
nand ( n3766 , n3678 , n3765 );
not ( n3767 , n3682 );
nand ( n3768 , n3767 , n3761 );
nand ( n3769 , n3766 , n3768 );
not ( n3770 , n3769 );
not ( n3771 , n3749 );
not ( n3772 , n3755 );
and ( n3773 , n3771 , n3772 );
xor ( n3774 , n3748 , n3733 );
and ( n3775 , n3774 , n3278 );
nor ( n3776 , n3773 , n3775 );
not ( n3777 , n2550 );
not ( n3778 , n40 );
not ( n3779 , n2660 );
or ( n3780 , n3778 , n3779 );
or ( n3781 , n2660 , n40 );
nand ( n3782 , n3780 , n3781 );
not ( n3783 , n3782 );
or ( n3784 , n3777 , n3783 );
and ( n3785 , n2782 , n41 );
not ( n3786 , n2782 );
and ( n3787 , n3786 , n424 );
nor ( n3788 , n3785 , n3787 );
nand ( n3789 , n3788 , n3043 );
nand ( n3790 , n3784 , n3789 );
not ( n3791 , n2982 );
not ( n3792 , n1924 );
or ( n3793 , n3791 , n3792 );
nand ( n3794 , n3037 , n3716 );
nand ( n3795 , n3793 , n3794 );
xor ( n3796 , n3790 , n3795 );
not ( n3797 , n3736 );
not ( n3798 , n2905 );
or ( n3799 , n3797 , n3798 );
not ( n3800 , n3607 );
nand ( n3801 , n3800 , n1890 );
nand ( n3802 , n3799 , n3801 );
not ( n3803 , n3743 );
and ( n3804 , n2533 , n40 );
not ( n3805 , n3804 );
nor ( n3806 , n3803 , n3805 );
nor ( n3807 , n3802 , n3806 );
not ( n3808 , n3807 );
nand ( n3809 , n3806 , n3802 );
nand ( n3810 , n3808 , n3809 );
not ( n3811 , n3810 );
and ( n3812 , n3796 , n3811 );
not ( n3813 , n3796 );
and ( n3814 , n3813 , n3810 );
nor ( n3815 , n3812 , n3814 );
and ( n3816 , n3776 , n3815 );
not ( n3817 , n3776 );
not ( n3818 , n3815 );
and ( n3819 , n3817 , n3818 );
nor ( n3820 , n3816 , n3819 );
not ( n3821 , n3820 );
not ( n3822 , n3700 );
not ( n3823 , n3707 );
and ( n3824 , n3822 , n3823 );
and ( n3825 , n3707 , n3700 );
nor ( n3826 , n3825 , n3718 );
nor ( n3827 , n3824 , n3826 );
not ( n3828 , n3748 );
not ( n3829 , n3733 );
and ( n3830 , n3828 , n3829 );
and ( n3831 , n3744 , n3735 , n3737 );
nor ( n3832 , n3830 , n3831 );
xor ( n3833 , n3827 , n3832 );
not ( n3834 , n2632 );
not ( n3835 , n1877 );
or ( n3836 , n3834 , n3835 );
not ( n3837 , n3731 );
or ( n3838 , n3837 , n2955 );
nand ( n3839 , n3836 , n3838 );
not ( n3840 , n2641 );
not ( n3841 , n3840 );
not ( n3842 , n3210 );
and ( n3843 , n3841 , n3842 );
and ( n3844 , n1916 , n51 );
nor ( n3845 , n3843 , n3844 );
not ( n3846 , n3845 );
not ( n3847 , n2715 );
not ( n3848 , n2024 );
or ( n3849 , n3847 , n3848 );
nand ( n3850 , n2722 , n3696 );
nand ( n3851 , n3849 , n3850 );
not ( n3852 , n3851 );
or ( n3853 , n3846 , n3852 );
or ( n3854 , n3845 , n3851 );
nand ( n3855 , n3853 , n3854 );
xor ( n3856 , n3839 , n3855 );
xor ( n3857 , n3833 , n3856 );
or ( n3858 , n3821 , n3857 );
buf ( n3859 , n3776 );
or ( n3860 , n3859 , n3815 );
nand ( n3861 , n3858 , n3860 );
not ( n3862 , n3861 );
or ( n3863 , n1876 , n2955 );
and ( n3864 , n675 , n968 );
and ( n3865 , n756 , n44 );
nor ( n3866 , n3864 , n3865 );
or ( n3867 , n3866 , n2633 );
nand ( n3868 , n3863 , n3867 );
not ( n3869 , n3868 );
not ( n3870 , n2562 );
nor ( n3871 , n2782 , n3870 );
not ( n3872 , n3871 );
not ( n3873 , n2005 );
not ( n3874 , n2747 );
or ( n3875 , n3873 , n3874 );
xor ( n3876 , n2645 , n48 );
nand ( n3877 , n3876 , n2732 );
nand ( n3878 , n3875 , n3877 );
not ( n3879 , n3878 );
not ( n3880 , n3879 );
or ( n3881 , n3872 , n3880 );
not ( n3882 , n3871 );
nand ( n3883 , n3878 , n3882 );
nand ( n3884 , n3881 , n3883 );
not ( n3885 , n3884 );
or ( n3886 , n3869 , n3885 );
or ( n3887 , n3868 , n3884 );
nand ( n3888 , n3886 , n3887 );
not ( n3889 , n3888 );
not ( n3890 , n3889 );
not ( n3891 , n3796 );
not ( n3892 , n3811 );
or ( n3893 , n3891 , n3892 );
nand ( n3894 , n3795 , n3790 );
nand ( n3895 , n3893 , n3894 );
not ( n3896 , n3895 );
not ( n3897 , n3896 );
or ( n3898 , n3890 , n3897 );
nand ( n3899 , n3888 , n3895 );
nand ( n3900 , n3898 , n3899 );
not ( n3901 , n2550 );
not ( n3902 , n3228 );
not ( n3903 , n40 );
and ( n3904 , n3902 , n3903 );
and ( n3905 , n3375 , n40 );
nor ( n3906 , n3904 , n3905 );
not ( n3907 , n3906 );
or ( n3908 , n3901 , n3907 );
nand ( n3909 , n3043 , n3782 );
nand ( n3910 , n3908 , n3909 );
and ( n3911 , n360 , n3705 );
not ( n3912 , n360 );
and ( n3913 , n3912 , n3216 );
nor ( n3914 , n3911 , n3913 );
nand ( n3915 , n409 , n2795 );
nand ( n3916 , n3914 , n3915 );
xor ( n3917 , n3910 , n3916 );
or ( n3918 , n2025 , n2986 );
xor ( n3919 , n42 , n2853 );
not ( n3920 , n3007 );
or ( n3921 , n3919 , n3920 );
nand ( n3922 , n3918 , n3921 );
xor ( n3923 , n3917 , n3922 );
xor ( n3924 , n3900 , n3923 );
not ( n3925 , n3924 );
and ( n3926 , n3833 , n3856 );
and ( n3927 , n3827 , n3832 );
nor ( n3928 , n3926 , n3927 );
not ( n3929 , n3839 );
not ( n3930 , n3855 );
or ( n3931 , n3929 , n3930 );
not ( n3932 , n3845 );
nand ( n3933 , n3932 , n3851 );
nand ( n3934 , n3931 , n3933 );
not ( n3935 , n3809 );
not ( n3936 , n1924 );
not ( n3937 , n2699 );
or ( n3938 , n3936 , n3937 );
and ( n3939 , n587 , n46 );
not ( n3940 , n587 );
and ( n3941 , n3940 , n916 );
nor ( n3942 , n3939 , n3941 );
or ( n3943 , n3942 , n2709 );
nand ( n3944 , n3938 , n3943 );
not ( n3945 , n3944 );
or ( n3946 , n3935 , n3945 );
or ( n3947 , n3944 , n3809 );
nand ( n3948 , n3946 , n3947 );
xnor ( n3949 , n3934 , n3948 );
and ( n3950 , n3928 , n3949 );
not ( n3951 , n3928 );
not ( n3952 , n3949 );
and ( n3953 , n3951 , n3952 );
nor ( n3954 , n3950 , n3953 );
not ( n3955 , n3954 );
not ( n3956 , n3955 );
or ( n3957 , n3925 , n3956 );
not ( n3958 , n3924 );
nand ( n3959 , n3958 , n3954 );
nand ( n3960 , n3957 , n3959 );
not ( n3961 , n3960 );
or ( n3962 , n3862 , n3961 );
or ( n3963 , n3861 , n3960 );
nand ( n3964 , n3962 , n3963 );
not ( n3965 , n3964 );
not ( n3966 , n3928 );
not ( n3967 , n3949 );
and ( n3968 , n3966 , n3967 );
and ( n3969 , n3954 , n3924 );
nor ( n3970 , n3968 , n3969 );
not ( n3971 , n3970 );
not ( n3972 , n3923 );
not ( n3973 , n3900 );
or ( n3974 , n3972 , n3973 );
not ( n3975 , n3896 );
nand ( n3976 , n3975 , n3889 );
nand ( n3977 , n3974 , n3976 );
not ( n3978 , n3922 );
not ( n3979 , n3917 );
or ( n3980 , n3978 , n3979 );
nand ( n3981 , n3910 , n3916 );
nand ( n3982 , n3980 , n3981 );
not ( n3983 , n2701 );
not ( n3984 , n3325 );
not ( n3985 , n3984 );
and ( n3986 , n3983 , n3985 );
and ( n3987 , n1636 , n51 );
nor ( n3988 , n3986 , n3987 );
not ( n3989 , n3988 );
nand ( n3990 , n39 , n40 );
and ( n3991 , n3990 , n38 );
not ( n3992 , n3991 );
nor ( n3993 , n3871 , n3992 );
nand ( n3994 , n3989 , n3993 );
not ( n3995 , n3993 );
nand ( n3996 , n3995 , n3988 );
and ( n3997 , n3994 , n3996 );
not ( n3998 , n3997 );
and ( n3999 , n3982 , n3998 );
not ( n4000 , n3982 );
and ( n4001 , n4000 , n3997 );
or ( n4002 , n3999 , n4001 );
not ( n4003 , n4002 );
not ( n4004 , n3882 );
not ( n4005 , n3879 );
or ( n4006 , n4004 , n4005 );
not ( n4007 , n3868 );
nand ( n4008 , n4007 , n3884 );
nand ( n4009 , n4006 , n4008 );
not ( n4010 , n4009 );
and ( n4011 , n4003 , n4010 );
and ( n4012 , n4002 , n4009 );
nor ( n4013 , n4011 , n4012 );
or ( n4014 , n3977 , n4013 );
not ( n4015 , n3923 );
not ( n4016 , n3900 );
or ( n4017 , n4015 , n4016 );
nand ( n4018 , n4017 , n3976 );
nand ( n4019 , n4018 , n4013 );
nand ( n4020 , n4014 , n4019 );
not ( n4021 , n4020 );
not ( n4022 , n3007 );
not ( n4023 , n1665 );
or ( n4024 , n4022 , n4023 );
xnor ( n4025 , n42 , n2853 );
nand ( n4026 , n4025 , n2722 );
nand ( n4027 , n4024 , n4026 );
not ( n4028 , n3593 );
not ( n4029 , n3876 );
not ( n4030 , n4029 );
and ( n4031 , n4028 , n4030 );
and ( n4032 , n2732 , n1626 );
nor ( n4033 , n4031 , n4032 );
xnor ( n4034 , n4027 , n4033 );
or ( n4035 , n3866 , n2955 );
or ( n4036 , n1792 , n2633 );
nand ( n4037 , n4035 , n4036 );
xnor ( n4038 , n4034 , n4037 );
not ( n4039 , n4038 );
or ( n4040 , n2868 , n3942 );
or ( n4041 , n1681 , n2709 );
nand ( n4042 , n4040 , n4041 );
not ( n4043 , n4042 );
not ( n4044 , n2573 );
not ( n4045 , n38 );
not ( n4046 , n2660 );
or ( n4047 , n4045 , n4046 );
or ( n4048 , n2660 , n38 );
nand ( n4049 , n4047 , n4048 );
not ( n4050 , n4049 );
or ( n4051 , n4044 , n4050 );
and ( n4052 , n38 , n3391 );
not ( n4053 , n38 );
and ( n4054 , n4053 , n3440 );
or ( n4055 , n4052 , n4054 );
nand ( n4056 , n4055 , n2564 );
nand ( n4057 , n4051 , n4056 );
not ( n4058 , n2550 );
not ( n4059 , n1770 );
or ( n4060 , n4058 , n4059 );
nand ( n4061 , n3906 , n3043 );
nand ( n4062 , n4060 , n4061 );
xor ( n4063 , n4057 , n4062 );
not ( n4064 , n4063 );
not ( n4065 , n4064 );
or ( n4066 , n4043 , n4065 );
not ( n4067 , n4042 );
nand ( n4068 , n4067 , n4063 );
nand ( n4069 , n4066 , n4068 );
not ( n4070 , n4069 );
or ( n4071 , n4039 , n4070 );
or ( n4072 , n4069 , n4038 );
nand ( n4073 , n4071 , n4072 );
not ( n4074 , n3948 );
not ( n4075 , n3934 );
or ( n4076 , n4074 , n4075 );
not ( n4077 , n3809 );
nand ( n4078 , n4077 , n3944 );
nand ( n4079 , n4076 , n4078 );
xnor ( n4080 , n4073 , n4079 );
not ( n4081 , n4080 );
or ( n4082 , n4021 , n4081 );
or ( n4083 , n4080 , n4020 );
nand ( n4084 , n4082 , n4083 );
nand ( n4085 , n3971 , n4084 );
or ( n4086 , n3723 , n3760 );
not ( n4087 , n3719 );
or ( n4088 , n3689 , n4087 );
nand ( n4089 , n4086 , n4088 );
not ( n4090 , n4089 );
xor ( n4091 , n3820 , n3857 );
not ( n4092 , n4091 );
or ( n4093 , n4090 , n4092 );
or ( n4094 , n4091 , n4089 );
nand ( n4095 , n4093 , n4094 );
nand ( n4096 , n4085 , n4095 );
nor ( n4097 , n3965 , n4096 );
not ( n4098 , n4097 );
or ( n4099 , n3770 , n4098 );
xor ( n4100 , n4084 , n3970 );
not ( n4101 , n3964 );
not ( n4102 , n4091 );
nand ( n4103 , n4102 , n4089 );
or ( n4104 , n4101 , n4103 );
not ( n4105 , n3960 );
nand ( n4106 , n4105 , n3861 );
nand ( n4107 , n4104 , n4106 );
or ( n4108 , n4100 , n4107 );
nand ( n4109 , n4108 , n4085 );
nand ( n4110 , n4099 , n4109 );
not ( n4111 , n4110 );
not ( n4112 , n4080 );
and ( n4113 , n4112 , n4020 );
not ( n4114 , n4013 );
and ( n4115 , n4018 , n4114 );
nor ( n4116 , n4113 , n4115 );
not ( n4117 , n4116 );
not ( n4118 , n4037 );
not ( n4119 , n4034 );
or ( n4120 , n4118 , n4119 );
not ( n4121 , n4033 );
nand ( n4122 , n4121 , n4027 );
nand ( n4123 , n4120 , n4122 );
not ( n4124 , n1626 );
not ( n4125 , n2905 );
or ( n4126 , n4124 , n4125 );
nand ( n4127 , n2830 , n2733 );
nand ( n4128 , n4126 , n4127 );
not ( n4129 , n4128 );
not ( n4130 , n2783 );
not ( n4131 , n4130 );
not ( n4132 , n2790 );
not ( n4133 , n50 );
and ( n4134 , n4132 , n4133 );
nor ( n4135 , n4134 , n1591 );
and ( n4136 , n3705 , n2790 );
nor ( n4137 , n4136 , n2314 );
and ( n4138 , n4135 , n4137 );
not ( n4139 , n4138 );
or ( n4140 , n4131 , n4139 );
not ( n4141 , n4130 );
nand ( n4142 , n4135 , n4137 );
nand ( n4143 , n4141 , n4142 );
nand ( n4144 , n4140 , n4143 );
not ( n4145 , n4144 );
not ( n4146 , n4145 );
or ( n4147 , n4129 , n4146 );
not ( n4148 , n4128 );
nand ( n4149 , n4148 , n4144 );
nand ( n4150 , n4147 , n4149 );
xor ( n4151 , n4123 , n4150 );
not ( n4152 , n4042 );
not ( n4153 , n4063 );
or ( n4154 , n4152 , n4153 );
nand ( n4155 , n4062 , n4057 );
nand ( n4156 , n4154 , n4155 );
xnor ( n4157 , n4151 , n4156 );
not ( n4158 , n4079 );
not ( n4159 , n4073 );
or ( n4160 , n4158 , n4159 );
not ( n4161 , n4038 );
nand ( n4162 , n4161 , n4069 );
nand ( n4163 , n4160 , n4162 );
xnor ( n4164 , n4157 , n4163 );
not ( n4165 , n4009 );
not ( n4166 , n4165 );
not ( n4167 , n4002 );
or ( n4168 , n4166 , n4167 );
nand ( n4169 , n3982 , n3997 );
nand ( n4170 , n4168 , n4169 );
not ( n4171 , n3043 );
not ( n4172 , n1770 );
or ( n4173 , n4171 , n4172 );
nand ( n4174 , n2550 , n2855 );
nand ( n4175 , n4173 , n4174 );
not ( n4176 , n4175 );
xor ( n4177 , n1377 , n38 );
not ( n4178 , n4177 );
not ( n4179 , n2926 );
and ( n4180 , n4178 , n4179 );
and ( n4181 , n2564 , n4049 );
nor ( n4182 , n4180 , n4181 );
not ( n4183 , n4182 );
or ( n4184 , n4176 , n4183 );
or ( n4185 , n4175 , n4182 );
nand ( n4186 , n4184 , n4185 );
not ( n4187 , n3994 );
and ( n4188 , n4186 , n4187 );
not ( n4189 , n4186 );
not ( n4190 , n4187 );
and ( n4191 , n4189 , n4190 );
nor ( n4192 , n4188 , n4191 );
not ( n4193 , n449 );
xor ( n4194 , n46 , n4193 );
not ( n4195 , n4194 );
not ( n4196 , n2699 );
or ( n4197 , n4195 , n4196 );
nand ( n4198 , n2866 , n3381 );
nand ( n4199 , n4197 , n4198 );
not ( n4200 , n2722 );
not ( n4201 , n1785 );
or ( n4202 , n4200 , n4201 );
nand ( n4203 , n2841 , n2713 );
nand ( n4204 , n4202 , n4203 );
xor ( n4205 , n4199 , n4204 );
or ( n4206 , n2955 , n1792 );
not ( n4207 , n2805 );
or ( n4208 , n4207 , n2633 );
nand ( n4209 , n4206 , n4208 );
and ( n4210 , n4205 , n4209 );
not ( n4211 , n4205 );
not ( n4212 , n4209 );
and ( n4213 , n4211 , n4212 );
nor ( n4214 , n4210 , n4213 );
xor ( n4215 , n4192 , n4214 );
buf ( n4216 , n4215 );
xor ( n4217 , n4170 , n4216 );
xor ( n4218 , n4164 , n4217 );
not ( n4219 , n4218 );
or ( n4220 , n4117 , n4219 );
or ( n4221 , n4218 , n4116 );
nand ( n4222 , n4220 , n4221 );
not ( n4223 , n4222 );
or ( n4224 , n4111 , n4223 );
and ( n4225 , n4164 , n4217 );
not ( n4226 , n4157 );
and ( n4227 , n4163 , n4226 );
nor ( n4228 , n4225 , n4227 );
not ( n4229 , n4228 );
not ( n4230 , n4214 );
not ( n4231 , n4192 );
or ( n4232 , n4230 , n4231 );
nand ( n4233 , n4170 , n4215 );
nand ( n4234 , n4232 , n4233 );
not ( n4235 , n2832 );
and ( n4236 , n2821 , n4235 );
not ( n4237 , n2821 );
and ( n4238 , n4237 , n2832 );
nor ( n4239 , n4236 , n4238 );
not ( n4240 , n4209 );
not ( n4241 , n4205 );
or ( n4242 , n4240 , n4241 );
nand ( n4243 , n4199 , n4204 );
nand ( n4244 , n4242 , n4243 );
and ( n4245 , n4239 , n4244 );
not ( n4246 , n4239 );
not ( n4247 , n4244 );
and ( n4248 , n4246 , n4247 );
or ( n4249 , n4245 , n4248 );
xor ( n4250 , n2874 , n2862 );
and ( n4251 , n4249 , n4250 );
not ( n4252 , n4249 );
not ( n4253 , n4250 );
and ( n4254 , n4252 , n4253 );
nor ( n4255 , n4251 , n4254 );
xor ( n4256 , n4234 , n4255 );
not ( n4257 , n4156 );
not ( n4258 , n4151 );
or ( n4259 , n4257 , n4258 );
nand ( n4260 , n4150 , n4123 );
nand ( n4261 , n4259 , n4260 );
buf ( n4262 , n4261 );
not ( n4263 , n4262 );
not ( n4264 , n4175 );
not ( n4265 , n4264 );
not ( n4266 , n4182 );
and ( n4267 , n4265 , n4266 );
and ( n4268 , n4186 , n4187 );
nor ( n4269 , n4267 , n4268 );
not ( n4270 , n4269 );
not ( n4271 , n4270 );
not ( n4272 , n4128 );
not ( n4273 , n4144 );
or ( n4274 , n4272 , n4273 );
not ( n4275 , n4130 );
nand ( n4276 , n4275 , n4138 );
nand ( n4277 , n4274 , n4276 );
not ( n4278 , n4277 );
nor ( n4279 , n2784 , n2797 );
not ( n4280 , n4279 );
nand ( n4281 , n4280 , n2798 );
not ( n4282 , n4281 );
not ( n4283 , n2564 );
not ( n4284 , n4177 );
not ( n4285 , n4284 );
or ( n4286 , n4283 , n4285 );
or ( n4287 , n1523 , n3870 );
nand ( n4288 , n4286 , n4287 );
not ( n4289 , n4288 );
and ( n4290 , n4282 , n4289 );
and ( n4291 , n4281 , n4288 );
nor ( n4292 , n4290 , n4291 );
not ( n4293 , n4292 );
or ( n4294 , n4278 , n4293 );
or ( n4295 , n4292 , n4277 );
nand ( n4296 , n4294 , n4295 );
not ( n4297 , n4296 );
not ( n4298 , n4297 );
or ( n4299 , n4271 , n4298 );
nand ( n4300 , n4296 , n4269 );
nand ( n4301 , n4299 , n4300 );
not ( n4302 , n4301 );
and ( n4303 , n4263 , n4302 );
and ( n4304 , n4301 , n4262 );
nor ( n4305 , n4303 , n4304 );
not ( n4306 , n4305 );
and ( n4307 , n4256 , n4306 );
not ( n4308 , n4256 );
and ( n4309 , n4308 , n4305 );
nor ( n4310 , n4307 , n4309 );
not ( n4311 , n4310 );
not ( n4312 , n4311 );
or ( n4313 , n4229 , n4312 );
not ( n4314 , n4228 );
nand ( n4315 , n4314 , n4310 );
nand ( n4316 , n4313 , n4315 );
not ( n4317 , n4218 );
nand ( n4318 , n4317 , n4116 );
and ( n4319 , n4316 , n4318 );
nand ( n4320 , n4224 , n4319 );
nand ( n4321 , n2875 , n2877 );
and ( n4322 , n2836 , n4321 );
not ( n4323 , n2836 );
and ( n4324 , n4323 , n2878 );
nor ( n4325 , n4322 , n4324 );
not ( n4326 , n4277 );
or ( n4327 , n4326 , n4292 );
not ( n4328 , n4288 );
or ( n4329 , n4281 , n4328 );
nand ( n4330 , n4327 , n4329 );
and ( n4331 , n4325 , n4330 );
not ( n4332 , n4325 );
not ( n4333 , n4330 );
and ( n4334 , n4332 , n4333 );
nor ( n4335 , n4331 , n4334 );
not ( n4336 , n4335 );
not ( n4337 , n4336 );
not ( n4338 , n4247 );
not ( n4339 , n4239 );
and ( n4340 , n4338 , n4339 );
and ( n4341 , n4249 , n4250 );
nor ( n4342 , n4340 , n4341 );
not ( n4343 , n4342 );
not ( n4344 , n4343 );
or ( n4345 , n4337 , n4344 );
nand ( n4346 , n4335 , n4342 );
nand ( n4347 , n4345 , n4346 );
xor ( n4348 , n3177 , n3172 );
not ( n4349 , n4348 );
not ( n4350 , n4270 );
not ( n4351 , n4350 );
not ( n4352 , n4297 );
or ( n4353 , n4351 , n4352 );
not ( n4354 , n4261 );
nand ( n4355 , n4354 , n4301 );
nand ( n4356 , n4353 , n4355 );
not ( n4357 , n4356 );
not ( n4358 , n4357 );
or ( n4359 , n4349 , n4358 );
not ( n4360 , n4348 );
nand ( n4361 , n4360 , n4356 );
nand ( n4362 , n4359 , n4361 );
xor ( n4363 , n4347 , n4362 );
not ( n4364 , n4363 );
and ( n4365 , n4305 , n4256 );
and ( n4366 , n4234 , n4255 );
nor ( n4367 , n4365 , n4366 );
buf ( n4368 , n4367 );
nand ( n4369 , n4364 , n4368 );
not ( n4370 , n3152 );
not ( n4371 , n3201 );
or ( n4372 , n4370 , n4371 );
or ( n4373 , n3152 , n3201 );
nand ( n4374 , n4372 , n4373 );
not ( n4375 , n4374 );
not ( n4376 , n4336 );
not ( n4377 , n4342 );
and ( n4378 , n4376 , n4377 );
and ( n4379 , n4325 , n4330 );
nor ( n4380 , n4378 , n4379 );
not ( n4381 , n4380 );
not ( n4382 , n4381 );
xor ( n4383 , n2881 , n2773 );
buf ( n4384 , n4383 );
not ( n4385 , n4384 );
xor ( n4386 , n3186 , n3179 );
not ( n4387 , n4386 );
not ( n4388 , n4387 );
or ( n4389 , n4385 , n4388 );
not ( n4390 , n4383 );
nand ( n4391 , n4390 , n4386 );
nand ( n4392 , n4389 , n4391 );
not ( n4393 , n4392 );
or ( n4394 , n4382 , n4393 );
nand ( n4395 , n4386 , n4384 );
nand ( n4396 , n4394 , n4395 );
not ( n4397 , n4396 );
nand ( n4398 , n4375 , n4397 );
xor ( n4399 , n4380 , n4392 );
and ( n4400 , n4347 , n4362 );
not ( n4401 , n4357 );
nor ( n4402 , n4401 , n4348 );
nor ( n4403 , n4400 , n4402 );
xor ( n4404 , n4399 , n4403 );
nand ( n4405 , n4369 , n4398 , n4404 );
or ( n4406 , n4320 , n4405 );
not ( n4407 , n4368 );
xor ( n4408 , n4363 , n4407 );
not ( n4409 , n4228 );
nand ( n4410 , n4409 , n4311 );
nand ( n4411 , n4408 , n4410 );
and ( n4412 , n4404 , n4398 , n4369 );
and ( n4413 , n4411 , n4412 );
not ( n4414 , n4403 );
and ( n4415 , n4392 , n4380 );
not ( n4416 , n4392 );
and ( n4417 , n4416 , n4381 );
or ( n4418 , n4415 , n4417 );
nand ( n4419 , n4414 , n4418 );
not ( n4420 , n4419 );
xor ( n4421 , n4374 , n4396 );
not ( n4422 , n4421 );
or ( n4423 , n4420 , n4422 );
nand ( n4424 , n4423 , n4398 );
not ( n4425 , n3205 );
not ( n4426 , n3150 );
or ( n4427 , n4425 , n4426 );
or ( n4428 , n3205 , n3150 );
nand ( n4429 , n4427 , n4428 );
nand ( n4430 , n4424 , n4429 );
nor ( n4431 , n4413 , n4430 );
nand ( n4432 , n4406 , n4431 );
nand ( n4433 , n3208 , n4432 );
and ( n4434 , n2966 , n3149 );
and ( n4435 , n2894 , n2961 );
nor ( n4436 , n4434 , n4435 );
not ( n4437 , n4436 );
not ( n4438 , n3148 );
not ( n4439 , n3093 );
and ( n4440 , n4438 , n4439 );
not ( n4441 , n3099 );
and ( n4442 , n3147 , n4441 );
nor ( n4443 , n4440 , n4442 );
xor ( n4444 , n2922 , n2944 );
and ( n4445 , n4444 , n2960 );
and ( n4446 , n2922 , n2944 );
nor ( n4447 , n4445 , n4446 );
and ( n4448 , n4443 , n4447 );
not ( n4449 , n4443 );
not ( n4450 , n4447 );
and ( n4451 , n4449 , n4450 );
nor ( n4452 , n4448 , n4451 );
not ( n4453 , n3118 );
not ( n4454 , n4453 );
not ( n4455 , n3143 );
or ( n4456 , n4454 , n4455 );
not ( n4457 , n3125 );
nand ( n4458 , n4457 , n3139 );
nand ( n4459 , n4456 , n4458 );
not ( n4460 , n2699 );
not ( n4461 , n922 );
or ( n4462 , n4460 , n4461 );
nand ( n4463 , n4462 , n3474 );
not ( n4464 , n4463 );
and ( n4465 , n2954 , n2959 );
and ( n4466 , n2946 , n2953 );
nor ( n4467 , n4465 , n4466 );
xnor ( n4468 , n4464 , n4467 );
not ( n4469 , n3117 );
not ( n4470 , n3113 );
or ( n4471 , n4469 , n4470 );
not ( n4472 , n3104 );
not ( n4473 , n3109 );
or ( n4474 , n4472 , n4473 );
nand ( n4475 , n4471 , n4474 );
xor ( n4476 , n4468 , n4475 );
xor ( n4477 , n4459 , n4476 );
not ( n4478 , n952 );
not ( n4479 , n2564 );
or ( n4480 , n4478 , n4479 );
not ( n4481 , n38 );
not ( n4482 , n587 );
or ( n4483 , n4481 , n4482 );
or ( n4484 , n38 , n587 );
nand ( n4485 , n4483 , n4484 );
nand ( n4486 , n4485 , n2927 );
nand ( n4487 , n4480 , n4486 );
not ( n4488 , n4487 );
and ( n4489 , n933 , n3043 );
not ( n4490 , n2640 );
not ( n4491 , n40 );
and ( n4492 , n4490 , n4491 );
and ( n4493 , n2646 , n40 );
nor ( n4494 , n4492 , n4493 );
and ( n4495 , n2550 , n4494 );
nor ( n4496 , n4489 , n4495 );
not ( n4497 , n4496 );
or ( n4498 , n4488 , n4497 );
or ( n4499 , n4487 , n4496 );
nand ( n4500 , n4498 , n4499 );
or ( n4501 , n971 , n2955 );
and ( n4502 , n968 , n2790 );
not ( n4503 , n968 );
not ( n4504 , n2790 );
and ( n4505 , n4503 , n4504 );
nor ( n4506 , n4502 , n4505 );
or ( n4507 , n4506 , n2633 );
nand ( n4508 , n4501 , n4507 );
xnor ( n4509 , n4500 , n4508 );
not ( n4510 , n4509 );
not ( n4511 , n961 );
not ( n4512 , n2722 );
or ( n4513 , n4511 , n4512 );
not ( n4514 , n42 );
not ( n4515 , n2595 );
or ( n4516 , n4514 , n4515 );
or ( n4517 , n2595 , n42 );
nand ( n4518 , n4516 , n4517 );
nand ( n4519 , n4518 , n2715 );
nand ( n4520 , n4513 , n4519 );
not ( n4521 , n4520 );
not ( n4522 , n2897 );
not ( n4523 , n4522 );
and ( n4524 , n4521 , n4523 );
and ( n4525 , n4520 , n4522 );
nor ( n4526 , n4524 , n4525 );
not ( n4527 , n4526 );
not ( n4528 , n2678 );
nand ( n4529 , n1101 , n4528 );
xor ( n4530 , n36 , n675 );
nand ( n4531 , n4530 , n3011 );
and ( n4532 , n4529 , n4531 );
not ( n4533 , n4532 );
or ( n4534 , n4527 , n4533 );
or ( n4535 , n4526 , n4532 );
nand ( n4536 , n4534 , n4535 );
not ( n4537 , n4536 );
not ( n4538 , n2939 );
not ( n4539 , n2934 );
or ( n4540 , n4538 , n4539 );
nand ( n4541 , n2929 , n2910 );
nand ( n4542 , n4540 , n4541 );
not ( n4543 , n4542 );
or ( n4544 , n4537 , n4543 );
or ( n4545 , n4536 , n4542 );
nand ( n4546 , n4544 , n4545 );
not ( n4547 , n4546 );
or ( n4548 , n4510 , n4547 );
or ( n4549 , n4546 , n4509 );
nand ( n4550 , n4548 , n4549 );
xor ( n4551 , n4477 , n4550 );
xor ( n4552 , n4452 , n4551 );
not ( n4553 , n4552 );
or ( n4554 , n4437 , n4553 );
or ( n4555 , n4552 , n4436 );
nand ( n4556 , n4554 , n4555 );
nor ( n4557 , n4433 , n4556 );
not ( n4558 , n4557 );
nand ( n4559 , n4433 , n4556 );
buf ( n4560 , n4559 );
nand ( n4561 , n4558 , n4560 );
nand ( n4562 , n1 , n2 );
not ( n4563 , n4562 );
nand ( n4564 , n4561 , n4563 );
or ( n4565 , n36 , n62 );
nand ( n4566 , n36 , n62 );
nand ( n4567 , n4565 , n4566 );
or ( n4568 , n2678 , n4567 );
or ( n4569 , n36 , n61 );
nand ( n4570 , n36 , n61 );
nand ( n4571 , n4569 , n4570 );
or ( n4572 , n2776 , n4571 );
nand ( n4573 , n4568 , n4572 );
not ( n4574 , n3920 );
and ( n4575 , n42 , n55 );
not ( n4576 , n42 );
not ( n4577 , n55 );
and ( n4578 , n4576 , n4577 );
nor ( n4579 , n4575 , n4578 );
not ( n4580 , n4579 );
not ( n4581 , n4580 );
and ( n4582 , n4574 , n4581 );
and ( n4583 , n42 , n56 );
not ( n4584 , n42 );
not ( n4585 , n56 );
and ( n4586 , n4584 , n4585 );
nor ( n4587 , n4583 , n4586 );
and ( n4588 , n2722 , n4587 );
nor ( n4589 , n4582 , n4588 );
and ( n4590 , n36 , n63 );
xnor ( n4591 , n4589 , n4590 );
xor ( n4592 , n4573 , n4591 );
and ( n4593 , n38 , n60 );
not ( n4594 , n38 );
not ( n4595 , n60 );
and ( n4596 , n4594 , n4595 );
nor ( n4597 , n4593 , n4596 );
and ( n4598 , n2564 , n4597 );
and ( n4599 , n38 , n59 );
nor ( n4600 , n38 , n59 );
nor ( n4601 , n4599 , n4600 );
and ( n4602 , n2573 , n4601 );
nor ( n4603 , n4598 , n4602 );
not ( n4604 , n4603 );
not ( n4605 , n44 );
not ( n4606 , n54 );
and ( n4607 , n4605 , n4606 );
and ( n4608 , n44 , n54 );
nor ( n4609 , n4607 , n4608 );
not ( n4610 , n4609 );
not ( n4611 , n2581 );
or ( n4612 , n4610 , n4611 );
and ( n4613 , n44 , n53 );
not ( n4614 , n44 );
not ( n4615 , n53 );
and ( n4616 , n4614 , n4615 );
nor ( n4617 , n4613 , n4616 );
nand ( n4618 , n2587 , n4617 );
nand ( n4619 , n4612 , n4618 );
not ( n4620 , n4619 );
or ( n4621 , n4604 , n4620 );
or ( n4622 , n4603 , n4619 );
nand ( n4623 , n4621 , n4622 );
not ( n4624 , n40 );
not ( n4625 , n58 );
and ( n4626 , n4624 , n4625 );
and ( n4627 , n40 , n58 );
nor ( n4628 , n4626 , n4627 );
and ( n4629 , n2951 , n4628 );
not ( n4630 , n57 );
and ( n4631 , n427 , n4630 );
and ( n4632 , n40 , n57 );
nor ( n4633 , n4631 , n4632 );
and ( n4634 , n2550 , n4633 );
nor ( n4635 , n4629 , n4634 );
not ( n4636 , n4635 );
and ( n4637 , n4623 , n4636 );
not ( n4638 , n4623 );
and ( n4639 , n4638 , n4635 );
nor ( n4640 , n4637 , n4639 );
not ( n4641 , n2901 );
nor ( n4642 , n36 , n63 );
or ( n4643 , n4590 , n4642 );
or ( n4644 , n4641 , n4643 );
or ( n4645 , n2776 , n4567 );
nand ( n4646 , n4644 , n4645 );
not ( n4647 , n4646 );
not ( n4648 , n2926 );
not ( n4649 , n4597 );
not ( n4650 , n4649 );
and ( n4651 , n4648 , n4650 );
not ( n4652 , n38 );
not ( n4653 , n61 );
and ( n4654 , n4652 , n4653 );
and ( n4655 , n38 , n61 );
nor ( n4656 , n4654 , n4655 );
and ( n4657 , n2564 , n4656 );
nor ( n4658 , n4651 , n4657 );
not ( n4659 , n4658 );
and ( n4660 , n4647 , n4659 );
buf ( n4661 , n4646 );
and ( n4662 , n4661 , n4658 );
nor ( n4663 , n4660 , n4662 );
and ( n4664 , n48 , n52 );
not ( n4665 , n48 );
not ( n4666 , n52 );
and ( n4667 , n4665 , n4666 );
nor ( n4668 , n4664 , n4667 );
not ( n4669 , n4668 );
not ( n4670 , n2748 );
or ( n4671 , n4669 , n4670 );
nand ( n4672 , n4671 , n2909 );
not ( n4673 , n4672 );
or ( n4674 , n4663 , n4673 );
not ( n4675 , n4661 );
or ( n4676 , n4675 , n4658 );
nand ( n4677 , n4674 , n4676 );
and ( n4678 , n4640 , n4677 );
not ( n4679 , n4640 );
not ( n4680 , n4677 );
and ( n4681 , n4679 , n4680 );
nor ( n4682 , n4678 , n4681 );
xnor ( n4683 , n4592 , n4682 );
and ( n4684 , n54 , n46 );
not ( n4685 , n54 );
and ( n4686 , n4685 , n916 );
nor ( n4687 , n4684 , n4686 );
not ( n4688 , n4687 );
not ( n4689 , n3037 );
or ( n4690 , n4688 , n4689 );
and ( n4691 , n46 , n53 );
not ( n4692 , n46 );
and ( n4693 , n4692 , n4615 );
nor ( n4694 , n4691 , n4693 );
nand ( n4695 , n3381 , n4694 );
nand ( n4696 , n4690 , n4695 );
nand ( n4697 , n36 , n65 );
xor ( n4698 , n4696 , n4697 );
not ( n4699 , n4698 );
not ( n4700 , n2986 );
not ( n4701 , n58 );
and ( n4702 , n42 , n4701 );
not ( n4703 , n42 );
and ( n4704 , n4703 , n58 );
nor ( n4705 , n4702 , n4704 );
not ( n4706 , n4705 );
and ( n4707 , n4700 , n4706 );
and ( n4708 , n1899 , n4630 );
and ( n4709 , n42 , n57 );
nor ( n4710 , n4708 , n4709 );
and ( n4711 , n3007 , n4710 );
nor ( n4712 , n4707 , n4711 );
and ( n4713 , n4699 , n4712 );
not ( n4714 , n4697 );
nor ( n4715 , n4714 , n4696 );
nor ( n4716 , n4713 , n4715 );
not ( n4717 , n4716 );
not ( n4718 , n38 );
not ( n4719 , n62 );
and ( n4720 , n4718 , n4719 );
and ( n4721 , n38 , n62 );
nor ( n4722 , n4720 , n4721 );
and ( n4723 , n2564 , n4722 );
and ( n4724 , n2573 , n4656 );
nor ( n4725 , n4723 , n4724 );
not ( n4726 , n4725 );
not ( n4727 , n2581 );
and ( n4728 , n44 , n56 );
not ( n4729 , n44 );
and ( n4730 , n4729 , n4585 );
nor ( n4731 , n4728 , n4730 );
not ( n4732 , n4731 );
or ( n4733 , n4727 , n4732 );
not ( n4734 , n2586 );
and ( n4735 , n44 , n55 );
not ( n4736 , n44 );
and ( n4737 , n4736 , n4577 );
nor ( n4738 , n4735 , n4737 );
nand ( n4739 , n4734 , n4738 );
nand ( n4740 , n4733 , n4739 );
not ( n4741 , n4740 );
and ( n4742 , n427 , n4595 );
and ( n4743 , n40 , n60 );
nor ( n4744 , n4742 , n4743 );
not ( n4745 , n4744 );
not ( n4746 , n3042 );
or ( n4747 , n4745 , n4746 );
and ( n4748 , n40 , n59 );
not ( n4749 , n40 );
not ( n4750 , n59 );
and ( n4751 , n4749 , n4750 );
nor ( n4752 , n4748 , n4751 );
nand ( n4753 , n2550 , n4752 );
nand ( n4754 , n4747 , n4753 );
not ( n4755 , n4754 );
not ( n4756 , n4755 );
or ( n4757 , n4741 , n4756 );
not ( n4758 , n4740 );
nand ( n4759 , n4758 , n4754 );
nand ( n4760 , n4757 , n4759 );
nand ( n4761 , n4726 , n4760 );
not ( n4762 , n4755 );
nand ( n4763 , n4762 , n4740 );
and ( n4764 , n4761 , n4763 );
not ( n4765 , n4764 );
and ( n4766 , n4717 , n4765 );
and ( n4767 , n4716 , n4764 );
nor ( n4768 , n4766 , n4767 );
not ( n4769 , n4768 );
and ( n4770 , n2870 , n4694 );
and ( n4771 , n46 , n52 );
not ( n4772 , n46 );
and ( n4773 , n4772 , n4666 );
nor ( n4774 , n4771 , n4773 );
and ( n4775 , n3381 , n4774 );
nor ( n4776 , n4770 , n4775 );
and ( n4777 , n2722 , n4710 );
and ( n4778 , n2715 , n4587 );
nor ( n4779 , n4777 , n4778 );
and ( n4780 , n4779 , n3109 );
not ( n4781 , n4779 );
and ( n4782 , n4781 , n3108 );
nor ( n4783 , n4780 , n4782 );
xor ( n4784 , n4776 , n4783 );
and ( n4785 , n4769 , n4784 );
not ( n4786 , n4764 );
and ( n4787 , n4716 , n4786 );
nor ( n4788 , n4785 , n4787 );
nand ( n4789 , n36 , n64 );
not ( n4790 , n4789 );
not ( n4791 , n4752 );
not ( n4792 , n2541 );
or ( n4793 , n4791 , n4792 );
nand ( n4794 , n2550 , n4628 );
nand ( n4795 , n4793 , n4794 );
not ( n4796 , n4795 );
or ( n4797 , n4790 , n4796 );
or ( n4798 , n4795 , n4789 );
nand ( n4799 , n4797 , n4798 );
not ( n4800 , n4799 );
and ( n4801 , n2581 , n4738 );
and ( n4802 , n2632 , n4609 );
nor ( n4803 , n4801 , n4802 );
not ( n4804 , n4803 );
not ( n4805 , n4804 );
or ( n4806 , n4800 , n4805 );
not ( n4807 , n4789 );
nand ( n4808 , n4807 , n4795 );
nand ( n4809 , n4806 , n4808 );
not ( n4810 , n4774 );
not ( n4811 , n2699 );
or ( n4812 , n4810 , n4811 );
nand ( n4813 , n4812 , n3474 );
not ( n4814 , n4813 );
and ( n4815 , n4809 , n4814 );
not ( n4816 , n4809 );
and ( n4817 , n4816 , n4813 );
nor ( n4818 , n4815 , n4817 );
not ( n4819 , n4818 );
not ( n4820 , n4819 );
or ( n4821 , n4783 , n4776 );
or ( n4822 , n4779 , n4473 );
nand ( n4823 , n4821 , n4822 );
not ( n4824 , n4823 );
and ( n4825 , n4820 , n4824 );
and ( n4826 , n4819 , n4823 );
nor ( n4827 , n4825 , n4826 );
not ( n4828 , n4827 );
and ( n4829 , n4788 , n4828 );
not ( n4830 , n4788 );
and ( n4831 , n4830 , n4827 );
nor ( n4832 , n4829 , n4831 );
xor ( n4833 , n4683 , n4832 );
not ( n4834 , n4833 );
and ( n4835 , n42 , n60 );
not ( n4836 , n42 );
and ( n4837 , n4836 , n4595 );
nor ( n4838 , n4835 , n4837 );
not ( n4839 , n4838 );
not ( n4840 , n43 );
not ( n4841 , n44 );
nor ( n4842 , n4841 , n42 );
not ( n4843 , n4842 );
or ( n4844 , n4840 , n4843 );
nand ( n4845 , n4844 , n2719 );
not ( n4846 , n4845 );
or ( n4847 , n4839 , n4846 );
and ( n4848 , n42 , n59 );
not ( n4849 , n42 );
and ( n4850 , n4849 , n4750 );
nor ( n4851 , n4848 , n4850 );
nand ( n4852 , n2713 , n4851 );
nand ( n4853 , n4847 , n4852 );
not ( n4854 , n4853 );
not ( n4855 , n4854 );
not ( n4856 , n3396 );
and ( n4857 , n44 , n58 );
not ( n4858 , n44 );
and ( n4859 , n4858 , n4701 );
nor ( n4860 , n4857 , n4859 );
not ( n4861 , n4860 );
or ( n4862 , n4856 , n4861 );
and ( n4863 , n44 , n57 );
not ( n4864 , n44 );
and ( n4865 , n4864 , n4630 );
nor ( n4866 , n4863 , n4865 );
nand ( n4867 , n2631 , n4866 );
nand ( n4868 , n4862 , n4867 );
not ( n4869 , n4868 );
not ( n4870 , n4869 );
or ( n4871 , n4855 , n4870 );
not ( n4872 , n4868 );
not ( n4873 , n4853 );
or ( n4874 , n4872 , n4873 );
xor ( n4875 , n36 , n66 );
not ( n4876 , n4875 );
not ( n4877 , n2818 );
or ( n4878 , n4876 , n4877 );
or ( n4879 , n36 , n65 );
nand ( n4880 , n4879 , n4697 );
not ( n4881 , n4880 );
nand ( n4882 , n4881 , n2681 );
nand ( n4883 , n4878 , n4882 );
not ( n4884 , n4883 );
nand ( n4885 , n4874 , n4884 );
nand ( n4886 , n4871 , n4885 );
not ( n4887 , n4886 );
nand ( n4888 , n36 , n67 );
not ( n4889 , n4888 );
not ( n4890 , n50 );
not ( n4891 , n4666 );
or ( n4892 , n4890 , n4891 );
nand ( n4893 , n4892 , n3060 );
nand ( n4894 , n4889 , n4893 );
not ( n4895 , n4893 );
nand ( n4896 , n4895 , n4888 );
and ( n4897 , n4894 , n4896 );
not ( n4898 , n4897 );
xor ( n4899 , n48 , n54 );
not ( n4900 , n4899 );
not ( n4901 , n2905 );
or ( n4902 , n4900 , n4901 );
and ( n4903 , n48 , n53 );
not ( n4904 , n48 );
and ( n4905 , n4904 , n4615 );
nor ( n4906 , n4903 , n4905 );
nand ( n4907 , n2732 , n4906 );
nand ( n4908 , n4902 , n4907 );
not ( n4909 , n4908 );
or ( n4910 , n4898 , n4909 );
nand ( n4911 , n4910 , n4894 );
not ( n4912 , n4911 );
not ( n4913 , n4912 );
and ( n4914 , n4887 , n4913 );
and ( n4915 , n4886 , n4911 );
not ( n4916 , n4886 );
and ( n4917 , n4916 , n4912 );
or ( n4918 , n4915 , n4917 );
and ( n4919 , n46 , n56 );
not ( n4920 , n46 );
and ( n4921 , n4920 , n4585 );
nor ( n4922 , n4919 , n4921 );
not ( n4923 , n4922 );
not ( n4924 , n2699 );
or ( n4925 , n4923 , n4924 );
and ( n4926 , n46 , n55 );
not ( n4927 , n46 );
and ( n4928 , n4927 , n4577 );
nor ( n4929 , n4926 , n4928 );
nand ( n4930 , n3381 , n4929 );
nand ( n4931 , n4925 , n4930 );
not ( n4932 , n4931 );
and ( n4933 , n40 , n62 );
not ( n4934 , n40 );
not ( n4935 , n62 );
and ( n4936 , n4934 , n4935 );
nor ( n4937 , n4933 , n4936 );
not ( n4938 , n4937 );
not ( n4939 , n3042 );
or ( n4940 , n4938 , n4939 );
not ( n4941 , n40 );
not ( n4942 , n61 );
and ( n4943 , n4941 , n4942 );
and ( n4944 , n40 , n61 );
nor ( n4945 , n4943 , n4944 );
nand ( n4946 , n3742 , n4945 );
nand ( n4947 , n4940 , n4946 );
nor ( n4948 , n2561 , n2562 );
and ( n4949 , n38 , n64 );
not ( n4950 , n38 );
not ( n4951 , n64 );
and ( n4952 , n4950 , n4951 );
nor ( n4953 , n4949 , n4952 );
and ( n4954 , n4948 , n4953 );
not ( n4955 , n38 );
not ( n4956 , n63 );
and ( n4957 , n4955 , n4956 );
and ( n4958 , n38 , n63 );
nor ( n4959 , n4957 , n4958 );
and ( n4960 , n2562 , n4959 );
nor ( n4961 , n4954 , n4960 );
not ( n4962 , n4961 );
and ( n4963 , n4947 , n4962 );
not ( n4964 , n4947 );
and ( n4965 , n4964 , n4961 );
nor ( n4966 , n4963 , n4965 );
not ( n4967 , n4966 );
or ( n4968 , n4932 , n4967 );
nand ( n4969 , n4947 , n4962 );
nand ( n4970 , n4968 , n4969 );
and ( n4971 , n4918 , n4970 );
nor ( n4972 , n4914 , n4971 );
buf ( n4973 , n4972 );
and ( n4974 , n4712 , n4698 );
not ( n4975 , n4712 );
and ( n4976 , n4975 , n4699 );
or ( n4977 , n4974 , n4976 );
or ( n4978 , n36 , n64 );
nand ( n4979 , n4978 , n4789 );
not ( n4980 , n4979 );
nand ( n4981 , n4980 , n2818 );
not ( n4982 , n4643 );
nand ( n4983 , n4982 , n2813 );
nand ( n4984 , n4981 , n4983 );
not ( n4985 , n4984 );
not ( n4986 , n4866 );
not ( n4987 , n3396 );
or ( n4988 , n4986 , n4987 );
nand ( n4989 , n2587 , n4731 );
nand ( n4990 , n4988 , n4989 );
not ( n4991 , n4990 );
not ( n4992 , n4991 );
or ( n4993 , n4985 , n4992 );
or ( n4994 , n4984 , n4991 );
nand ( n4995 , n4993 , n4994 );
not ( n4996 , n4995 );
not ( n4997 , n4672 );
and ( n4998 , n4996 , n4997 );
and ( n4999 , n4995 , n4672 );
nor ( n5000 , n4998 , n4999 );
xnor ( n5001 , n4977 , n5000 );
or ( n5002 , n4973 , n5001 );
or ( n5003 , n4977 , n5000 );
nand ( n5004 , n5002 , n5003 );
not ( n5005 , n5004 );
and ( n5006 , n2699 , n4929 );
and ( n5007 , n2982 , n4687 );
nor ( n5008 , n5006 , n5007 );
not ( n5009 , n5008 );
not ( n5010 , n5009 );
not ( n5011 , n2714 );
not ( n5012 , n4705 );
and ( n5013 , n5011 , n5012 );
and ( n5014 , n4845 , n4851 );
nor ( n5015 , n5013 , n5014 );
not ( n5016 , n5015 );
not ( n5017 , n5016 );
not ( n5018 , n4906 );
not ( n5019 , n2905 );
or ( n5020 , n5018 , n5019 );
nand ( n5021 , n2824 , n4668 );
nand ( n5022 , n5020 , n5021 );
not ( n5023 , n5022 );
not ( n5024 , n5023 );
or ( n5025 , n5017 , n5024 );
nand ( n5026 , n5015 , n5022 );
nand ( n5027 , n5025 , n5026 );
not ( n5028 , n5027 );
or ( n5029 , n5010 , n5028 );
nand ( n5030 , n5022 , n5016 );
nand ( n5031 , n5029 , n5030 );
not ( n5032 , n5031 );
not ( n5033 , n5032 );
xor ( n5034 , n4725 , n4760 );
nand ( n5035 , n36 , n66 );
not ( n5036 , n5035 );
not ( n5037 , n50 );
and ( n5038 , n5036 , n5037 );
not ( n5039 , n2818 );
or ( n5040 , n5039 , n4880 );
or ( n5041 , n2814 , n4979 );
nand ( n5042 , n5040 , n5041 );
xor ( n5043 , n5035 , n50 );
and ( n5044 , n5042 , n5043 );
nor ( n5045 , n5038 , n5044 );
xor ( n5046 , n5034 , n5045 );
not ( n5047 , n5046 );
or ( n5048 , n5033 , n5047 );
or ( n5049 , n4760 , n4725 );
nand ( n5050 , n4760 , n4725 );
nand ( n5051 , n5049 , n5050 , n5045 );
nand ( n5052 , n5048 , n5051 );
not ( n5053 , n5052 );
not ( n5054 , n4784 );
not ( n5055 , n4768 );
or ( n5056 , n5054 , n5055 );
or ( n5057 , n4784 , n4768 );
nand ( n5058 , n5056 , n5057 );
xor ( n5059 , n5053 , n5058 );
not ( n5060 , n5059 );
or ( n5061 , n5005 , n5060 );
nand ( n5062 , n5058 , n5053 );
nand ( n5063 , n5061 , n5062 );
and ( n5064 , n4799 , n4804 );
not ( n5065 , n4799 );
and ( n5066 , n5065 , n4803 );
nor ( n5067 , n5064 , n5066 );
and ( n5068 , n4995 , n4673 );
and ( n5069 , n4990 , n4984 );
nor ( n5070 , n5068 , n5069 );
xnor ( n5071 , n5067 , n5070 );
and ( n5072 , n4663 , n4673 );
not ( n5073 , n4663 );
and ( n5074 , n5073 , n4672 );
nor ( n5075 , n5072 , n5074 );
and ( n5076 , n5071 , n5075 );
not ( n5077 , n5070 );
and ( n5078 , n5077 , n5067 );
nor ( n5079 , n5076 , n5078 );
not ( n5080 , n5079 );
and ( n5081 , n5063 , n5080 );
not ( n5082 , n5063 );
and ( n5083 , n5082 , n5079 );
or ( n5084 , n5081 , n5083 );
not ( n5085 , n5084 );
or ( n5086 , n4834 , n5085 );
or ( n5087 , n5084 , n4833 );
nand ( n5088 , n5086 , n5087 );
xor ( n5089 , n5059 , n5004 );
not ( n5090 , n5089 );
xnor ( n5091 , n5008 , n5027 );
and ( n5092 , n5042 , n5043 );
not ( n5093 , n5042 );
not ( n5094 , n5043 );
and ( n5095 , n5093 , n5094 );
nor ( n5096 , n5092 , n5095 );
xnor ( n5097 , n5091 , n5096 );
not ( n5098 , n5097 );
and ( n5099 , n44 , n59 );
not ( n5100 , n44 );
and ( n5101 , n5100 , n4750 );
nor ( n5102 , n5099 , n5101 );
and ( n5103 , n3396 , n5102 );
and ( n5104 , n2587 , n4860 );
nor ( n5105 , n5103 , n5104 );
not ( n5106 , n5105 );
and ( n5107 , n48 , n55 );
not ( n5108 , n48 );
and ( n5109 , n5108 , n4577 );
nor ( n5110 , n5107 , n5109 );
not ( n5111 , n5110 );
not ( n5112 , n50 );
nand ( n5113 , n5112 , n48 , n1363 );
nand ( n5114 , n5113 , n2744 );
not ( n5115 , n5114 );
or ( n5116 , n5111 , n5115 );
nand ( n5117 , n2823 , n4899 );
nand ( n5118 , n5116 , n5117 );
not ( n5119 , n4875 );
not ( n5120 , n2675 );
and ( n5121 , n5119 , n5120 );
nand ( n5122 , n2673 , n2674 );
and ( n5123 , n38 , n67 );
not ( n5124 , n38 );
not ( n5125 , n67 );
and ( n5126 , n5124 , n5125 );
nor ( n5127 , n5123 , n5126 );
not ( n5128 , n5127 );
nand ( n5129 , n5128 , n2676 );
and ( n5130 , n5122 , n5129 );
nor ( n5131 , n5121 , n5130 );
xor ( n5132 , n5118 , n5131 );
nand ( n5133 , n5106 , n5132 );
nand ( n5134 , n5118 , n5131 );
nand ( n5135 , n5133 , n5134 );
not ( n5136 , n5135 );
not ( n5137 , n5136 );
nand ( n5138 , n2813 , n67 );
nand ( n5139 , n5138 , n2774 );
not ( n5140 , n52 );
not ( n5141 , n3061 );
or ( n5142 , n5140 , n5141 );
not ( n5143 , n51 );
and ( n5144 , n5143 , n53 );
nor ( n5145 , n50 , n52 );
nor ( n5146 , n5144 , n2314 , n5145 );
nand ( n5147 , n5142 , n5146 );
nor ( n5148 , n5139 , n5147 );
not ( n5149 , n5148 );
not ( n5150 , n5149 );
and ( n5151 , n5137 , n5150 );
not ( n5152 , n5148 );
not ( n5153 , n5136 );
or ( n5154 , n5152 , n5153 );
nand ( n5155 , n5149 , n5135 );
nand ( n5156 , n5154 , n5155 );
and ( n5157 , n42 , n61 );
not ( n5158 , n42 );
and ( n5159 , n5158 , n4653 );
nor ( n5160 , n5157 , n5159 );
and ( n5161 , n2722 , n5160 );
and ( n5162 , n2715 , n4838 );
nor ( n5163 , n5161 , n5162 );
not ( n5164 , n5163 );
not ( n5165 , n40 );
not ( n5166 , n63 );
and ( n5167 , n5165 , n5166 );
and ( n5168 , n40 , n63 );
nor ( n5169 , n5167 , n5168 );
and ( n5170 , n3042 , n5169 );
and ( n5171 , n3742 , n4937 );
nor ( n5172 , n5170 , n5171 );
not ( n5173 , n5172 );
and ( n5174 , n46 , n57 );
not ( n5175 , n46 );
and ( n5176 , n5175 , n4630 );
nor ( n5177 , n5174 , n5176 );
not ( n5178 , n5177 );
not ( n5179 , n48 );
not ( n5180 , n2694 );
or ( n5181 , n5179 , n5180 );
nand ( n5182 , n2121 , n1624 , n46 );
nand ( n5183 , n5181 , n5182 );
not ( n5184 , n5183 );
or ( n5185 , n5178 , n5184 );
nand ( n5186 , n3381 , n4922 );
nand ( n5187 , n5185 , n5186 );
not ( n5188 , n5187 );
or ( n5189 , n5173 , n5188 );
or ( n5190 , n5187 , n5172 );
nand ( n5191 , n5189 , n5190 );
nand ( n5192 , n5164 , n5191 );
not ( n5193 , n5172 );
nand ( n5194 , n5193 , n5187 );
nand ( n5195 , n5192 , n5194 );
and ( n5196 , n5156 , n5195 );
nor ( n5197 , n5151 , n5196 );
not ( n5198 , n5197 );
and ( n5199 , n5098 , n5198 );
and ( n5200 , n5091 , n5096 );
nor ( n5201 , n5199 , n5200 );
not ( n5202 , n5201 );
nand ( n5203 , n4948 , n4959 );
nand ( n5204 , n2562 , n4722 );
and ( n5205 , n5203 , n5204 );
xor ( n5206 , n5205 , n4990 );
and ( n5207 , n2951 , n4945 );
and ( n5208 , n2550 , n4744 );
nor ( n5209 , n5207 , n5208 );
and ( n5210 , n5206 , n5209 );
and ( n5211 , n5205 , n4990 );
nor ( n5212 , n5210 , n5211 );
xor ( n5213 , n5031 , n5212 );
not ( n5214 , n5046 );
xnor ( n5215 , n5213 , n5214 );
not ( n5216 , n5215 );
or ( n5217 , n5202 , n5216 );
and ( n5218 , n5214 , n5032 );
and ( n5219 , n5046 , n5031 );
nor ( n5220 , n5218 , n5219 );
or ( n5221 , n5220 , n5212 );
nand ( n5222 , n5217 , n5221 );
xnor ( n5223 , n5071 , n5075 );
xor ( n5224 , n5222 , n5223 );
not ( n5225 , n5224 );
or ( n5226 , n5090 , n5225 );
or ( n5227 , n5222 , n5223 );
nand ( n5228 , n5226 , n5227 );
nor ( n5229 , n5088 , n5228 );
not ( n5230 , n5229 );
nand ( n5231 , n5228 , n5088 );
nand ( n5232 , n5230 , n5231 );
not ( n5233 , n5232 );
xnor ( n5234 , n5224 , n5089 );
not ( n5235 , n5201 );
and ( n5236 , n5215 , n5235 );
not ( n5237 , n5215 );
and ( n5238 , n5237 , n5201 );
nor ( n5239 , n5236 , n5238 );
xor ( n5240 , n4966 , n4931 );
not ( n5241 , n5240 );
not ( n5242 , n4869 );
not ( n5243 , n4853 );
or ( n5244 , n5242 , n5243 );
nand ( n5245 , n4854 , n4868 );
nand ( n5246 , n5244 , n5245 );
buf ( n5247 , n4883 );
xnor ( n5248 , n5246 , n5247 );
xor ( n5249 , n4897 , n4908 );
not ( n5250 , n5249 );
and ( n5251 , n5248 , n5250 );
not ( n5252 , n5248 );
and ( n5253 , n5252 , n5249 );
nor ( n5254 , n5251 , n5253 );
not ( n5255 , n5254 );
or ( n5256 , n5241 , n5255 );
not ( n5257 , n5248 );
nand ( n5258 , n5257 , n5249 );
nand ( n5259 , n5256 , n5258 );
xor ( n5260 , n5205 , n4990 );
xor ( n5261 , n5260 , n5209 );
not ( n5262 , n5261 );
xor ( n5263 , n4918 , n4970 );
not ( n5264 , n5263 );
or ( n5265 , n5262 , n5264 );
or ( n5266 , n5261 , n5263 );
nand ( n5267 , n5265 , n5266 );
nand ( n5268 , n5259 , n5267 );
not ( n5269 , n5261 );
nand ( n5270 , n5269 , n5263 );
and ( n5271 , n5268 , n5270 );
xor ( n5272 , n5001 , n4973 );
not ( n5273 , n5272 );
and ( n5274 , n5271 , n5273 );
not ( n5275 , n5271 );
and ( n5276 , n5275 , n5272 );
nor ( n5277 , n5274 , n5276 );
and ( n5278 , n5239 , n5277 );
not ( n5279 , n5271 );
and ( n5280 , n5279 , n5272 );
nor ( n5281 , n5278 , n5280 );
buf ( n5282 , n5281 );
or ( n5283 , n5234 , n5282 );
not ( n5284 , n5282 );
not ( n5285 , n5234 );
or ( n5286 , n5284 , n5285 );
not ( n5287 , n66 );
and ( n5288 , n916 , n5287 );
and ( n5289 , n46 , n66 );
nor ( n5290 , n5288 , n5289 );
not ( n5291 , n5290 );
not ( n5292 , n2869 );
or ( n5293 , n5291 , n5292 );
not ( n5294 , n65 );
and ( n5295 , n916 , n5294 );
and ( n5296 , n46 , n65 );
nor ( n5297 , n5295 , n5296 );
nand ( n5298 , n2982 , n5297 );
nand ( n5299 , n5293 , n5298 );
not ( n5300 , n63 );
not ( n5301 , n5300 );
not ( n5302 , n3325 );
or ( n5303 , n5301 , n5302 );
and ( n5304 , n3216 , n62 );
and ( n5305 , n3061 , n4935 );
nor ( n5306 , n5304 , n5305 );
nand ( n5307 , n5303 , n5306 );
or ( n5308 , n3474 , n67 );
nand ( n5309 , n5308 , n3477 );
nand ( n5310 , n5307 , n5309 );
xor ( n5311 , n5299 , n5310 );
and ( n5312 , n4653 , n3061 );
not ( n5313 , n4653 );
and ( n5314 , n5313 , n3216 );
nor ( n5315 , n5312 , n5314 );
nand ( n5316 , n3471 , n4935 );
nand ( n5317 , n5315 , n5316 );
and ( n5318 , n2587 , n67 );
nor ( n5319 , n5317 , n5318 );
not ( n5320 , n5319 );
nand ( n5321 , n5317 , n5318 );
nand ( n5322 , n5320 , n5321 );
not ( n5323 , n5322 );
not ( n5324 , n48 );
not ( n5325 , n64 );
and ( n5326 , n5324 , n5325 );
and ( n5327 , n48 , n64 );
nor ( n5328 , n5326 , n5327 );
and ( n5329 , n2747 , n5328 );
and ( n5330 , n48 , n63 );
not ( n5331 , n48 );
and ( n5332 , n5331 , n5300 );
nor ( n5333 , n5330 , n5332 );
and ( n5334 , n2733 , n5333 );
nor ( n5335 , n5329 , n5334 );
not ( n5336 , n5335 );
not ( n5337 , n5336 );
and ( n5338 , n5323 , n5337 );
and ( n5339 , n5322 , n5336 );
nor ( n5340 , n5338 , n5339 );
or ( n5341 , n5311 , n5340 );
not ( n5342 , n5299 );
or ( n5343 , n5342 , n5310 );
nand ( n5344 , n5341 , n5343 );
not ( n5345 , n5344 );
not ( n5346 , n5345 );
not ( n5347 , n5322 );
not ( n5348 , n5335 );
and ( n5349 , n5347 , n5348 );
not ( n5350 , n5321 );
nor ( n5351 , n5349 , n5350 );
nand ( n5352 , n2585 , n44 );
not ( n5353 , n5352 );
not ( n5354 , n67 );
and ( n5355 , n5353 , n5354 );
not ( n5356 , n3332 );
nor ( n5357 , n5355 , n5356 );
not ( n5358 , n5357 );
not ( n5359 , n4653 );
not ( n5360 , n2795 );
or ( n5361 , n5359 , n5360 );
and ( n5362 , n3216 , n60 );
and ( n5363 , n3061 , n4595 );
nor ( n5364 , n5362 , n5363 );
nand ( n5365 , n5361 , n5364 );
not ( n5366 , n5365 );
not ( n5367 , n5366 );
or ( n5368 , n5358 , n5367 );
not ( n5369 , n5357 );
nand ( n5370 , n5369 , n5365 );
nand ( n5371 , n5368 , n5370 );
not ( n5372 , n5371 );
and ( n5373 , n5351 , n5372 );
not ( n5374 , n5351 );
and ( n5375 , n5374 , n5371 );
nor ( n5376 , n5373 , n5375 );
not ( n5377 , n5376 );
not ( n5378 , n5297 );
not ( n5379 , n5183 );
or ( n5380 , n5378 , n5379 );
and ( n5381 , n46 , n64 );
not ( n5382 , n46 );
and ( n5383 , n5382 , n4951 );
nor ( n5384 , n5381 , n5383 );
nand ( n5385 , n3381 , n5384 );
nand ( n5386 , n5380 , n5385 );
not ( n5387 , n5333 );
not ( n5388 , n2747 );
or ( n5389 , n5387 , n5388 );
and ( n5390 , n48 , n62 );
not ( n5391 , n48 );
and ( n5392 , n5391 , n4935 );
nor ( n5393 , n5390 , n5392 );
nand ( n5394 , n2733 , n5393 );
nand ( n5395 , n5389 , n5394 );
xor ( n5396 , n5386 , n5395 );
not ( n5397 , n44 );
not ( n5398 , n67 );
and ( n5399 , n5397 , n5398 );
and ( n5400 , n44 , n67 );
nor ( n5401 , n5399 , n5400 );
and ( n5402 , n2581 , n5401 );
and ( n5403 , n968 , n5287 );
and ( n5404 , n44 , n66 );
nor ( n5405 , n5403 , n5404 );
and ( n5406 , n2587 , n5405 );
nor ( n5407 , n5402 , n5406 );
not ( n5408 , n5407 );
and ( n5409 , n5396 , n5408 );
not ( n5410 , n5396 );
and ( n5411 , n5410 , n5407 );
nor ( n5412 , n5409 , n5411 );
not ( n5413 , n5412 );
and ( n5414 , n5377 , n5413 );
not ( n5415 , n5412 );
not ( n5416 , n5415 );
and ( n5417 , n5416 , n5376 );
nor ( n5418 , n5414 , n5417 );
not ( n5419 , n5418 );
or ( n5420 , n5346 , n5419 );
xor ( n5421 , n5418 , n5345 );
or ( n5422 , n5309 , n5307 );
nand ( n5423 , n5422 , n5310 );
not ( n5424 , n5423 );
not ( n5425 , n5424 );
and ( n5426 , n48 , n67 );
not ( n5427 , n48 );
and ( n5428 , n5427 , n5125 );
nor ( n5429 , n5426 , n5428 );
not ( n5430 , n5429 );
not ( n5431 , n5430 );
not ( n5432 , n5183 );
or ( n5433 , n5431 , n5432 );
nand ( n5434 , n3381 , n5290 );
nand ( n5435 , n5433 , n5434 );
not ( n5436 , n5435 );
and ( n5437 , n48 , n65 );
not ( n5438 , n48 );
and ( n5439 , n5438 , n5294 );
nor ( n5440 , n5437 , n5439 );
and ( n5441 , n2905 , n5440 );
and ( n5442 , n2732 , n5328 );
nor ( n5443 , n5441 , n5442 );
not ( n5444 , n5443 );
or ( n5445 , n5436 , n5444 );
or ( n5446 , n5435 , n5443 );
nand ( n5447 , n5445 , n5446 );
not ( n5448 , n5447 );
or ( n5449 , n5425 , n5448 );
not ( n5450 , n5443 );
nand ( n5451 , n5450 , n5435 );
nand ( n5452 , n5449 , n5451 );
xnor ( n5453 , n5299 , n5310 );
not ( n5454 , n5453 );
not ( n5455 , n5340 );
or ( n5456 , n5454 , n5455 );
or ( n5457 , n5453 , n5340 );
nand ( n5458 , n5456 , n5457 );
or ( n5459 , n5452 , n5458 );
xor ( n5460 , n48 , n66 );
not ( n5461 , n5460 );
not ( n5462 , n2745 );
or ( n5463 , n5461 , n5462 );
nand ( n5464 , n2732 , n5440 );
nand ( n5465 , n5463 , n5464 );
not ( n5466 , n5465 );
not ( n5467 , n51 );
nor ( n5468 , n5467 , n50 );
nand ( n5469 , n5468 , n63 );
not ( n5470 , n51 );
nand ( n5471 , n5470 , n50 , n4951 );
nand ( n5472 , n3430 , n5300 );
nand ( n5473 , n5469 , n5471 , n5472 );
and ( n5474 , n2980 , n67 );
nor ( n5475 , n5473 , n5474 );
not ( n5476 , n5475 );
nand ( n5477 , n5473 , n5474 );
nand ( n5478 , n5476 , n5477 );
or ( n5479 , n5466 , n5478 );
nand ( n5480 , n5479 , n5477 );
not ( n5481 , n5424 );
not ( n5482 , n5447 );
not ( n5483 , n5482 );
or ( n5484 , n5481 , n5483 );
nand ( n5485 , n5423 , n5447 );
nand ( n5486 , n5484 , n5485 );
xor ( n5487 , n5480 , n5486 );
and ( n5488 , n64 , n5468 );
not ( n5489 , n64 );
and ( n5490 , n5489 , n3430 );
nor ( n5491 , n5488 , n5490 );
nand ( n5492 , n2794 , n5294 );
and ( n5493 , n5491 , n5492 );
not ( n5494 , n67 );
nand ( n5495 , n1363 , n1490 );
not ( n5496 , n5495 );
or ( n5497 , n5494 , n5496 );
nand ( n5498 , n5497 , n3108 );
nor ( n5499 , n5493 , n5498 );
buf ( n5500 , n5499 );
not ( n5501 , n5500 );
not ( n5502 , n5478 );
not ( n5503 , n5465 );
and ( n5504 , n5502 , n5503 );
and ( n5505 , n5465 , n5478 );
nor ( n5506 , n5504 , n5505 );
not ( n5507 , n5506 );
not ( n5508 , n5507 );
or ( n5509 , n5501 , n5508 );
not ( n5510 , n5500 );
not ( n5511 , n5506 );
or ( n5512 , n5510 , n5511 );
or ( n5513 , n5500 , n5506 );
nand ( n5514 , n5512 , n5513 );
and ( n5515 , n2905 , n5429 );
and ( n5516 , n48 , n66 );
nor ( n5517 , n48 , n66 );
nor ( n5518 , n5516 , n5517 );
and ( n5519 , n2732 , n5518 );
nor ( n5520 , n5515 , n5519 );
not ( n5521 , n67 );
not ( n5522 , n3607 );
or ( n5523 , n5521 , n5522 );
not ( n5524 , n5294 );
not ( n5525 , n51 );
nor ( n5526 , n5525 , n50 );
not ( n5527 , n5526 );
or ( n5528 , n5524 , n5527 );
not ( n5529 , n67 );
not ( n5530 , n51 );
or ( n5531 , n5529 , n5530 );
not ( n5532 , n66 );
nand ( n5533 , n5532 , n50 );
nand ( n5534 , n5531 , n5533 );
nand ( n5535 , n5528 , n5534 );
nor ( n5536 , n3060 , n5294 );
nor ( n5537 , n5535 , n5536 );
nand ( n5538 , n5523 , n5537 );
and ( n5539 , n5520 , n5538 );
not ( n5540 , n5499 );
nand ( n5541 , n5498 , n5493 );
nand ( n5542 , n5540 , n5541 );
or ( n5543 , n5539 , n5542 );
buf ( n5544 , n5538 );
or ( n5545 , n5520 , n5544 );
nand ( n5546 , n5543 , n5545 );
nand ( n5547 , n5514 , n5546 );
nand ( n5548 , n5509 , n5547 );
and ( n5549 , n5487 , n5548 );
and ( n5550 , n5480 , n5486 );
or ( n5551 , n5549 , n5550 );
not ( n5552 , n5551 );
xor ( n5553 , n5452 , n5458 );
nand ( n5554 , n5552 , n5553 );
nand ( n5555 , n5459 , n5554 );
nand ( n5556 , n5421 , n5555 );
nand ( n5557 , n5420 , n5556 );
not ( n5558 , n5557 );
not ( n5559 , n5376 );
and ( n5560 , n5559 , n5416 );
nor ( n5561 , n5371 , n5351 );
nor ( n5562 , n5560 , n5561 );
not ( n5563 , n5562 );
not ( n5564 , n3363 );
and ( n5565 , n5564 , n5393 );
and ( n5566 , n48 , n61 );
not ( n5567 , n48 );
and ( n5568 , n5567 , n4653 );
nor ( n5569 , n5566 , n5568 );
and ( n5570 , n2824 , n5569 );
nor ( n5571 , n5565 , n5570 );
not ( n5572 , n5384 );
not ( n5573 , n2699 );
or ( n5574 , n5572 , n5573 );
and ( n5575 , n916 , n5300 );
and ( n5576 , n46 , n63 );
nor ( n5577 , n5575 , n5576 );
nand ( n5578 , n3381 , n5577 );
nand ( n5579 , n5574 , n5578 );
not ( n5580 , n5579 );
not ( n5581 , n5370 );
or ( n5582 , n5580 , n5581 );
or ( n5583 , n5579 , n5370 );
nand ( n5584 , n5582 , n5583 );
xnor ( n5585 , n5571 , n5584 );
not ( n5586 , n5585 );
nand ( n5587 , n3216 , n59 );
nand ( n5588 , n2794 , n4595 );
nand ( n5589 , n3061 , n4750 );
and ( n5590 , n5587 , n5588 , n5589 );
not ( n5591 , n5590 );
and ( n5592 , n2713 , n67 );
not ( n5593 , n5592 );
and ( n5594 , n5591 , n5593 );
and ( n5595 , n5590 , n5592 );
nor ( n5596 , n5594 , n5595 );
and ( n5597 , n2581 , n5405 );
and ( n5598 , n44 , n65 );
nor ( n5599 , n44 , n65 );
nor ( n5600 , n5598 , n5599 );
and ( n5601 , n2587 , n5600 );
nor ( n5602 , n5597 , n5601 );
and ( n5603 , n5596 , n5602 );
not ( n5604 , n5596 );
not ( n5605 , n5602 );
and ( n5606 , n5604 , n5605 );
nor ( n5607 , n5603 , n5606 );
not ( n5608 , n5408 );
not ( n5609 , n5396 );
or ( n5610 , n5608 , n5609 );
nand ( n5611 , n5386 , n5395 );
nand ( n5612 , n5610 , n5611 );
xor ( n5613 , n5607 , n5612 );
not ( n5614 , n5613 );
not ( n5615 , n5614 );
or ( n5616 , n5586 , n5615 );
not ( n5617 , n5585 );
nand ( n5618 , n5617 , n5613 );
nand ( n5619 , n5616 , n5618 );
not ( n5620 , n5619 );
or ( n5621 , n5563 , n5620 );
or ( n5622 , n5619 , n5562 );
nand ( n5623 , n5621 , n5622 );
and ( n5624 , n5613 , n5585 );
and ( n5625 , n5607 , n5612 );
nor ( n5626 , n5624 , n5625 );
not ( n5627 , n5626 );
not ( n5628 , n5584 );
or ( n5629 , n5628 , n5571 );
not ( n5630 , n5579 );
or ( n5631 , n5630 , n5370 );
nand ( n5632 , n5629 , n5631 );
not ( n5633 , n5632 );
not ( n5634 , n5633 );
or ( n5635 , n5596 , n5602 );
not ( n5636 , n5590 );
nand ( n5637 , n5636 , n5592 );
nand ( n5638 , n5635 , n5637 );
not ( n5639 , n5638 );
not ( n5640 , n5569 );
not ( n5641 , n5114 );
or ( n5642 , n5640 , n5641 );
and ( n5643 , n48 , n60 );
not ( n5644 , n48 );
and ( n5645 , n5644 , n4595 );
nor ( n5646 , n5643 , n5645 );
nand ( n5647 , n2732 , n5646 );
nand ( n5648 , n5642 , n5647 );
not ( n5649 , n5125 );
not ( n5650 , n3273 );
or ( n5651 , n5649 , n5650 );
nand ( n5652 , n5651 , n2719 );
nor ( n5653 , n5648 , n5652 );
not ( n5654 , n5653 );
nand ( n5655 , n5648 , n5652 );
nand ( n5656 , n5654 , n5655 );
not ( n5657 , n5656 );
not ( n5658 , n5577 );
not ( n5659 , n2869 );
or ( n5660 , n5658 , n5659 );
and ( n5661 , n916 , n4935 );
and ( n5662 , n46 , n62 );
nor ( n5663 , n5661 , n5662 );
nand ( n5664 , n2982 , n5663 );
nand ( n5665 , n5660 , n5664 );
not ( n5666 , n5665 );
and ( n5667 , n5657 , n5666 );
and ( n5668 , n5656 , n5665 );
nor ( n5669 , n5667 , n5668 );
not ( n5670 , n5669 );
or ( n5671 , n5639 , n5670 );
or ( n5672 , n5638 , n5669 );
nand ( n5673 , n5671 , n5672 );
not ( n5674 , n5673 );
not ( n5675 , n4750 );
not ( n5676 , n2795 );
or ( n5677 , n5675 , n5676 );
and ( n5678 , n58 , n3216 );
not ( n5679 , n58 );
and ( n5680 , n5679 , n3061 );
nor ( n5681 , n5678 , n5680 );
nand ( n5682 , n5677 , n5681 );
not ( n5683 , n5401 );
not ( n5684 , n5683 );
not ( n5685 , n4845 );
or ( n5686 , n5684 , n5685 );
not ( n5687 , n42 );
not ( n5688 , n66 );
and ( n5689 , n5687 , n5688 );
and ( n5690 , n42 , n66 );
nor ( n5691 , n5689 , n5690 );
nand ( n5692 , n2713 , n5691 );
nand ( n5693 , n5686 , n5692 );
xor ( n5694 , n5682 , n5693 );
not ( n5695 , n5694 );
and ( n5696 , n2581 , n5600 );
and ( n5697 , n44 , n64 );
not ( n5698 , n44 );
and ( n5699 , n5698 , n4951 );
nor ( n5700 , n5697 , n5699 );
and ( n5701 , n2632 , n5700 );
nor ( n5702 , n5696 , n5701 );
not ( n5703 , n5702 );
and ( n5704 , n5695 , n5703 );
and ( n5705 , n5694 , n5702 );
nor ( n5706 , n5704 , n5705 );
not ( n5707 , n5706 );
and ( n5708 , n5674 , n5707 );
and ( n5709 , n5673 , n5706 );
nor ( n5710 , n5708 , n5709 );
not ( n5711 , n5710 );
not ( n5712 , n5711 );
or ( n5713 , n5634 , n5712 );
nand ( n5714 , n5710 , n5632 );
nand ( n5715 , n5713 , n5714 );
nand ( n5716 , n5627 , n5715 );
and ( n5717 , n5623 , n5716 );
not ( n5718 , n5717 );
or ( n5719 , n5558 , n5718 );
not ( n5720 , n5716 );
not ( n5721 , n5619 );
nand ( n5722 , n5721 , n5562 );
nor ( n5723 , n5720 , n5722 );
not ( n5724 , n5626 );
nor ( n5725 , n5724 , n5715 );
nor ( n5726 , n5723 , n5725 );
nand ( n5727 , n5719 , n5726 );
not ( n5728 , n5663 );
not ( n5729 , n5183 );
or ( n5730 , n5728 , n5729 );
not ( n5731 , n46 );
not ( n5732 , n61 );
and ( n5733 , n5731 , n5732 );
and ( n5734 , n46 , n61 );
nor ( n5735 , n5733 , n5734 );
nand ( n5736 , n3381 , n5735 );
nand ( n5737 , n5730 , n5736 );
not ( n5738 , n5737 );
buf ( n5739 , n5526 );
and ( n5740 , n5739 , n57 );
and ( n5741 , n3705 , n4630 );
nor ( n5742 , n5740 , n5741 );
nand ( n5743 , n2795 , n4701 );
and ( n5744 , n5742 , n5743 );
not ( n5745 , n5744 );
or ( n5746 , n5738 , n5745 );
or ( n5747 , n5737 , n5744 );
nand ( n5748 , n5746 , n5747 );
and ( n5749 , n2722 , n5691 );
and ( n5750 , n42 , n65 );
not ( n5751 , n42 );
and ( n5752 , n5751 , n5294 );
nor ( n5753 , n5750 , n5752 );
and ( n5754 , n2715 , n5753 );
nor ( n5755 , n5749 , n5754 );
not ( n5756 , n5755 );
and ( n5757 , n5748 , n5756 );
not ( n5758 , n5748 );
and ( n5759 , n5758 , n5755 );
nor ( n5760 , n5757 , n5759 );
not ( n5761 , n5638 );
not ( n5762 , n5669 );
not ( n5763 , n5762 );
or ( n5764 , n5761 , n5763 );
not ( n5765 , n5656 );
nand ( n5766 , n5765 , n5665 );
nand ( n5767 , n5764 , n5766 );
xor ( n5768 , n5760 , n5767 );
not ( n5769 , n5768 );
not ( n5770 , n5646 );
not ( n5771 , n2905 );
or ( n5772 , n5770 , n5771 );
not ( n5773 , n48 );
not ( n5774 , n59 );
and ( n5775 , n5773 , n5774 );
and ( n5776 , n48 , n59 );
nor ( n5777 , n5775 , n5776 );
nand ( n5778 , n2732 , n5777 );
nand ( n5779 , n5772 , n5778 );
xor ( n5780 , n5655 , n5779 );
not ( n5781 , n5700 );
not ( n5782 , n3396 );
or ( n5783 , n5781 , n5782 );
and ( n5784 , n44 , n63 );
not ( n5785 , n44 );
and ( n5786 , n5785 , n5300 );
nor ( n5787 , n5784 , n5786 );
nand ( n5788 , n2585 , n5787 );
nand ( n5789 , n5783 , n5788 );
not ( n5790 , n5789 );
nand ( n5791 , n3742 , n67 );
not ( n5792 , n5791 );
and ( n5793 , n5790 , n5792 );
and ( n5794 , n5789 , n5791 );
nor ( n5795 , n5793 , n5794 );
xor ( n5796 , n5780 , n5795 );
not ( n5797 , n5693 );
not ( n5798 , n5682 );
or ( n5799 , n5797 , n5798 );
not ( n5800 , n5702 );
nand ( n5801 , n5800 , n5694 );
nand ( n5802 , n5799 , n5801 );
not ( n5803 , n5802 );
and ( n5804 , n5796 , n5803 );
not ( n5805 , n5796 );
and ( n5806 , n5805 , n5802 );
nor ( n5807 , n5804 , n5806 );
not ( n5808 , n5807 );
and ( n5809 , n5769 , n5808 );
buf ( n5810 , n5807 );
and ( n5811 , n5768 , n5810 );
nor ( n5812 , n5809 , n5811 );
not ( n5813 , n5673 );
not ( n5814 , n5813 );
not ( n5815 , n5706 );
and ( n5816 , n5814 , n5815 );
and ( n5817 , n5711 , n5632 );
nor ( n5818 , n5816 , n5817 );
xor ( n5819 , n5812 , n5818 );
nand ( n5820 , n5727 , n5819 );
not ( n5821 , n5779 );
or ( n5822 , n5795 , n5821 );
not ( n5823 , n5791 );
nand ( n5824 , n5823 , n5789 );
nand ( n5825 , n5822 , n5824 );
not ( n5826 , n5756 );
not ( n5827 , n5748 );
or ( n5828 , n5826 , n5827 );
not ( n5829 , n5744 );
nand ( n5830 , n5829 , n5737 );
nand ( n5831 , n5828 , n5830 );
xor ( n5832 , n5825 , n5831 );
and ( n5833 , n56 , n3216 );
not ( n5834 , n4630 );
not ( n5835 , n2795 );
or ( n5836 , n5834 , n5835 );
nand ( n5837 , n3705 , n4585 );
nand ( n5838 , n5836 , n5837 );
nor ( n5839 , n5833 , n5838 );
not ( n5840 , n5839 );
not ( n5841 , n5787 );
not ( n5842 , n2581 );
or ( n5843 , n5841 , n5842 );
and ( n5844 , n44 , n62 );
not ( n5845 , n44 );
and ( n5846 , n5845 , n4935 );
nor ( n5847 , n5844 , n5846 );
nand ( n5848 , n2587 , n5847 );
nand ( n5849 , n5843 , n5848 );
not ( n5850 , n5849 );
and ( n5851 , n5840 , n5850 );
and ( n5852 , n5839 , n5849 );
nor ( n5853 , n5851 , n5852 );
and ( n5854 , n2722 , n5753 );
and ( n5855 , n42 , n64 );
not ( n5856 , n42 );
and ( n5857 , n5856 , n4951 );
nor ( n5858 , n5855 , n5857 );
and ( n5859 , n3007 , n5858 );
nor ( n5860 , n5854 , n5859 );
xor ( n5861 , n5853 , n5860 );
xnor ( n5862 , n5832 , n5861 );
not ( n5863 , n5802 );
not ( n5864 , n5796 );
or ( n5865 , n5863 , n5864 );
not ( n5866 , n5655 );
and ( n5867 , n5795 , n5821 );
not ( n5868 , n5795 );
and ( n5869 , n5868 , n5779 );
nor ( n5870 , n5867 , n5869 );
nand ( n5871 , n5866 , n5870 );
nand ( n5872 , n5865 , n5871 );
not ( n5873 , n5872 );
and ( n5874 , n5125 , n40 );
and ( n5875 , n42 , n67 );
nor ( n5876 , n5874 , n5875 );
not ( n5877 , n5876 );
nand ( n5878 , n5877 , n2541 );
and ( n5879 , n5287 , n427 );
and ( n5880 , n40 , n66 );
nor ( n5881 , n5879 , n5880 );
nand ( n5882 , n2550 , n5881 );
and ( n5883 , n5878 , n5882 );
not ( n5884 , n5735 );
not ( n5885 , n3037 );
or ( n5886 , n5884 , n5885 );
not ( n5887 , n46 );
not ( n5888 , n60 );
and ( n5889 , n5887 , n5888 );
and ( n5890 , n46 , n60 );
nor ( n5891 , n5889 , n5890 );
nand ( n5892 , n3381 , n5891 );
nand ( n5893 , n5886 , n5892 );
xnor ( n5894 , n5883 , n5893 );
not ( n5895 , n5777 );
not ( n5896 , n2747 );
or ( n5897 , n5895 , n5896 );
and ( n5898 , n48 , n58 );
not ( n5899 , n48 );
and ( n5900 , n5899 , n4701 );
nor ( n5901 , n5898 , n5900 );
nand ( n5902 , n2732 , n5901 );
nand ( n5903 , n5897 , n5902 );
not ( n5904 , n5903 );
and ( n5905 , n5791 , n3804 );
not ( n5906 , n5905 );
and ( n5907 , n5904 , n5906 );
and ( n5908 , n5903 , n5905 );
nor ( n5909 , n5907 , n5908 );
xnor ( n5910 , n5894 , n5909 );
not ( n5911 , n5910 );
and ( n5912 , n5873 , n5911 );
and ( n5913 , n5872 , n5910 );
nor ( n5914 , n5912 , n5913 );
xnor ( n5915 , n5862 , n5914 );
not ( n5916 , n5810 );
and ( n5917 , n5916 , n5768 );
and ( n5918 , n5767 , n5760 );
nor ( n5919 , n5917 , n5918 );
and ( n5920 , n5915 , n5919 );
nand ( n5921 , n5812 , n5818 );
not ( n5922 , n5921 );
nor ( n5923 , n5920 , n5922 );
nand ( n5924 , n5820 , n5923 );
or ( n5925 , n5914 , n5862 );
not ( n5926 , n5872 );
or ( n5927 , n5926 , n5910 );
nand ( n5928 , n5925 , n5927 );
not ( n5929 , n5928 );
nand ( n5930 , n5832 , n5861 );
nand ( n5931 , n5831 , n5825 );
and ( n5932 , n5930 , n5931 );
or ( n5933 , n5853 , n5860 );
not ( n5934 , n5849 );
or ( n5935 , n5934 , n5839 );
nand ( n5936 , n5933 , n5935 );
and ( n5937 , n2870 , n5891 );
and ( n5938 , n916 , n4750 );
and ( n5939 , n46 , n59 );
nor ( n5940 , n5938 , n5939 );
and ( n5941 , n3381 , n5940 );
nor ( n5942 , n5937 , n5941 );
xnor ( n5943 , n5942 , n5908 );
not ( n5944 , n5943 );
and ( n5945 , n5936 , n5944 );
not ( n5946 , n5936 );
and ( n5947 , n5946 , n5943 );
nor ( n5948 , n5945 , n5947 );
and ( n5949 , n5932 , n5948 );
not ( n5950 , n5932 );
not ( n5951 , n5948 );
and ( n5952 , n5950 , n5951 );
nor ( n5953 , n5949 , n5952 );
nand ( n5954 , n2562 , n67 );
and ( n5955 , n2905 , n5901 );
and ( n5956 , n48 , n57 );
not ( n5957 , n48 );
and ( n5958 , n5957 , n4630 );
nor ( n5959 , n5956 , n5958 );
and ( n5960 , n2823 , n5959 );
nor ( n5961 , n5955 , n5960 );
xor ( n5962 , n5954 , n5961 );
and ( n5963 , n2581 , n5847 );
and ( n5964 , n968 , n4653 );
and ( n5965 , n44 , n61 );
nor ( n5966 , n5964 , n5965 );
and ( n5967 , n2587 , n5966 );
nor ( n5968 , n5963 , n5967 );
not ( n5969 , n5968 );
and ( n5970 , n5962 , n5969 );
not ( n5971 , n5962 );
and ( n5972 , n5971 , n5968 );
nor ( n5973 , n5970 , n5972 );
and ( n5974 , n2541 , n5881 );
and ( n5975 , n40 , n65 );
not ( n5976 , n40 );
and ( n5977 , n5976 , n5294 );
nor ( n5978 , n5975 , n5977 );
and ( n5979 , n2550 , n5978 );
nor ( n5980 , n5974 , n5979 );
nand ( n5981 , n5739 , n55 );
nand ( n5982 , n3325 , n4585 );
nand ( n5983 , n3061 , n4577 );
and ( n5984 , n5981 , n5982 , n5983 );
not ( n5985 , n5984 );
not ( n5986 , n5858 );
not ( n5987 , n4845 );
or ( n5988 , n5986 , n5987 );
xor ( n5989 , n63 , n42 );
nand ( n5990 , n2713 , n5989 );
nand ( n5991 , n5988 , n5990 );
not ( n5992 , n5991 );
or ( n5993 , n5985 , n5992 );
or ( n5994 , n5991 , n5984 );
nand ( n5995 , n5993 , n5994 );
xnor ( n5996 , n5980 , n5995 );
xor ( n5997 , n5973 , n5996 );
not ( n5998 , n5909 );
not ( n5999 , n5894 );
or ( n6000 , n5998 , n5999 );
not ( n6001 , n5893 );
or ( n6002 , n6001 , n5883 );
nand ( n6003 , n6000 , n6002 );
xnor ( n6004 , n5997 , n6003 );
xor ( n6005 , n5953 , n6004 );
not ( n6006 , n6005 );
or ( n6007 , n5929 , n6006 );
or ( n6008 , n5928 , n6005 );
nand ( n6009 , n6007 , n6008 );
or ( n6010 , n5915 , n5919 );
nand ( n6011 , n5924 , n6009 , n6010 );
not ( n6012 , n6004 );
not ( n6013 , n5953 );
or ( n6014 , n6012 , n6013 );
nand ( n6015 , n5932 , n5948 );
nand ( n6016 , n6014 , n6015 );
nand ( n6017 , n5954 , n3991 );
not ( n6018 , n6017 );
nand ( n6019 , n5739 , n54 );
nand ( n6020 , n3471 , n4577 );
not ( n6021 , n54 );
nand ( n6022 , n3061 , n6021 );
nand ( n6023 , n6019 , n6020 , n6022 );
not ( n6024 , n6023 );
not ( n6025 , n6024 );
or ( n6026 , n6018 , n6025 );
not ( n6027 , n6017 );
nand ( n6028 , n6027 , n6023 );
nand ( n6029 , n6026 , n6028 );
and ( n6030 , n5962 , n5968 );
and ( n6031 , n5954 , n5961 );
nor ( n6032 , n6030 , n6031 );
xnor ( n6033 , n6029 , n6032 );
not ( n6034 , n5991 );
or ( n6035 , n6034 , n5984 );
not ( n6036 , n5980 );
nand ( n6037 , n6036 , n5995 );
nand ( n6038 , n6035 , n6037 );
not ( n6039 , n6038 );
and ( n6040 , n6033 , n6039 );
not ( n6041 , n6033 );
and ( n6042 , n6041 , n6038 );
nor ( n6043 , n6040 , n6042 );
and ( n6044 , n6003 , n5997 );
and ( n6045 , n5973 , n5996 );
nor ( n6046 , n6044 , n6045 );
xor ( n6047 , n6043 , n6046 );
not ( n6048 , n5940 );
not ( n6049 , n2869 );
or ( n6050 , n6048 , n6049 );
and ( n6051 , n916 , n4701 );
and ( n6052 , n46 , n58 );
nor ( n6053 , n6051 , n6052 );
nand ( n6054 , n2982 , n6053 );
nand ( n6055 , n6050 , n6054 );
not ( n6056 , n6055 );
nand ( n6057 , n3042 , n5978 );
and ( n6058 , n40 , n64 );
not ( n6059 , n40 );
and ( n6060 , n6059 , n4951 );
nor ( n6061 , n6058 , n6060 );
nand ( n6062 , n2549 , n6061 );
and ( n6063 , n6057 , n6062 );
not ( n6064 , n6063 );
and ( n6065 , n6056 , n6064 );
and ( n6066 , n6055 , n6063 );
nor ( n6067 , n6065 , n6066 );
and ( n6068 , n2564 , n5127 );
not ( n6069 , n3870 );
not ( n6070 , n38 );
not ( n6071 , n66 );
and ( n6072 , n6070 , n6071 );
and ( n6073 , n38 , n66 );
nor ( n6074 , n6072 , n6073 );
and ( n6075 , n6069 , n6074 );
nor ( n6076 , n6068 , n6075 );
and ( n6077 , n6067 , n6076 );
not ( n6078 , n6067 );
not ( n6079 , n6076 );
and ( n6080 , n6078 , n6079 );
nor ( n6081 , n6077 , n6080 );
not ( n6082 , n6081 );
and ( n6083 , n2905 , n5959 );
and ( n6084 , n48 , n56 );
not ( n6085 , n48 );
and ( n6086 , n6085 , n4585 );
nor ( n6087 , n6084 , n6086 );
and ( n6088 , n2732 , n6087 );
nor ( n6089 , n6083 , n6088 );
and ( n6090 , n4845 , n5989 );
and ( n6091 , n42 , n62 );
nor ( n6092 , n42 , n62 );
nor ( n6093 , n6091 , n6092 );
and ( n6094 , n2713 , n6093 );
nor ( n6095 , n6090 , n6094 );
and ( n6096 , n6089 , n6095 );
not ( n6097 , n6089 );
not ( n6098 , n6095 );
and ( n6099 , n6097 , n6098 );
nor ( n6100 , n6096 , n6099 );
and ( n6101 , n2581 , n5966 );
xor ( n6102 , n44 , n60 );
and ( n6103 , n2631 , n6102 );
nor ( n6104 , n6101 , n6103 );
not ( n6105 , n6104 );
and ( n6106 , n6100 , n6105 );
not ( n6107 , n6100 );
and ( n6108 , n6107 , n6104 );
or ( n6109 , n6106 , n6108 );
not ( n6110 , n6109 );
or ( n6111 , n6082 , n6110 );
or ( n6112 , n6081 , n6109 );
nand ( n6113 , n6111 , n6112 );
not ( n6114 , n5943 );
not ( n6115 , n5936 );
or ( n6116 , n6114 , n6115 );
not ( n6117 , n5942 );
nand ( n6118 , n6117 , n5908 );
nand ( n6119 , n6116 , n6118 );
xnor ( n6120 , n6113 , n6119 );
xor ( n6121 , n6047 , n6120 );
nand ( n6122 , n6016 , n6121 );
xor ( n6123 , n6043 , n6046 );
and ( n6124 , n6123 , n6120 );
and ( n6125 , n6043 , n6046 );
nor ( n6126 , n6124 , n6125 );
not ( n6127 , n6126 );
not ( n6128 , n5138 );
nand ( n6129 , n3705 , n4615 );
nand ( n6130 , n6021 , n3471 );
nand ( n6131 , n53 , n3216 );
nand ( n6132 , n6129 , n6130 , n6131 );
not ( n6133 , n6132 );
or ( n6134 , n6128 , n6133 );
not ( n6135 , n6132 );
not ( n6136 , n5138 );
nand ( n6137 , n6135 , n6136 );
nand ( n6138 , n6134 , n6137 );
and ( n6139 , n6087 , n2905 );
and ( n6140 , n2732 , n5110 );
nor ( n6141 , n6139 , n6140 );
xor ( n6142 , n6138 , n6141 );
not ( n6143 , n6142 );
not ( n6144 , n6100 );
not ( n6145 , n6105 );
or ( n6146 , n6144 , n6145 );
not ( n6147 , n6089 );
nand ( n6148 , n6147 , n6098 );
nand ( n6149 , n6146 , n6148 );
not ( n6150 , n6149 );
or ( n6151 , n6143 , n6150 );
or ( n6152 , n6142 , n6149 );
nand ( n6153 , n6151 , n6152 );
or ( n6154 , n6067 , n6076 );
not ( n6155 , n6055 );
or ( n6156 , n6155 , n6063 );
nand ( n6157 , n6154 , n6156 );
and ( n6158 , n6153 , n6157 );
not ( n6159 , n6153 );
not ( n6160 , n6157 );
and ( n6161 , n6159 , n6160 );
or ( n6162 , n6158 , n6161 );
nand ( n6163 , n6113 , n6119 );
not ( n6164 , n6109 );
nand ( n6165 , n6164 , n6081 );
and ( n6166 , n6163 , n6165 );
xor ( n6167 , n6162 , n6166 );
not ( n6168 , n6038 );
not ( n6169 , n6033 );
or ( n6170 , n6168 , n6169 );
not ( n6171 , n6029 );
nand ( n6172 , n6171 , n6032 );
nand ( n6173 , n6170 , n6172 );
not ( n6174 , n5169 );
not ( n6175 , n2549 );
or ( n6176 , n6174 , n6175 );
nand ( n6177 , n3042 , n6061 );
nand ( n6178 , n6176 , n6177 );
not ( n6179 , n6178 );
and ( n6180 , n4948 , n6074 );
not ( n6181 , n38 );
not ( n6182 , n65 );
and ( n6183 , n6181 , n6182 );
and ( n6184 , n38 , n65 );
nor ( n6185 , n6183 , n6184 );
and ( n6186 , n6069 , n6185 );
nor ( n6187 , n6180 , n6186 );
not ( n6188 , n6187 );
and ( n6189 , n6179 , n6188 );
and ( n6190 , n6178 , n6187 );
nor ( n6191 , n6189 , n6190 );
xor ( n6192 , n6028 , n6191 );
and ( n6193 , n2581 , n6102 );
and ( n6194 , n2631 , n5102 );
nor ( n6195 , n6193 , n6194 );
not ( n6196 , n6195 );
not ( n6197 , n6053 );
not ( n6198 , n5183 );
or ( n6199 , n6197 , n6198 );
nand ( n6200 , n2982 , n5177 );
nand ( n6201 , n6199 , n6200 );
not ( n6202 , n6201 );
or ( n6203 , n6196 , n6202 );
or ( n6204 , n6201 , n6195 );
nand ( n6205 , n6203 , n6204 );
not ( n6206 , n6205 );
and ( n6207 , n2987 , n6093 );
and ( n6208 , n2715 , n5160 );
nor ( n6209 , n6207 , n6208 );
not ( n6210 , n6209 );
and ( n6211 , n6206 , n6210 );
and ( n6212 , n6205 , n6209 );
nor ( n6213 , n6211 , n6212 );
xnor ( n6214 , n6192 , n6213 );
xor ( n6215 , n6173 , n6214 );
not ( n6216 , n6215 );
xor ( n6217 , n6167 , n6216 );
nand ( n6218 , n6127 , n6217 );
not ( n6219 , n5928 );
nand ( n6220 , n6219 , n6005 );
and ( n6221 , n6122 , n6218 , n6220 );
nand ( n6222 , n6011 , n6221 );
not ( n6223 , n6126 );
not ( n6224 , n6217 );
or ( n6225 , n6223 , n6224 );
buf ( n6226 , n6126 );
or ( n6227 , n6217 , n6226 );
nand ( n6228 , n6225 , n6227 );
not ( n6229 , n6121 );
not ( n6230 , n6016 );
nand ( n6231 , n6229 , n6230 );
nand ( n6232 , n6228 , n6231 );
buf ( n6233 , n6218 );
and ( n6234 , n6232 , n6233 );
not ( n6235 , n6173 );
not ( n6236 , n6214 );
or ( n6237 , n6235 , n6236 );
not ( n6238 , n6213 );
nand ( n6239 , n6238 , n6192 );
nand ( n6240 , n6237 , n6239 );
not ( n6241 , n6201 );
or ( n6242 , n6241 , n6195 );
not ( n6243 , n6209 );
nand ( n6244 , n6243 , n6205 );
nand ( n6245 , n6242 , n6244 );
not ( n6246 , n5163 );
not ( n6247 , n5191 );
or ( n6248 , n6246 , n6247 );
or ( n6249 , n5191 , n5163 );
nand ( n6250 , n6248 , n6249 );
xor ( n6251 , n5132 , n5105 );
nor ( n6252 , n6250 , n6251 );
not ( n6253 , n6252 );
nand ( n6254 , n6250 , n6251 );
nand ( n6255 , n6253 , n6254 );
xor ( n6256 , n6245 , n6255 );
and ( n6257 , n6240 , n6256 );
not ( n6258 , n6240 );
not ( n6259 , n6256 );
and ( n6260 , n6258 , n6259 );
nor ( n6261 , n6257 , n6260 );
not ( n6262 , n6136 );
not ( n6263 , n6132 );
or ( n6264 , n6262 , n6263 );
not ( n6265 , n6141 );
nand ( n6266 , n6265 , n6138 );
nand ( n6267 , n6264 , n6266 );
not ( n6268 , n6267 );
not ( n6269 , n6268 );
not ( n6270 , n5148 );
nand ( n6271 , n5139 , n5147 );
nand ( n6272 , n6270 , n6271 );
not ( n6273 , n6272 );
and ( n6274 , n38 , n64 );
not ( n6275 , n38 );
and ( n6276 , n6275 , n4951 );
or ( n6277 , n6274 , n6276 );
or ( n6278 , n6277 , n2926 );
nand ( n6279 , n4948 , n6185 );
nand ( n6280 , n6278 , n6279 );
not ( n6281 , n6280 );
and ( n6282 , n6273 , n6281 );
and ( n6283 , n6272 , n6280 );
nor ( n6284 , n6282 , n6283 );
not ( n6285 , n6284 );
not ( n6286 , n6285 );
or ( n6287 , n6269 , n6286 );
nand ( n6288 , n6284 , n6267 );
nand ( n6289 , n6287 , n6288 );
or ( n6290 , n6191 , n6028 );
not ( n6291 , n6178 );
or ( n6292 , n6291 , n6187 );
nand ( n6293 , n6290 , n6292 );
and ( n6294 , n6289 , n6293 );
not ( n6295 , n6289 );
not ( n6296 , n6293 );
and ( n6297 , n6295 , n6296 );
nor ( n6298 , n6294 , n6297 );
not ( n6299 , n6157 );
not ( n6300 , n6153 );
or ( n6301 , n6299 , n6300 );
not ( n6302 , n6142 );
nand ( n6303 , n6302 , n6149 );
nand ( n6304 , n6301 , n6303 );
not ( n6305 , n6304 );
and ( n6306 , n6298 , n6305 );
not ( n6307 , n6298 );
and ( n6308 , n6307 , n6304 );
nor ( n6309 , n6306 , n6308 );
not ( n6310 , n6309 );
and ( n6311 , n6261 , n6310 );
not ( n6312 , n6261 );
and ( n6313 , n6312 , n6309 );
nor ( n6314 , n6311 , n6313 );
not ( n6315 , n6162 );
nor ( n6316 , n6315 , n6215 );
or ( n6317 , n6316 , n6166 );
or ( n6318 , n6216 , n6162 );
nand ( n6319 , n6317 , n6318 );
and ( n6320 , n6314 , n6319 );
nor ( n6321 , n6234 , n6320 );
nand ( n6322 , n6222 , n6321 );
not ( n6323 , n5277 );
and ( n6324 , n5239 , n6323 );
not ( n6325 , n5239 );
and ( n6326 , n6325 , n5277 );
nor ( n6327 , n6324 , n6326 );
xor ( n6328 , n5197 , n5097 );
not ( n6329 , n6250 );
not ( n6330 , n6329 );
not ( n6331 , n6251 );
and ( n6332 , n6330 , n6331 );
and ( n6333 , n6255 , n6245 );
nor ( n6334 , n6332 , n6333 );
not ( n6335 , n6334 );
not ( n6336 , n6335 );
or ( n6337 , n6268 , n6284 );
not ( n6338 , n6280 );
or ( n6339 , n6272 , n6338 );
nand ( n6340 , n6337 , n6339 );
buf ( n6341 , n6340 );
not ( n6342 , n6341 );
xor ( n6343 , n5156 , n5195 );
not ( n6344 , n6343 );
not ( n6345 , n6344 );
or ( n6346 , n6342 , n6345 );
not ( n6347 , n6340 );
nand ( n6348 , n6347 , n6343 );
nand ( n6349 , n6346 , n6348 );
not ( n6350 , n6349 );
or ( n6351 , n6336 , n6350 );
not ( n6352 , n6344 );
nand ( n6353 , n6352 , n6341 );
nand ( n6354 , n6351 , n6353 );
xor ( n6355 , n6328 , n6354 );
xor ( n6356 , n5259 , n5267 );
and ( n6357 , n6355 , n6356 );
and ( n6358 , n6328 , n6354 );
nor ( n6359 , n6357 , n6358 );
nand ( n6360 , n6327 , n6359 );
or ( n6361 , n6319 , n6314 );
nand ( n6362 , n6360 , n6361 );
and ( n6363 , n6349 , n6335 );
not ( n6364 , n6349 );
and ( n6365 , n6364 , n6334 );
or ( n6366 , n6363 , n6365 );
not ( n6367 , n6366 );
not ( n6368 , n6367 );
not ( n6369 , n6304 );
not ( n6370 , n6298 );
or ( n6371 , n6369 , n6370 );
nand ( n6372 , n6289 , n6293 );
nand ( n6373 , n6371 , n6372 );
xnor ( n6374 , n5254 , n5240 );
xnor ( n6375 , n6373 , n6374 );
not ( n6376 , n6375 );
or ( n6377 , n6368 , n6376 );
not ( n6378 , n6374 );
nand ( n6379 , n6378 , n6373 );
nand ( n6380 , n6377 , n6379 );
not ( n6381 , n6380 );
not ( n6382 , n6381 );
xnor ( n6383 , n6356 , n6355 );
not ( n6384 , n6383 );
or ( n6385 , n6382 , n6384 );
not ( n6386 , n6375 );
not ( n6387 , n6366 );
and ( n6388 , n6386 , n6387 );
and ( n6389 , n6375 , n6366 );
nor ( n6390 , n6388 , n6389 );
not ( n6391 , n6309 );
not ( n6392 , n6261 );
or ( n6393 , n6391 , n6392 );
or ( n6394 , n6240 , n6256 );
nand ( n6395 , n6393 , n6394 );
nand ( n6396 , n6390 , n6395 );
nand ( n6397 , n6385 , n6396 );
nor ( n6398 , n6362 , n6397 );
nand ( n6399 , n6322 , n6398 );
buf ( n6400 , n6360 );
xor ( n6401 , n6390 , n6395 );
or ( n6402 , n6397 , n6401 );
or ( n6403 , n6383 , n6381 );
nand ( n6404 , n6402 , n6403 );
and ( n6405 , n6400 , n6404 );
nor ( n6406 , n6327 , n6359 );
nor ( n6407 , n6405 , n6406 );
nand ( n6408 , n6399 , n6407 );
nand ( n6409 , n5286 , n6408 );
nand ( n6410 , n5283 , n6409 );
not ( n6411 , n6410 );
or ( n6412 , n5233 , n6411 );
or ( n6413 , n6410 , n5232 );
nand ( n6414 , n6412 , n6413 );
not ( n6415 , n2 );
and ( n6416 , n6415 , n1 );
nand ( n6417 , n6414 , n6416 );
or ( n6418 , n96 , n95 );
nand ( n6419 , n95 , n96 );
nand ( n6420 , n6418 , n6419 );
xor ( n6421 , n94 , n95 );
nand ( n6422 , n6420 , n6421 );
not ( n6423 , n6422 );
not ( n6424 , n94 );
not ( n6425 , n74 );
and ( n6426 , n6424 , n6425 );
and ( n6427 , n74 , n94 );
nor ( n6428 , n6426 , n6427 );
and ( n6429 , n6423 , n6428 );
not ( n6430 , n6420 );
not ( n6431 , n73 );
and ( n6432 , n6424 , n6431 );
and ( n6433 , n73 , n94 );
nor ( n6434 , n6432 , n6433 );
and ( n6435 , n6430 , n6434 );
nor ( n6436 , n6429 , n6435 );
xor ( n6437 , n86 , n87 );
not ( n6438 , n88 );
not ( n6439 , n6438 );
not ( n6440 , n87 );
not ( n6441 , n6440 );
or ( n6442 , n6439 , n6441 );
nand ( n6443 , n87 , n88 );
nand ( n6444 , n6442 , n6443 );
and ( n6445 , n6437 , n6444 );
not ( n6446 , n86 );
not ( n6447 , n82 );
and ( n6448 , n6446 , n6447 );
and ( n6449 , n82 , n86 );
nor ( n6450 , n6448 , n6449 );
and ( n6451 , n6445 , n6450 );
not ( n6452 , n6444 );
not ( n6453 , n81 );
and ( n6454 , n6453 , n6446 );
and ( n6455 , n81 , n86 );
nor ( n6456 , n6454 , n6455 );
and ( n6457 , n6452 , n6456 );
nor ( n6458 , n6451 , n6457 );
xor ( n6459 , n6436 , n6458 );
not ( n6460 , n93 );
not ( n6461 , n92 );
or ( n6462 , n6460 , n6461 );
or ( n6463 , n92 , n93 );
nand ( n6464 , n6462 , n6463 );
xor ( n6465 , n93 , n94 );
or ( n6466 , n6464 , n6465 );
not ( n6467 , n6466 );
not ( n6468 , n92 );
not ( n6469 , n76 );
and ( n6470 , n6468 , n6469 );
and ( n6471 , n76 , n92 );
nor ( n6472 , n6470 , n6471 );
and ( n6473 , n6467 , n6472 );
buf ( n6474 , n6465 );
not ( n6475 , n92 );
not ( n6476 , n75 );
and ( n6477 , n6475 , n6476 );
and ( n6478 , n75 , n92 );
nor ( n6479 , n6477 , n6478 );
and ( n6480 , n6474 , n6479 );
nor ( n6481 , n6473 , n6480 );
xor ( n6482 , n6459 , n6481 );
not ( n6483 , n96 );
nand ( n6484 , n6483 , n97 );
not ( n6485 , n6484 );
not ( n6486 , n97 );
nand ( n6487 , n6486 , n96 );
not ( n6488 , n6487 );
or ( n6489 , n6485 , n6488 );
and ( n6490 , n98 , n6486 );
not ( n6491 , n98 );
and ( n6492 , n6491 , n97 );
nor ( n6493 , n6490 , n6492 );
nand ( n6494 , n6489 , n6493 );
not ( n6495 , n6494 );
not ( n6496 , n72 );
and ( n6497 , n6483 , n6496 );
and ( n6498 , n72 , n96 );
nor ( n6499 , n6497 , n6498 );
and ( n6500 , n6495 , n6499 );
not ( n6501 , n6493 );
not ( n6502 , n71 );
and ( n6503 , n6483 , n6502 );
and ( n6504 , n71 , n96 );
nor ( n6505 , n6503 , n6504 );
and ( n6506 , n6501 , n6505 );
nor ( n6507 , n6500 , n6506 );
not ( n6508 , n6437 );
not ( n6509 , n6444 );
or ( n6510 , n6508 , n6509 );
nand ( n6511 , n6510 , n83 );
and ( n6512 , n6443 , n86 );
and ( n6513 , n6511 , n6512 );
nand ( n6514 , n6513 , n6 );
xor ( n6515 , n6507 , n6514 );
not ( n6516 , n91 );
nand ( n6517 , n6516 , n90 );
not ( n6518 , n6517 );
not ( n6519 , n90 );
nand ( n6520 , n6519 , n91 );
not ( n6521 , n6520 );
or ( n6522 , n6518 , n6521 );
xor ( n6523 , n91 , n92 );
buf ( n6524 , n6523 );
not ( n6525 , n6524 );
nand ( n6526 , n6522 , n6525 );
not ( n6527 , n6526 );
not ( n6528 , n90 );
not ( n6529 , n78 );
and ( n6530 , n6528 , n6529 );
and ( n6531 , n78 , n90 );
nor ( n6532 , n6530 , n6531 );
and ( n6533 , n6527 , n6532 );
not ( n6534 , n6525 );
not ( n6535 , n77 );
and ( n6536 , n6528 , n6535 );
and ( n6537 , n77 , n90 );
nor ( n6538 , n6536 , n6537 );
and ( n6539 , n6534 , n6538 );
nor ( n6540 , n6533 , n6539 );
xor ( n6541 , n6515 , n6540 );
xor ( n6542 , n6482 , n6541 );
or ( n6543 , n6513 , n6 );
nand ( n6544 , n6543 , n6514 );
not ( n6545 , n6544 );
not ( n6546 , n99 );
nand ( n6547 , n6546 , n98 );
or ( n6548 , n6547 , n71 );
nand ( n6549 , n98 , n99 );
or ( n6550 , n6549 , n70 );
not ( n6551 , n99 );
nor ( n6552 , n6551 , n98 );
not ( n6553 , n6552 );
not ( n6554 , n70 );
or ( n6555 , n6553 , n6554 );
nand ( n6556 , n6548 , n6550 , n6555 );
not ( n6557 , n6556 );
and ( n6558 , n6545 , n6557 );
and ( n6559 , n6544 , n6556 );
nor ( n6560 , n6558 , n6559 );
not ( n6561 , n83 );
and ( n6562 , n6561 , n6446 );
and ( n6563 , n83 , n86 );
nor ( n6564 , n6562 , n6563 );
and ( n6565 , n6445 , n6564 );
and ( n6566 , n6452 , n6450 );
nor ( n6567 , n6565 , n6566 );
or ( n6568 , n6560 , n6567 );
not ( n6569 , n6556 );
or ( n6570 , n6544 , n6569 );
nand ( n6571 , n6568 , n6570 );
not ( n6572 , n6571 );
and ( n6573 , n6542 , n6572 );
and ( n6574 , n6541 , n6482 );
nor ( n6575 , n6573 , n6574 );
or ( n6576 , n6547 , n70 );
or ( n6577 , n6549 , n69 );
not ( n6578 , n69 );
or ( n6579 , n6553 , n6578 );
nand ( n6580 , n6576 , n6577 , n6579 );
xor ( n6581 , n85 , n86 );
nand ( n6582 , n6581 , n83 );
not ( n6583 , n6582 );
xor ( n6584 , n6583 , n5 );
and ( n6585 , n6580 , n6584 );
and ( n6586 , n6583 , n5 );
nor ( n6587 , n6585 , n6586 );
not ( n6588 , n6587 );
xor ( n6589 , n6507 , n6514 );
and ( n6590 , n6589 , n6540 );
and ( n6591 , n6507 , n6514 );
nor ( n6592 , n6590 , n6591 );
not ( n6593 , n6592 );
or ( n6594 , n6588 , n6593 );
or ( n6595 , n6592 , n6587 );
nand ( n6596 , n6594 , n6595 );
xor ( n6597 , n6436 , n6458 );
and ( n6598 , n6597 , n6481 );
and ( n6599 , n6436 , n6458 );
nor ( n6600 , n6598 , n6599 );
xor ( n6601 , n6596 , n6600 );
xor ( n6602 , n6575 , n6601 );
xor ( n6603 , n6580 , n6584 );
not ( n6604 , n6603 );
and ( n6605 , n6424 , n6476 );
and ( n6606 , n75 , n94 );
nor ( n6607 , n6605 , n6606 );
and ( n6608 , n6423 , n6607 );
and ( n6609 , n6430 , n6428 );
nor ( n6610 , n6608 , n6609 );
and ( n6611 , n6475 , n6535 );
and ( n6612 , n77 , n92 );
nor ( n6613 , n6611 , n6612 );
and ( n6614 , n6467 , n6613 );
and ( n6615 , n6474 , n6472 );
nor ( n6616 , n6614 , n6615 );
xor ( n6617 , n6610 , n6616 );
and ( n6618 , n6483 , n6431 );
and ( n6619 , n73 , n96 );
nor ( n6620 , n6618 , n6619 );
and ( n6621 , n6495 , n6620 );
and ( n6622 , n6501 , n6499 );
nor ( n6623 , n6621 , n6622 );
and ( n6624 , n6617 , n6623 );
and ( n6625 , n6610 , n6616 );
nor ( n6626 , n6624 , n6625 );
not ( n6627 , n6626 );
or ( n6628 , n6604 , n6627 );
xnor ( n6629 , n6626 , n6603 );
not ( n6630 , n88 );
nand ( n6631 , n6630 , n89 );
not ( n6632 , n89 );
nand ( n6633 , n6632 , n88 );
and ( n6634 , n6631 , n6633 );
xor ( n6635 , n89 , n90 );
nor ( n6636 , n6634 , n6635 );
buf ( n6637 , n6636 );
buf ( n6638 , n6637 );
not ( n6639 , n80 );
and ( n6640 , n6639 , n6630 );
and ( n6641 , n80 , n88 );
nor ( n6642 , n6640 , n6641 );
and ( n6643 , n6638 , n6642 );
buf ( n6644 , n6635 );
not ( n6645 , n79 );
and ( n6646 , n6645 , n6630 );
and ( n6647 , n79 , n88 );
nor ( n6648 , n6646 , n6647 );
and ( n6649 , n6644 , n6648 );
nor ( n6650 , n6643 , n6649 );
or ( n6651 , n6629 , n6650 );
nand ( n6652 , n6628 , n6651 );
and ( n6653 , n6602 , n6652 );
and ( n6654 , n6575 , n6601 );
nor ( n6655 , n6653 , n6654 );
and ( n6656 , n6483 , n6554 );
and ( n6657 , n70 , n96 );
nor ( n6658 , n6656 , n6657 );
and ( n6659 , n6495 , n6658 );
and ( n6660 , n6483 , n6578 );
and ( n6661 , n69 , n96 );
nor ( n6662 , n6660 , n6661 );
and ( n6663 , n6501 , n6662 );
nor ( n6664 , n6659 , n6663 );
not ( n6665 , n6581 );
and ( n6666 , n85 , n84 );
not ( n6667 , n85 );
not ( n6668 , n84 );
and ( n6669 , n6667 , n6668 );
nor ( n6670 , n6666 , n6669 );
nand ( n6671 , n6665 , n6670 );
or ( n6672 , n82 , n84 );
nand ( n6673 , n82 , n84 );
nand ( n6674 , n6672 , n6673 );
or ( n6675 , n6671 , n6674 );
or ( n6676 , n81 , n84 );
nand ( n6677 , n81 , n84 );
nand ( n6678 , n6676 , n6677 );
or ( n6679 , n6678 , n6665 );
nand ( n6680 , n6675 , n6679 );
and ( n6681 , n6664 , n6680 );
not ( n6682 , n6664 );
not ( n6683 , n6680 );
and ( n6684 , n6682 , n6683 );
nor ( n6685 , n6681 , n6684 );
and ( n6686 , n6468 , n6425 );
and ( n6687 , n74 , n92 );
nor ( n6688 , n6686 , n6687 );
and ( n6689 , n6467 , n6688 );
and ( n6690 , n6468 , n6431 );
and ( n6691 , n73 , n92 );
nor ( n6692 , n6690 , n6691 );
and ( n6693 , n6474 , n6692 );
nor ( n6694 , n6689 , n6693 );
xnor ( n6695 , n6685 , n6694 );
nand ( n6696 , n85 , n86 );
and ( n6697 , n6696 , n84 );
and ( n6698 , n6582 , n6697 );
nand ( n6699 , n6698 , n4 );
and ( n6700 , n6424 , n6496 );
and ( n6701 , n72 , n94 );
nor ( n6702 , n6700 , n6701 );
and ( n6703 , n6423 , n6702 );
and ( n6704 , n6424 , n6502 );
and ( n6705 , n71 , n94 );
nor ( n6706 , n6704 , n6705 );
and ( n6707 , n6430 , n6706 );
nor ( n6708 , n6703 , n6707 );
xor ( n6709 , n6699 , n6708 );
and ( n6710 , n6528 , n6469 );
and ( n6711 , n76 , n90 );
nor ( n6712 , n6710 , n6711 );
and ( n6713 , n6527 , n6712 );
and ( n6714 , n6528 , n6476 );
and ( n6715 , n75 , n90 );
nor ( n6716 , n6714 , n6715 );
and ( n6717 , n6534 , n6716 );
nor ( n6718 , n6713 , n6717 );
xor ( n6719 , n6709 , n6718 );
xor ( n6720 , n6695 , n6719 );
and ( n6721 , n6639 , n6446 );
and ( n6722 , n80 , n86 );
nor ( n6723 , n6721 , n6722 );
and ( n6724 , n6445 , n6723 );
and ( n6725 , n6446 , n6645 );
and ( n6726 , n79 , n86 );
nor ( n6727 , n6725 , n6726 );
and ( n6728 , n6452 , n6727 );
nor ( n6729 , n6724 , n6728 );
and ( n6730 , n78 , n88 );
nor ( n6731 , n78 , n88 );
nor ( n6732 , n6730 , n6731 );
and ( n6733 , n6637 , n6732 );
not ( n6734 , n88 );
and ( n6735 , n6734 , n6535 );
and ( n6736 , n77 , n88 );
nor ( n6737 , n6735 , n6736 );
and ( n6738 , n6644 , n6737 );
nor ( n6739 , n6733 , n6738 );
xor ( n6740 , n6729 , n6739 );
not ( n6741 , n68 );
and ( n6742 , n6741 , n98 );
not ( n6743 , n6549 );
nor ( n6744 , n6742 , n6743 );
nand ( n6745 , n83 , n84 );
and ( n6746 , n6744 , n6745 );
nor ( n6747 , n6744 , n6745 );
nor ( n6748 , n6746 , n6747 );
xnor ( n6749 , n6740 , n6748 );
xor ( n6750 , n6720 , n6749 );
xnor ( n6751 , n6655 , n6750 );
or ( n6752 , n4 , n6698 );
nand ( n6753 , n6752 , n6699 );
not ( n6754 , n68 );
not ( n6755 , n6743 );
or ( n6756 , n6754 , n6755 );
not ( n6757 , n98 );
and ( n6758 , n6757 , n6741 );
and ( n6759 , n6578 , n98 );
nor ( n6760 , n6759 , n99 );
nor ( n6761 , n6758 , n6760 );
nand ( n6762 , n6756 , n6761 );
xor ( n6763 , n6753 , n6762 );
and ( n6764 , n6467 , n6479 );
and ( n6765 , n6474 , n6688 );
nor ( n6766 , n6764 , n6765 );
xor ( n6767 , n6763 , n6766 );
and ( n6768 , n6527 , n6538 );
and ( n6769 , n6524 , n6712 );
nor ( n6770 , n6768 , n6769 );
and ( n6771 , n6636 , n6648 );
and ( n6772 , n6644 , n6732 );
nor ( n6773 , n6771 , n6772 );
xor ( n6774 , n6770 , n6773 );
and ( n6775 , n6495 , n6505 );
and ( n6776 , n6501 , n6658 );
nor ( n6777 , n6775 , n6776 );
xor ( n6778 , n6774 , n6777 );
xor ( n6779 , n6767 , n6778 );
and ( n6780 , n6445 , n6456 );
and ( n6781 , n6452 , n6723 );
nor ( n6782 , n6780 , n6781 );
or ( n6783 , n6671 , n6564 );
or ( n6784 , n6665 , n6674 );
nand ( n6785 , n6783 , n6784 );
and ( n6786 , n6782 , n6785 );
not ( n6787 , n6782 );
not ( n6788 , n6785 );
and ( n6789 , n6787 , n6788 );
nor ( n6790 , n6786 , n6789 );
and ( n6791 , n6423 , n6434 );
not ( n6792 , n6420 );
and ( n6793 , n6792 , n6702 );
nor ( n6794 , n6791 , n6793 );
xnor ( n6795 , n6790 , n6794 );
and ( n6796 , n6779 , n6795 );
and ( n6797 , n6767 , n6778 );
nor ( n6798 , n6796 , n6797 );
and ( n6799 , n6596 , n6600 );
not ( n6800 , n6587 );
and ( n6801 , n6592 , n6800 );
nor ( n6802 , n6799 , n6801 );
and ( n6803 , n6798 , n6802 );
not ( n6804 , n6798 );
not ( n6805 , n6802 );
and ( n6806 , n6804 , n6805 );
nor ( n6807 , n6803 , n6806 );
xor ( n6808 , n6753 , n6762 );
and ( n6809 , n6808 , n6766 );
and ( n6810 , n6753 , n6762 );
nor ( n6811 , n6809 , n6810 );
xor ( n6812 , n6770 , n6773 );
and ( n6813 , n6812 , n6777 );
and ( n6814 , n6770 , n6773 );
nor ( n6815 , n6813 , n6814 );
xor ( n6816 , n6811 , n6815 );
or ( n6817 , n6790 , n6794 );
or ( n6818 , n6782 , n6788 );
nand ( n6819 , n6817 , n6818 );
xor ( n6820 , n6816 , n6819 );
xor ( n6821 , n6807 , n6820 );
or ( n6822 , n6751 , n6821 );
or ( n6823 , n6655 , n6750 );
nand ( n6824 , n6822 , n6823 );
nand ( n6825 , n6824 , n2526 );
and ( n6826 , n4564 , n6417 , n6825 );
not ( n6827 , n6826 );
not ( n6828 , n6827 );
or ( n6829 , n6807 , n6820 );
or ( n6830 , n6805 , n6798 );
nand ( n6831 , n6829 , n6830 );
and ( n6832 , n6495 , n6662 );
and ( n6833 , n6483 , n6741 );
and ( n6834 , n68 , n96 );
nor ( n6835 , n6833 , n6834 );
and ( n6836 , n6501 , n6835 );
nor ( n6837 , n6832 , n6836 );
and ( n6838 , n6637 , n6737 );
and ( n6839 , n6734 , n6469 );
and ( n6840 , n76 , n88 );
nor ( n6841 , n6839 , n6840 );
and ( n6842 , n6644 , n6841 );
nor ( n6843 , n6838 , n6842 );
xor ( n6844 , n6837 , n6843 );
and ( n6845 , n6423 , n6706 );
and ( n6846 , n6424 , n6554 );
and ( n6847 , n70 , n94 );
nor ( n6848 , n6846 , n6847 );
and ( n6849 , n6792 , n6848 );
nor ( n6850 , n6845 , n6849 );
xor ( n6851 , n6844 , n6850 );
not ( n6852 , n6729 );
not ( n6853 , n6739 );
and ( n6854 , n6852 , n6853 );
and ( n6855 , n6740 , n6748 );
nor ( n6856 , n6854 , n6855 );
xor ( n6857 , n6851 , n6856 );
and ( n6858 , n6816 , n6819 );
and ( n6859 , n6811 , n6815 );
nor ( n6860 , n6858 , n6859 );
xor ( n6861 , n6857 , n6860 );
xor ( n6862 , n6831 , n6861 );
xor ( n6863 , n6695 , n6719 );
and ( n6864 , n6863 , n6749 );
and ( n6865 , n6695 , n6719 );
nor ( n6866 , n6864 , n6865 );
xor ( n6867 , n6699 , n6708 );
and ( n6868 , n6867 , n6718 );
and ( n6869 , n6699 , n6708 );
nor ( n6870 , n6868 , n6869 );
xor ( n6871 , n6870 , n6747 );
and ( n6872 , n6445 , n6727 );
and ( n6873 , n6529 , n6446 );
and ( n6874 , n78 , n86 );
nor ( n6875 , n6873 , n6874 );
and ( n6876 , n6452 , n6875 );
nor ( n6877 , n6872 , n6876 );
not ( n6878 , n6877 );
xor ( n6879 , n6871 , n6878 );
xor ( n6880 , n6866 , n6879 );
or ( n6881 , n6671 , n6678 );
or ( n6882 , n80 , n84 );
nand ( n6883 , n80 , n84 );
nand ( n6884 , n6882 , n6883 );
or ( n6885 , n6665 , n6884 );
nand ( n6886 , n6881 , n6885 );
not ( n6887 , n6673 );
xor ( n6888 , n6886 , n6887 );
and ( n6889 , n6467 , n6692 );
and ( n6890 , n92 , n72 );
not ( n6891 , n92 );
and ( n6892 , n6891 , n6496 );
nor ( n6893 , n6890 , n6892 );
and ( n6894 , n6474 , n6893 );
nor ( n6895 , n6889 , n6894 );
not ( n6896 , n6895 );
and ( n6897 , n6888 , n6896 );
not ( n6898 , n6888 );
and ( n6899 , n6898 , n6895 );
nor ( n6900 , n6897 , n6899 );
and ( n6901 , n6527 , n6716 );
and ( n6902 , n6528 , n6425 );
and ( n6903 , n74 , n90 );
nor ( n6904 , n6902 , n6903 );
and ( n6905 , n6534 , n6904 );
nor ( n6906 , n6901 , n6905 );
or ( n6907 , n6906 , n98 );
nand ( n6908 , n6906 , n98 );
nand ( n6909 , n6907 , n6908 );
xor ( n6910 , n6900 , n6909 );
or ( n6911 , n6685 , n6694 );
or ( n6912 , n6664 , n6683 );
nand ( n6913 , n6911 , n6912 );
xor ( n6914 , n6910 , n6913 );
xor ( n6915 , n6880 , n6914 );
nand ( n6916 , n6862 , n6915 );
not ( n6917 , n6916 );
or ( n6918 , n6862 , n6915 );
nand ( n6919 , n6918 , n2526 );
nor ( n6920 , n6917 , n6919 );
not ( n6921 , n6920 );
or ( n6922 , n6828 , n6921 );
xor ( n6923 , n6751 , n6821 );
xnor ( n6924 , n6560 , n6567 );
and ( n6925 , n6452 , n83 );
xor ( n6926 , n7 , n6925 );
or ( n6927 , n6547 , n72 );
or ( n6928 , n6549 , n71 );
or ( n6929 , n6553 , n6502 );
nand ( n6930 , n6927 , n6928 , n6929 );
and ( n6931 , n6926 , n6930 );
and ( n6932 , n7 , n6925 );
nor ( n6933 , n6931 , n6932 );
not ( n6934 , n6423 );
not ( n6935 , n6934 );
and ( n6936 , n6424 , n76 );
and ( n6937 , n6469 , n94 );
nor ( n6938 , n6936 , n6937 );
not ( n6939 , n6938 );
and ( n6940 , n6935 , n6939 );
and ( n6941 , n6792 , n6607 );
nor ( n6942 , n6940 , n6941 );
not ( n6943 , n88 );
not ( n6944 , n6528 );
or ( n6945 , n6943 , n6944 );
nand ( n6946 , n6945 , n6633 );
nand ( n6947 , n6635 , n83 );
nand ( n6948 , n6946 , n6947 );
not ( n6949 , n6948 );
nand ( n6950 , n6949 , n8 );
xor ( n6951 , n6942 , n6950 );
and ( n6952 , n6475 , n6529 );
and ( n6953 , n78 , n92 );
nor ( n6954 , n6952 , n6953 );
and ( n6955 , n6467 , n6954 );
and ( n6956 , n6474 , n6613 );
nor ( n6957 , n6955 , n6956 );
and ( n6958 , n6951 , n6957 );
and ( n6959 , n6942 , n6950 );
nor ( n6960 , n6958 , n6959 );
and ( n6961 , n6933 , n6960 );
not ( n6962 , n6933 );
not ( n6963 , n6960 );
and ( n6964 , n6962 , n6963 );
nor ( n6965 , n6961 , n6964 );
or ( n6966 , n6924 , n6965 );
or ( n6967 , n6963 , n6933 );
nand ( n6968 , n6966 , n6967 );
and ( n6969 , n6528 , n6645 );
and ( n6970 , n79 , n90 );
nor ( n6971 , n6969 , n6970 );
and ( n6972 , n6527 , n6971 );
and ( n6973 , n6534 , n6532 );
nor ( n6974 , n6972 , n6973 );
and ( n6975 , n6453 , n6630 );
and ( n6976 , n81 , n88 );
nor ( n6977 , n6975 , n6976 );
and ( n6978 , n6638 , n6977 );
and ( n6979 , n6644 , n6642 );
nor ( n6980 , n6978 , n6979 );
xor ( n6981 , n6974 , n6980 );
not ( n6982 , n6981 );
and ( n6983 , n6483 , n6425 );
and ( n6984 , n74 , n96 );
nor ( n6985 , n6983 , n6984 );
and ( n6986 , n6495 , n6985 );
and ( n6987 , n6501 , n6620 );
nor ( n6988 , n6986 , n6987 );
and ( n6989 , n6438 , n6447 );
and ( n6990 , n82 , n88 );
nor ( n6991 , n6989 , n6990 );
and ( n6992 , n6637 , n6991 );
and ( n6993 , n6644 , n6977 );
nor ( n6994 , n6992 , n6993 );
xor ( n6995 , n6988 , n6994 );
and ( n6996 , n6528 , n6639 );
and ( n6997 , n80 , n90 );
nor ( n6998 , n6996 , n6997 );
and ( n6999 , n6527 , n6998 );
and ( n7000 , n6534 , n6971 );
nor ( n7001 , n6999 , n7000 );
and ( n7002 , n6995 , n7001 );
and ( n7003 , n6988 , n6994 );
nor ( n7004 , n7002 , n7003 );
not ( n7005 , n7004 );
or ( n7006 , n6982 , n7005 );
or ( n7007 , n6974 , n6980 );
nand ( n7008 , n7006 , n7007 );
xor ( n7009 , n6968 , n7008 );
xor ( n7010 , n6629 , n6650 );
and ( n7011 , n7009 , n7010 );
and ( n7012 , n6968 , n7008 );
nor ( n7013 , n7011 , n7012 );
xor ( n7014 , n6779 , n6795 );
or ( n7015 , n7013 , n7014 );
xor ( n7016 , n7013 , n7014 );
xor ( n7017 , n6575 , n6601 );
xor ( n7018 , n7017 , n6652 );
nand ( n7019 , n7016 , n7018 );
nand ( n7020 , n7015 , n7019 );
nand ( n7021 , n6923 , n7020 , n2526 );
nand ( n7022 , n6922 , n7021 );
or ( n7023 , n6831 , n6861 );
nand ( n7024 , n7023 , n6916 );
and ( n7025 , n6880 , n6914 );
and ( n7026 , n6866 , n6879 );
nor ( n7027 , n7025 , n7026 );
and ( n7028 , n6637 , n6841 );
and ( n7029 , n6734 , n6476 );
and ( n7030 , n75 , n88 );
nor ( n7031 , n7029 , n7030 );
and ( n7032 , n6644 , n7031 );
nor ( n7033 , n7028 , n7032 );
xor ( n7034 , n7033 , n6677 );
and ( n7035 , n6527 , n6904 );
and ( n7036 , n6528 , n6431 );
and ( n7037 , n73 , n90 );
nor ( n7038 , n7036 , n7037 );
and ( n7039 , n6534 , n7038 );
nor ( n7040 , n7035 , n7039 );
xor ( n7041 , n7034 , n7040 );
not ( n7042 , n7041 );
xor ( n7043 , n6870 , n6747 );
not ( n7044 , n6877 );
and ( n7045 , n7043 , n7044 );
and ( n7046 , n6870 , n6747 );
or ( n7047 , n7045 , n7046 );
xor ( n7048 , n7042 , n7047 );
buf ( n7049 , n6671 );
or ( n7050 , n7049 , n6884 );
or ( n7051 , n79 , n84 );
nand ( n7052 , n79 , n84 );
nand ( n7053 , n7051 , n7052 );
or ( n7054 , n6665 , n7053 );
nand ( n7055 , n7050 , n7054 );
xor ( n7056 , n6908 , n7055 );
not ( n7057 , n7056 );
and ( n7058 , n6888 , n6896 );
and ( n7059 , n6886 , n6887 );
nor ( n7060 , n7058 , n7059 );
not ( n7061 , n7060 );
or ( n7062 , n7057 , n7061 );
or ( n7063 , n7060 , n7056 );
nand ( n7064 , n7062 , n7063 );
xnor ( n7065 , n7048 , n7064 );
xnor ( n7066 , n7027 , n7065 );
and ( n7067 , n6860 , n6857 );
and ( n7068 , n6851 , n6856 );
nor ( n7069 , n7067 , n7068 );
and ( n7070 , n6495 , n6835 );
and ( n7071 , n6757 , n6486 );
not ( n7072 , n96 );
not ( n7073 , n6757 );
or ( n7074 , n7072 , n7073 );
nand ( n7075 , n7074 , n6487 );
not ( n7076 , n7075 );
nor ( n7077 , n7071 , n7076 );
nor ( n7078 , n7070 , n7077 );
and ( n7079 , n6423 , n6848 );
and ( n7080 , n6424 , n6578 );
and ( n7081 , n69 , n94 );
nor ( n7082 , n7080 , n7081 );
and ( n7083 , n6430 , n7082 );
nor ( n7084 , n7079 , n7083 );
or ( n7085 , n7078 , n7084 );
nand ( n7086 , n7078 , n7084 );
nand ( n7087 , n7085 , n7086 );
and ( n7088 , n6467 , n6893 );
and ( n7089 , n6475 , n6502 );
and ( n7090 , n71 , n92 );
nor ( n7091 , n7089 , n7090 );
and ( n7092 , n6474 , n7091 );
nor ( n7093 , n7088 , n7092 );
and ( n7094 , n6445 , n6875 );
and ( n7095 , n6535 , n6446 );
and ( n7096 , n77 , n86 );
nor ( n7097 , n7095 , n7096 );
and ( n7098 , n6452 , n7097 );
nor ( n7099 , n7094 , n7098 );
and ( n7100 , n7093 , n7099 );
nor ( n7101 , n7093 , n7099 );
nor ( n7102 , n7100 , n7101 );
xor ( n7103 , n7087 , n7102 );
xor ( n7104 , n6837 , n6843 );
and ( n7105 , n7104 , n6850 );
and ( n7106 , n6837 , n6843 );
nor ( n7107 , n7105 , n7106 );
xnor ( n7108 , n7103 , n7107 );
and ( n7109 , n6910 , n6913 );
and ( n7110 , n6900 , n6909 );
nor ( n7111 , n7109 , n7110 );
xor ( n7112 , n7108 , n7111 );
xnor ( n7113 , n7069 , n7112 );
xor ( n7114 , n7066 , n7113 );
nand ( n7115 , n7024 , n7114 , n2526 );
xor ( n7116 , n7033 , n6677 );
and ( n7117 , n7116 , n7040 );
and ( n7118 , n7033 , n6677 );
nor ( n7119 , n7117 , n7118 );
xor ( n7120 , n7119 , n7086 );
and ( n7121 , n6527 , n7038 );
and ( n7122 , n6528 , n6496 );
and ( n7123 , n72 , n90 );
nor ( n7124 , n7122 , n7123 );
and ( n7125 , n6534 , n7124 );
nor ( n7126 , n7121 , n7125 );
xnor ( n7127 , n7126 , n7075 );
and ( n7128 , n6423 , n7082 );
and ( n7129 , n6424 , n6741 );
and ( n7130 , n68 , n94 );
nor ( n7131 , n7129 , n7130 );
and ( n7132 , n6792 , n7131 );
nor ( n7133 , n7128 , n7132 );
xor ( n7134 , n7127 , n7133 );
xnor ( n7135 , n7120 , n7134 );
and ( n7136 , n7103 , n7107 );
and ( n7137 , n7087 , n7102 );
nor ( n7138 , n7136 , n7137 );
xnor ( n7139 , n7135 , n7138 );
and ( n7140 , n7048 , n7064 );
and ( n7141 , n7047 , n7042 );
nor ( n7142 , n7140 , n7141 );
xor ( n7143 , n7139 , n7142 );
and ( n7144 , n6637 , n7031 );
and ( n7145 , n6438 , n6425 );
and ( n7146 , n74 , n88 );
nor ( n7147 , n7145 , n7146 );
and ( n7148 , n6644 , n7147 );
nor ( n7149 , n7144 , n7148 );
xnor ( n7150 , n7149 , n6883 );
and ( n7151 , n6467 , n7091 );
buf ( n7152 , n6474 );
and ( n7153 , n92 , n70 );
not ( n7154 , n92 );
and ( n7155 , n7154 , n6554 );
nor ( n7156 , n7153 , n7155 );
and ( n7157 , n7152 , n7156 );
nor ( n7158 , n7151 , n7157 );
xor ( n7159 , n7150 , n7158 );
not ( n7160 , n7159 );
not ( n7161 , n7060 );
and ( n7162 , n7161 , n7056 );
and ( n7163 , n6908 , n7055 );
nor ( n7164 , n7162 , n7163 );
not ( n7165 , n7164 );
or ( n7166 , n7160 , n7165 );
or ( n7167 , n7164 , n7159 );
nand ( n7168 , n7166 , n7167 );
or ( n7169 , n7049 , n7053 );
not ( n7170 , n6665 );
not ( n7171 , n7170 );
or ( n7172 , n78 , n84 );
nand ( n7173 , n78 , n84 );
nand ( n7174 , n7172 , n7173 );
or ( n7175 , n7171 , n7174 );
nand ( n7176 , n7169 , n7175 );
and ( n7177 , n6445 , n7097 );
and ( n7178 , n6446 , n6469 );
and ( n7179 , n76 , n86 );
nor ( n7180 , n7178 , n7179 );
and ( n7181 , n6452 , n7180 );
nor ( n7182 , n7177 , n7181 );
not ( n7183 , n7182 );
and ( n7184 , n7176 , n7183 );
not ( n7185 , n7176 );
and ( n7186 , n7185 , n7182 );
nor ( n7187 , n7184 , n7186 );
xor ( n7188 , n7187 , n7101 );
xor ( n7189 , n7168 , n7188 );
not ( n7190 , n7112 );
not ( n7191 , n7069 );
or ( n7192 , n7190 , n7191 );
or ( n7193 , n7108 , n7111 );
nand ( n7194 , n7192 , n7193 );
xor ( n7195 , n7189 , n7194 );
xor ( n7196 , n7143 , n7195 );
or ( n7197 , n7066 , n7113 );
or ( n7198 , n7027 , n7065 );
nand ( n7199 , n7197 , n7198 );
nand ( n7200 , n7196 , n7199 , n2526 );
nand ( n7201 , n7115 , n7200 );
nor ( n7202 , n7022 , n7201 );
not ( n7203 , n7202 );
nand ( n7204 , n4110 , n4222 );
nand ( n7205 , n7204 , n4319 );
and ( n7206 , n7205 , n4410 );
buf ( n7207 , n4408 );
xnor ( n7208 , n7206 , n7207 );
not ( n7209 , n7208 );
not ( n7210 , n4563 );
or ( n7211 , n7209 , n7210 );
buf ( n7212 , n6401 );
not ( n7213 , n7212 );
nand ( n7214 , n6322 , n6361 );
not ( n7215 , n7214 );
or ( n7216 , n7213 , n7215 );
or ( n7217 , n7214 , n7212 );
nand ( n7218 , n7216 , n7217 );
and ( n7219 , n7218 , n6416 );
not ( n7220 , n90 );
not ( n7221 , n6475 );
or ( n7222 , n7220 , n7221 );
nand ( n7223 , n7222 , n6517 );
nand ( n7224 , n6523 , n83 );
and ( n7225 , n7223 , n7224 );
nor ( n7226 , n7225 , n10 );
not ( n7227 , n7226 );
nand ( n7228 , n7225 , n10 );
nand ( n7229 , n7227 , n7228 );
and ( n7230 , n6743 , n6425 );
or ( n7231 , n6547 , n75 );
or ( n7232 , n6553 , n6425 );
nand ( n7233 , n7231 , n7232 );
nor ( n7234 , n7230 , n7233 );
xnor ( n7235 , n7229 , n7234 );
and ( n7236 , n6424 , n6645 );
and ( n7237 , n79 , n94 );
nor ( n7238 , n7236 , n7237 );
and ( n7239 , n6423 , n7238 );
and ( n7240 , n94 , n78 );
not ( n7241 , n94 );
and ( n7242 , n7241 , n6529 );
nor ( n7243 , n7240 , n7242 );
and ( n7244 , n6792 , n7243 );
nor ( n7245 , n7239 , n7244 );
or ( n7246 , n7235 , n7245 );
or ( n7247 , n7229 , n7234 );
nand ( n7248 , n7246 , n7247 );
not ( n7249 , n7248 );
and ( n7250 , n6483 , n6469 );
and ( n7251 , n76 , n96 );
nor ( n7252 , n7250 , n7251 );
and ( n7253 , n6495 , n7252 );
and ( n7254 , n6483 , n6476 );
and ( n7255 , n75 , n96 );
nor ( n7256 , n7254 , n7255 );
and ( n7257 , n6501 , n7256 );
nor ( n7258 , n7253 , n7257 );
and ( n7259 , n6528 , n6447 );
and ( n7260 , n82 , n90 );
nor ( n7261 , n7259 , n7260 );
and ( n7262 , n6527 , n7261 );
and ( n7263 , n6453 , n6528 );
and ( n7264 , n81 , n90 );
nor ( n7265 , n7263 , n7264 );
and ( n7266 , n6534 , n7265 );
nor ( n7267 , n7262 , n7266 );
xor ( n7268 , n7258 , n7267 );
not ( n7269 , n7268 );
or ( n7270 , n7249 , n7269 );
or ( n7271 , n7258 , n7267 );
nand ( n7272 , n7270 , n7271 );
and ( n7273 , n6468 , n6645 );
and ( n7274 , n79 , n92 );
nor ( n7275 , n7273 , n7274 );
and ( n7276 , n6467 , n7275 );
and ( n7277 , n6474 , n6954 );
nor ( n7278 , n7276 , n7277 );
and ( n7279 , n6527 , n7265 );
and ( n7280 , n6524 , n6998 );
nor ( n7281 , n7279 , n7280 );
xnor ( n7282 , n7278 , n7281 );
and ( n7283 , n6495 , n7256 );
and ( n7284 , n6501 , n6985 );
nor ( n7285 , n7283 , n7284 );
xor ( n7286 , n7282 , n7285 );
xor ( n7287 , n7272 , n7286 );
not ( n7288 , n8 );
nand ( n7289 , n7288 , n6948 );
nand ( n7290 , n6950 , n7289 );
and ( n7291 , n6743 , n6496 );
or ( n7292 , n6547 , n73 );
or ( n7293 , n6553 , n6496 );
nand ( n7294 , n7292 , n7293 );
nor ( n7295 , n7291 , n7294 );
xnor ( n7296 , n7290 , n7295 );
and ( n7297 , n94 , n77 );
not ( n7298 , n94 );
and ( n7299 , n7298 , n6535 );
nor ( n7300 , n7297 , n7299 );
and ( n7301 , n6423 , n7300 );
not ( n7302 , n6938 );
and ( n7303 , n6792 , n7302 );
nor ( n7304 , n7301 , n7303 );
xor ( n7305 , n7296 , n7304 );
and ( n7306 , n7287 , n7305 );
and ( n7307 , n7272 , n7286 );
nor ( n7308 , n7306 , n7307 );
or ( n7309 , n7304 , n7296 );
or ( n7310 , n7290 , n7295 );
nand ( n7311 , n7309 , n7310 );
xor ( n7312 , n7 , n6925 );
xor ( n7313 , n7312 , n6930 );
xor ( n7314 , n7311 , n7313 );
or ( n7315 , n7282 , n7285 );
or ( n7316 , n7278 , n7281 );
nand ( n7317 , n7315 , n7316 );
xor ( n7318 , n7314 , n7317 );
not ( n7319 , n7318 );
or ( n7320 , n7308 , n7319 , n1 );
xnor ( n7321 , n7308 , n7319 );
not ( n7322 , n6422 );
and ( n7323 , n7322 , n7243 );
and ( n7324 , n6430 , n7300 );
nor ( n7325 , n7323 , n7324 );
xor ( n7326 , n7325 , n7228 );
and ( n7327 , n6475 , n6639 );
and ( n7328 , n80 , n92 );
nor ( n7329 , n7327 , n7328 );
and ( n7330 , n6467 , n7329 );
and ( n7331 , n6474 , n7275 );
nor ( n7332 , n7330 , n7331 );
and ( n7333 , n7326 , n7332 );
and ( n7334 , n7325 , n7228 );
nor ( n7335 , n7333 , n7334 );
not ( n7336 , n6991 );
not ( n7337 , n6644 );
or ( n7338 , n7336 , n7337 );
not ( n7339 , n6633 );
and ( n7340 , n6561 , n7339 );
not ( n7341 , n6631 );
and ( n7342 , n7341 , n83 );
nor ( n7343 , n7340 , n7342 );
or ( n7344 , n7343 , n6644 );
nand ( n7345 , n7338 , n7344 );
not ( n7346 , n9 );
not ( n7347 , n6947 );
or ( n7348 , n7346 , n7347 );
or ( n7349 , n6947 , n9 );
nand ( n7350 , n7348 , n7349 );
not ( n7351 , n7350 );
or ( n7352 , n6547 , n74 );
or ( n7353 , n6549 , n73 );
or ( n7354 , n6553 , n6431 );
nand ( n7355 , n7352 , n7353 , n7354 );
not ( n7356 , n7355 );
or ( n7357 , n7351 , n7356 );
not ( n7358 , n6947 );
nand ( n7359 , n7358 , n9 );
nand ( n7360 , n7357 , n7359 );
xor ( n7361 , n7345 , n7360 );
and ( n7362 , n7335 , n7361 );
and ( n7363 , n7345 , n7360 );
nor ( n7364 , n7362 , n7363 );
xor ( n7365 , n6942 , n6950 );
xor ( n7366 , n7365 , n6957 );
xor ( n7367 , n7364 , n7366 );
xor ( n7368 , n6988 , n6994 );
xor ( n7369 , n7368 , n7001 );
xor ( n7370 , n7367 , n7369 );
or ( n7371 , n7370 , n1 );
or ( n7372 , n7321 , n7371 );
nand ( n7373 , n7320 , n7372 );
nor ( n7374 , n7219 , n7373 );
nand ( n7375 , n7211 , n7374 );
and ( n7376 , n6446 , n1 );
xor ( n7377 , n6965 , n6924 );
not ( n7378 , n7377 );
xor ( n7379 , n7364 , n7366 );
and ( n7380 , n7379 , n7369 );
and ( n7381 , n7364 , n7366 );
nor ( n7382 , n7380 , n7381 );
not ( n7383 , n7382 );
or ( n7384 , n7378 , n7383 );
or ( n7385 , n7382 , n7377 );
nand ( n7386 , n7384 , n7385 );
xor ( n7387 , n7311 , n7313 );
and ( n7388 , n7387 , n7317 );
and ( n7389 , n7311 , n7313 );
nor ( n7390 , n7388 , n7389 );
xor ( n7391 , n6610 , n6616 );
xor ( n7392 , n7391 , n6623 );
xor ( n7393 , n7390 , n7392 );
xnor ( n7394 , n7004 , n6981 );
xor ( n7395 , n7393 , n7394 );
nor ( n7396 , n7386 , n7395 , n1 );
not ( n7397 , n7386 );
not ( n7398 , n7395 );
nor ( n7399 , n7397 , n7398 , n1 );
nor ( n7400 , n7376 , n7396 , n7399 );
nand ( n7401 , n7375 , n7400 );
not ( n7402 , n7401 );
not ( n7403 , n4316 );
nand ( n7404 , n7204 , n4318 );
not ( n7405 , n7404 );
or ( n7406 , n7403 , n7405 );
or ( n7407 , n7404 , n4316 );
nand ( n7408 , n7406 , n7407 );
nand ( n7409 , n7408 , n4563 );
not ( n7410 , n6222 );
and ( n7411 , n6232 , n6233 );
nor ( n7412 , n7410 , n7411 );
not ( n7413 , n6320 );
nand ( n7414 , n7413 , n6361 );
xor ( n7415 , n7412 , n7414 );
nand ( n7416 , n7415 , n6416 );
xor ( n7417 , n7325 , n7228 );
xor ( n7418 , n7417 , n7332 );
xnor ( n7419 , n7355 , n7350 );
and ( n7420 , n7418 , n7419 );
xor ( n7421 , n7419 , n7418 );
not ( n7422 , n7421 );
or ( n7423 , n6517 , n83 );
or ( n7424 , n6520 , n6561 );
nand ( n7425 , n7423 , n7424 );
and ( n7426 , n6525 , n7425 );
and ( n7427 , n6524 , n7261 );
nor ( n7428 , n7426 , n7427 );
and ( n7429 , n6483 , n6535 );
and ( n7430 , n77 , n96 );
nor ( n7431 , n7429 , n7430 );
and ( n7432 , n6495 , n7431 );
and ( n7433 , n6501 , n7252 );
nor ( n7434 , n7432 , n7433 );
xor ( n7435 , n7428 , n7434 );
and ( n7436 , n6475 , n6453 );
and ( n7437 , n81 , n92 );
nor ( n7438 , n7436 , n7437 );
and ( n7439 , n6467 , n7438 );
and ( n7440 , n6474 , n7329 );
nor ( n7441 , n7439 , n7440 );
and ( n7442 , n7435 , n7441 );
and ( n7443 , n7428 , n7434 );
nor ( n7444 , n7442 , n7443 );
nor ( n7445 , n7422 , n7444 );
nor ( n7446 , n7420 , n7445 );
xor ( n7447 , n7335 , n7361 );
and ( n7448 , n7446 , n7447 , n2526 );
xor ( n7449 , n7287 , n7305 );
xor ( n7450 , n7446 , n7447 );
nand ( n7451 , n7449 , n7450 , n2526 );
not ( n7452 , n7451 );
nor ( n7453 , n7448 , n7452 );
and ( n7454 , n7416 , n7453 );
or ( n7455 , n2526 , n87 );
nand ( n7456 , n7321 , n7370 , n2526 );
nand ( n7457 , n7455 , n7456 );
nor ( n7458 , n7321 , n7371 );
or ( n7459 , n7457 , n7458 );
nand ( n7460 , n7409 , n7454 , n7459 );
not ( n7461 , n7460 );
or ( n7462 , n2526 , n90 );
or ( n7463 , n6549 , n76 );
or ( n7464 , n6547 , n77 );
or ( n7465 , n6553 , n6469 );
nand ( n7466 , n7463 , n7464 , n7465 );
not ( n7467 , n7466 );
not ( n7468 , n512 );
nand ( n7469 , n83 , n6465 );
not ( n7470 , n93 );
not ( n7471 , n94 );
or ( n7472 , n7470 , n7471 );
nand ( n7473 , n7472 , n92 );
not ( n7474 , n7473 );
nand ( n7475 , n7469 , n7474 );
not ( n7476 , n7475 );
or ( n7477 , n7468 , n7476 );
or ( n7478 , n7475 , n512 );
nand ( n7479 , n7477 , n7478 );
not ( n7480 , n7479 );
or ( n7481 , n7467 , n7480 );
or ( n7482 , n7479 , n7466 );
nand ( n7483 , n7481 , n7482 );
not ( n7484 , n94 );
not ( n7485 , n81 );
or ( n7486 , n7484 , n7485 );
or ( n7487 , n81 , n94 );
nand ( n7488 , n7486 , n7487 );
or ( n7489 , n6934 , n7488 );
and ( n7490 , n6424 , n80 );
and ( n7491 , n6639 , n94 );
nor ( n7492 , n7490 , n7491 );
or ( n7493 , n6420 , n7492 );
nand ( n7494 , n7489 , n7493 );
and ( n7495 , n7483 , n7494 );
not ( n7496 , n7479 );
and ( n7497 , n7496 , n7466 );
nor ( n7498 , n7495 , n7497 );
or ( n7499 , n6549 , n75 );
not ( n7500 , n6547 );
nand ( n7501 , n7500 , n6469 );
nand ( n7502 , n6552 , n75 );
nand ( n7503 , n7499 , n7501 , n7502 );
not ( n7504 , n7503 );
and ( n7505 , n11 , n7224 );
not ( n7506 , n11 );
not ( n7507 , n7224 );
and ( n7508 , n7506 , n7507 );
nor ( n7509 , n7505 , n7508 );
not ( n7510 , n7509 );
and ( n7511 , n7504 , n7510 );
and ( n7512 , n7503 , n7509 );
nor ( n7513 , n7511 , n7512 );
and ( n7514 , n6483 , n6529 );
and ( n7515 , n78 , n96 );
nor ( n7516 , n7514 , n7515 );
and ( n7517 , n6495 , n7516 );
and ( n7518 , n6501 , n7431 );
nor ( n7519 , n7517 , n7518 );
xor ( n7520 , n7513 , n7519 );
and ( n7521 , n7498 , n7520 );
and ( n7522 , n7513 , n7519 );
nor ( n7523 , n7521 , n7522 );
not ( n7524 , n7523 );
xor ( n7525 , n7428 , n7434 );
xor ( n7526 , n7525 , n7441 );
not ( n7527 , n7526 );
not ( n7528 , n7527 );
and ( n7529 , n7524 , n7528 );
and ( n7530 , n7523 , n7527 );
nor ( n7531 , n7529 , n7530 );
xor ( n7532 , n7235 , n7245 );
and ( n7533 , n6475 , n6447 );
and ( n7534 , n82 , n92 );
nor ( n7535 , n7533 , n7534 );
and ( n7536 , n6467 , n7535 );
and ( n7537 , n6474 , n7438 );
nor ( n7538 , n7536 , n7537 );
xor ( n7539 , n7538 , n7478 );
not ( n7540 , n7492 );
and ( n7541 , n6423 , n7540 );
and ( n7542 , n6792 , n7238 );
nor ( n7543 , n7541 , n7542 );
and ( n7544 , n7539 , n7543 );
and ( n7545 , n7538 , n7478 );
nor ( n7546 , n7544 , n7545 );
xnor ( n7547 , n7532 , n7546 );
not ( n7548 , n7509 );
and ( n7549 , n7503 , n7548 );
and ( n7550 , n7507 , n11 );
nor ( n7551 , n7549 , n7550 );
xor ( n7552 , n7547 , n7551 );
nand ( n7553 , n7531 , n7552 , n2526 );
not ( n7554 , n7531 );
not ( n7555 , n7552 );
nand ( n7556 , n7554 , n7555 , n2526 );
nand ( n7557 , n7462 , n7553 , n7556 );
not ( n7558 , n7557 );
not ( n7559 , n3768 );
not ( n7560 , n3766 );
or ( n7561 , n7559 , n7560 );
nand ( n7562 , n7561 , n4095 );
nand ( n7563 , n7562 , n4103 );
not ( n7564 , n4101 );
or ( n7565 , n7563 , n7564 );
not ( n7566 , n4103 );
not ( n7567 , n7562 );
or ( n7568 , n7566 , n7567 );
nand ( n7569 , n7568 , n7564 );
nand ( n7570 , n7565 , n7569 );
not ( n7571 , n7570 );
not ( n7572 , n4563 );
or ( n7573 , n7571 , n7572 );
and ( n7574 , n5924 , n6010 );
nor ( n7575 , n7574 , n6009 );
not ( n7576 , n6011 );
or ( n7577 , n7575 , n7576 );
and ( n7578 , n7577 , n6416 );
xor ( n7579 , n7498 , n7520 );
xor ( n7580 , n7539 , n7543 );
xor ( n7581 , n7579 , n7580 );
and ( n7582 , n6483 , n6645 );
and ( n7583 , n79 , n96 );
nor ( n7584 , n7582 , n7583 );
and ( n7585 , n6495 , n7584 );
and ( n7586 , n6501 , n7516 );
nor ( n7587 , n7585 , n7586 );
and ( n7588 , n6424 , n6561 );
and ( n7589 , n83 , n94 );
nor ( n7590 , n7588 , n7589 );
not ( n7591 , n7590 );
and ( n7592 , n6467 , n7591 );
and ( n7593 , n6474 , n7535 );
nor ( n7594 , n7592 , n7593 );
xnor ( n7595 , n7587 , n7594 );
and ( n7596 , n6424 , n6447 );
and ( n7597 , n82 , n94 );
nor ( n7598 , n7596 , n7597 );
and ( n7599 , n6423 , n7598 );
not ( n7600 , n7488 );
and ( n7601 , n6792 , n7600 );
nor ( n7602 , n7599 , n7601 );
not ( n7603 , n7602 );
not ( n7604 , n7469 );
xor ( n7605 , n7604 , n13 );
and ( n7606 , n7603 , n7605 );
and ( n7607 , n7604 , n13 );
nor ( n7608 , n7606 , n7607 );
or ( n7609 , n7595 , n7608 );
or ( n7610 , n7587 , n7594 );
nand ( n7611 , n7609 , n7610 );
not ( n7612 , n7611 );
and ( n7613 , n7581 , n7612 );
and ( n7614 , n7579 , n7580 );
nor ( n7615 , n7613 , n7614 , n1 );
nor ( n7616 , n7578 , n7615 );
nand ( n7617 , n7573 , n7616 );
not ( n7618 , n7617 );
or ( n7619 , n7558 , n7618 );
or ( n7620 , n7617 , n7557 );
nand ( n7621 , n7619 , n7620 );
not ( n7622 , n7621 );
xor ( n7623 , n7595 , n7608 );
not ( n7624 , n7623 );
nand ( n7625 , n7624 , n2526 );
xnor ( n7626 , n7483 , n7494 );
not ( n7627 , n83 );
not ( n7628 , n6422 );
or ( n7629 , n7627 , n7628 );
and ( n7630 , n6419 , n94 );
nand ( n7631 , n7629 , n7630 );
not ( n7632 , n14 );
nor ( n7633 , n7631 , n7632 );
or ( n7634 , n6547 , n78 );
or ( n7635 , n6549 , n77 );
or ( n7636 , n6553 , n6535 );
nand ( n7637 , n7634 , n7635 , n7636 );
xnor ( n7638 , n7633 , n7637 );
not ( n7639 , n7638 );
and ( n7640 , n6483 , n6639 );
and ( n7641 , n80 , n96 );
nor ( n7642 , n7640 , n7641 );
and ( n7643 , n6495 , n7642 );
and ( n7644 , n6501 , n7584 );
nor ( n7645 , n7643 , n7644 );
not ( n7646 , n7645 );
and ( n7647 , n7639 , n7646 );
and ( n7648 , n7633 , n7637 );
nor ( n7649 , n7647 , n7648 );
xor ( n7650 , n7626 , n7649 );
or ( n7651 , n7625 , n7650 );
or ( n7652 , n92 , n2526 );
nand ( n7653 , n7650 , n7623 , n2526 );
nand ( n7654 , n7651 , n7652 , n7653 );
not ( n7655 , n7654 );
not ( n7656 , n4563 );
not ( n7657 , n3765 );
not ( n7658 , n7657 );
not ( n7659 , n3678 );
not ( n7660 , n7659 );
or ( n7661 , n7658 , n7660 );
nand ( n7662 , n7661 , n3766 );
not ( n7663 , n7662 );
or ( n7664 , n7656 , n7663 );
or ( n7665 , n5727 , n5819 );
nand ( n7666 , n7665 , n5820 );
and ( n7667 , n7666 , n6416 );
xnor ( n7668 , n7638 , n7645 );
and ( n7669 , n7605 , n7602 );
not ( n7670 , n7605 );
and ( n7671 , n7670 , n7603 );
nor ( n7672 , n7669 , n7671 );
and ( n7673 , n7668 , n7672 );
not ( n7674 , n7633 );
not ( n7675 , n14 );
nand ( n7676 , n7675 , n7631 );
nand ( n7677 , n7674 , n7676 );
not ( n7678 , n7677 );
or ( n7679 , n6547 , n79 );
or ( n7680 , n6549 , n78 );
or ( n7681 , n6553 , n6529 );
nand ( n7682 , n7679 , n7680 , n7681 );
not ( n7683 , n7682 );
and ( n7684 , n7678 , n7683 );
and ( n7685 , n7677 , n7682 );
nor ( n7686 , n7684 , n7685 );
not ( n7687 , n7686 );
and ( n7688 , n6423 , n7590 );
and ( n7689 , n6792 , n7598 );
nor ( n7690 , n7688 , n7689 );
not ( n7691 , n7690 );
and ( n7692 , n7687 , n7691 );
not ( n7693 , n7677 );
and ( n7694 , n7693 , n7682 );
nor ( n7695 , n7692 , n7694 );
xor ( n7696 , n7668 , n7672 );
and ( n7697 , n7695 , n7696 );
nor ( n7698 , n7673 , n7697 , n1 );
nor ( n7699 , n7667 , n7698 );
nand ( n7700 , n7664 , n7699 );
nand ( n7701 , n7655 , n7700 );
not ( n7702 , n7701 );
nand ( n7703 , n5820 , n5921 );
xor ( n7704 , n5915 , n5919 );
xnor ( n7705 , n7703 , n7704 );
and ( n7706 , n7705 , n6416 );
or ( n7707 , n7626 , n7649 , n1 );
nand ( n7708 , n7707 , n7653 );
nor ( n7709 , n7706 , n7708 );
or ( n7710 , n3769 , n4095 );
nand ( n7711 , n7710 , n7562 );
nand ( n7712 , n7711 , n4563 );
nand ( n7713 , n7709 , n7712 );
not ( n7714 , n7713 );
and ( n7715 , n7581 , n7611 );
not ( n7716 , n7581 );
and ( n7717 , n7716 , n7612 );
nor ( n7718 , n7715 , n7717 );
or ( n7719 , n7718 , n1 );
or ( n7720 , n2526 , n91 );
nand ( n7721 , n7719 , n7720 );
nor ( n7722 , n7714 , n7721 );
nor ( n7723 , n7702 , n7722 );
not ( n7724 , n7723 );
and ( n7725 , n6483 , n1 );
or ( n7726 , n6547 , n81 );
or ( n7727 , n6549 , n80 );
or ( n7728 , n6553 , n6639 );
nand ( n7729 , n7726 , n7727 , n7728 );
not ( n7730 , n7075 );
and ( n7731 , n6501 , n83 );
nor ( n7732 , n7730 , n7731 );
or ( n7733 , n7732 , n16 );
nor ( n7734 , n7076 , n7731 );
nand ( n7735 , n7734 , n16 );
nand ( n7736 , n7733 , n7735 );
and ( n7737 , n7729 , n7736 );
not ( n7738 , n7729 );
not ( n7739 , n7736 );
and ( n7740 , n7738 , n7739 );
nor ( n7741 , n7737 , n7740 );
and ( n7742 , n96 , n82 );
not ( n7743 , n96 );
and ( n7744 , n7743 , n6447 );
nor ( n7745 , n7742 , n7744 );
and ( n7746 , n6501 , n7745 );
not ( n7747 , n6501 );
or ( n7748 , n6487 , n83 );
or ( n7749 , n6484 , n6561 );
nand ( n7750 , n7748 , n7749 );
and ( n7751 , n7747 , n7750 );
nor ( n7752 , n7746 , n7751 );
nor ( n7753 , n7741 , n7752 , n1 );
not ( n7754 , n7741 );
not ( n7755 , n7752 );
nor ( n7756 , n7754 , n7755 , n1 );
nor ( n7757 , n7725 , n7753 , n7756 );
not ( n7758 , n5553 );
and ( n7759 , n7758 , n5551 );
not ( n7760 , n5554 );
nor ( n7761 , n7759 , n7760 );
not ( n7762 , n6416 );
or ( n7763 , n7761 , n7762 );
and ( n7764 , n7731 , n2526 , n17 );
nand ( n7765 , n6561 , n98 );
nand ( n7766 , n6547 , n7765 );
nand ( n7767 , n7766 , n18 );
nor ( n7768 , n7767 , n1 );
and ( n7769 , n7731 , n17 );
not ( n7770 , n7731 );
not ( n7771 , n17 );
and ( n7772 , n7770 , n7771 );
nor ( n7773 , n7769 , n7772 );
and ( n7774 , n7768 , n7773 );
nor ( n7775 , n7764 , n7774 );
nand ( n7776 , n7763 , n7775 );
not ( n7777 , n7776 );
not ( n7778 , n3639 );
not ( n7779 , n3631 );
and ( n7780 , n7778 , n7779 );
and ( n7781 , n3639 , n3631 );
nor ( n7782 , n7780 , n7781 );
not ( n7783 , n7782 );
nand ( n7784 , n3634 , n3621 );
nand ( n7785 , n7783 , n7784 );
not ( n7786 , n7785 );
not ( n7787 , n7784 );
nand ( n7788 , n7787 , n7782 );
not ( n7789 , n7788 );
or ( n7790 , n7786 , n7789 );
nand ( n7791 , n7790 , n4563 );
nand ( n7792 , n7777 , n7791 );
xor ( n7793 , n7757 , n7792 );
and ( n7794 , n6486 , n1 );
not ( n7795 , n7767 );
nor ( n7796 , n7795 , n7773 , n1 );
nor ( n7797 , n7794 , n7774 , n7796 );
xor ( n7798 , n5480 , n5486 );
xor ( n7799 , n7798 , n5548 );
and ( n7800 , n7799 , n6416 );
or ( n7801 , n6547 , n82 );
or ( n7802 , n81 , n6549 );
or ( n7803 , n6453 , n6553 );
nand ( n7804 , n7801 , n7802 , n7803 );
and ( n7805 , n7804 , n2526 );
nor ( n7806 , n7800 , n7805 );
not ( n7807 , n3574 );
not ( n7808 , n3620 );
nand ( n7809 , n7807 , n7808 );
not ( n7810 , n7809 );
not ( n7811 , n3621 );
or ( n7812 , n7810 , n7811 );
nand ( n7813 , n7812 , n4563 );
nand ( n7814 , n7806 , n7813 );
xor ( n7815 , n7797 , n7814 );
xor ( n7816 , n3595 , n3610 );
xor ( n7817 , n7816 , n3613 );
and ( n7818 , n7817 , n4563 );
not ( n7819 , n19 );
not ( n7820 , n2526 );
or ( n7821 , n7819 , n7820 );
xor ( n7822 , n5538 , n5520 );
xor ( n7823 , n7822 , n5542 );
or ( n7824 , n7823 , n7762 );
nand ( n7825 , n7821 , n7824 );
nor ( n7826 , n7818 , n7825 );
or ( n7827 , n1 , n83 );
nand ( n7828 , n7827 , n99 );
nor ( n7829 , n7826 , n7828 );
and ( n7830 , n6757 , n1 );
nor ( n7831 , n7766 , n1 , n18 );
nor ( n7832 , n7830 , n7768 , n7831 );
xor ( n7833 , n7829 , n7832 );
xor ( n7834 , n3587 , n3588 );
xor ( n7835 , n7834 , n3617 );
or ( n7836 , n7835 , n4562 );
xnor ( n7837 , n5514 , n5546 );
or ( n7838 , n7837 , n7762 );
and ( n7839 , n82 , n99 );
not ( n7840 , n7765 );
nor ( n7841 , n7839 , n7840 );
and ( n7842 , n6549 , n7841 );
not ( n7843 , n6549 );
and ( n7844 , n7843 , n82 );
nor ( n7845 , n7842 , n7844 );
nand ( n7846 , n7845 , n2526 );
nand ( n7847 , n7836 , n7838 , n7846 );
and ( n7848 , n7833 , n7847 );
and ( n7849 , n7829 , n7832 );
or ( n7850 , n7848 , n7849 );
and ( n7851 , n7815 , n7850 );
and ( n7852 , n7797 , n7814 );
or ( n7853 , n7851 , n7852 );
and ( n7854 , n7793 , n7853 );
and ( n7855 , n7757 , n7792 );
or ( n7856 , n7854 , n7855 );
not ( n7857 , n7856 );
and ( n7858 , n6792 , n83 );
or ( n7859 , n7858 , n15 );
nand ( n7860 , n7858 , n15 );
nand ( n7861 , n7859 , n7860 );
xor ( n7862 , n7861 , n7735 );
not ( n7863 , n7862 );
nand ( n7864 , n7863 , n2526 );
or ( n7865 , n6547 , n80 );
or ( n7866 , n79 , n6549 );
or ( n7867 , n6645 , n6553 );
nand ( n7868 , n7865 , n7866 , n7867 );
not ( n7869 , n7868 );
and ( n7870 , n6495 , n7745 );
and ( n7871 , n96 , n81 );
not ( n7872 , n96 );
and ( n7873 , n7872 , n6453 );
nor ( n7874 , n7871 , n7873 );
and ( n7875 , n6501 , n7874 );
nor ( n7876 , n7870 , n7875 );
not ( n7877 , n7876 );
or ( n7878 , n7869 , n7877 );
or ( n7879 , n7876 , n7868 );
nand ( n7880 , n7878 , n7879 );
or ( n7881 , n7864 , n7880 );
or ( n7882 , n95 , n2526 );
nand ( n7883 , n7862 , n7880 , n2526 );
nand ( n7884 , n7881 , n7882 , n7883 );
buf ( n7885 , n7884 );
not ( n7886 , n7885 );
not ( n7887 , n3642 );
not ( n7888 , n7887 );
nand ( n7889 , n7785 , n3503 , n3632 );
not ( n7890 , n7889 );
or ( n7891 , n7888 , n7890 );
nand ( n7892 , n7891 , n4563 );
or ( n7893 , n5421 , n5555 );
nand ( n7894 , n7893 , n5556 );
nand ( n7895 , n7894 , n6416 );
and ( n7896 , n7739 , n7729 , n2526 );
nor ( n7897 , n7896 , n7753 );
nand ( n7898 , n7892 , n7895 , n7897 );
not ( n7899 , n7898 );
or ( n7900 , n7886 , n7899 );
or ( n7901 , n7898 , n7885 );
nand ( n7902 , n7900 , n7901 );
not ( n7903 , n7902 );
or ( n7904 , n7857 , n7903 );
not ( n7905 , n7885 );
nand ( n7906 , n7905 , n7898 );
nand ( n7907 , n7904 , n7906 );
not ( n7908 , n7907 );
xor ( n7909 , n7686 , n7690 );
and ( n7910 , n6495 , n7874 );
and ( n7911 , n6501 , n7642 );
nor ( n7912 , n7910 , n7911 );
not ( n7913 , n7912 );
and ( n7914 , n7909 , n7913 );
not ( n7915 , n7909 );
and ( n7916 , n7915 , n7912 );
nor ( n7917 , n7914 , n7916 );
or ( n7918 , n7861 , n7735 );
nand ( n7919 , n7918 , n7860 );
or ( n7920 , n7917 , n7919 , n1 );
or ( n7921 , n2526 , n94 );
nand ( n7922 , n7920 , n7921 );
and ( n7923 , n7917 , n7919 , n2526 );
nor ( n7924 , n7922 , n7923 );
not ( n7925 , n7924 );
not ( n7926 , n3661 );
not ( n7927 , n3644 );
nor ( n7928 , n7926 , n7927 );
or ( n7929 , n7928 , n3662 );
nand ( n7930 , n7929 , n4563 );
or ( n7931 , n5557 , n5623 );
nand ( n7932 , n5557 , n5623 );
nand ( n7933 , n7931 , n7932 );
nand ( n7934 , n7933 , n6416 );
not ( n7935 , n7883 );
not ( n7936 , n7868 );
nor ( n7937 , n7876 , n7936 , n1 );
nor ( n7938 , n7935 , n7937 );
and ( n7939 , n7930 , n7934 , n7938 );
not ( n7940 , n7939 );
or ( n7941 , n7925 , n7940 );
or ( n7942 , n7924 , n7939 );
nand ( n7943 , n7941 , n7942 );
not ( n7944 , n7943 );
or ( n7945 , n7908 , n7944 );
not ( n7946 , n7939 );
nand ( n7947 , n7946 , n7924 );
nand ( n7948 , n7945 , n7947 );
not ( n7949 , n3665 );
nor ( n7950 , n7949 , n3662 );
buf ( n7951 , n3673 );
xor ( n7952 , n7950 , n7951 );
nand ( n7953 , n7952 , n4563 );
not ( n7954 , n5626 );
not ( n7955 , n5715 );
or ( n7956 , n7954 , n7955 );
or ( n7957 , n5715 , n5626 );
nand ( n7958 , n7956 , n7957 );
not ( n7959 , n7958 );
nand ( n7960 , n5722 , n7932 );
not ( n7961 , n7960 );
or ( n7962 , n7959 , n7961 );
or ( n7963 , n7960 , n7958 );
nand ( n7964 , n7962 , n7963 );
nand ( n7965 , n7964 , n6416 );
and ( n7966 , n7909 , n7913 , n2526 );
nor ( n7967 , n7966 , n7923 );
nand ( n7968 , n7953 , n7965 , n7967 );
xor ( n7969 , n7695 , n7696 );
and ( n7970 , n7969 , n2526 );
not ( n7971 , n93 );
and ( n7972 , n7971 , n1 );
nor ( n7973 , n7970 , n7972 );
nor ( n7974 , n7968 , n7973 );
not ( n7975 , n7974 );
nand ( n7976 , n7968 , n7973 );
nand ( n7977 , n7975 , n7976 );
nor ( n7978 , n7948 , n7977 );
buf ( n7979 , n7974 );
nor ( n7980 , n7978 , n7979 );
xnor ( n7981 , n7654 , n7700 );
nand ( n7982 , n7980 , n7981 );
not ( n7983 , n7982 );
or ( n7984 , n7724 , n7983 );
not ( n7985 , n7713 );
nand ( n7986 , n7985 , n7721 );
nand ( n7987 , n7984 , n7986 );
not ( n7988 , n7987 );
or ( n7989 , n7622 , n7988 );
not ( n7990 , n7617 );
nand ( n7991 , n7990 , n7557 );
nand ( n7992 , n7989 , n7991 );
not ( n7993 , n4563 );
nand ( n7994 , n7569 , n4106 );
xor ( n7995 , n7994 , n4100 );
not ( n7996 , n7995 );
or ( n7997 , n7993 , n7996 );
not ( n7998 , n6220 );
nor ( n7999 , n7576 , n7998 );
not ( n8000 , n7999 );
xnor ( n8001 , n6230 , n6229 );
not ( n8002 , n8001 );
or ( n8003 , n8000 , n8002 );
or ( n8004 , n8001 , n7999 );
nand ( n8005 , n8003 , n8004 );
and ( n8006 , n6416 , n8005 );
nand ( n8007 , n7523 , n7527 , n2526 );
nand ( n8008 , n7553 , n8007 );
nor ( n8009 , n8006 , n8008 );
nand ( n8010 , n7997 , n8009 );
not ( n8011 , n7444 );
not ( n8012 , n7421 );
and ( n8013 , n8011 , n8012 );
and ( n8014 , n7421 , n7444 );
nor ( n8015 , n8013 , n8014 );
xor ( n8016 , n7248 , n7268 );
xor ( n8017 , n8015 , n8016 );
not ( n8018 , n7546 );
not ( n8019 , n7532 );
or ( n8020 , n8018 , n8019 );
or ( n8021 , n7547 , n7551 );
nand ( n8022 , n8020 , n8021 );
or ( n8023 , n8017 , n8022 );
nand ( n8024 , n8017 , n8022 );
nand ( n8025 , n8023 , n8024 );
and ( n8026 , n8025 , n2526 );
and ( n8027 , n6632 , n1 );
nor ( n8028 , n8026 , n8027 );
or ( n8029 , n8010 , n8028 );
or ( n8030 , n4110 , n4222 );
nand ( n8031 , n8030 , n7204 );
not ( n8032 , n8031 );
not ( n8033 , n4563 );
or ( n8034 , n8032 , n8033 );
not ( n8035 , n6122 );
nor ( n8036 , n6228 , n8035 , n7762 );
nand ( n8037 , n7999 , n8036 );
not ( n8038 , n8037 );
and ( n8039 , n6228 , n6231 , n6416 );
not ( n8040 , n8039 );
not ( n8041 , n7999 );
not ( n8042 , n8041 );
or ( n8043 , n8040 , n8042 );
and ( n8044 , n8039 , n8035 );
or ( n8045 , n6228 , n6231 , n7762 );
and ( n8046 , n8015 , n8016 );
not ( n8047 , n8024 );
nor ( n8048 , n8046 , n8047 );
or ( n8049 , n8048 , n1 );
nand ( n8050 , n8045 , n8049 );
nor ( n8051 , n8044 , n8050 );
nand ( n8052 , n8043 , n8051 );
nor ( n8053 , n8038 , n8052 );
nand ( n8054 , n8034 , n8053 );
or ( n8055 , n2526 , n88 );
not ( n8056 , n7449 );
not ( n8057 , n7450 );
nand ( n8058 , n8056 , n8057 , n2526 );
nand ( n8059 , n8055 , n7451 , n8058 );
xor ( n8060 , n8054 , n8059 );
not ( n8061 , n8060 );
nand ( n8062 , n8029 , n8061 );
nor ( n8063 , n7461 , n7992 , n8062 );
nand ( n8064 , n8010 , n8028 );
or ( n8065 , n8060 , n8064 );
not ( n8066 , n8059 );
nand ( n8067 , n8066 , n8054 );
nand ( n8068 , n8065 , n8067 );
not ( n8069 , n8068 );
not ( n8070 , n7460 );
or ( n8071 , n8069 , n8070 );
not ( n8072 , n7459 );
nand ( n8073 , n7409 , n7454 );
nand ( n8074 , n8072 , n8073 );
nand ( n8075 , n8071 , n8074 );
nor ( n8076 , n8063 , n8075 );
not ( n8077 , n8076 );
or ( n8078 , n7402 , n8077 );
xor ( n8079 , n7009 , n7010 );
not ( n8080 , n8079 );
nand ( n8081 , n8080 , n2526 );
xor ( n8082 , n7390 , n7392 );
and ( n8083 , n8082 , n7394 );
and ( n8084 , n7390 , n7392 );
nor ( n8085 , n8083 , n8084 );
not ( n8086 , n6542 );
not ( n8087 , n6571 );
and ( n8088 , n8086 , n8087 );
and ( n8089 , n6542 , n6571 );
nor ( n8090 , n8088 , n8089 );
xor ( n8091 , n8085 , n8090 );
or ( n8092 , n8081 , n8091 );
or ( n8093 , n85 , n2526 );
nand ( n8094 , n8091 , n2526 , n8079 );
nand ( n8095 , n8092 , n8093 , n8094 );
xnor ( n8096 , n6383 , n6381 );
not ( n8097 , n8096 );
not ( n8098 , n7212 );
not ( n8099 , n7214 );
or ( n8100 , n8098 , n8099 );
nand ( n8101 , n8100 , n6396 );
not ( n8102 , n8101 );
or ( n8103 , n8097 , n8102 );
not ( n8104 , n8101 );
not ( n8105 , n8096 );
and ( n8106 , n8104 , n8105 );
nor ( n8107 , n8106 , n7762 );
nand ( n8108 , n8103 , n8107 );
nand ( n8109 , n8095 , n8108 );
not ( n8110 , n8109 );
not ( n8111 , n7206 );
not ( n8112 , n7207 );
or ( n8113 , n8111 , n8112 );
buf ( n8114 , n4369 );
nand ( n8115 , n8113 , n8114 );
not ( n8116 , n4404 );
xnor ( n8117 , n8115 , n8116 );
nor ( n8118 , n8117 , n4562 );
not ( n8119 , n8118 );
and ( n8120 , n7382 , n7377 , n2526 );
nor ( n8121 , n8120 , n7396 );
and ( n8122 , n8110 , n8119 , n8121 );
nor ( n8123 , n7375 , n7400 );
nor ( n8124 , n8122 , n8123 );
nand ( n8125 , n8078 , n8124 );
buf ( n8126 , n4421 );
not ( n8127 , n8115 );
not ( n8128 , n8116 );
and ( n8129 , n8127 , n8128 );
not ( n8130 , n4419 );
nor ( n8131 , n8129 , n8130 );
xnor ( n8132 , n8126 , n8131 );
not ( n8133 , n8132 );
not ( n8134 , n4563 );
or ( n8135 , n8133 , n8134 );
not ( n8136 , n6404 );
or ( n8137 , n7214 , n6397 );
nand ( n8138 , n8136 , n8137 );
not ( n8139 , n6406 );
nand ( n8140 , n8139 , n6400 );
xnor ( n8141 , n8138 , n8140 );
nand ( n8142 , n8141 , n6416 );
and ( n8143 , n8085 , n8090 , n2526 );
not ( n8144 , n8094 );
nor ( n8145 , n8143 , n8144 );
and ( n8146 , n8142 , n8145 );
nand ( n8147 , n8135 , n8146 );
or ( n8148 , n7016 , n7018 );
nand ( n8149 , n8148 , n7019 );
and ( n8150 , n8149 , n2526 );
and ( n8151 , n6668 , n1 );
nor ( n8152 , n8150 , n8151 );
buf ( n8153 , n8152 );
and ( n8154 , n8147 , n8153 );
not ( n8155 , n8121 );
nor ( n8156 , n8155 , n8118 );
buf ( n8157 , n8108 );
and ( n8158 , n8156 , n8157 );
buf ( n8159 , n8095 );
nor ( n8160 , n8158 , n8159 );
nor ( n8161 , n8154 , n8160 );
nand ( n8162 , n8125 , n8161 );
not ( n8163 , n2 );
not ( n8164 , n8131 );
not ( n8165 , n8126 );
or ( n8166 , n8164 , n8165 );
buf ( n8167 , n4398 );
nand ( n8168 , n8166 , n8167 );
xor ( n8169 , n8168 , n4429 );
not ( n8170 , n8169 );
or ( n8171 , n8163 , n8170 );
not ( n8172 , n6408 );
xnor ( n8173 , n5234 , n5282 );
or ( n8174 , n8172 , n8173 );
and ( n8175 , n8172 , n8173 );
nor ( n8176 , n8175 , n2526 );
nand ( n8177 , n8174 , n8176 );
nand ( n8178 , n8177 , n4562 );
nand ( n8179 , n8171 , n8178 );
or ( n8180 , n6923 , n7020 );
nand ( n8181 , n8180 , n2526 );
nand ( n8182 , n8179 , n8181 );
not ( n8183 , n8147 );
not ( n8184 , n8153 );
nand ( n8185 , n8183 , n8184 );
nand ( n8186 , n8162 , n8182 , n8185 );
not ( n8187 , n8186 );
or ( n8188 , n7203 , n8187 );
not ( n8189 , n4552 );
nand ( n8190 , n8189 , n4436 );
not ( n8191 , n8190 );
not ( n8192 , n4559 );
or ( n8193 , n8191 , n8192 );
nand ( n8194 , n2121 , n46 );
and ( n8195 , n3474 , n8194 );
not ( n8196 , n710 );
not ( n8197 , n2632 );
or ( n8198 , n8196 , n8197 );
not ( n8199 , n4506 );
nand ( n8200 , n8199 , n2581 );
nand ( n8201 , n8198 , n8200 );
xor ( n8202 , n8195 , n8201 );
buf ( n8203 , n2541 );
not ( n8204 , n8203 );
not ( n8205 , n4494 );
or ( n8206 , n8204 , n8205 );
not ( n8207 , n788 );
nand ( n8208 , n8207 , n2550 );
nand ( n8209 , n8206 , n8208 );
xor ( n8210 , n8202 , n8209 );
not ( n8211 , n4526 );
and ( n8212 , n8211 , n4532 );
not ( n8213 , n4522 );
nor ( n8214 , n8213 , n4520 );
nor ( n8215 , n8212 , n8214 );
not ( n8216 , n8215 );
and ( n8217 , n8210 , n8216 );
not ( n8218 , n8210 );
and ( n8219 , n8218 , n8215 );
nor ( n8220 , n8217 , n8219 );
not ( n8221 , n4518 );
or ( n8222 , n2986 , n8221 );
or ( n8223 , n2714 , n721 );
nand ( n8224 , n8222 , n8223 );
not ( n8225 , n8224 );
and ( n8226 , n752 , n374 );
nor ( n8227 , n8226 , n2776 );
and ( n8228 , n749 , n8227 );
not ( n8229 , n4530 );
nor ( n8230 , n8229 , n5039 );
nor ( n8231 , n8228 , n8230 );
not ( n8232 , n8231 );
or ( n8233 , n8225 , n8232 );
or ( n8234 , n8224 , n8231 );
nand ( n8235 , n8233 , n8234 );
not ( n8236 , n4485 );
not ( n8237 , n2564 );
or ( n8238 , n8236 , n8237 );
not ( n8239 , n6069 );
or ( n8240 , n769 , n8239 );
nand ( n8241 , n8238 , n8240 );
xnor ( n8242 , n8235 , n8241 );
xnor ( n8243 , n8220 , n8242 );
not ( n8244 , n4475 );
not ( n8245 , n4468 );
or ( n8246 , n8244 , n8245 );
not ( n8247 , n4467 );
nand ( n8248 , n8247 , n4464 );
nand ( n8249 , n8246 , n8248 );
not ( n8250 , n4487 );
not ( n8251 , n8250 );
not ( n8252 , n4496 );
and ( n8253 , n8251 , n8252 );
and ( n8254 , n4500 , n4508 );
nor ( n8255 , n8253 , n8254 );
and ( n8256 , n1002 , n4463 );
not ( n8257 , n1002 );
and ( n8258 , n8257 , n4464 );
nor ( n8259 , n8256 , n8258 );
and ( n8260 , n8255 , n8259 );
not ( n8261 , n8255 );
not ( n8262 , n8259 );
and ( n8263 , n8261 , n8262 );
nor ( n8264 , n8260 , n8263 );
xor ( n8265 , n8249 , n8264 );
not ( n8266 , n8265 );
not ( n8267 , n4509 );
nand ( n8268 , n8267 , n4546 );
not ( n8269 , n4536 );
nand ( n8270 , n8269 , n4542 );
and ( n8271 , n8268 , n8270 );
not ( n8272 , n8271 );
and ( n8273 , n8266 , n8272 );
and ( n8274 , n8265 , n8271 );
nor ( n8275 , n8273 , n8274 );
xor ( n8276 , n8243 , n8275 );
xor ( n8277 , n4459 , n4476 );
and ( n8278 , n8277 , n4550 );
and ( n8279 , n4459 , n4476 );
nor ( n8280 , n8278 , n8279 );
xor ( n8281 , n8276 , n8280 );
not ( n8282 , n8281 );
not ( n8283 , n4551 );
not ( n8284 , n4452 );
or ( n8285 , n8283 , n8284 );
not ( n8286 , n4443 );
nand ( n8287 , n8286 , n4450 );
nand ( n8288 , n8285 , n8287 );
not ( n8289 , n8288 );
or ( n8290 , n8282 , n8289 );
or ( n8291 , n8281 , n8288 );
nand ( n8292 , n8290 , n8291 );
not ( n8293 , n8292 );
not ( n8294 , n8293 );
nand ( n8295 , n8193 , n8294 );
buf ( n8296 , n8295 );
not ( n8297 , n8288 );
nand ( n8298 , n8297 , n8281 );
nand ( n8299 , n8296 , n8298 );
xor ( n8300 , n8243 , n8275 );
and ( n8301 , n8300 , n8280 );
and ( n8302 , n8243 , n8275 );
nor ( n8303 , n8301 , n8302 );
not ( n8304 , n8220 );
not ( n8305 , n8242 );
and ( n8306 , n8304 , n8305 );
and ( n8307 , n8210 , n8215 );
nor ( n8308 , n8306 , n8307 );
not ( n8309 , n40 );
not ( n8310 , n2595 );
or ( n8311 , n8309 , n8310 );
or ( n8312 , n2595 , n40 );
nand ( n8313 , n8311 , n8312 );
not ( n8314 , n8313 );
not ( n8315 , n2550 );
or ( n8316 , n8314 , n8315 );
not ( n8317 , n788 );
nand ( n8318 , n8317 , n8203 );
nand ( n8319 , n8316 , n8318 );
and ( n8320 , n36 , n675 );
not ( n8321 , n8320 );
not ( n8322 , n720 );
not ( n8323 , n2722 );
or ( n8324 , n8322 , n8323 );
xor ( n8325 , n42 , n2790 );
nand ( n8326 , n8325 , n2713 );
nand ( n8327 , n8324 , n8326 );
not ( n8328 , n8327 );
or ( n8329 , n8321 , n8328 );
or ( n8330 , n8327 , n8320 );
nand ( n8331 , n8329 , n8330 );
xnor ( n8332 , n8319 , n8331 );
or ( n8333 , n8259 , n8255 );
or ( n8334 , n4464 , n1002 );
nand ( n8335 , n8333 , n8334 );
xor ( n8336 , n8332 , n8335 );
xnor ( n8337 , n8308 , n8336 );
not ( n8338 , n8268 );
not ( n8339 , n8270 );
or ( n8340 , n8338 , n8339 );
nand ( n8341 , n8340 , n8265 );
nand ( n8342 , n8249 , n8264 );
and ( n8343 , n8341 , n8342 );
not ( n8344 , n8231 );
not ( n8345 , n8224 );
not ( n8346 , n8345 );
and ( n8347 , n8344 , n8346 );
and ( n8348 , n8235 , n8241 );
nor ( n8349 , n8347 , n8348 );
xor ( n8350 , n8195 , n8201 );
and ( n8351 , n8350 , n8209 );
and ( n8352 , n8195 , n8201 );
nor ( n8353 , n8351 , n8352 );
xor ( n8354 , n8349 , n8353 );
or ( n8355 , n769 , n8237 );
and ( n8356 , n38 , n2646 );
not ( n8357 , n38 );
and ( n8358 , n8357 , n2641 );
or ( n8359 , n8356 , n8358 );
or ( n8360 , n8239 , n8359 );
nand ( n8361 , n8355 , n8360 );
not ( n8362 , n8361 );
not ( n8363 , n869 );
not ( n8364 , n5039 );
and ( n8365 , n8363 , n8364 );
not ( n8366 , n587 );
not ( n8367 , n374 );
or ( n8368 , n8366 , n8367 );
nand ( n8369 , n2555 , n36 );
nand ( n8370 , n8368 , n8369 );
not ( n8371 , n8370 );
and ( n8372 , n8371 , n2682 );
nor ( n8373 , n8365 , n8372 );
not ( n8374 , n8373 );
or ( n8375 , n8362 , n8374 );
or ( n8376 , n8373 , n8361 );
nand ( n8377 , n8375 , n8376 );
or ( n8378 , n711 , n2955 );
nand ( n8379 , n8378 , n5352 );
xnor ( n8380 , n8377 , n8379 );
xor ( n8381 , n8354 , n8380 );
and ( n8382 , n8343 , n8381 );
not ( n8383 , n8343 );
not ( n8384 , n8381 );
and ( n8385 , n8383 , n8384 );
nor ( n8386 , n8382 , n8385 );
xnor ( n8387 , n8337 , n8386 );
xor ( n8388 , n8303 , n8387 );
nor ( n8389 , n8299 , n8388 );
not ( n8390 , n8389 );
not ( n8391 , n8298 );
not ( n8392 , n8295 );
or ( n8393 , n8391 , n8392 );
nand ( n8394 , n8393 , n8388 );
buf ( n8395 , n8394 );
nand ( n8396 , n8390 , n8395 );
nand ( n8397 , n8396 , n4563 );
and ( n8398 , n4818 , n4823 );
and ( n8399 , n4809 , n4814 );
nor ( n8400 , n8398 , n8399 );
not ( n8401 , n4636 );
not ( n8402 , n4623 );
or ( n8403 , n8401 , n8402 );
not ( n8404 , n4603 );
nand ( n8405 , n8404 , n4619 );
nand ( n8406 , n8403 , n8405 );
and ( n8407 , n4566 , n4814 );
not ( n8408 , n4566 );
and ( n8409 , n8408 , n4813 );
nor ( n8410 , n8407 , n8409 );
xnor ( n8411 , n8406 , n8410 );
xor ( n8412 , n8400 , n8411 );
and ( n8413 , n4682 , n4592 );
not ( n8414 , n4680 );
and ( n8415 , n4640 , n8414 );
nor ( n8416 , n8413 , n8415 );
and ( n8417 , n8412 , n8416 );
and ( n8418 , n8400 , n8411 );
nor ( n8419 , n8417 , n8418 );
and ( n8420 , n4617 , n2581 );
and ( n8421 , n44 , n52 );
not ( n8422 , n44 );
and ( n8423 , n8422 , n4666 );
nor ( n8424 , n8421 , n8423 );
and ( n8425 , n2587 , n8424 );
nor ( n8426 , n8420 , n8425 );
not ( n8427 , n8426 );
not ( n8428 , n8195 );
and ( n8429 , n8427 , n8428 );
and ( n8430 , n8426 , n8195 );
nor ( n8431 , n8429 , n8430 );
and ( n8432 , n8203 , n4633 );
not ( n8433 , n40 );
not ( n8434 , n56 );
and ( n8435 , n8433 , n8434 );
and ( n8436 , n40 , n56 );
nor ( n8437 , n8435 , n8436 );
and ( n8438 , n2550 , n8437 );
nor ( n8439 , n8432 , n8438 );
or ( n8440 , n8431 , n8439 );
not ( n8441 , n8195 );
or ( n8442 , n8426 , n8441 );
nand ( n8443 , n8440 , n8442 );
and ( n8444 , n304 , n4701 );
and ( n8445 , n38 , n58 );
nor ( n8446 , n8444 , n8445 );
and ( n8447 , n2564 , n8446 );
and ( n8448 , n38 , n57 );
nor ( n8449 , n38 , n57 );
nor ( n8450 , n8448 , n8449 );
and ( n8451 , n6069 , n8450 );
nor ( n8452 , n8447 , n8451 );
not ( n8453 , n8452 );
not ( n8454 , n8424 );
not ( n8455 , n2581 );
or ( n8456 , n8454 , n8455 );
nand ( n8457 , n8456 , n5352 );
or ( n8458 , n36 , n60 );
nand ( n8459 , n36 , n60 );
nand ( n8460 , n8458 , n8459 );
not ( n8461 , n8460 );
not ( n8462 , n8461 );
not ( n8463 , n4528 );
or ( n8464 , n8462 , n8463 );
or ( n8465 , n36 , n59 );
nand ( n8466 , n36 , n59 );
nand ( n8467 , n8465 , n8466 );
not ( n8468 , n8467 );
nand ( n8469 , n8468 , n2682 );
nand ( n8470 , n8464 , n8469 );
xor ( n8471 , n8457 , n8470 );
not ( n8472 , n8471 );
or ( n8473 , n8453 , n8472 );
or ( n8474 , n8471 , n8452 );
nand ( n8475 , n8473 , n8474 );
xor ( n8476 , n8443 , n8475 );
and ( n8477 , n2564 , n4601 );
and ( n8478 , n6069 , n8446 );
nor ( n8479 , n8477 , n8478 );
or ( n8480 , n2678 , n4571 );
not ( n8481 , n2682 );
or ( n8482 , n8481 , n8460 );
nand ( n8483 , n8480 , n8482 );
and ( n8484 , n8479 , n8483 );
not ( n8485 , n8479 );
not ( n8486 , n8483 );
and ( n8487 , n8485 , n8486 );
nor ( n8488 , n8484 , n8487 );
and ( n8489 , n2722 , n4579 );
xor ( n8490 , n42 , n54 );
and ( n8491 , n2715 , n8490 );
nor ( n8492 , n8489 , n8491 );
or ( n8493 , n8488 , n8492 );
or ( n8494 , n8486 , n8479 );
nand ( n8495 , n8493 , n8494 );
xor ( n8496 , n8476 , n8495 );
xor ( n8497 , n8419 , n8496 );
xor ( n8498 , n8488 , n8492 );
not ( n8499 , n8498 );
xnor ( n8500 , n8431 , n8439 );
not ( n8501 , n8500 );
not ( n8502 , n4573 );
not ( n8503 , n4591 );
or ( n8504 , n8502 , n8503 );
not ( n8505 , n4589 );
nand ( n8506 , n8505 , n4590 );
nand ( n8507 , n8504 , n8506 );
not ( n8508 , n8507 );
or ( n8509 , n8501 , n8508 );
or ( n8510 , n8507 , n8500 );
nand ( n8511 , n8509 , n8510 );
not ( n8512 , n8511 );
or ( n8513 , n8499 , n8512 );
not ( n8514 , n8500 );
nand ( n8515 , n8514 , n8507 );
nand ( n8516 , n8513 , n8515 );
not ( n8517 , n2540 );
not ( n8518 , n8437 );
not ( n8519 , n8518 );
and ( n8520 , n8517 , n8519 );
and ( n8521 , n427 , n4577 );
and ( n8522 , n40 , n55 );
nor ( n8523 , n8521 , n8522 );
and ( n8524 , n2550 , n8523 );
nor ( n8525 , n8520 , n8524 );
xor ( n8526 , n8525 , n4570 );
and ( n8527 , n2722 , n8490 );
and ( n8528 , n42 , n53 );
not ( n8529 , n42 );
and ( n8530 , n8529 , n4615 );
nor ( n8531 , n8528 , n8530 );
and ( n8532 , n2713 , n8531 );
nor ( n8533 , n8527 , n8532 );
xor ( n8534 , n8526 , n8533 );
not ( n8535 , n8534 );
not ( n8536 , n4566 );
not ( n8537 , n4814 );
or ( n8538 , n8536 , n8537 );
not ( n8539 , n8406 );
nand ( n8540 , n8539 , n8410 );
nand ( n8541 , n8538 , n8540 );
not ( n8542 , n8541 );
or ( n8543 , n8535 , n8542 );
or ( n8544 , n8541 , n8534 );
nand ( n8545 , n8543 , n8544 );
xnor ( n8546 , n8516 , n8545 );
not ( n8547 , n8546 );
xor ( n8548 , n8497 , n8547 );
not ( n8549 , n8548 );
xor ( n8550 , n8400 , n8411 );
xor ( n8551 , n8550 , n8416 );
not ( n8552 , n8551 );
xor ( n8553 , n8498 , n8511 );
xor ( n8554 , n8552 , n8553 );
or ( n8555 , n4832 , n4683 );
or ( n8556 , n4788 , n4827 );
nand ( n8557 , n8555 , n8556 );
and ( n8558 , n8554 , n8557 );
and ( n8559 , n8552 , n8553 );
nor ( n8560 , n8558 , n8559 );
not ( n8561 , n8560 );
and ( n8562 , n8549 , n8561 );
and ( n8563 , n8560 , n8548 );
nor ( n8564 , n8562 , n8563 );
not ( n8565 , n8564 );
xor ( n8566 , n8552 , n8553 );
xor ( n8567 , n8566 , n8557 );
not ( n8568 , n8567 );
nand ( n8569 , n6409 , n5283 );
nor ( n8570 , n8569 , n5232 );
buf ( n8571 , n5229 );
nor ( n8572 , n8570 , n8571 );
not ( n8573 , n8572 );
or ( n8574 , n8568 , n8573 );
not ( n8575 , n8571 );
not ( n8576 , n8575 );
not ( n8577 , n8569 );
or ( n8578 , n8576 , n8577 );
not ( n8579 , n5231 );
nor ( n8580 , n8579 , n8567 );
nand ( n8581 , n8578 , n8580 );
not ( n8582 , n4833 );
not ( n8583 , n5084 );
not ( n8584 , n8583 );
or ( n8585 , n8582 , n8584 );
not ( n8586 , n5063 );
not ( n8587 , n5080 );
or ( n8588 , n8586 , n8587 );
nand ( n8589 , n8585 , n8588 );
nand ( n8590 , n8581 , n8589 );
nand ( n8591 , n8574 , n8590 );
buf ( n8592 , n8591 );
not ( n8593 , n8592 );
or ( n8594 , n8565 , n8593 );
or ( n8595 , n8592 , n8564 );
nand ( n8596 , n8594 , n8595 );
nand ( n8597 , n8596 , n6416 );
or ( n8598 , n7199 , n7196 );
nand ( n8599 , n8598 , n2526 );
nand ( n8600 , n8397 , n8597 , n8599 );
not ( n8601 , n6920 );
nand ( n8602 , n8601 , n6826 );
not ( n8603 , n8602 );
nand ( n8604 , n4560 , n8190 , n8293 );
nand ( n8605 , n8604 , n8296 , n2 );
not ( n8606 , n8605 );
not ( n8607 , n1 );
xnor ( n8608 , n8567 , n8589 );
xnor ( n8609 , n8608 , n8572 );
not ( n8610 , n8609 );
or ( n8611 , n8607 , n8610 );
nand ( n8612 , n8611 , n4562 );
not ( n8613 , n8612 );
or ( n8614 , n8606 , n8613 );
or ( n8615 , n7024 , n7114 );
nand ( n8616 , n8615 , n2526 );
nand ( n8617 , n8614 , n8616 );
not ( n8618 , n8617 );
or ( n8619 , n8603 , n8618 );
not ( n8620 , n7201 );
nand ( n8621 , n8619 , n8620 );
nand ( n8622 , n8600 , n8621 );
not ( n8623 , n8622 );
nand ( n8624 , n8188 , n8623 );
not ( n8625 , n8624 );
not ( n8626 , n8625 );
or ( n8627 , n7142 , n7139 );
or ( n8628 , n7135 , n7138 );
nand ( n8629 , n8627 , n8628 );
and ( n8630 , n7187 , n7101 );
and ( n8631 , n7183 , n7176 );
nor ( n8632 , n8630 , n8631 );
or ( n8633 , n7049 , n7174 );
or ( n8634 , n77 , n84 );
nand ( n8635 , n77 , n84 );
nand ( n8636 , n8634 , n8635 );
or ( n8637 , n6665 , n8636 );
nand ( n8638 , n8633 , n8637 );
not ( n8639 , n8638 );
not ( n8640 , n7052 );
and ( n8641 , n8639 , n8640 );
and ( n8642 , n8638 , n7052 );
nor ( n8643 , n8641 , n8642 );
and ( n8644 , n6527 , n7124 );
and ( n8645 , n6528 , n6502 );
and ( n8646 , n71 , n90 );
nor ( n8647 , n8645 , n8646 );
and ( n8648 , n6534 , n8647 );
nor ( n8649 , n8644 , n8648 );
xnor ( n8650 , n8643 , n8649 );
xnor ( n8651 , n8632 , n8650 );
and ( n8652 , n6638 , n7147 );
and ( n8653 , n6630 , n6431 );
and ( n8654 , n73 , n88 );
nor ( n8655 , n8653 , n8654 );
and ( n8656 , n6644 , n8655 );
nor ( n8657 , n8652 , n8656 );
and ( n8658 , n6445 , n7180 );
and ( n8659 , n6446 , n6476 );
and ( n8660 , n75 , n86 );
nor ( n8661 , n8659 , n8660 );
and ( n8662 , n6452 , n8661 );
nor ( n8663 , n8658 , n8662 );
xor ( n8664 , n8657 , n8663 );
and ( n8665 , n6467 , n7156 );
and ( n8666 , n92 , n69 );
not ( n8667 , n92 );
and ( n8668 , n8667 , n6578 );
nor ( n8669 , n8666 , n8668 );
and ( n8670 , n7152 , n8669 );
nor ( n8671 , n8665 , n8670 );
xor ( n8672 , n8664 , n8671 );
xor ( n8673 , n8651 , n8672 );
xor ( n8674 , n8629 , n8673 );
and ( n8675 , n7120 , n7134 );
and ( n8676 , n7119 , n7086 );
nor ( n8677 , n8675 , n8676 );
or ( n8678 , n7150 , n7158 );
or ( n8679 , n7149 , n6883 );
nand ( n8680 , n8678 , n8679 );
and ( n8681 , n6423 , n7131 );
and ( n8682 , n6792 , n94 );
nor ( n8683 , n8681 , n8682 );
xor ( n8684 , n8680 , n8683 );
or ( n8685 , n7127 , n7133 );
or ( n8686 , n7126 , n7075 );
nand ( n8687 , n8685 , n8686 );
xnor ( n8688 , n8684 , n8687 );
xnor ( n8689 , n8677 , n8688 );
and ( n8690 , n7168 , n7188 );
not ( n8691 , n7164 );
and ( n8692 , n8691 , n7159 );
nor ( n8693 , n8690 , n8692 );
xor ( n8694 , n8689 , n8693 );
or ( n8695 , n8674 , n8694 );
nand ( n8696 , n8674 , n8694 );
nand ( n8697 , n8695 , n8696 , n2526 );
and ( n8698 , n8476 , n8495 );
and ( n8699 , n8475 , n8443 );
nor ( n8700 , n8698 , n8699 );
not ( n8701 , n8700 );
not ( n8702 , n8545 );
not ( n8703 , n8516 );
or ( n8704 , n8702 , n8703 );
not ( n8705 , n8541 );
nand ( n8706 , n8705 , n8534 );
nand ( n8707 , n8704 , n8706 );
not ( n8708 , n8707 );
or ( n8709 , n8701 , n8708 );
or ( n8710 , n8707 , n8700 );
nand ( n8711 , n8709 , n8710 );
or ( n8712 , n2678 , n8467 );
or ( n8713 , n36 , n58 );
nand ( n8714 , n36 , n58 );
nand ( n8715 , n8713 , n8714 );
or ( n8716 , n2776 , n8715 );
nand ( n8717 , n8712 , n8716 );
not ( n8718 , n8459 );
xor ( n8719 , n8717 , n8718 );
and ( n8720 , n3043 , n8523 );
and ( n8721 , n54 , n40 );
not ( n8722 , n54 );
and ( n8723 , n8722 , n427 );
nor ( n8724 , n8721 , n8723 );
and ( n8725 , n2550 , n8724 );
nor ( n8726 , n8720 , n8725 );
not ( n8727 , n8726 );
and ( n8728 , n8719 , n8727 );
not ( n8729 , n8719 );
and ( n8730 , n8729 , n8726 );
nor ( n8731 , n8728 , n8730 );
not ( n8732 , n8731 );
not ( n8733 , n8457 );
not ( n8734 , n8470 );
or ( n8735 , n8733 , n8734 );
not ( n8736 , n8452 );
nand ( n8737 , n8736 , n8471 );
nand ( n8738 , n8735 , n8737 );
not ( n8739 , n8738 );
not ( n8740 , n8533 );
and ( n8741 , n8739 , n8740 );
and ( n8742 , n8738 , n8533 );
nor ( n8743 , n8741 , n8742 );
not ( n8744 , n8743 );
or ( n8745 , n8732 , n8744 );
or ( n8746 , n8731 , n8743 );
nand ( n8747 , n8745 , n8746 );
not ( n8748 , n8533 );
not ( n8749 , n8526 );
or ( n8750 , n8748 , n8749 );
or ( n8751 , n8525 , n4570 );
nand ( n8752 , n8750 , n8751 );
not ( n8753 , n8752 );
and ( n8754 , n2564 , n8450 );
and ( n8755 , n304 , n4585 );
and ( n8756 , n38 , n56 );
nor ( n8757 , n8755 , n8756 );
and ( n8758 , n2573 , n8757 );
nor ( n8759 , n8754 , n8758 );
nand ( n8760 , n5352 , n3328 );
not ( n8761 , n8760 );
and ( n8762 , n8759 , n8761 );
not ( n8763 , n8759 );
and ( n8764 , n8763 , n8760 );
nor ( n8765 , n8762 , n8764 );
and ( n8766 , n2722 , n8531 );
and ( n8767 , n42 , n52 );
not ( n8768 , n42 );
and ( n8769 , n8768 , n4666 );
nor ( n8770 , n8767 , n8769 );
and ( n8771 , n2715 , n8770 );
nor ( n8772 , n8766 , n8771 );
xnor ( n8773 , n8765 , n8772 );
not ( n8774 , n8773 );
or ( n8775 , n8753 , n8774 );
or ( n8776 , n8752 , n8773 );
nand ( n8777 , n8775 , n8776 );
xnor ( n8778 , n8747 , n8777 );
xnor ( n8779 , n8711 , n8778 );
xor ( n8780 , n8419 , n8496 );
not ( n8781 , n8546 );
and ( n8782 , n8780 , n8781 );
and ( n8783 , n8419 , n8496 );
or ( n8784 , n8782 , n8783 );
xor ( n8785 , n8779 , n8784 );
nor ( n8786 , n8591 , n8564 );
not ( n8787 , n8560 );
nor ( n8788 , n8787 , n8548 );
nor ( n8789 , n8786 , n8788 );
xor ( n8790 , n8785 , n8789 );
nand ( n8791 , n8790 , n6416 );
or ( n8792 , n8387 , n8303 );
not ( n8793 , n8792 );
not ( n8794 , n8394 );
or ( n8795 , n8793 , n8794 );
not ( n8796 , n8386 );
or ( n8797 , n8796 , n8337 );
or ( n8798 , n8343 , n8381 );
nand ( n8799 , n8797 , n8798 );
not ( n8800 , n8799 );
or ( n8801 , n8336 , n8308 );
not ( n8802 , n8335 );
or ( n8803 , n8802 , n8332 );
nand ( n8804 , n8801 , n8803 );
not ( n8805 , n8379 );
not ( n8806 , n8377 );
or ( n8807 , n8805 , n8806 );
not ( n8808 , n8373 );
nand ( n8809 , n8808 , n8361 );
nand ( n8810 , n8807 , n8809 );
not ( n8811 , n8810 );
not ( n8812 , n8327 );
not ( n8813 , n8812 );
and ( n8814 , n8811 , n8813 );
and ( n8815 , n8810 , n8812 );
nor ( n8816 , n8814 , n8815 );
not ( n8817 , n8816 );
and ( n8818 , n596 , n2682 );
nor ( n8819 , n8370 , n2678 );
nor ( n8820 , n8818 , n8819 );
not ( n8821 , n8313 );
not ( n8822 , n2951 );
or ( n8823 , n8821 , n8822 );
nand ( n8824 , n640 , n2550 );
nand ( n8825 , n8823 , n8824 );
not ( n8826 , n8825 );
not ( n8827 , n749 );
and ( n8828 , n8826 , n8827 );
and ( n8829 , n8825 , n749 );
nor ( n8830 , n8828 , n8829 );
xor ( n8831 , n8820 , n8830 );
not ( n8832 , n8831 );
and ( n8833 , n8817 , n8832 );
and ( n8834 , n8831 , n8816 );
nor ( n8835 , n8833 , n8834 );
not ( n8836 , n8761 );
not ( n8837 , n8325 );
not ( n8838 , n2722 );
or ( n8839 , n8837 , n8838 );
nand ( n8840 , n570 , n2715 );
nand ( n8841 , n8839 , n8840 );
not ( n8842 , n8841 );
not ( n8843 , n8842 );
or ( n8844 , n8836 , n8843 );
nand ( n8845 , n8841 , n8760 );
nand ( n8846 , n8844 , n8845 );
not ( n8847 , n8846 );
not ( n8848 , n561 );
not ( n8849 , n8239 );
and ( n8850 , n8848 , n8849 );
not ( n8851 , n8359 );
buf ( n8852 , n2564 );
and ( n8853 , n8851 , n8852 );
nor ( n8854 , n8850 , n8853 );
not ( n8855 , n8854 );
and ( n8856 , n8847 , n8855 );
and ( n8857 , n8846 , n8854 );
nor ( n8858 , n8856 , n8857 );
and ( n8859 , n8319 , n8331 );
and ( n8860 , n8812 , n8320 );
nor ( n8861 , n8859 , n8860 );
xor ( n8862 , n8858 , n8861 );
not ( n8863 , n8862 );
and ( n8864 , n8835 , n8863 );
not ( n8865 , n8835 );
and ( n8866 , n8865 , n8862 );
nor ( n8867 , n8864 , n8866 );
xor ( n8868 , n8349 , n8353 );
and ( n8869 , n8868 , n8380 );
and ( n8870 , n8349 , n8353 );
nor ( n8871 , n8869 , n8870 );
xor ( n8872 , n8867 , n8871 );
xnor ( n8873 , n8804 , n8872 );
nand ( n8874 , n8800 , n8873 );
not ( n8875 , n8873 );
nand ( n8876 , n8875 , n8799 );
nand ( n8877 , n8874 , n8876 );
nand ( n8878 , n8795 , n8877 );
and ( n8879 , n8874 , n8792 );
and ( n8880 , n8879 , n8298 );
and ( n8881 , n8880 , n8190 );
not ( n8882 , n8881 );
not ( n8883 , n4559 );
or ( n8884 , n8882 , n8883 );
not ( n8885 , n8293 );
not ( n8886 , n8298 );
or ( n8887 , n8885 , n8886 );
nand ( n8888 , n8887 , n8388 );
nand ( n8889 , n8888 , n8879 );
nand ( n8890 , n8884 , n8889 );
nand ( n8891 , n8876 , n8890 );
nand ( n8892 , n8878 , n8891 , n4563 );
and ( n8893 , n7143 , n7195 );
and ( n8894 , n7189 , n7194 );
or ( n8895 , n8893 , n8894 );
nand ( n8896 , n8895 , n2526 );
nand ( n8897 , n8791 , n8892 , n8896 );
xnor ( n8898 , n8697 , n8897 );
not ( n8899 , n8898 );
not ( n8900 , n8899 );
or ( n8901 , n8626 , n8900 );
nand ( n8902 , n8624 , n8898 );
nand ( n8903 , n8901 , n8902 );
not ( n8904 , n8903 );
buf ( n8905 , n7115 );
not ( n8906 , n8905 );
nand ( n8907 , n8600 , n7200 );
not ( n8908 , n8907 );
or ( n8909 , n8906 , n8908 );
or ( n8910 , n8907 , n8905 );
nand ( n8911 , n8909 , n8910 );
and ( n8912 , n8162 , n8185 );
not ( n8913 , n8912 );
and ( n8914 , n8182 , n7021 );
and ( n8915 , n8913 , n8914 );
not ( n8916 , n8913 );
not ( n8917 , n8914 );
and ( n8918 , n8916 , n8917 );
nor ( n8919 , n8915 , n8918 );
nor ( n8920 , n8911 , n8919 );
not ( n8921 , n8912 );
not ( n8922 , n8914 );
or ( n8923 , n8921 , n8922 );
nand ( n8924 , n8923 , n7021 );
not ( n8925 , n8924 );
and ( n8926 , n6920 , n6827 );
not ( n8927 , n6920 );
and ( n8928 , n8927 , n6826 );
nor ( n8929 , n8926 , n8928 );
not ( n8930 , n8929 );
and ( n8931 , n8925 , n8930 );
and ( n8932 , n8924 , n8929 );
nor ( n8933 , n8931 , n8932 );
not ( n8934 , n7022 );
not ( n8935 , n8934 );
not ( n8936 , n8186 );
or ( n8937 , n8935 , n8936 );
nand ( n8938 , n8937 , n8602 );
nand ( n8939 , n8617 , n8905 );
nand ( n8940 , n8938 , n8939 );
nand ( n8941 , n8920 , n8933 , n8940 );
nor ( n8942 , n8904 , n8941 );
nand ( n8943 , n7982 , n7701 );
not ( n8944 , n8943 );
xnor ( n8945 , n7985 , n7721 );
not ( n8946 , n8945 );
and ( n8947 , n8944 , n8946 );
and ( n8948 , n8943 , n8945 );
nor ( n8949 , n8947 , n8948 );
not ( n8950 , n8949 );
not ( n8951 , n16 );
or ( n8952 , n8950 , n8951 );
or ( n8953 , n8949 , n16 );
nand ( n8954 , n8952 , n8953 );
not ( n8955 , n8954 );
not ( n8956 , n17 );
not ( n8957 , n7980 );
xor ( n8958 , n8957 , n7981 );
not ( n8959 , n8958 );
or ( n8960 , n8956 , n8959 );
or ( n8961 , n17 , n8958 );
nand ( n8962 , n8960 , n8961 );
not ( n8963 , n18 );
not ( n8964 , n8963 );
xor ( n8965 , n7943 , n7907 );
nand ( n8966 , n8965 , n19 );
not ( n8967 , n8966 );
and ( n8968 , n8964 , n8967 );
not ( n8969 , n18 );
not ( n8970 , n8966 );
or ( n8971 , n8969 , n8970 );
or ( n8972 , n8966 , n18 );
nand ( n8973 , n8971 , n8972 );
not ( n8974 , n7978 );
nand ( n8975 , n7977 , n7948 );
nand ( n8976 , n8974 , n8975 );
and ( n8977 , n8973 , n8976 );
nor ( n8978 , n8968 , n8977 );
nand ( n8979 , n8962 , n8978 );
nand ( n8980 , n8958 , n7771 );
and ( n8981 , n8979 , n8980 );
not ( n8982 , n8981 );
or ( n8983 , n8955 , n8982 );
not ( n8984 , n8949 );
nand ( n8985 , n16 , n8984 );
nand ( n8986 , n8983 , n8985 );
buf ( n8987 , n7987 );
xnor ( n8988 , n7621 , n8987 );
and ( n8989 , n8986 , n8988 );
not ( n8990 , n8989 );
not ( n8991 , n7621 );
not ( n8992 , n7987 );
or ( n8993 , n8991 , n8992 );
nand ( n8994 , n8993 , n7991 );
nor ( n8995 , n8010 , n8028 );
not ( n8996 , n8995 );
nand ( n8997 , n8996 , n8064 );
xor ( n8998 , n8994 , n8997 );
or ( n8999 , n8997 , n8994 );
buf ( n9000 , n8064 );
nand ( n9001 , n8999 , n9000 );
buf ( n9002 , n8061 );
and ( n9003 , n9001 , n9002 );
not ( n9004 , n9001 );
not ( n9005 , n9002 );
and ( n9006 , n9004 , n9005 );
nor ( n9007 , n9003 , n9006 );
nand ( n9008 , n8998 , n9007 );
nor ( n9009 , n8990 , n9008 );
xor ( n9010 , n7400 , n7375 );
not ( n9011 , n9010 );
buf ( n9012 , n8076 );
not ( n9013 , n9012 );
not ( n9014 , n9013 );
or ( n9015 , n9011 , n9014 );
nand ( n9016 , n9015 , n7401 );
nand ( n9017 , n8119 , n8110 , n8121 );
not ( n9018 , n8160 );
nand ( n9019 , n9017 , n9018 );
not ( n9020 , n9019 );
and ( n9021 , n9016 , n9020 );
not ( n9022 , n9016 );
and ( n9023 , n9022 , n9019 );
nor ( n9024 , n9021 , n9023 );
not ( n9025 , n9002 );
not ( n9026 , n9001 );
or ( n9027 , n9025 , n9026 );
nand ( n9028 , n9027 , n8067 );
not ( n9029 , n9028 );
nand ( n9030 , n7460 , n8074 );
not ( n9031 , n9030 );
or ( n9032 , n9029 , n9031 );
or ( n9033 , n9028 , n9030 );
nand ( n9034 , n9032 , n9033 );
xnor ( n9035 , n9012 , n9010 );
nand ( n9036 , n9009 , n9024 , n9034 , n9035 );
nand ( n9037 , n8125 , n9018 );
and ( n9038 , n8183 , n8153 );
not ( n9039 , n8183 );
and ( n9040 , n9039 , n8184 );
nor ( n9041 , n9038 , n9040 );
xor ( n9042 , n9037 , n9041 );
nor ( n9043 , n9036 , n9042 );
not ( n9044 , n9043 );
not ( n9045 , n9044 );
not ( n9046 , n8897 );
nand ( n9047 , n9046 , n8697 );
nand ( n9048 , n8902 , n9047 );
and ( n9049 , n8684 , n8687 );
and ( n9050 , n8680 , n8683 );
nor ( n9051 , n9049 , n9050 );
xor ( n9052 , n8657 , n8663 );
and ( n9053 , n9052 , n8671 );
and ( n9054 , n8657 , n8663 );
nor ( n9055 , n9053 , n9054 );
xor ( n9056 , n8683 , n7173 );
xnor ( n9057 , n9055 , n9056 );
xnor ( n9058 , n9051 , n9057 );
and ( n9059 , n6527 , n8647 );
and ( n9060 , n6528 , n6554 );
and ( n9061 , n70 , n90 );
nor ( n9062 , n9060 , n9061 );
and ( n9063 , n6534 , n9062 );
nor ( n9064 , n9059 , n9063 );
and ( n9065 , n6445 , n8661 );
and ( n9066 , n6446 , n6425 );
and ( n9067 , n74 , n86 );
nor ( n9068 , n9066 , n9067 );
and ( n9069 , n6452 , n9068 );
nor ( n9070 , n9065 , n9069 );
xor ( n9071 , n9064 , n9070 );
or ( n9072 , n7049 , n8636 );
or ( n9073 , n76 , n84 );
and ( n9074 , n76 , n84 );
not ( n9075 , n9074 );
nand ( n9076 , n9073 , n9075 );
or ( n9077 , n7171 , n9076 );
nand ( n9078 , n9072 , n9077 );
xor ( n9079 , n9071 , n9078 );
or ( n9080 , n8643 , n8649 );
not ( n9081 , n8638 );
or ( n9082 , n9081 , n7052 );
nand ( n9083 , n9080 , n9082 );
xor ( n9084 , n9079 , n9083 );
and ( n9085 , n6638 , n8655 );
and ( n9086 , n6734 , n6496 );
and ( n9087 , n72 , n88 );
nor ( n9088 , n9086 , n9087 );
and ( n9089 , n6644 , n9088 );
nor ( n9090 , n9085 , n9089 );
xnor ( n9091 , n9090 , n7630 );
and ( n9092 , n6467 , n8669 );
and ( n9093 , n92 , n68 );
not ( n9094 , n92 );
and ( n9095 , n9094 , n6741 );
nor ( n9096 , n9093 , n9095 );
and ( n9097 , n7152 , n9096 );
nor ( n9098 , n9092 , n9097 );
xor ( n9099 , n9091 , n9098 );
xnor ( n9100 , n9084 , n9099 );
xor ( n9101 , n9058 , n9100 );
or ( n9102 , n8651 , n8672 );
or ( n9103 , n8632 , n8650 );
nand ( n9104 , n9102 , n9103 );
xor ( n9105 , n9101 , n9104 );
or ( n9106 , n8689 , n8693 );
or ( n9107 , n8677 , n8688 );
nand ( n9108 , n9106 , n9107 );
xnor ( n9109 , n9105 , n9108 );
and ( n9110 , n8674 , n8694 );
and ( n9111 , n8629 , n8673 );
nor ( n9112 , n9110 , n9111 );
or ( n9113 , n9109 , n9112 , n1 );
not ( n9114 , n4562 );
xor ( n9115 , n8779 , n8784 );
and ( n9116 , n9115 , n8789 );
and ( n9117 , n8779 , n8784 );
or ( n9118 , n9116 , n9117 );
and ( n9119 , n8711 , n8778 );
not ( n9120 , n8700 );
nor ( n9121 , n9120 , n8707 );
nor ( n9122 , n9119 , n9121 );
not ( n9123 , n8718 );
not ( n9124 , n8717 );
or ( n9125 , n9123 , n9124 );
nand ( n9126 , n8719 , n8727 );
nand ( n9127 , n9125 , n9126 );
not ( n9128 , n8724 );
not ( n9129 , n2541 );
or ( n9130 , n9128 , n9129 );
and ( n9131 , n40 , n53 );
not ( n9132 , n40 );
and ( n9133 , n9132 , n4615 );
nor ( n9134 , n9131 , n9133 );
nand ( n9135 , n2550 , n9134 );
nand ( n9136 , n9130 , n9135 );
not ( n9137 , n9136 );
and ( n9138 , n2564 , n8757 );
and ( n9139 , n304 , n4577 );
and ( n9140 , n38 , n55 );
nor ( n9141 , n9139 , n9140 );
and ( n9142 , n6069 , n9141 );
nor ( n9143 , n9138 , n9142 );
not ( n9144 , n9143 );
and ( n9145 , n9137 , n9144 );
not ( n9146 , n9137 );
and ( n9147 , n9146 , n9143 );
nor ( n9148 , n9145 , n9147 );
xor ( n9149 , n9127 , n9148 );
not ( n9150 , n8770 );
not ( n9151 , n2722 );
or ( n9152 , n9150 , n9151 );
nand ( n9153 , n42 , n2715 );
nand ( n9154 , n9152 , n9153 );
xnor ( n9155 , n9154 , n8466 );
or ( n9156 , n2678 , n8715 );
or ( n9157 , n36 , n57 );
nand ( n9158 , n36 , n57 );
nand ( n9159 , n9157 , n9158 );
or ( n9160 , n2776 , n9159 );
nand ( n9161 , n9156 , n9160 );
xor ( n9162 , n9155 , n9161 );
or ( n9163 , n8765 , n8772 );
or ( n9164 , n8759 , n8760 );
nand ( n9165 , n9163 , n9164 );
xor ( n9166 , n9162 , n9165 );
xor ( n9167 , n9149 , n9166 );
not ( n9168 , n9167 );
not ( n9169 , n8777 );
not ( n9170 , n8747 );
or ( n9171 , n9169 , n9170 );
not ( n9172 , n8773 );
nand ( n9173 , n9172 , n8752 );
nand ( n9174 , n9171 , n9173 );
not ( n9175 , n8738 );
not ( n9176 , n9175 );
not ( n9177 , n8533 );
and ( n9178 , n9176 , n9177 );
not ( n9179 , n8743 );
and ( n9180 , n9179 , n8731 );
nor ( n9181 , n9178 , n9180 );
xor ( n9182 , n9174 , n9181 );
not ( n9183 , n9182 );
or ( n9184 , n9168 , n9183 );
or ( n9185 , n9182 , n9167 );
nand ( n9186 , n9184 , n9185 );
nand ( n9187 , n9122 , n9186 );
or ( n9188 , n9122 , n9186 );
and ( n9189 , n9187 , n9188 );
xnor ( n9190 , n9118 , n9189 );
not ( n9191 , n9190 );
or ( n9192 , n9114 , n9191 );
not ( n9193 , n2722 );
not ( n9194 , n570 );
or ( n9195 , n9193 , n9194 );
nand ( n9196 , n9195 , n9153 );
xor ( n9197 , n9196 , n8369 );
and ( n9198 , n663 , n4528 );
and ( n9199 , n2641 , n374 );
and ( n9200 , n3840 , n36 );
nor ( n9201 , n9199 , n9200 );
and ( n9202 , n9201 , n2682 );
nor ( n9203 , n9198 , n9202 );
xor ( n9204 , n9197 , n9203 );
not ( n9205 , n8846 );
or ( n9206 , n9205 , n8854 );
or ( n9207 , n8842 , n8760 );
nand ( n9208 , n9206 , n9207 );
xor ( n9209 , n9204 , n9208 );
or ( n9210 , n8830 , n8820 );
not ( n9211 , n8825 );
or ( n9212 , n9211 , n749 );
nand ( n9213 , n9210 , n9212 );
not ( n9214 , n8852 );
or ( n9215 , n561 , n9214 );
xnor ( n9216 , n2701 , n38 );
or ( n9217 , n9216 , n8239 );
nand ( n9218 , n9215 , n9217 );
not ( n9219 , n9218 );
not ( n9220 , n8203 );
not ( n9221 , n9220 );
not ( n9222 , n641 );
and ( n9223 , n9221 , n9222 );
and ( n9224 , n4504 , n427 );
not ( n9225 , n4504 );
and ( n9226 , n9225 , n40 );
nor ( n9227 , n9224 , n9226 );
and ( n9228 , n9227 , n2550 );
nor ( n9229 , n9223 , n9228 );
not ( n9230 , n9229 );
not ( n9231 , n9230 );
or ( n9232 , n9219 , n9231 );
or ( n9233 , n9230 , n9218 );
nand ( n9234 , n9232 , n9233 );
xor ( n9235 , n9213 , n9234 );
xnor ( n9236 , n9209 , n9235 );
not ( n9237 , n8816 );
and ( n9238 , n9237 , n8831 );
and ( n9239 , n8810 , n8327 );
nor ( n9240 , n9238 , n9239 );
xor ( n9241 , n9236 , n9240 );
and ( n9242 , n8835 , n8862 );
and ( n9243 , n8858 , n8861 );
nor ( n9244 , n9242 , n9243 );
not ( n9245 , n9244 );
xor ( n9246 , n9241 , n9245 );
and ( n9247 , n8872 , n8804 );
and ( n9248 , n8867 , n8871 );
nor ( n9249 , n9247 , n9248 );
xor ( n9250 , n9246 , n9249 );
not ( n9251 , n8876 );
nor ( n9252 , n9251 , n8890 );
xor ( n9253 , n9250 , n9252 );
and ( n9254 , n9253 , n2 );
nor ( n9255 , n9254 , n2526 );
nand ( n9256 , n9192 , n9255 );
not ( n9257 , n9109 );
not ( n9258 , n9112 );
or ( n9259 , n9257 , n9258 );
nand ( n9260 , n9259 , n2526 );
nand ( n9261 , n9256 , n9260 );
nand ( n9262 , n9113 , n9261 );
and ( n9263 , n9048 , n9262 );
not ( n9264 , n9048 );
not ( n9265 , n9262 );
and ( n9266 , n9264 , n9265 );
nor ( n9267 , n9263 , n9266 );
nor ( n9268 , n8938 , n8939 );
not ( n9269 , n9268 );
nand ( n9270 , n8942 , n9045 , n9267 , n9269 );
xor ( n9271 , n9236 , n9240 );
not ( n9272 , n9244 );
and ( n9273 , n9271 , n9272 );
and ( n9274 , n9236 , n9240 );
or ( n9275 , n9273 , n9274 );
and ( n9276 , n4528 , n9201 );
and ( n9277 , n460 , n2682 );
nor ( n9278 , n9276 , n9277 );
buf ( n9279 , n3274 );
and ( n9280 , n9278 , n9279 );
not ( n9281 , n9278 );
not ( n9282 , n9279 );
and ( n9283 , n9281 , n9282 );
nor ( n9284 , n9280 , n9283 );
not ( n9285 , n9220 );
and ( n9286 , n9285 , n9227 );
and ( n9287 , n429 , n2550 );
nor ( n9288 , n9286 , n9287 );
xor ( n9289 , n9284 , n9288 );
or ( n9290 , n9197 , n9203 );
not ( n9291 , n2986 );
not ( n9292 , n624 );
and ( n9293 , n9291 , n9292 );
not ( n9294 , n9153 );
nor ( n9295 , n9293 , n9294 );
or ( n9296 , n9295 , n8369 );
nand ( n9297 , n9290 , n9296 );
xnor ( n9298 , n9289 , n9297 );
and ( n9299 , n36 , n595 );
and ( n9300 , n9299 , n9230 );
not ( n9301 , n9299 );
and ( n9302 , n9301 , n9229 );
nor ( n9303 , n9300 , n9302 );
or ( n9304 , n9216 , n9214 );
or ( n9305 , n419 , n8239 );
nand ( n9306 , n9304 , n9305 );
xor ( n9307 , n9303 , n9306 );
xor ( n9308 , n9298 , n9307 );
and ( n9309 , n9213 , n9234 );
and ( n9310 , n9218 , n9229 );
nor ( n9311 , n9309 , n9310 );
xnor ( n9312 , n9308 , n9311 );
and ( n9313 , n9209 , n9235 );
and ( n9314 , n9204 , n9208 );
nor ( n9315 , n9313 , n9314 );
xor ( n9316 , n9312 , n9315 );
xor ( n9317 , n9275 , n9316 );
not ( n9318 , n9317 );
not ( n9319 , n9318 );
xor ( n9320 , n9246 , n9249 );
and ( n9321 , n9320 , n9252 );
and ( n9322 , n9246 , n9249 );
or ( n9323 , n9321 , n9322 );
buf ( n9324 , n9323 );
not ( n9325 , n9324 );
or ( n9326 , n9319 , n9325 );
or ( n9327 , n9324 , n9318 );
nand ( n9328 , n9326 , n9327 );
and ( n9329 , n9328 , n2 );
nor ( n9330 , n9329 , n2526 );
not ( n9331 , n9330 );
not ( n9332 , n9167 );
or ( n9333 , n9332 , n9182 );
not ( n9334 , n9174 );
or ( n9335 , n9334 , n9181 );
nand ( n9336 , n9333 , n9335 );
not ( n9337 , n9154 );
not ( n9338 , n9337 );
not ( n9339 , n8466 );
and ( n9340 , n9338 , n9339 );
and ( n9341 , n9155 , n9161 );
nor ( n9342 , n9340 , n9341 );
and ( n9343 , n2564 , n9141 );
xor ( n9344 , n38 , n54 );
and ( n9345 , n6069 , n9344 );
nor ( n9346 , n9343 , n9345 );
not ( n9347 , n9346 );
not ( n9348 , n9347 );
and ( n9349 , n8714 , n9136 );
not ( n9350 , n8714 );
and ( n9351 , n9350 , n9137 );
or ( n9352 , n9349 , n9351 );
not ( n9353 , n9352 );
or ( n9354 , n9348 , n9353 );
or ( n9355 , n9352 , n9347 );
nand ( n9356 , n9354 , n9355 );
xor ( n9357 , n9342 , n9356 );
not ( n9358 , n9159 );
not ( n9359 , n9358 );
not ( n9360 , n2818 );
or ( n9361 , n9359 , n9360 );
or ( n9362 , n36 , n56 );
nand ( n9363 , n36 , n56 );
and ( n9364 , n9362 , n9363 );
nand ( n9365 , n3011 , n9364 );
nand ( n9366 , n9361 , n9365 );
and ( n9367 , n9366 , n9282 );
not ( n9368 , n9366 );
and ( n9369 , n9368 , n9279 );
nor ( n9370 , n9367 , n9369 );
and ( n9371 , n3043 , n9134 );
and ( n9372 , n427 , n4666 );
and ( n9373 , n40 , n52 );
nor ( n9374 , n9372 , n9373 );
and ( n9375 , n2550 , n9374 );
nor ( n9376 , n9371 , n9375 );
xnor ( n9377 , n9370 , n9376 );
xor ( n9378 , n9357 , n9377 );
and ( n9379 , n9127 , n9148 );
and ( n9380 , n9137 , n9144 );
nor ( n9381 , n9379 , n9380 );
xor ( n9382 , n9378 , n9381 );
and ( n9383 , n9149 , n9166 );
and ( n9384 , n9162 , n9165 );
nor ( n9385 , n9383 , n9384 );
xnor ( n9386 , n9382 , n9385 );
xnor ( n9387 , n9336 , n9386 );
not ( n9388 , n9387 );
nand ( n9389 , n9118 , n9188 );
nand ( n9390 , n9389 , n9187 );
not ( n9391 , n9390 );
or ( n9392 , n9388 , n9391 );
or ( n9393 , n9390 , n9387 );
nand ( n9394 , n9392 , n9393 );
nand ( n9395 , n9394 , n4562 );
not ( n9396 , n9395 );
or ( n9397 , n9331 , n9396 );
or ( n9398 , n9058 , n9100 );
or ( n9399 , n9051 , n9057 );
nand ( n9400 , n9398 , n9399 );
not ( n9401 , n9056 );
not ( n9402 , n9055 );
or ( n9403 , n9401 , n9402 );
or ( n9404 , n8683 , n7173 );
nand ( n9405 , n9403 , n9404 );
and ( n9406 , n6638 , n9088 );
and ( n9407 , n6630 , n6502 );
and ( n9408 , n71 , n88 );
nor ( n9409 , n9407 , n9408 );
and ( n9410 , n6644 , n9409 );
nor ( n9411 , n9406 , n9410 );
xnor ( n9412 , n9411 , n8635 );
and ( n9413 , n6527 , n9062 );
and ( n9414 , n6528 , n6578 );
and ( n9415 , n69 , n90 );
nor ( n9416 , n9414 , n9415 );
and ( n9417 , n6534 , n9416 );
nor ( n9418 , n9413 , n9417 );
not ( n9419 , n9418 );
and ( n9420 , n9412 , n9419 );
not ( n9421 , n9412 );
and ( n9422 , n9421 , n9418 );
nor ( n9423 , n9420 , n9422 );
xor ( n9424 , n9405 , n9423 );
not ( n9425 , n9424 );
and ( n9426 , n9084 , n9099 );
and ( n9427 , n9079 , n9083 );
nor ( n9428 , n9426 , n9427 );
not ( n9429 , n9428 );
or ( n9430 , n9425 , n9429 );
or ( n9431 , n9428 , n9424 );
nand ( n9432 , n9430 , n9431 );
xnor ( n9433 , n9400 , n9432 );
not ( n9434 , n9078 );
not ( n9435 , n9071 );
or ( n9436 , n9434 , n9435 );
or ( n9437 , n9064 , n9070 );
nand ( n9438 , n9436 , n9437 );
and ( n9439 , n6445 , n9068 );
and ( n9440 , n6446 , n6431 );
and ( n9441 , n73 , n86 );
nor ( n9442 , n9440 , n9441 );
and ( n9443 , n6452 , n9442 );
nor ( n9444 , n9439 , n9443 );
not ( n9445 , n9444 );
or ( n9446 , n7049 , n9076 );
or ( n9447 , n75 , n84 );
nand ( n9448 , n75 , n84 );
nand ( n9449 , n9447 , n9448 );
or ( n9450 , n6665 , n9449 );
nand ( n9451 , n9446 , n9450 );
not ( n9452 , n9451 );
and ( n9453 , n9445 , n9452 );
and ( n9454 , n9444 , n9451 );
nor ( n9455 , n9453 , n9454 );
and ( n9456 , n6467 , n9096 );
and ( n9457 , n7152 , n92 );
nor ( n9458 , n9456 , n9457 );
xor ( n9459 , n9455 , n9458 );
xor ( n9460 , n9438 , n9459 );
or ( n9461 , n9091 , n9098 );
or ( n9462 , n9090 , n7630 );
nand ( n9463 , n9461 , n9462 );
xor ( n9464 , n9460 , n9463 );
and ( n9465 , n9433 , n9464 );
or ( n9466 , n9433 , n9464 );
nand ( n9467 , n9466 , n2526 );
nor ( n9468 , n9465 , n9467 );
and ( n9469 , n9105 , n9108 );
and ( n9470 , n9101 , n9104 );
nor ( n9471 , n9469 , n9470 );
and ( n9472 , n9468 , n9471 );
nor ( n9473 , n9468 , n9471 , n1 );
nor ( n9474 , n9472 , n9473 );
nand ( n9475 , n9397 , n9474 );
not ( n9476 , n9475 );
not ( n9477 , n9476 );
and ( n9478 , n9261 , n9047 );
not ( n9479 , n9478 );
not ( n9480 , n8902 );
or ( n9481 , n9479 , n9480 );
nand ( n9482 , n9481 , n9113 );
not ( n9483 , n9482 );
or ( n9484 , n9477 , n9483 );
or ( n9485 , n9476 , n9482 );
nand ( n9486 , n9484 , n9485 );
nor ( n9487 , n9270 , n9486 );
not ( n9488 , n9478 );
not ( n9489 , n8902 );
or ( n9490 , n9488 , n9489 );
not ( n9491 , n9473 );
and ( n9492 , n9491 , n9113 );
nand ( n9493 , n9490 , n9492 );
or ( n9494 , n9455 , n9458 );
not ( n9495 , n9451 );
or ( n9496 , n9444 , n9495 );
nand ( n9497 , n9494 , n9496 );
and ( n9498 , n9497 , n9419 );
not ( n9499 , n9497 );
and ( n9500 , n9499 , n9418 );
nor ( n9501 , n9498 , n9500 );
or ( n9502 , n7049 , n9449 );
or ( n9503 , n74 , n84 );
nand ( n9504 , n74 , n84 );
nand ( n9505 , n9503 , n9504 );
or ( n9506 , n7171 , n9505 );
nand ( n9507 , n9502 , n9506 );
xnor ( n9508 , n9507 , n9074 );
and ( n9509 , n6638 , n9409 );
and ( n9510 , n6630 , n6554 );
and ( n9511 , n70 , n88 );
nor ( n9512 , n9510 , n9511 );
and ( n9513 , n6644 , n9512 );
nor ( n9514 , n9509 , n9513 );
xor ( n9515 , n9508 , n9514 );
xor ( n9516 , n9501 , n9515 );
and ( n9517 , n6527 , n9416 );
and ( n9518 , n6528 , n6741 );
and ( n9519 , n68 , n90 );
nor ( n9520 , n9518 , n9519 );
and ( n9521 , n6534 , n9520 );
nor ( n9522 , n9517 , n9521 );
xor ( n9523 , n9522 , n7473 );
and ( n9524 , n6445 , n9442 );
and ( n9525 , n6446 , n6496 );
and ( n9526 , n72 , n86 );
nor ( n9527 , n9525 , n9526 );
and ( n9528 , n6452 , n9527 );
nor ( n9529 , n9524 , n9528 );
xor ( n9530 , n9523 , n9529 );
or ( n9531 , n9412 , n9419 );
or ( n9532 , n9411 , n8635 );
nand ( n9533 , n9531 , n9532 );
xor ( n9534 , n9530 , n9533 );
xnor ( n9535 , n9516 , n9534 );
xor ( n9536 , n9438 , n9459 );
and ( n9537 , n9536 , n9463 );
and ( n9538 , n9438 , n9459 );
nor ( n9539 , n9537 , n9538 );
xnor ( n9540 , n9535 , n9539 );
not ( n9541 , n9428 );
and ( n9542 , n9541 , n9424 );
and ( n9543 , n9405 , n9423 );
nor ( n9544 , n9542 , n9543 );
xnor ( n9545 , n9540 , n9544 );
not ( n9546 , n9545 );
or ( n9547 , n9400 , n9432 );
not ( n9548 , n9467 );
nand ( n9549 , n9547 , n9548 );
nor ( n9550 , n9546 , n9549 );
not ( n9551 , n9550 );
not ( n9552 , n6416 );
or ( n9553 , n9336 , n9386 );
not ( n9554 , n9553 );
not ( n9555 , n9389 );
not ( n9556 , n9555 );
or ( n9557 , n9554 , n9556 );
not ( n9558 , n9386 );
not ( n9559 , n9336 );
or ( n9560 , n9558 , n9559 );
nand ( n9561 , n9560 , n9187 );
nand ( n9562 , n9553 , n9561 );
nand ( n9563 , n9557 , n9562 );
and ( n9564 , n9382 , n9385 );
and ( n9565 , n9378 , n9381 );
nor ( n9566 , n9564 , n9565 );
and ( n9567 , n2564 , n9344 );
and ( n9568 , n4652 , n4615 );
and ( n9569 , n38 , n53 );
nor ( n9570 , n9568 , n9569 );
and ( n9571 , n2573 , n9570 );
nor ( n9572 , n9567 , n9571 );
xor ( n9573 , n9158 , n9572 );
not ( n9574 , n9364 );
not ( n9575 , n2901 );
or ( n9576 , n9574 , n9575 );
not ( n9577 , n36 );
not ( n9578 , n55 );
and ( n9579 , n9577 , n9578 );
nand ( n9580 , n36 , n55 );
not ( n9581 , n9580 );
nor ( n9582 , n9579 , n9581 );
nand ( n9583 , n2682 , n9582 );
nand ( n9584 , n9576 , n9583 );
not ( n9585 , n9584 );
xor ( n9586 , n9573 , n9585 );
and ( n9587 , n8203 , n9374 );
nor ( n9588 , n2551 , n427 );
nor ( n9589 , n9587 , n9588 );
not ( n9590 , n9589 );
and ( n9591 , n9586 , n9590 );
not ( n9592 , n9586 );
and ( n9593 , n9592 , n9589 );
nor ( n9594 , n9591 , n9593 );
not ( n9595 , n9370 );
not ( n9596 , n9376 );
and ( n9597 , n9595 , n9596 );
and ( n9598 , n9366 , n9279 );
nor ( n9599 , n9597 , n9598 );
xnor ( n9600 , n9594 , n9599 );
and ( n9601 , n9352 , n9346 );
and ( n9602 , n9137 , n8714 );
nor ( n9603 , n9601 , n9602 );
xor ( n9604 , n9600 , n9603 );
xor ( n9605 , n9342 , n9356 );
and ( n9606 , n9605 , n9377 );
and ( n9607 , n9342 , n9356 );
nor ( n9608 , n9606 , n9607 );
xor ( n9609 , n9604 , n9608 );
nor ( n9610 , n9566 , n9609 );
and ( n9611 , n9566 , n9609 );
nor ( n9612 , n9610 , n9611 );
and ( n9613 , n9563 , n9612 );
not ( n9614 , n9563 );
not ( n9615 , n9612 );
and ( n9616 , n9614 , n9615 );
nor ( n9617 , n9613 , n9616 );
not ( n9618 , n9617 );
or ( n9619 , n9552 , n9618 );
or ( n9620 , n9323 , n9317 );
not ( n9621 , n9275 );
nand ( n9622 , n9621 , n9316 );
nand ( n9623 , n9620 , n9622 );
or ( n9624 , n9312 , n9315 );
or ( n9625 , n9308 , n9311 );
nand ( n9626 , n9624 , n9625 );
not ( n9627 , n9626 );
or ( n9628 , n9284 , n9288 );
or ( n9629 , n9278 , n9282 );
nand ( n9630 , n9628 , n9629 );
and ( n9631 , n429 , n9285 );
nor ( n9632 , n9631 , n9588 );
not ( n9633 , n9632 );
xnor ( n9634 , n9630 , n9633 );
and ( n9635 , n4528 , n509 );
and ( n9636 , n2595 , n374 );
nor ( n9637 , n2595 , n374 );
nor ( n9638 , n9636 , n9637 );
and ( n9639 , n9638 , n2682 );
nor ( n9640 , n9635 , n9639 );
not ( n9641 , n9640 );
and ( n9642 , n9200 , n9641 );
not ( n9643 , n9200 );
and ( n9644 , n9643 , n9640 );
nor ( n9645 , n9642 , n9644 );
not ( n9646 , n8239 );
not ( n9647 , n9646 );
or ( n9648 , n4504 , n38 );
not ( n9649 , n4504 );
or ( n9650 , n9649 , n304 );
nand ( n9651 , n9648 , n9650 );
not ( n9652 , n9651 );
or ( n9653 , n9647 , n9652 );
or ( n9654 , n419 , n9214 );
nand ( n9655 , n9653 , n9654 );
xor ( n9656 , n9645 , n9655 );
xnor ( n9657 , n9634 , n9656 );
and ( n9658 , n9303 , n9306 );
and ( n9659 , n9230 , n9299 );
nor ( n9660 , n9658 , n9659 );
xor ( n9661 , n9657 , n9660 );
or ( n9662 , n9298 , n9307 );
or ( n9663 , n9289 , n9297 );
nand ( n9664 , n9662 , n9663 );
xor ( n9665 , n9661 , n9664 );
not ( n9666 , n9665 );
or ( n9667 , n9627 , n9666 );
or ( n9668 , n9665 , n9626 );
nand ( n9669 , n9667 , n9668 );
xor ( n9670 , n9623 , n9669 );
and ( n9671 , n9670 , n4563 );
nor ( n9672 , n9545 , n1 );
nor ( n9673 , n9671 , n9672 );
nand ( n9674 , n9619 , n9673 );
nand ( n9675 , n9674 , n9549 );
nand ( n9676 , n9551 , n9675 );
nand ( n9677 , n9475 , n9491 );
nand ( n9678 , n9493 , n9676 , n9677 );
not ( n9679 , n9678 );
and ( n9680 , n9476 , n9482 );
not ( n9681 , n9676 );
nand ( n9682 , n9681 , n9491 );
nor ( n9683 , n9680 , n9682 );
nor ( n9684 , n9679 , n9683 );
and ( n9685 , n9487 , n9684 );
and ( n9686 , n9516 , n9534 );
and ( n9687 , n9530 , n9533 );
nor ( n9688 , n9686 , n9687 );
or ( n9689 , n7049 , n9505 );
or ( n9690 , n73 , n84 );
nand ( n9691 , n73 , n84 );
nand ( n9692 , n9690 , n9691 );
or ( n9693 , n7171 , n9692 );
nand ( n9694 , n9689 , n9693 );
not ( n9695 , n9448 );
xnor ( n9696 , n9694 , n9695 );
and ( n9697 , n6527 , n9520 );
and ( n9698 , n6534 , n90 );
nor ( n9699 , n9697 , n9698 );
xor ( n9700 , n9696 , n9699 );
or ( n9701 , n9523 , n9529 );
or ( n9702 , n9522 , n7474 );
nand ( n9703 , n9701 , n9702 );
xor ( n9704 , n9700 , n9703 );
not ( n9705 , n9508 );
not ( n9706 , n9514 );
and ( n9707 , n9705 , n9706 );
and ( n9708 , n9507 , n9074 );
nor ( n9709 , n9707 , n9708 );
and ( n9710 , n6445 , n9527 );
and ( n9711 , n6446 , n6502 );
and ( n9712 , n71 , n86 );
nor ( n9713 , n9711 , n9712 );
and ( n9714 , n6452 , n9713 );
nor ( n9715 , n9710 , n9714 );
and ( n9716 , n6638 , n9512 );
and ( n9717 , n6630 , n6578 );
and ( n9718 , n69 , n88 );
nor ( n9719 , n9717 , n9718 );
and ( n9720 , n6644 , n9719 );
nor ( n9721 , n9716 , n9720 );
and ( n9722 , n9715 , n9721 );
not ( n9723 , n9715 );
not ( n9724 , n9721 );
and ( n9725 , n9723 , n9724 );
nor ( n9726 , n9722 , n9725 );
xor ( n9727 , n9709 , n9726 );
xnor ( n9728 , n9704 , n9727 );
xnor ( n9729 , n9688 , n9728 );
and ( n9730 , n9501 , n9515 );
and ( n9731 , n9497 , n9419 );
nor ( n9732 , n9730 , n9731 );
and ( n9733 , n9729 , n9732 );
nor ( n9734 , n9729 , n9732 );
nor ( n9735 , n9733 , n9734 , n1 );
not ( n9736 , n9735 );
not ( n9737 , n9736 );
not ( n9738 , n9669 );
not ( n9739 , n9623 );
or ( n9740 , n9738 , n9739 );
not ( n9741 , n9665 );
nand ( n9742 , n9741 , n9626 );
nand ( n9743 , n9740 , n9742 );
xor ( n9744 , n9657 , n9660 );
and ( n9745 , n9744 , n9664 );
and ( n9746 , n9657 , n9660 );
nor ( n9747 , n9745 , n9746 );
and ( n9748 , n9634 , n9656 );
and ( n9749 , n9630 , n9632 );
nor ( n9750 , n9748 , n9749 );
and ( n9751 , n9651 , n8852 );
and ( n9752 , n307 , n9646 );
nor ( n9753 , n9751 , n9752 );
nand ( n9754 , n1914 , n36 );
and ( n9755 , n9754 , n3804 );
not ( n9756 , n9754 );
and ( n9757 , n9756 , n3805 );
nor ( n9758 , n9755 , n9757 );
xor ( n9759 , n9753 , n9758 );
xor ( n9760 , n9750 , n9759 );
and ( n9761 , n9645 , n9655 );
and ( n9762 , n9641 , n9200 );
nor ( n9763 , n9761 , n9762 );
and ( n9764 , n9638 , n4528 );
and ( n9765 , n377 , n2682 );
nor ( n9766 , n9764 , n9765 );
and ( n9767 , n9766 , n9633 );
not ( n9768 , n9766 );
and ( n9769 , n9768 , n9632 );
nor ( n9770 , n9767 , n9769 );
xnor ( n9771 , n9763 , n9770 );
xor ( n9772 , n9760 , n9771 );
xor ( n9773 , n9747 , n9772 );
and ( n9774 , n9743 , n9773 );
not ( n9775 , n9743 );
not ( n9776 , n9773 );
and ( n9777 , n9775 , n9776 );
nor ( n9778 , n9774 , n9777 );
nand ( n9779 , n9778 , n4563 );
not ( n9780 , n9553 );
nor ( n9781 , n9780 , n9610 );
not ( n9782 , n9781 );
not ( n9783 , n9555 );
or ( n9784 , n9782 , n9783 );
not ( n9785 , n9562 );
not ( n9786 , n9610 );
and ( n9787 , n9785 , n9786 );
nor ( n9788 , n9787 , n9611 );
nand ( n9789 , n9784 , n9788 );
and ( n9790 , n9604 , n9608 );
and ( n9791 , n9600 , n9603 );
nor ( n9792 , n9790 , n9791 );
xor ( n9793 , n9158 , n9572 );
not ( n9794 , n9584 );
and ( n9795 , n9793 , n9794 );
and ( n9796 , n9158 , n9572 );
or ( n9797 , n9795 , n9796 );
and ( n9798 , n4528 , n9582 );
and ( n9799 , n374 , n6021 );
nor ( n9800 , n374 , n6021 );
nor ( n9801 , n9799 , n9800 );
and ( n9802 , n2682 , n9801 );
nor ( n9803 , n9798 , n9802 );
and ( n9804 , n9803 , n9589 );
not ( n9805 , n9803 );
and ( n9806 , n9805 , n9590 );
nor ( n9807 , n9804 , n9806 );
xnor ( n9808 , n9797 , n9807 );
and ( n9809 , n8852 , n9570 );
and ( n9810 , n304 , n4666 );
and ( n9811 , n38 , n52 );
nor ( n9812 , n9810 , n9811 );
and ( n9813 , n9646 , n9812 );
nor ( n9814 , n9809 , n9813 );
xnor ( n9815 , n9814 , n9363 );
or ( n9816 , n9815 , n3805 );
nand ( n9817 , n9815 , n3805 );
nand ( n9818 , n9816 , n9817 );
xor ( n9819 , n9808 , n9818 );
and ( n9820 , n9594 , n9599 );
and ( n9821 , n9590 , n9586 );
nor ( n9822 , n9820 , n9821 );
xnor ( n9823 , n9819 , n9822 );
xnor ( n9824 , n9792 , n9823 );
and ( n9825 , n9789 , n9824 );
not ( n9826 , n9789 );
not ( n9827 , n9824 );
and ( n9828 , n9826 , n9827 );
nor ( n9829 , n9825 , n9828 );
nand ( n9830 , n9829 , n6416 );
or ( n9831 , n9540 , n9544 );
or ( n9832 , n9539 , n9535 );
nand ( n9833 , n9831 , n9832 , n2526 );
nand ( n9834 , n9779 , n9830 , n9833 );
not ( n9835 , n9834 );
not ( n9836 , n9835 );
or ( n9837 , n9737 , n9836 );
nand ( n9838 , n9834 , n9735 );
nand ( n9839 , n9837 , n9838 );
not ( n9840 , n9839 );
or ( n9841 , n9549 , n9545 );
nand ( n9842 , n9678 , n9841 );
not ( n9843 , n9842 );
or ( n9844 , n9840 , n9843 );
nand ( n9845 , n9835 , n9735 );
nand ( n9846 , n9844 , n9845 );
or ( n9847 , n9688 , n9728 );
not ( n9848 , n9734 );
nand ( n9849 , n9847 , n9848 );
and ( n9850 , n6638 , n9719 );
and ( n9851 , n6438 , n6741 );
and ( n9852 , n68 , n88 );
nor ( n9853 , n9851 , n9852 );
and ( n9854 , n6644 , n9853 );
nor ( n9855 , n9850 , n9854 );
xor ( n9856 , n9855 , n7223 );
or ( n9857 , n7049 , n9692 );
or ( n9858 , n72 , n84 );
nand ( n9859 , n72 , n84 );
nand ( n9860 , n9858 , n9859 );
or ( n9861 , n7171 , n9860 );
nand ( n9862 , n9857 , n9861 );
xnor ( n9863 , n9856 , n9862 );
not ( n9864 , n9696 );
not ( n9865 , n9699 );
and ( n9866 , n9864 , n9865 );
and ( n9867 , n9694 , n9695 );
nor ( n9868 , n9866 , n9867 );
xor ( n9869 , n9863 , n9868 );
not ( n9870 , n9724 );
not ( n9871 , n9504 );
and ( n9872 , n9870 , n9871 );
and ( n9873 , n9724 , n9504 );
nor ( n9874 , n9872 , n9873 );
and ( n9875 , n6445 , n9713 );
and ( n9876 , n6446 , n6554 );
and ( n9877 , n70 , n86 );
nor ( n9878 , n9876 , n9877 );
and ( n9879 , n6452 , n9878 );
nor ( n9880 , n9875 , n9879 );
xnor ( n9881 , n9874 , n9880 );
xnor ( n9882 , n9869 , n9881 );
or ( n9883 , n9709 , n9726 );
or ( n9884 , n9715 , n9724 );
nand ( n9885 , n9883 , n9884 );
xor ( n9886 , n9882 , n9885 );
and ( n9887 , n9704 , n9727 );
and ( n9888 , n9700 , n9703 );
nor ( n9889 , n9887 , n9888 );
not ( n9890 , n9889 );
xor ( n9891 , n9886 , n9890 );
nand ( n9892 , n9849 , n9891 , n2526 );
not ( n9893 , n9637 );
and ( n9894 , n307 , n8852 );
nor ( n9895 , n8239 , n304 );
nor ( n9896 , n9894 , n9895 );
and ( n9897 , n9893 , n9896 );
not ( n9898 , n9893 );
not ( n9899 , n9896 );
and ( n9900 , n9898 , n9899 );
nor ( n9901 , n9897 , n9900 );
and ( n9902 , n393 , n4528 );
xor ( n9903 , n36 , n9649 );
and ( n9904 , n9903 , n2682 );
nor ( n9905 , n9902 , n9904 );
xnor ( n9906 , n9901 , n9905 );
not ( n9907 , n9906 );
and ( n9908 , n9753 , n9758 );
and ( n9909 , n9754 , n3804 );
nor ( n9910 , n9908 , n9909 );
not ( n9911 , n9910 );
and ( n9912 , n9907 , n9911 );
and ( n9913 , n9906 , n9910 );
nor ( n9914 , n9912 , n9913 );
or ( n9915 , n9763 , n9770 );
or ( n9916 , n9766 , n9632 );
nand ( n9917 , n9915 , n9916 );
xor ( n9918 , n9914 , n9917 );
xor ( n9919 , n9750 , n9759 );
and ( n9920 , n9919 , n9771 );
and ( n9921 , n9750 , n9759 );
nor ( n9922 , n9920 , n9921 );
xor ( n9923 , n9918 , n9922 );
or ( n9924 , n9743 , n9773 );
not ( n9925 , n9747 );
nand ( n9926 , n9925 , n9772 );
nand ( n9927 , n9924 , n9926 );
xor ( n9928 , n9923 , n9927 );
nand ( n9929 , n9928 , n4563 );
and ( n9930 , n9819 , n9822 );
and ( n9931 , n9808 , n9818 );
nor ( n9932 , n9930 , n9931 );
and ( n9933 , n9797 , n9807 );
and ( n9934 , n9803 , n9589 );
nor ( n9935 , n9933 , n9934 );
and ( n9936 , n8852 , n9812 );
nor ( n9937 , n9936 , n9895 );
not ( n9938 , n9937 );
not ( n9939 , n9801 );
or ( n9940 , n2678 , n9939 );
and ( n9941 , n4615 , n36 );
and ( n9942 , n374 , n53 );
nor ( n9943 , n9941 , n9942 );
or ( n9944 , n8481 , n9943 );
nand ( n9945 , n9940 , n9944 );
not ( n9946 , n9945 );
not ( n9947 , n9580 );
and ( n9948 , n9946 , n9947 );
and ( n9949 , n9945 , n9580 );
nor ( n9950 , n9948 , n9949 );
not ( n9951 , n9950 );
or ( n9952 , n9938 , n9951 );
or ( n9953 , n9950 , n9937 );
nand ( n9954 , n9952 , n9953 );
xor ( n9955 , n9935 , n9954 );
or ( n9956 , n9815 , n3804 );
or ( n9957 , n9814 , n9363 );
nand ( n9958 , n9956 , n9957 );
xnor ( n9959 , n9955 , n9958 );
nor ( n9960 , n9932 , n9959 );
not ( n9961 , n9960 );
nand ( n9962 , n9932 , n9959 );
nand ( n9963 , n9961 , n9962 );
not ( n9964 , n9963 );
nand ( n9965 , n9792 , n9823 );
and ( n9966 , n9118 , n9781 , n9188 , n9965 );
not ( n9967 , n9966 );
or ( n9968 , n9792 , n9823 );
nand ( n9969 , n9968 , n9788 );
nand ( n9970 , n9965 , n9969 );
nand ( n9971 , n9967 , n9970 );
not ( n9972 , n9971 );
or ( n9973 , n9964 , n9972 );
not ( n9974 , n9970 );
nor ( n9975 , n9974 , n9960 );
nand ( n9976 , n9967 , n9975 );
nand ( n9977 , n9973 , n9976 );
or ( n9978 , n9962 , n9971 );
nand ( n9979 , n9977 , n9978 , n6416 );
or ( n9980 , n9849 , n9891 );
nand ( n9981 , n9980 , n2526 );
nand ( n9982 , n9929 , n9979 , n9981 );
nand ( n9983 , n9892 , n9982 );
buf ( n9984 , n9983 );
not ( n9985 , n9984 );
and ( n9986 , n9846 , n9985 );
not ( n9987 , n9846 );
and ( n9988 , n9987 , n9984 );
nor ( n9989 , n9986 , n9988 );
buf ( n9990 , n9842 );
and ( n9991 , n9990 , n9839 );
not ( n9992 , n9990 );
not ( n9993 , n9839 );
and ( n9994 , n9992 , n9993 );
nor ( n9995 , n9991 , n9994 );
nand ( n9996 , n9685 , n9989 , n9995 );
and ( n9997 , n9835 , n9735 );
nand ( n9998 , n9841 , n9892 );
nor ( n9999 , n9997 , n9998 );
not ( n10000 , n9999 );
not ( n10001 , n9678 );
or ( n10002 , n10000 , n10001 );
nand ( n10003 , n9834 , n9892 , n9736 );
and ( n10004 , n9982 , n10003 );
nand ( n10005 , n10002 , n10004 );
buf ( n10006 , n10005 );
not ( n10007 , n9918 );
not ( n10008 , n9922 );
or ( n10009 , n10007 , n10008 );
or ( n10010 , n9922 , n9918 );
nand ( n10011 , n10009 , n10010 );
not ( n10012 , n10011 );
not ( n10013 , n9927 );
or ( n10014 , n10012 , n10013 );
not ( n10015 , n9922 );
nand ( n10016 , n10015 , n9918 );
nand ( n10017 , n10014 , n10016 );
not ( n10018 , n9914 );
nand ( n10019 , n10018 , n9917 );
not ( n10020 , n9906 );
nand ( n10021 , n10020 , n9910 );
and ( n10022 , n10019 , n10021 );
or ( n10023 , n9901 , n9905 );
or ( n10024 , n9899 , n9893 );
nand ( n10025 , n10023 , n10024 );
not ( n10026 , n9903 );
not ( n10027 , n4528 );
or ( n10028 , n10026 , n10027 );
or ( n10029 , n475 , n8481 );
nand ( n10030 , n10028 , n10029 );
and ( n10031 , n376 , n3992 );
not ( n10032 , n376 );
and ( n10033 , n10032 , n3991 );
nor ( n10034 , n10031 , n10033 );
xor ( n10035 , n10030 , n10034 );
or ( n10036 , n10035 , n9896 );
nand ( n10037 , n10035 , n9896 );
nand ( n10038 , n10036 , n10037 );
xnor ( n10039 , n10025 , n10038 );
xnor ( n10040 , n10022 , n10039 );
not ( n10041 , n10040 );
xor ( n10042 , n10017 , n10041 );
or ( n10043 , n10042 , n4562 );
and ( n10044 , n9955 , n9958 );
and ( n10045 , n9935 , n9954 );
nor ( n10046 , n10044 , n10045 );
or ( n10047 , n2678 , n9943 );
and ( n10048 , n4666 , n36 );
and ( n10049 , n374 , n52 );
nor ( n10050 , n10048 , n10049 );
or ( n10051 , n8481 , n10050 );
nand ( n10052 , n10047 , n10051 );
xor ( n10053 , n10052 , n9800 );
xnor ( n10054 , n10053 , n3991 );
not ( n10055 , n9945 );
and ( n10056 , n10055 , n9937 , n9580 );
nor ( n10057 , n10055 , n9937 , n9580 );
nor ( n10058 , n10056 , n10057 );
xnor ( n10059 , n10054 , n10058 );
nor ( n10060 , n10046 , n10059 );
not ( n10061 , n10060 );
nand ( n10062 , n10046 , n10059 );
and ( n10063 , n10062 , n9962 );
nand ( n10064 , n10061 , n10063 );
and ( n10065 , n10064 , n6416 );
nand ( n10066 , n9976 , n10065 , n9962 );
nand ( n10067 , n10043 , n10066 );
not ( n10068 , n10060 );
nand ( n10069 , n10068 , n10062 );
or ( n10070 , n9976 , n10069 , n7762 );
xor ( n10071 , n9882 , n9885 );
not ( n10072 , n9889 );
and ( n10073 , n10071 , n10072 );
and ( n10074 , n9882 , n9885 );
or ( n10075 , n10073 , n10074 );
not ( n10076 , n10075 );
nor ( n10077 , n10076 , n1 );
not ( n10078 , n9862 );
not ( n10079 , n9856 );
or ( n10080 , n10078 , n10079 );
or ( n10081 , n9855 , n7223 );
nand ( n10082 , n10080 , n10081 );
and ( n10083 , n6638 , n9853 );
and ( n10084 , n6644 , n88 );
nor ( n10085 , n10083 , n10084 );
and ( n10086 , n10082 , n10085 );
not ( n10087 , n10082 );
not ( n10088 , n10085 );
and ( n10089 , n10087 , n10088 );
nor ( n10090 , n10086 , n10089 );
or ( n10091 , n7049 , n9860 );
or ( n10092 , n71 , n84 );
nand ( n10093 , n71 , n84 );
nand ( n10094 , n10092 , n10093 );
or ( n10095 , n7171 , n10094 );
nand ( n10096 , n10091 , n10095 );
not ( n10097 , n10096 );
not ( n10098 , n9691 );
and ( n10099 , n10097 , n10098 );
and ( n10100 , n10096 , n9691 );
nor ( n10101 , n10099 , n10100 );
and ( n10102 , n6445 , n9878 );
and ( n10103 , n6446 , n6578 );
and ( n10104 , n69 , n86 );
nor ( n10105 , n10103 , n10104 );
and ( n10106 , n6452 , n10105 );
nor ( n10107 , n10102 , n10106 );
xor ( n10108 , n10101 , n10107 );
xor ( n10109 , n10090 , n10108 );
or ( n10110 , n9874 , n9880 );
or ( n10111 , n9721 , n9504 );
nand ( n10112 , n10110 , n10111 );
xnor ( n10113 , n10109 , n10112 );
and ( n10114 , n9869 , n9881 );
and ( n10115 , n9868 , n9863 );
nor ( n10116 , n10114 , n10115 );
xor ( n10117 , n10113 , n10116 );
and ( n10118 , n10077 , n10117 );
not ( n10119 , n10064 );
nor ( n10120 , n10119 , n10069 , n7762 );
nor ( n10121 , n10077 , n10117 , n1 );
nor ( n10122 , n10118 , n10120 , n10121 );
nand ( n10123 , n10070 , n10122 );
nor ( n10124 , n10067 , n10123 );
buf ( n10125 , n10124 );
not ( n10126 , n10125 );
and ( n10127 , n10006 , n10126 );
not ( n10128 , n10006 );
and ( n10129 , n10128 , n10125 );
nor ( n10130 , n10127 , n10129 );
nor ( n10131 , n9996 , n10130 );
or ( n10132 , n10005 , n10124 );
not ( n10133 , n10117 );
nand ( n10134 , n10133 , n10077 );
nand ( n10135 , n10132 , n10134 );
buf ( n10136 , n10135 );
not ( n10137 , n10136 );
or ( n10138 , n10113 , n10116 );
or ( n10139 , n10112 , n10109 );
nand ( n10140 , n10138 , n10139 , n2526 );
not ( n10141 , n10140 );
and ( n10142 , n10090 , n10108 );
and ( n10143 , n10082 , n10085 );
nor ( n10144 , n10142 , n10143 );
or ( n10145 , n10101 , n10107 );
not ( n10146 , n10096 );
or ( n10147 , n10146 , n9691 );
nand ( n10148 , n10145 , n10147 );
or ( n10149 , n7049 , n10094 );
or ( n10150 , n70 , n84 );
nand ( n10151 , n70 , n84 );
nand ( n10152 , n10150 , n10151 );
or ( n10153 , n7171 , n10152 );
nand ( n10154 , n10149 , n10153 );
and ( n10155 , n10154 , n10088 );
not ( n10156 , n10154 );
and ( n10157 , n10156 , n10085 );
nor ( n10158 , n10155 , n10157 );
xnor ( n10159 , n10148 , n10158 );
and ( n10160 , n6445 , n10105 );
and ( n10161 , n6446 , n6741 );
and ( n10162 , n68 , n86 );
nor ( n10163 , n10161 , n10162 );
and ( n10164 , n6452 , n10163 );
nor ( n10165 , n10160 , n10164 );
xor ( n10166 , n6946 , n9859 );
xor ( n10167 , n10165 , n10166 );
xor ( n10168 , n10159 , n10167 );
xor ( n10169 , n10144 , n10168 );
nand ( n10170 , n10141 , n10169 );
or ( n10171 , n10017 , n10040 );
or ( n10172 , n10022 , n10039 );
nand ( n10173 , n10171 , n10172 );
or ( n10174 , n2678 , n475 );
nand ( n10175 , n2682 , n36 );
nand ( n10176 , n10174 , n10175 );
and ( n10177 , n36 , n9649 );
nor ( n10178 , n10176 , n10177 );
not ( n10179 , n10178 );
nand ( n10180 , n10176 , n10177 );
nand ( n10181 , n10179 , n10180 );
not ( n10182 , n10181 );
and ( n10183 , n10030 , n10034 );
and ( n10184 , n376 , n3992 );
nor ( n10185 , n10183 , n10184 );
not ( n10186 , n10185 );
or ( n10187 , n10182 , n10186 );
or ( n10188 , n10185 , n10181 );
nand ( n10189 , n10187 , n10188 );
and ( n10190 , n10025 , n10038 );
and ( n10191 , n10035 , n9899 );
nor ( n10192 , n10190 , n10191 );
xnor ( n10193 , n10189 , n10192 );
xnor ( n10194 , n10173 , n10193 );
or ( n10195 , n10194 , n4562 );
and ( n10196 , n10053 , n3992 );
and ( n10197 , n10052 , n9800 );
nor ( n10198 , n10196 , n10197 );
not ( n10199 , n10198 );
or ( n10200 , n2678 , n10050 );
nand ( n10201 , n10200 , n10175 );
not ( n10202 , n10201 );
nand ( n10203 , n36 , n53 );
nor ( n10204 , n10202 , n10203 );
not ( n10205 , n10203 );
nor ( n10206 , n10205 , n10201 );
nor ( n10207 , n10204 , n10206 );
not ( n10208 , n10207 );
and ( n10209 , n10199 , n10208 );
and ( n10210 , n10198 , n10207 );
nor ( n10211 , n10209 , n10210 );
not ( n10212 , n10211 );
and ( n10213 , n10054 , n10058 );
nor ( n10214 , n10213 , n10057 );
not ( n10215 , n10214 );
and ( n10216 , n10212 , n10215 );
and ( n10217 , n10211 , n10214 );
nor ( n10218 , n10216 , n10217 );
not ( n10219 , n10063 );
not ( n10220 , n9966 );
or ( n10221 , n10219 , n10220 );
not ( n10222 , n9975 );
not ( n10223 , n10064 );
and ( n10224 , n10222 , n10223 );
nor ( n10225 , n10224 , n10060 );
nand ( n10226 , n10221 , n10225 );
xnor ( n10227 , n10218 , n10226 );
and ( n10228 , n10227 , n6416 );
nor ( n10229 , n10169 , n1 );
nor ( n10230 , n10228 , n10229 );
nand ( n10231 , n10195 , n10230 );
nand ( n10232 , n10231 , n10140 );
nand ( n10233 , n10170 , n10232 );
buf ( n10234 , n10233 );
not ( n10235 , n10234 );
not ( n10236 , n10235 );
or ( n10237 , n10137 , n10236 );
or ( n10238 , n10235 , n10136 );
nand ( n10239 , n10237 , n10238 );
nand ( n10240 , n10131 , n10239 );
and ( n10241 , n10144 , n10168 );
and ( n10242 , n10159 , n10167 );
nor ( n10243 , n10241 , n10242 , n1 );
and ( n10244 , n10148 , n10158 );
and ( n10245 , n10088 , n10154 );
nor ( n10246 , n10244 , n10245 );
and ( n10247 , n6445 , n10163 );
and ( n10248 , n6452 , n86 );
nor ( n10249 , n10247 , n10248 );
not ( n10250 , n10249 );
or ( n10251 , n7049 , n10152 );
or ( n10252 , n69 , n84 );
nand ( n10253 , n69 , n84 );
nand ( n10254 , n10252 , n10253 );
or ( n10255 , n7171 , n10254 );
nand ( n10256 , n10251 , n10255 );
not ( n10257 , n10256 );
not ( n10258 , n10093 );
and ( n10259 , n10257 , n10258 );
and ( n10260 , n10256 , n10093 );
nor ( n10261 , n10259 , n10260 );
not ( n10262 , n10261 );
or ( n10263 , n10250 , n10262 );
or ( n10264 , n10261 , n10249 );
nand ( n10265 , n10263 , n10264 );
and ( n10266 , n10165 , n10166 );
and ( n10267 , n6946 , n9859 );
nor ( n10268 , n10266 , n10267 );
xnor ( n10269 , n10265 , n10268 );
xnor ( n10270 , n10246 , n10269 );
nor ( n10271 , n10270 , n1 );
nand ( n10272 , n10243 , n10271 );
not ( n10273 , n10272 );
not ( n10274 , n10185 );
not ( n10275 , n10180 );
and ( n10276 , n10274 , n10275 );
and ( n10277 , n10185 , n10178 );
nor ( n10278 , n10276 , n10277 );
not ( n10279 , n10278 );
and ( n10280 , n10198 , n10206 );
not ( n10281 , n10198 );
and ( n10282 , n10281 , n10204 );
nor ( n10283 , n10280 , n10282 );
nor ( n10284 , n374 , n2674 );
and ( n10285 , n10284 , n52 );
and ( n10286 , n2774 , n4666 );
nor ( n10287 , n10285 , n10286 );
xor ( n10288 , n10283 , n10287 );
not ( n10289 , n10218 );
not ( n10290 , n10289 );
not ( n10291 , n10226 );
or ( n10292 , n10290 , n10291 );
not ( n10293 , n10214 );
nand ( n10294 , n10293 , n10211 );
nand ( n10295 , n10292 , n10294 );
xnor ( n10296 , n10288 , n10295 );
nand ( n10297 , n10296 , n4562 );
not ( n10298 , n10193 );
not ( n10299 , n10173 );
or ( n10300 , n10298 , n10299 );
not ( n10301 , n10192 );
nand ( n10302 , n10301 , n10189 );
nand ( n10303 , n10300 , n10302 );
and ( n10304 , n335 , n10284 );
not ( n10305 , n335 );
and ( n10306 , n10305 , n2774 );
nor ( n10307 , n10304 , n10306 );
and ( n10308 , n10303 , n10307 );
not ( n10309 , n10303 );
not ( n10310 , n10307 );
and ( n10311 , n10309 , n10310 );
nor ( n10312 , n10308 , n10311 );
nand ( n10313 , n10279 , n10297 , n10312 , n1 );
nand ( n10314 , n10278 , n1 );
nor ( n10315 , n10312 , n10314 );
nand ( n10316 , n10315 , n10297 );
nand ( n10317 , n10297 , n6416 );
nor ( n10318 , n10243 , n10271 );
nand ( n10319 , n10313 , n10316 , n10317 , n10318 );
not ( n10320 , n10319 );
or ( n10321 , n10273 , n10320 );
nand ( n10322 , n10135 , n10233 );
or ( n10323 , n10140 , n10169 );
nand ( n10324 , n10322 , n10323 );
nand ( n10325 , n10321 , n10324 );
and ( n10326 , n10323 , n10272 );
nand ( n10327 , n10319 , n10326 , n10322 );
and ( n10328 , n10325 , n10327 );
nor ( n10329 , n10240 , n10328 );
not ( n10330 , n10326 );
not ( n10331 , n10322 );
or ( n10332 , n10330 , n10331 );
nand ( n10333 , n10332 , n10319 );
not ( n10334 , n10268 );
not ( n10335 , n10265 );
or ( n10336 , n10334 , n10335 );
or ( n10337 , n10246 , n10269 );
nand ( n10338 , n10336 , n10337 );
not ( n10339 , n7049 );
not ( n10340 , n10254 );
and ( n10341 , n10339 , n10340 );
and ( n10342 , n6668 , n68 );
and ( n10343 , n6741 , n84 );
nor ( n10344 , n10342 , n10343 );
not ( n10345 , n10344 );
and ( n10346 , n7170 , n10345 );
nor ( n10347 , n10341 , n10346 );
xnor ( n10348 , n10347 , n10151 );
xor ( n10349 , n10348 , n6512 );
not ( n10350 , n10256 );
and ( n10351 , n10249 , n10350 , n10093 );
nor ( n10352 , n10249 , n10350 , n10093 );
nor ( n10353 , n10351 , n10352 );
xor ( n10354 , n10349 , n10353 );
or ( n10355 , n10338 , n10354 );
nand ( n10356 , n10338 , n10354 , n2526 );
and ( n10357 , n10355 , n10356 , n2526 );
xnor ( n10358 , n10333 , n10357 );
and ( n10359 , n10329 , n10358 );
or ( n10360 , n10348 , n6512 );
or ( n10361 , n10347 , n10151 );
nand ( n10362 , n10360 , n10361 );
or ( n10363 , n7049 , n10344 );
or ( n10364 , n7171 , n6668 );
nand ( n10365 , n10363 , n10364 );
and ( n10366 , n10365 , n10253 );
not ( n10367 , n10365 );
not ( n10368 , n10253 );
and ( n10369 , n10367 , n10368 );
nor ( n10370 , n10366 , n10369 );
xnor ( n10371 , n10362 , n10370 );
and ( n10372 , n10353 , n10349 );
nor ( n10373 , n10372 , n10352 );
and ( n10374 , n10371 , n10373 );
nor ( n10375 , n10374 , n1 );
not ( n10376 , n10373 );
not ( n10377 , n10371 );
nand ( n10378 , n10376 , n10377 , n2526 );
nand ( n10379 , n10375 , n10378 );
not ( n10380 , n10379 );
not ( n10381 , n10357 );
not ( n10382 , n10333 );
not ( n10383 , n10382 );
or ( n10384 , n10381 , n10383 );
nand ( n10385 , n10384 , n10356 );
not ( n10386 , n10385 );
or ( n10387 , n10380 , n10386 );
or ( n10388 , n10379 , n10385 );
nand ( n10389 , n10387 , n10388 );
and ( n10390 , n10359 , n10389 );
and ( n10391 , n10362 , n10370 );
and ( n10392 , n10365 , n10253 );
nor ( n10393 , n10391 , n10392 );
or ( n10394 , n6668 , n10368 , n6741 );
or ( n10395 , n10253 , n68 );
nand ( n10396 , n10394 , n10395 );
not ( n10397 , n6697 );
or ( n10398 , n10396 , n10397 );
nand ( n10399 , n10396 , n10397 );
nand ( n10400 , n10398 , n10399 );
nor ( n10401 , n10393 , n10400 );
not ( n10402 , n10401 );
and ( n10403 , n10393 , n10400 );
nor ( n10404 , n10403 , n1 );
nand ( n10405 , n10402 , n10404 );
not ( n10406 , n10405 );
not ( n10407 , n10356 );
not ( n10408 , n10333 );
or ( n10409 , n10407 , n10408 );
and ( n10410 , n10355 , n10375 );
nand ( n10411 , n10409 , n10410 );
nand ( n10412 , n10411 , n10378 );
not ( n10413 , n10412 );
or ( n10414 , n10406 , n10413 );
or ( n10415 , n10405 , n10412 );
nand ( n10416 , n10414 , n10415 );
and ( n10417 , n10416 , n2531 );
or ( n10418 , n10401 , n10412 );
nand ( n10419 , n10418 , n10404 );
and ( n10420 , n10368 , n68 );
not ( n10421 , n10399 );
nor ( n10422 , n10420 , n10421 , n1 );
nand ( n10423 , n10419 , n10422 );
not ( n10424 , n10423 );
nand ( n10425 , n10390 , n10417 , n10424 );
nand ( n10426 , n2532 , n10425 );
xnor ( n10427 , n10379 , n10385 );
and ( n10428 , n10329 , n10358 );
or ( n10429 , n10427 , n10428 );
nand ( n10430 , n10429 , n2530 );
or ( n10431 , n10430 , n10390 );
xnor ( n10432 , n2486 , n615 );
or ( n10433 , n10432 , n2531 );
nand ( n10434 , n10431 , n10433 );
nand ( n10435 , n10416 , n10389 , n10359 );
nand ( n10436 , n10435 , n2531 );
buf ( n10437 , n10329 );
or ( n10438 , n10437 , n10358 );
nand ( n10439 , n10438 , n2530 );
or ( n10440 , n10439 , n10428 );
xnor ( n10441 , n2481 , n708 );
or ( n10442 , n10441 , n2530 );
nand ( n10443 , n10440 , n10442 );
buf ( n10444 , n10131 );
buf ( n10445 , n10239 );
and ( n10446 , n10444 , n10445 );
not ( n10447 , n10328 );
or ( n10448 , n10446 , n10447 );
nand ( n10449 , n10448 , n2530 );
or ( n10450 , n10449 , n10437 );
xnor ( n10451 , n2476 , n818 );
or ( n10452 , n10451 , n2530 );
nand ( n10453 , n10450 , n10452 );
not ( n10454 , n10444 );
not ( n10455 , n10445 );
and ( n10456 , n10454 , n10455 );
not ( n10457 , n2530 );
nor ( n10458 , n10456 , n10457 );
nand ( n10459 , n10240 , n10458 );
xor ( n10460 , n2471 , n1030 );
nand ( n10461 , n10460 , n10457 );
nand ( n10462 , n10459 , n10461 );
not ( n10463 , n10457 );
xor ( n10464 , n1128 , n2466 );
not ( n10465 , n10464 );
or ( n10466 , n10463 , n10465 );
buf ( n10467 , n9996 );
and ( n10468 , n10467 , n10130 );
not ( n10469 , n2530 );
nor ( n10470 , n10468 , n10469 );
nand ( n10471 , n10454 , n10470 );
nand ( n10472 , n10466 , n10471 );
not ( n10473 , n10469 );
xor ( n10474 , n2461 , n1261 );
not ( n10475 , n10474 );
or ( n10476 , n10473 , n10475 );
not ( n10477 , n9989 );
not ( n10478 , n9685 );
not ( n10479 , n10478 );
nand ( n10480 , n10479 , n9995 );
nand ( n10481 , n10477 , n10480 );
nand ( n10482 , n10481 , n2530 , n10467 );
nand ( n10483 , n10476 , n10482 );
xnor ( n10484 , n1357 , n2456 );
and ( n10485 , n10469 , n10484 );
not ( n10486 , n10469 );
and ( n10487 , n10478 , n9995 );
not ( n10488 , n10478 );
not ( n10489 , n9995 );
and ( n10490 , n10488 , n10489 );
nor ( n10491 , n10487 , n10490 );
and ( n10492 , n10486 , n10491 );
nor ( n10493 , n10485 , n10492 );
xnor ( n10494 , n2451 , n1482 );
and ( n10495 , n10469 , n10494 );
not ( n10496 , n10469 );
buf ( n10497 , n9487 );
not ( n10498 , n10497 );
not ( n10499 , n9684 );
not ( n10500 , n10499 );
and ( n10501 , n10498 , n10500 );
and ( n10502 , n10497 , n10499 );
nor ( n10503 , n10501 , n10502 );
and ( n10504 , n10496 , n10503 );
nor ( n10505 , n10495 , n10504 );
not ( n10506 , n2519 );
not ( n10507 , n10506 );
not ( n10508 , n2501 );
or ( n10509 , n10507 , n10508 );
not ( n10510 , n2515 );
nand ( n10511 , n10510 , n2505 );
nand ( n10512 , n10509 , n10511 );
not ( n10513 , n10512 );
or ( n10514 , n323 , n2676 );
and ( n10515 , n323 , n2676 );
nor ( n10516 , n10515 , n303 );
nand ( n10517 , n10514 , n10516 );
not ( n10518 , n10517 );
or ( n10519 , n2509 , n2514 );
or ( n10520 , n2513 , n338 );
nand ( n10521 , n10519 , n10520 );
not ( n10522 , n10521 );
or ( n10523 , n10518 , n10522 );
or ( n10524 , n10521 , n10517 );
nand ( n10525 , n10523 , n10524 );
not ( n10526 , n10525 );
and ( n10527 , n10513 , n10526 );
and ( n10528 , n10512 , n10525 );
nor ( n10529 , n10527 , n10528 );
nor ( n10530 , n10529 , n2530 );
not ( n10531 , n10130 );
xnor ( n10532 , n2446 , n1617 );
or ( n10533 , n10532 , n2530 );
not ( n10534 , n8941 );
nand ( n10535 , n10534 , n9045 , n9269 );
not ( n10536 , n8903 );
nor ( n10537 , n10535 , n10536 );
and ( n10538 , n10537 , n9267 );
not ( n10539 , n9486 );
or ( n10540 , n10538 , n10539 );
not ( n10541 , n10497 );
nand ( n10542 , n10540 , n10541 , n2530 );
nand ( n10543 , n10533 , n10542 );
not ( n10544 , n490 );
buf ( n10545 , n2496 );
not ( n10546 , n10545 );
or ( n10547 , n10544 , n10546 );
or ( n10548 , n10545 , n490 );
nand ( n10549 , n10547 , n10548 );
not ( n10550 , n2531 );
nand ( n10551 , n10549 , n10550 );
or ( n10552 , n10537 , n9267 );
nand ( n10553 , n10552 , n2530 );
or ( n10554 , n10553 , n10538 );
xnor ( n10555 , n2441 , n1721 );
or ( n10556 , n10555 , n2530 );
nand ( n10557 , n10554 , n10556 );
not ( n10558 , n10535 );
or ( n10559 , n10558 , n8903 );
nand ( n10560 , n10559 , n2530 );
or ( n10561 , n10560 , n10537 );
xnor ( n10562 , n2436 , n1813 );
or ( n10563 , n10562 , n2530 );
nand ( n10564 , n10561 , n10563 );
xnor ( n10565 , n2431 , n1870 );
or ( n10566 , n10565 , n2530 );
buf ( n10567 , n8933 );
not ( n10568 , n8919 );
and ( n10569 , n9043 , n10568 );
nand ( n10570 , n10567 , n10569 );
nand ( n10571 , n9269 , n8940 );
nor ( n10572 , n10570 , n10571 );
not ( n10573 , n8905 );
nor ( n10574 , n9268 , n10573 );
and ( n10575 , n10574 , n8907 );
not ( n10576 , n10574 );
not ( n10577 , n8907 );
and ( n10578 , n10576 , n10577 );
nor ( n10579 , n10575 , n10578 );
or ( n10580 , n10572 , n10579 );
nand ( n10581 , n10580 , n10535 , n2530 );
nand ( n10582 , n10566 , n10581 );
not ( n10583 , n10570 );
not ( n10584 , n10571 );
or ( n10585 , n10583 , n10584 );
nand ( n10586 , n10585 , n2530 );
or ( n10587 , n10586 , n10572 );
xnor ( n10588 , n2426 , n1950 );
or ( n10589 , n10588 , n2530 );
nand ( n10590 , n10587 , n10589 );
not ( n10591 , n10469 );
xor ( n10592 , n2411 , n2423 );
not ( n10593 , n10592 );
or ( n10594 , n10591 , n10593 );
not ( n10595 , n10569 );
not ( n10596 , n10567 );
and ( n10597 , n10595 , n10596 );
nor ( n10598 , n10597 , n10469 );
nand ( n10599 , n10598 , n10570 );
nand ( n10600 , n10594 , n10599 );
not ( n10601 , n10469 );
xor ( n10602 , n2406 , n2394 );
not ( n10603 , n10602 );
not ( n10604 , n2390 );
or ( n10605 , n10603 , n10604 );
or ( n10606 , n2390 , n10602 );
nand ( n10607 , n10605 , n10606 );
not ( n10608 , n10607 );
or ( n10609 , n10601 , n10608 );
and ( n10610 , n9044 , n8919 );
nor ( n10611 , n10610 , n10469 );
nand ( n10612 , n10611 , n10595 );
nand ( n10613 , n10609 , n10612 );
not ( n10614 , n10469 );
xor ( n10615 , n2108 , n2385 );
not ( n10616 , n10615 );
or ( n10617 , n10614 , n10616 );
buf ( n10618 , n9036 );
not ( n10619 , n9042 );
not ( n10620 , n10619 );
and ( n10621 , n10618 , n10620 );
not ( n10622 , n2530 );
nor ( n10623 , n10621 , n10622 );
nand ( n10624 , n10623 , n9044 );
nand ( n10625 , n10617 , n10624 );
not ( n10626 , n10469 );
xor ( n10627 , n2380 , n2156 );
not ( n10628 , n10627 );
or ( n10629 , n10626 , n10628 );
buf ( n10630 , n9009 );
buf ( n10631 , n9034 );
nand ( n10632 , n10630 , n10631 , n9035 );
not ( n10633 , n9024 );
and ( n10634 , n10632 , n10633 );
not ( n10635 , n2530 );
nor ( n10636 , n10634 , n10635 );
nand ( n10637 , n10618 , n10636 );
nand ( n10638 , n10629 , n10637 );
xor ( n10639 , n2198 , n2376 );
nand ( n10640 , n10639 , n10469 );
nand ( n10641 , n10630 , n10631 );
not ( n10642 , n9035 );
and ( n10643 , n10641 , n10642 );
nor ( n10644 , n10643 , n10622 );
nand ( n10645 , n10644 , n10632 );
nand ( n10646 , n10640 , n10645 );
not ( n10647 , n10469 );
xor ( n10648 , n2372 , n2232 );
not ( n10649 , n10648 );
or ( n10650 , n10647 , n10649 );
not ( n10651 , n10630 );
not ( n10652 , n10631 );
and ( n10653 , n10651 , n10652 );
nor ( n10654 , n10653 , n10635 );
nand ( n10655 , n10654 , n10641 );
nand ( n10656 , n10650 , n10655 );
buf ( n10657 , n8989 );
and ( n10658 , n10657 , n8998 );
or ( n10659 , n10658 , n9007 );
nand ( n10660 , n10659 , n2530 );
or ( n10661 , n10660 , n10630 );
not ( n10662 , n2356 );
not ( n10663 , n2367 );
and ( n10664 , n10662 , n10663 );
and ( n10665 , n2356 , n2367 );
nor ( n10666 , n10664 , n10665 );
or ( n10667 , n10666 , n2530 );
nand ( n10668 , n10661 , n10667 );
or ( n10669 , n10657 , n8998 );
nand ( n10670 , n10669 , n2530 );
or ( n10671 , n10670 , n10658 );
xnor ( n10672 , n2352 , n2288 );
or ( n10673 , n10672 , n2530 );
nand ( n10674 , n10671 , n10673 );
or ( n10675 , n8986 , n8988 );
nand ( n10676 , n10675 , n2530 );
or ( n10677 , n10657 , n10676 );
xnor ( n10678 , n2311 , n2348 );
or ( n10679 , n10678 , n2530 );
nand ( n10680 , n10677 , n10679 );
xnor ( n10681 , n8981 , n8954 );
or ( n10682 , n10681 , n10469 );
xnor ( n10683 , n2343 , n2330 );
or ( n10684 , n10683 , n2530 );
nand ( n10685 , n10682 , n10684 );
and ( n10686 , n2329 , n2320 );
or ( n10687 , n2330 , n10686 , n2530 );
or ( n10688 , n8962 , n8978 );
nand ( n10689 , n10688 , n8979 );
not ( n10690 , n10689 );
not ( n10691 , n2530 );
or ( n10692 , n10690 , n10691 );
nand ( n10693 , n10687 , n10692 );
and ( n10694 , n3581 , n1379 );
and ( n10695 , n1179 , n1788 );
nor ( n10696 , n10694 , n10695 , n1382 );
or ( n10697 , n10696 , n2319 , n2529 );
xnor ( n10698 , n8973 , n8976 );
or ( n10699 , n10698 , n10691 );
nand ( n10700 , n10697 , n10699 );
not ( n10701 , n8958 );
or ( n10702 , n2529 , n1524 , n1788 );
or ( n10703 , n19 , n8965 );
nand ( n10704 , n10703 , n8966 , n2529 );
nand ( n10705 , n10702 , n10704 );
xor ( n10706 , n7757 , n7792 );
xor ( n10707 , n10706 , n7853 );
xor ( n10708 , n7797 , n7814 );
xor ( n10709 , n10708 , n7850 );
xor ( n10710 , n7829 , n7832 );
xor ( n10711 , n10710 , n7847 );
and ( n10712 , n7826 , n7828 );
nor ( n10713 , n10712 , n7829 );
xnor ( n10714 , n2491 , n546 );
and ( n10715 , n10359 , n10389 );
nor ( n10716 , n10715 , n10416 );
or ( n10717 , n10436 , n10716 );
or ( n10718 , n10714 , n2531 );
nand ( n10719 , n10717 , n10718 );
xor ( n10720 , n7902 , n7856 );
not ( n10721 , n10435 );
nor ( n10722 , n10423 , n10550 );
not ( n10723 , n10722 );
or ( n10724 , n10721 , n10723 );
nand ( n10725 , n10724 , n10551 );
endmodule

