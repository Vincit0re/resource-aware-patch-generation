module top ( g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 );
input g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 ;
output g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 ;

wire n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , 
     n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , 
     n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , 
     n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , 
     n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , 
     n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , 
     n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , 
     n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , 
     n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , 
     n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , 
     n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , 
     n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , 
     n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , 
     n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , 
     n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , 
     n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , 
     n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , 
     n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , 
     n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , 
     n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , 
     n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , 
     n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , 
     n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , 
     n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , 
     n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , 
     n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , 
     n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , 
     n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , 
     n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , 
     n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , 
     n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , 
     n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , 
     n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , 
     n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , 
     n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , 
     n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , 
     n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , 
     n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , 
     n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , 
     n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , 
     n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , 
     n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , 
     n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , 
     n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , 
     n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , 
     n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , 
     n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , 
     n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , 
     n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , 
     n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , 
     n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , 
     n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , 
     n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , 
     n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , 
     n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , 
     n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , 
     n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , 
     n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , 
     n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , 
     n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , 
     n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , 
     n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , 
     n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , 
     n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , 
     n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , 
     n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , 
     n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , 
     n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , 
     n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , 
     n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , 
     n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , 
     n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , 
     n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , 
     n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , 
     n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , 
     n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , 
     n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , 
     n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , 
     n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , 
     n790 , n791 , n792 , n793 , n794 , n795 , n796 ;
buf ( n1 , g0 );
buf ( n2 , g1 );
buf ( n3 , g2 );
buf ( n4 , g3 );
buf ( n5 , g4 );
buf ( n6 , g5 );
buf ( n7 , g6 );
buf ( n8 , g7 );
buf ( n9 , g8 );
buf ( n10 , g9 );
buf ( n11 , g10 );
buf ( n12 , g11 );
buf ( n13 , g12 );
buf ( n14 , g13 );
buf ( n15 , g14 );
buf ( n16 , g15 );
buf ( n17 , g16 );
buf ( n18 , g17 );
buf ( n19 , g18 );
buf ( n20 , g19 );
buf ( n21 , g20 );
buf ( n22 , g21 );
buf ( n23 , g22 );
buf ( n24 , g23 );
buf ( n25 , g24 );
buf ( n26 , g25 );
buf ( n27 , g26 );
buf ( n28 , g27 );
buf ( n29 , g28 );
buf ( n30 , g29 );
buf ( n31 , g30 );
buf ( n32 , g31 );
buf ( n33 , g32 );
buf ( n34 , g33 );
buf ( n35 , g34 );
buf ( n36 , g35 );
buf ( n37 , g36 );
buf ( n38 , g37 );
buf ( n39 , g38 );
buf ( n40 , g39 );
buf ( n41 , g40 );
buf ( n42 , g41 );
buf ( n43 , g42 );
buf ( n44 , g43 );
buf ( n45 , g44 );
buf ( n46 , g45 );
buf ( g46 , n47 );
buf ( g47 , n48 );
buf ( g48 , n49 );
buf ( g49 , n50 );
buf ( g50 , n51 );
buf ( g51 , n52 );
buf ( g52 , n53 );
buf ( g53 , n54 );
buf ( g54 , n55 );
buf ( g55 , n56 );
buf ( g56 , n57 );
buf ( g57 , n58 );
buf ( g58 , n59 );
buf ( g59 , n60 );
buf ( g60 , n61 );
buf ( g61 , n62 );
buf ( g62 , n63 );
buf ( g63 , n64 );
buf ( g64 , n65 );
buf ( g65 , n66 );
buf ( g66 , n67 );
buf ( g67 , n68 );
buf ( g68 , n69 );
buf ( g69 , n70 );
buf ( g70 , n71 );
buf ( g71 , n72 );
buf ( g72 , n73 );
buf ( n47 , n383 );
buf ( n48 , n237 );
buf ( n49 , n606 );
buf ( n50 , n505 );
buf ( n51 , n569 );
buf ( n52 , n793 );
buf ( n53 , n624 );
buf ( n54 , n521 );
buf ( n55 , n316 );
buf ( n56 , n325 );
buf ( n57 , n693 );
buf ( n58 , n631 );
buf ( n59 , n796 );
buf ( n60 , n729 );
buf ( n61 , n636 );
buf ( n62 , n640 );
buf ( n63 , n686 );
buf ( n64 , n659 );
buf ( n65 , n744 );
buf ( n66 , n709 );
buf ( n67 , n784 );
buf ( n68 , n792 );
buf ( n69 , n766 );
buf ( n70 , n531 );
buf ( n71 , n755 );
buf ( n72 , n725 );
buf ( n73 , n776 );
nor ( n76 , n6 , n7 );
not ( n77 , n31 );
nand ( n78 , n76 , n77 );
not ( n79 , n78 );
not ( n80 , n79 );
not ( n81 , n2 );
not ( n82 , n81 );
not ( n83 , n41 );
nor ( n84 , n83 , n40 );
not ( n85 , n84 );
or ( n86 , n82 , n85 );
or ( n87 , n84 , n11 );
nand ( n88 , n86 , n87 );
and ( n89 , n88 , n24 );
not ( n90 , n38 );
nor ( n91 , n90 , n39 );
and ( n92 , n91 , n4 );
not ( n93 , n91 );
and ( n94 , n93 , n5 );
or ( n95 , n92 , n94 );
nor ( n96 , n95 , n24 );
or ( n97 , n8 , n9 , n10 );
not ( n98 , n97 );
nor ( n99 , n89 , n96 , n98 );
not ( n100 , n5 );
nor ( n101 , n100 , n24 );
not ( n102 , n38 );
nor ( n103 , n102 , n39 );
nand ( n104 , n101 , n103 );
not ( n105 , n24 );
not ( n106 , n39 );
nand ( n107 , n106 , n38 );
nand ( n108 , n105 , n107 , n4 );
not ( n109 , n40 );
not ( n110 , n11 );
nand ( n111 , n109 , n110 , n41 );
not ( n112 , n24 );
nor ( n113 , n2 , n41 );
nor ( n114 , n112 , n113 );
not ( n115 , n2 );
nand ( n116 , n115 , n40 );
nand ( n117 , n111 , n114 , n116 );
nand ( n118 , n104 , n108 , n117 );
not ( n119 , n38 );
not ( n120 , n39 );
nand ( n121 , n119 , n120 );
not ( n122 , n121 );
and ( n123 , n122 , n1 );
not ( n124 , n1 );
nand ( n125 , n124 , n38 );
not ( n126 , n24 );
nand ( n127 , n125 , n126 );
nor ( n128 , n123 , n127 );
not ( n129 , n1 );
and ( n130 , n129 , n39 );
nor ( n131 , n130 , n3 );
and ( n132 , n128 , n131 );
not ( n133 , n13 );
nand ( n134 , n133 , n40 );
not ( n135 , n24 );
nor ( n136 , n135 , n12 );
not ( n137 , n13 );
nand ( n138 , n137 , n41 );
nand ( n139 , n134 , n136 , n138 );
not ( n140 , n13 );
nor ( n141 , n140 , n40 , n41 );
nor ( n142 , n139 , n141 );
nor ( n143 , n132 , n142 );
nor ( n144 , n118 , n143 );
and ( n145 , n99 , n144 );
not ( n146 , n145 );
or ( n147 , n80 , n146 );
nand ( n148 , n147 , n23 );
not ( n149 , n126 );
not ( n150 , n12 );
nand ( n151 , n150 , n13 );
not ( n152 , n151 );
nor ( n153 , n2 , n11 );
nand ( n154 , n152 , n153 );
not ( n155 , n154 );
not ( n156 , n155 );
or ( n157 , n149 , n156 );
not ( n158 , n4 );
nor ( n159 , n3 , n5 );
nand ( n160 , n158 , n159 );
not ( n161 , n160 );
nand ( n162 , n161 , n24 , n1 );
nand ( n163 , n157 , n162 );
not ( n164 , n160 );
and ( n165 , n164 , n24 , n42 );
or ( n166 , n163 , n165 );
not ( n167 , n33 );
nand ( n168 , n167 , n16 );
nand ( n169 , n19 , n33 );
nand ( n170 , n168 , n169 );
not ( n171 , n170 );
not ( n172 , n171 );
xor ( n173 , n14 , n36 );
not ( n174 , n173 );
not ( n175 , n174 );
or ( n176 , n172 , n175 );
nor ( n177 , n30 , n34 );
nand ( n178 , n176 , n177 );
xor ( n179 , n14 , n37 );
not ( n180 , n179 );
and ( n181 , n35 , n19 );
not ( n182 , n35 );
and ( n183 , n182 , n16 );
nor ( n184 , n181 , n183 );
not ( n185 , n32 );
nand ( n186 , n180 , n184 , n185 );
not ( n187 , n18 );
and ( n188 , n187 , n32 );
nor ( n189 , n188 , n25 );
nand ( n190 , n186 , n189 );
nand ( n191 , n20 , n34 );
or ( n192 , n191 , n30 );
nand ( n193 , n178 , n190 , n192 );
nand ( n194 , n166 , n193 );
not ( n195 , n194 );
not ( n196 , n25 );
nand ( n197 , n196 , n26 );
not ( n198 , n197 );
not ( n199 , n30 );
nand ( n200 , n199 , n29 );
buf ( n201 , n200 );
not ( n202 , n201 );
nor ( n203 , n198 , n202 );
not ( n204 , n203 );
or ( n205 , n195 , n204 );
nor ( n206 , n27 , n28 );
not ( n207 , n23 );
and ( n208 , n206 , n207 , n15 , n17 );
not ( n209 , n22 );
and ( n210 , n76 , n209 , n77 );
nand ( n211 , n208 , n210 );
not ( n212 , n211 );
nand ( n213 , n205 , n212 );
not ( n214 , n27 );
nand ( n215 , n214 , n15 );
not ( n216 , n28 );
nand ( n217 , n216 , n17 );
nor ( n218 , n215 , n217 );
not ( n219 , n218 );
nor ( n220 , n219 , n24 );
not ( n221 , n220 );
nand ( n222 , n164 , n1 );
nor ( n223 , n222 , n21 );
not ( n224 , n160 );
and ( n225 , n224 , n129 , n42 );
nor ( n226 , n223 , n225 );
not ( n227 , n226 );
not ( n228 , n227 );
or ( n229 , n221 , n228 );
not ( n230 , n21 );
nand ( n231 , n155 , n230 );
nand ( n232 , n24 , n218 );
or ( n233 , n231 , n232 );
nand ( n234 , n229 , n233 );
and ( n235 , n193 , n79 , n209 );
nand ( n236 , n234 , n235 );
nand ( n237 , n148 , n213 , n236 );
not ( n238 , n77 );
nand ( n239 , n12 , n13 );
buf ( n240 , n239 );
nand ( n241 , n24 , n240 , n153 );
nor ( n242 , n4 , n5 );
nand ( n243 , n1 , n3 );
nand ( n244 , n242 , n126 , n243 );
nor ( n245 , n207 , n7 );
nand ( n246 , n241 , n244 , n245 );
not ( n247 , n246 );
or ( n248 , n238 , n247 );
not ( n249 , n7 );
and ( n250 , n249 , n31 );
nor ( n251 , n250 , n6 );
nand ( n252 , n248 , n251 );
not ( n253 , n252 );
not ( n254 , n144 );
nor ( n255 , n8 , n31 );
nand ( n256 , n254 , n255 );
and ( n257 , n22 , n34 );
not ( n258 , n22 );
and ( n259 , n258 , n32 );
nor ( n260 , n257 , n259 );
or ( n261 , n260 , n77 );
nand ( n262 , n261 , n23 );
not ( n263 , n8 );
and ( n264 , n262 , n263 );
nand ( n265 , n263 , n31 , n9 );
not ( n266 , n265 );
nor ( n267 , n264 , n266 );
nand ( n268 , n253 , n256 , n267 );
nand ( n269 , n268 , n10 );
not ( n270 , n118 );
not ( n271 , n1 );
not ( n272 , n120 );
or ( n273 , n271 , n272 );
nand ( n274 , n273 , n131 );
and ( n275 , n274 , n101 );
not ( n276 , n40 );
nand ( n277 , n276 , n13 );
not ( n278 , n12 );
and ( n279 , n134 , n277 , n278 );
nand ( n280 , n11 , n24 );
nor ( n281 , n279 , n280 );
nor ( n282 , n275 , n281 );
nor ( n283 , n243 , n24 );
not ( n284 , n283 );
not ( n285 , n239 );
nand ( n286 , n285 , n24 );
nand ( n287 , n284 , n286 );
not ( n288 , n13 );
nand ( n289 , n288 , n2 );
and ( n290 , n24 , n289 );
not ( n291 , n24 );
not ( n292 , n1 );
nand ( n293 , n292 , n4 );
and ( n294 , n291 , n293 );
nor ( n295 , n290 , n294 );
nor ( n296 , n287 , n295 );
nand ( n297 , n270 , n282 , n296 );
nand ( n298 , n79 , n23 );
not ( n299 , n298 );
nand ( n300 , n297 , n299 );
not ( n301 , n300 );
not ( n302 , n10 );
and ( n303 , n302 , n8 );
and ( n304 , n301 , n303 );
not ( n305 , n303 );
not ( n306 , n6 );
nand ( n307 , n306 , n31 , n7 );
nor ( n308 , n305 , n307 );
not ( n309 , n308 );
nand ( n310 , n9 , n23 );
or ( n311 , n260 , n310 );
or ( n312 , n9 , n23 );
nand ( n313 , n311 , n312 );
nor ( n314 , n309 , n313 );
nor ( n315 , n304 , n314 );
nand ( n316 , n269 , n315 );
not ( n317 , n10 );
nor ( n318 , n317 , n9 );
and ( n319 , n318 , n260 , n23 );
nor ( n320 , n319 , n307 );
nor ( n321 , n301 , n320 );
or ( n322 , n321 , n8 );
not ( n323 , n252 );
or ( n324 , n323 , n263 );
nand ( n325 , n322 , n324 );
nor ( n326 , n18 , n26 );
not ( n327 , n326 );
not ( n328 , n32 );
or ( n329 , n327 , n328 );
not ( n330 , n25 );
nand ( n331 , n329 , n330 );
not ( n332 , n331 );
not ( n333 , n34 );
not ( n334 , n333 );
not ( n335 , n170 );
or ( n336 , n334 , n335 );
nand ( n337 , n336 , n191 );
nor ( n338 , n174 , n34 );
nor ( n339 , n337 , n338 );
not ( n340 , n339 );
not ( n341 , n340 );
or ( n342 , n332 , n341 );
not ( n343 , n35 );
nor ( n344 , n343 , n19 );
not ( n345 , n344 );
not ( n346 , n168 );
not ( n347 , n346 );
or ( n348 , n345 , n347 );
not ( n349 , n169 );
not ( n350 , n16 );
not ( n351 , n35 );
nand ( n352 , n349 , n350 , n351 );
nand ( n353 , n348 , n352 );
and ( n354 , n353 , n180 , n333 );
or ( n355 , n191 , n179 );
xor ( n356 , n36 , n37 );
or ( n357 , n14 , n36 );
nand ( n358 , n14 , n36 );
nand ( n359 , n356 , n357 , n333 , n358 );
nand ( n360 , n355 , n359 );
and ( n361 , n360 , n184 );
nor ( n362 , n354 , n361 );
not ( n363 , n362 );
nor ( n364 , n26 , n32 );
nand ( n365 , n363 , n364 );
nand ( n366 , n342 , n365 );
not ( n367 , n163 );
nand ( n368 , n367 , n226 , n231 );
not ( n369 , n217 );
nand ( n370 , n79 , n369 , n207 );
nor ( n371 , n370 , n30 );
nand ( n372 , n366 , n368 , n371 );
not ( n373 , n145 );
and ( n374 , n373 , n22 );
or ( n375 , n299 , n209 );
not ( n376 , n200 );
and ( n377 , n376 , n197 );
or ( n378 , n377 , n215 );
not ( n379 , n370 );
nand ( n380 , n378 , n379 );
nand ( n381 , n375 , n380 );
nor ( n382 , n374 , n381 );
nand ( n383 , n372 , n382 );
nor ( n384 , n25 , n26 );
not ( n385 , n184 );
not ( n386 , n32 );
and ( n387 , n385 , n386 );
and ( n388 , n18 , n32 );
nor ( n389 , n387 , n388 );
not ( n390 , n389 );
and ( n391 , n384 , n390 );
nand ( n392 , n185 , n37 );
nor ( n393 , n392 , n14 , n25 );
nor ( n394 , n391 , n393 );
nor ( n395 , n1 , n42 );
not ( n396 , n395 );
not ( n397 , n224 );
or ( n398 , n396 , n397 );
not ( n399 , n43 );
nand ( n400 , n398 , n399 );
not ( n401 , n400 );
nor ( n402 , n394 , n401 );
nor ( n403 , n211 , n154 );
buf ( n404 , n403 );
and ( n405 , n402 , n404 , n201 );
nor ( n406 , n22 , n23 );
nand ( n407 , n79 , n406 );
not ( n408 , n407 );
not ( n409 , n14 );
nor ( n410 , n409 , n28 );
nand ( n411 , n408 , n410 );
nor ( n412 , n411 , n27 );
nor ( n413 , n29 , n30 );
nor ( n414 , n34 , n36 );
nand ( n415 , n197 , n413 , n414 );
nor ( n416 , n32 , n37 );
nand ( n417 , n200 , n384 , n416 );
nand ( n418 , n415 , n417 );
nand ( n419 , n400 , n418 , n155 );
nand ( n420 , n15 , n419 );
and ( n421 , n412 , n420 );
nor ( n422 , n405 , n421 );
and ( n423 , n337 , n413 );
not ( n424 , n36 );
nor ( n425 , n424 , n14 );
and ( n426 , n425 , n177 );
nor ( n427 , n423 , n426 );
nand ( n428 , n197 , n400 );
nor ( n429 , n427 , n428 );
and ( n430 , n429 , n404 );
nor ( n431 , n424 , n34 );
not ( n432 , n431 );
not ( n433 , n33 );
not ( n434 , n344 );
or ( n435 , n433 , n434 );
not ( n436 , n16 );
or ( n437 , n35 , n33 );
nand ( n438 , n437 , n19 );
nand ( n439 , n436 , n438 );
nand ( n440 , n435 , n439 );
not ( n441 , n440 );
or ( n442 , n432 , n441 );
not ( n443 , n20 );
nand ( n444 , n443 , n34 );
or ( n445 , n444 , n29 );
nand ( n446 , n445 , n199 );
nand ( n447 , n446 , n184 );
nand ( n448 , n442 , n447 );
not ( n449 , n392 );
and ( n450 , n448 , n449 );
nand ( n451 , n326 , n32 );
nand ( n452 , n451 , n330 );
and ( n453 , n452 , n171 , n431 );
nor ( n454 , n450 , n453 );
not ( n455 , n27 );
nand ( n456 , n455 , n410 , n24 );
nor ( n457 , n454 , n456 );
nor ( n458 , n430 , n457 );
not ( n459 , n446 );
not ( n460 , n459 );
not ( n461 , n29 );
and ( n462 , n414 , n461 );
nand ( n463 , n171 , n462 , n409 );
not ( n464 , n463 );
or ( n465 , n460 , n464 );
nand ( n466 , n465 , n452 );
not ( n467 , n278 );
not ( n468 , n153 );
or ( n469 , n467 , n468 );
nand ( n470 , n469 , n43 );
not ( n471 , n470 );
nor ( n472 , n160 , n395 );
not ( n473 , n472 );
or ( n474 , n471 , n473 );
or ( n475 , n198 , n29 );
or ( n476 , n199 , n26 );
nand ( n477 , n475 , n476 );
nand ( n478 , n474 , n477 );
and ( n479 , n466 , n478 );
nor ( n480 , n479 , n232 );
nor ( n481 , n411 , n17 );
not ( n482 , n24 );
not ( n483 , n407 );
or ( n484 , n482 , n483 );
and ( n485 , n369 , n27 , n45 );
and ( n486 , n28 , n44 );
nor ( n487 , n485 , n486 );
or ( n488 , n407 , n487 );
nand ( n489 , n484 , n488 );
nor ( n490 , n480 , n481 , n489 );
not ( n491 , n37 );
nand ( n492 , n364 , n409 , n491 );
nor ( n493 , n232 , n492 );
not ( n494 , n440 );
not ( n495 , n462 );
or ( n496 , n494 , n495 );
nand ( n497 , n496 , n447 );
and ( n498 , n493 , n497 );
not ( n499 , n377 );
or ( n500 , n499 , n424 );
or ( n501 , n197 , n491 );
nand ( n502 , n500 , n501 );
and ( n503 , n502 , n212 );
nor ( n504 , n498 , n503 );
nand ( n505 , n422 , n458 , n490 , n504 );
or ( n506 , n10 , n31 );
nand ( n507 , n506 , n8 );
and ( n508 , n254 , n507 );
nor ( n509 , n508 , n252 );
not ( n510 , n9 );
or ( n511 , n509 , n510 );
nand ( n512 , n318 , n8 );
or ( n513 , n300 , n512 );
not ( n514 , n260 );
or ( n515 , n514 , n77 );
nand ( n516 , n515 , n23 );
and ( n517 , n516 , n302 , n9 );
or ( n518 , n512 , n307 );
nand ( n519 , n518 , n265 );
nor ( n520 , n517 , n519 );
nand ( n521 , n511 , n513 , n520 );
not ( n522 , n23 );
nor ( n523 , n522 , n22 );
not ( n524 , n523 );
not ( n525 , n413 );
nor ( n526 , n219 , n524 , n525 );
not ( n527 , n526 );
not ( n528 , n340 );
or ( n529 , n527 , n528 );
nor ( n530 , n6 , n7 );
buf ( n531 , n530 );
not ( n532 , n531 );
not ( n533 , n532 );
not ( n534 , n533 );
not ( n535 , n534 );
nand ( n536 , n529 , n535 );
and ( n537 , n536 , n21 );
not ( n538 , n185 );
not ( n539 , n179 );
or ( n540 , n538 , n539 );
nand ( n541 , n540 , n389 );
nand ( n542 , n22 , n23 );
not ( n543 , n542 );
nand ( n544 , n543 , n384 , n21 );
nor ( n545 , n219 , n544 );
and ( n546 , n541 , n545 );
nor ( n547 , n537 , n546 );
nor ( n548 , n198 , n525 );
not ( n549 , n548 );
not ( n550 , n340 );
or ( n551 , n549 , n550 );
not ( n552 , n384 );
nor ( n553 , n202 , n552 );
nand ( n554 , n541 , n553 );
nand ( n555 , n551 , n554 );
not ( n556 , n403 );
and ( n557 , n472 , n212 );
and ( n558 , n22 , n217 );
not ( n559 , n22 );
and ( n560 , n559 , n215 );
nor ( n561 , n558 , n560 );
nand ( n562 , n561 , n31 );
and ( n563 , n562 , n219 );
nand ( n564 , n207 , n21 );
nor ( n565 , n563 , n564 );
nor ( n566 , n557 , n565 );
nand ( n567 , n556 , n566 );
nand ( n568 , n555 , n567 );
nand ( n569 , n547 , n568 );
and ( n570 , n226 , n162 );
nand ( n571 , n212 , n399 );
nor ( n572 , n570 , n571 );
not ( n573 , n572 );
not ( n574 , n555 );
or ( n575 , n573 , n574 );
nand ( n576 , n171 , n174 );
or ( n577 , n576 , n189 );
nor ( n578 , n14 , n36 );
not ( n579 , n578 );
not ( n580 , n416 );
or ( n581 , n579 , n580 );
or ( n582 , n392 , n358 );
nand ( n583 , n581 , n582 );
and ( n584 , n440 , n583 );
nand ( n585 , n21 , n24 );
nand ( n586 , n197 , n585 );
nor ( n587 , n584 , n586 );
nand ( n588 , n577 , n587 );
not ( n589 , n586 );
nand ( n590 , n589 , n34 );
and ( n591 , n588 , n590 , n43 );
not ( n592 , n190 );
not ( n593 , n199 );
not ( n594 , n444 );
or ( n595 , n593 , n594 );
nand ( n596 , n595 , n43 );
or ( n597 , n592 , n596 );
not ( n598 , n201 );
not ( n599 , n399 );
and ( n600 , n598 , n599 );
and ( n601 , n154 , n43 );
nor ( n602 , n600 , n601 );
nand ( n603 , n211 , n43 );
nand ( n604 , n597 , n602 , n603 );
nor ( n605 , n591 , n604 );
nand ( n606 , n575 , n605 );
and ( n607 , n24 , n153 );
not ( n608 , n24 );
and ( n609 , n608 , n242 );
nor ( n610 , n607 , n609 );
not ( n611 , n610 );
nor ( n612 , n298 , n97 );
nand ( n613 , n611 , n612 , n287 );
nor ( n614 , n613 , n209 );
not ( n615 , n33 );
or ( n616 , n614 , n615 );
and ( n617 , n283 , n242 , n38 );
not ( n618 , n286 );
and ( n619 , n618 , n41 , n153 );
nor ( n620 , n617 , n619 );
not ( n621 , n620 );
buf ( n622 , n612 );
nand ( n623 , n621 , n622 , n22 );
nand ( n624 , n616 , n623 );
or ( n625 , n614 , n333 );
and ( n626 , n283 , n242 , n39 );
and ( n627 , n618 , n153 , n40 );
nor ( n628 , n626 , n627 );
not ( n629 , n628 );
nand ( n630 , n629 , n622 , n22 );
nand ( n631 , n625 , n630 );
nor ( n632 , n613 , n22 );
or ( n633 , n632 , n185 );
not ( n634 , n628 );
nand ( n635 , n634 , n622 , n209 );
nand ( n636 , n633 , n635 );
or ( n637 , n632 , n351 );
not ( n638 , n620 );
nand ( n639 , n638 , n622 , n209 );
nand ( n640 , n637 , n639 );
or ( n641 , n384 , n23 );
nand ( n642 , n641 , n524 );
and ( n643 , n642 , n29 );
nor ( n644 , n542 , n31 );
and ( n645 , n644 , n552 );
nor ( n646 , n643 , n645 );
or ( n647 , n646 , n356 );
not ( n648 , n46 );
nor ( n649 , n648 , n19 );
nor ( n650 , n615 , n34 );
nand ( n651 , n649 , n650 , n174 );
not ( n652 , n651 );
not ( n653 , n444 );
or ( n654 , n652 , n653 );
nor ( n655 , n199 , n29 );
nand ( n656 , n654 , n655 );
nand ( n657 , n656 , n201 );
nand ( n658 , n657 , n542 );
nand ( n659 , n647 , n658 );
not ( n660 , n24 );
nand ( n661 , n308 , n313 );
nor ( n662 , n307 , n8 );
nand ( n663 , n319 , n662 );
nand ( n664 , n661 , n663 );
not ( n665 , n664 );
or ( n666 , n660 , n665 );
not ( n667 , n116 );
not ( n668 , n667 );
and ( n669 , n530 , n11 );
not ( n670 , n669 );
or ( n671 , n668 , n670 );
and ( n672 , n530 , n110 );
not ( n673 , n40 );
nand ( n674 , n673 , n41 );
nor ( n675 , n674 , n81 );
nand ( n676 , n672 , n675 );
nand ( n677 , n671 , n676 );
and ( n678 , n677 , n152 );
not ( n679 , n13 );
nand ( n680 , n679 , n11 );
not ( n681 , n680 );
nor ( n682 , n40 , n41 );
and ( n683 , n681 , n682 , n81 , n278 );
and ( n684 , n683 , n533 );
nor ( n685 , n678 , n684 );
nand ( n686 , n666 , n685 );
not ( n687 , n461 );
not ( n688 , n339 );
or ( n689 , n687 , n688 );
nor ( n690 , n543 , n199 );
nand ( n691 , n689 , n690 );
not ( n692 , n644 );
nand ( n693 , n691 , n692 );
not ( n694 , n26 );
not ( n695 , n207 );
or ( n696 , n694 , n695 );
nand ( n697 , n523 , n77 );
nand ( n698 , n696 , n697 );
and ( n699 , n698 , n525 );
and ( n700 , n543 , n26 );
nor ( n701 , n699 , n700 );
or ( n702 , n701 , n356 );
and ( n703 , n198 , n524 );
nand ( n704 , n180 , n344 , n364 , n46 );
and ( n705 , n704 , n451 );
nand ( n706 , n524 , n25 );
nor ( n707 , n705 , n706 );
nor ( n708 , n703 , n707 );
nand ( n709 , n702 , n708 );
and ( n710 , n532 , n1 );
nor ( n711 , n710 , n223 );
not ( n712 , n531 );
not ( n713 , n712 );
and ( n714 , n121 , n5 );
not ( n715 , n42 );
or ( n716 , n715 , n5 );
not ( n717 , n3 );
nand ( n718 , n716 , n717 );
nor ( n719 , n714 , n718 );
or ( n720 , n719 , n1 );
nand ( n721 , n720 , n293 );
and ( n722 , n713 , n721 );
not ( n723 , n162 );
nor ( n724 , n722 , n723 );
nand ( n725 , n711 , n724 );
or ( n726 , n541 , n26 );
not ( n727 , n706 );
nand ( n728 , n726 , n727 );
nand ( n729 , n728 , n697 );
and ( n730 , n40 , n11 );
not ( n731 , n40 );
and ( n732 , n731 , n2 );
or ( n733 , n730 , n732 );
or ( n734 , n733 , n585 );
nand ( n735 , n674 , n2 );
nand ( n736 , n734 , n735 );
and ( n737 , n533 , n736 );
and ( n738 , n669 , n673 );
nor ( n739 , n737 , n738 );
or ( n740 , n739 , n151 );
not ( n741 , n13 );
or ( n742 , n712 , n741 );
nand ( n743 , n742 , n12 );
nand ( n744 , n740 , n743 );
and ( n745 , n107 , n4 );
nor ( n746 , n4 , n24 );
and ( n747 , n746 , n21 );
nor ( n748 , n747 , n5 );
nor ( n749 , n39 , n748 );
nor ( n750 , n120 , n230 , n24 , n5 );
nor ( n751 , n745 , n749 , n750 );
nand ( n752 , n531 , n1 );
or ( n753 , n751 , n752 , n3 );
nand ( n754 , n752 , n3 );
nand ( n755 , n753 , n754 );
or ( n756 , n674 , n12 );
or ( n757 , n151 , n40 );
nand ( n758 , n756 , n757 , n531 );
nand ( n759 , n758 , n11 );
not ( n760 , n240 );
nand ( n761 , n672 , n760 );
or ( n762 , n12 , n40 );
nand ( n763 , n762 , n681 );
not ( n764 , n12 );
nand ( n765 , n764 , n2 , n11 );
nand ( n766 , n759 , n761 , n763 , n765 );
and ( n767 , n717 , n5 );
not ( n768 , n107 );
and ( n769 , n768 , n717 );
nor ( n770 , n769 , n5 );
nor ( n771 , n767 , n770 , n752 );
not ( n772 , n4 );
or ( n773 , n771 , n772 );
not ( n774 , n243 );
nand ( n775 , n713 , n774 , n772 , n5 );
nand ( n776 , n773 , n775 );
or ( n777 , n680 , n682 );
or ( n778 , n278 , n13 );
nand ( n779 , n777 , n778 , n289 );
and ( n780 , n533 , n779 );
and ( n781 , n532 , n13 );
nor ( n782 , n780 , n781 );
nand ( n783 , n155 , n585 );
nand ( n784 , n782 , n783 );
nand ( n785 , n110 , n12 );
and ( n786 , n531 , n785 );
nor ( n787 , n786 , n81 );
nor ( n788 , n735 , n12 );
nand ( n789 , n765 , n289 );
nor ( n790 , n787 , n788 , n789 );
nand ( n791 , n669 , n81 , n760 );
nand ( n792 , n790 , n791 );
nor ( n793 , n783 , n534 );
or ( n794 , n692 , n126 );
or ( n795 , n424 , n644 );
nand ( n796 , n794 , n795 );
endmodule
