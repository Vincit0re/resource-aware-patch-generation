// Benchmark "top_top_miter" written by ABC on Tue Jul 05 22:48:42 2022

module top_top_miter ( 
    g0, g1, g10, g11, g12, g13, g14, g15, g16, g17, g18, g19, g2, g20, g21,
    g22, g23, g24, g25, g26, g27, g28, g29, g3, g30, g31, g32, g33, g34,
    g35, g36, g37, g38, g39, g4, g40, g41, g42, g43, g44, g45, g46, g47,
    g48, g49, g5, g50, g51, g52, g53, g54, g55, g56, g57, g58, g59, g6,
    g60, g61, g62, g63, g64, g65, g66, g67, g68, g69, g7, g70, g71, g72,
    g73, g74, g75, g76, g77, g78, g79, g8, g80, g81, g82, g83, g84, g85,
    g86, g87, g88, g89, g9, g90, g91, g92, g93, g94, g95, g96, g97, g98,
    miter  );
  input  g0, g1, g10, g11, g12, g13, g14, g15, g16, g17, g18, g19, g2,
    g20, g21, g22, g23, g24, g25, g26, g27, g28, g29, g3, g30, g31, g32,
    g33, g34, g35, g36, g37, g38, g39, g4, g40, g41, g42, g43, g44, g45,
    g46, g47, g48, g49, g5, g50, g51, g52, g53, g54, g55, g56, g57, g58,
    g59, g6, g60, g61, g62, g63, g64, g65, g66, g67, g68, g69, g7, g70,
    g71, g72, g73, g74, g75, g76, g77, g78, g79, g8, g80, g81, g82, g83,
    g84, g85, g86, g87, g88, g89, g9, g90, g91, g92, g93, g94, g95, g96,
    g97, g98;
  output miter;
  wire n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
    n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
    n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
    n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
    n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
    n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
    n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
    n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
    n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
    n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
    n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
    n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
    n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
    n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
    n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
    n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
    n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
    n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
    n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
    n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
    n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
    n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
    n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
    n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
    n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
    n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
    n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
    n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
    n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
    n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
    n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
    n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
    n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
    n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
    n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
    n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
    n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
    n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
    n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
    n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
    n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
    n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
    n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
    n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
    n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
    n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
    n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
    n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
    n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
    n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
    n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
    n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
    n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
    n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
    n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
    n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
    n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
    n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
    n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
    n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
    n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
    n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
    n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
    n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
    n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
    n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
    n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
    n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
    n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
    n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
    n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
    n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
    n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
    n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
    n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
    n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
    n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
    n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
    n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
    n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
    n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
    n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
    n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
    n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
    n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
    n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
    n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
    n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
    n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
    n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
    n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
    n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
    n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
    n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
    n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
    n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
    n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
    n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
    n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
    n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
    n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
    n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
    n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
    n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
    n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
    n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
    n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
    n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
    n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
    n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
    n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
    n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
    n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
    n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
    n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
    n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
    n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
    n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
    n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
    n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
    n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
    n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
    n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
    n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
    n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
    n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
    n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
    n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
    n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
    n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
    n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
    n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
    n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
    n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
    n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
    n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
    n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
    n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
    n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
    n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
    n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
    n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
    n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
    n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
    n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
    n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
    n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
    n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
    n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
    n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
    n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
    n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
    n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
    n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
    n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
    n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
    n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
    n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
    n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
    n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
    n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
    n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
    n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
    n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
    n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
    n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
    n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
    n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
    n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
    n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
    n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
    n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
    n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
    n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
    n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
    n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
    n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
    n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
    n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
    n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
    n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
    n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
    n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
    n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
    n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
    n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
    n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
    n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
    n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
    n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
    n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
    n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
    n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
    n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
    n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
    n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
    n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
    n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
    n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
    n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
    n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
    n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
    n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
    n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
    n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
    n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
    n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
    n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
    n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
    n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
    n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
    n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
    n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
    n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
    n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
    n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
    n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
    n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
    n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
    n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
    n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
    n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
    n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
    n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
    n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
    n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
    n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
    n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
    n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
    n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
    n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
    n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
    n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
    n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
    n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
    n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
    n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
    n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
    n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
    n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
    n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
    n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
    n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
    n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
    n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
    n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
    n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
    n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
    n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
    n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
    n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
    n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
    n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
    n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
    n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
    n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
    n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
    n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
    n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
    n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
    n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
    n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
    n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
    n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
    n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
    n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
    n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
    n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
    n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
    n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
    n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
    n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
    n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
    n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
    n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
    n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
    n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
    n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
    n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
    n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
    n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
    n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
    n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
    n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
    n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
    n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
    n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
    n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
    n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
    n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
    n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
    n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
    n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
    n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
    n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
    n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
    n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
    n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
    n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
    n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
    n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
    n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
    n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
    n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
    n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
    n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
    n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
    n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
    n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
    n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
    n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
    n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
    n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
    n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
    n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
    n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
    n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
    n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
    n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
    n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
    n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
    n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
    n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
    n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
    n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
    n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
    n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
    n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
    n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
    n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
    n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
    n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
    n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
    n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
    n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
    n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
    n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
    n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
    n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
    n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
    n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
    n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
    n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
    n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
    n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
    n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
    n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
    n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
    n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
    n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
    n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
    n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
    n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
    n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
    n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
    n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
    n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
    n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
    n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
    n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
    n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
    n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
    n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
    n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
    n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
    n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
    n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
    n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
    n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
    n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
    n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
    n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
    n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
    n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
    n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
    n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
    n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
    n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
    n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
    n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
    n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
    n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
    n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
    n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089,
    n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099,
    n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
    n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119,
    n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129,
    n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
    n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
    n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
    n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169,
    n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
    n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
    n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
    n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
    n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
    n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229,
    n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239,
    n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249,
    n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259,
    n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
    n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
    n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
    n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
    n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
    n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
    n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
    n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
    n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
    n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
    n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
    n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
    n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
    n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
    n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
    n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
    n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
    n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
    n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
    n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
    n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
    n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
    n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
    n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
    n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
    n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
    n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
    n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
    n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
    n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
    n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
    n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
    n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
    n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
    n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
    n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
    n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
    n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
    n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
    n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
    n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
    n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
    n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
    n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
    n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
    n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
    n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
    n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
    n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
    n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
    n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
    n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
    n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
    n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
    n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
    n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
    n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
    n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
    n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
    n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
    n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
    n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
    n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
    n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
    n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
    n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
    n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
    n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
    n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
    n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
    n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
    n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
    n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
    n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
    n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
    n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
    n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
    n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
    n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
    n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
    n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
    n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
    n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
    n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
    n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
    n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
    n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
    n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
    n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
    n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
    n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
    n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
    n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
    n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
    n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
    n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
    n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
    n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
    n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
    n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
    n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
    n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
    n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
    n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
    n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
    n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
    n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
    n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
    n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
    n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
    n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
    n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
    n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
    n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
    n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
    n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
    n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
    n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
    n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
    n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
    n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
    n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
    n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
    n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
    n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
    n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
    n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
    n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
    n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
    n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
    n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
    n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
    n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
    n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
    n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
    n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
    n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
    n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
    n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
    n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
    n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
    n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
    n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
    n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
    n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
    n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
    n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
    n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
    n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
    n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
    n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
    n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
    n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
    n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
    n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
    n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
    n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
    n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
    n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
    n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
    n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
    n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
    n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
    n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
    n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
    n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
    n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
    n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
    n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
    n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
    n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
    n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
    n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
    n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
    n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
    n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
    n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
    n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
    n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
    n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
    n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
    n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
    n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
    n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
    n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
    n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
    n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
    n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
    n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
    n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
    n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
    n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
    n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
    n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
    n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
    n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
    n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
    n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
    n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
    n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
    n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
    n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
    n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
    n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
    n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
    n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
    n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
    n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
    n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
    n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
    n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
    n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
    n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
    n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
    n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
    n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
    n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
    n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
    n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
    n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
    n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
    n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
    n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
    n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
    n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
    n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
    n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
    n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
    n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
    n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
    n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
    n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
    n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
    n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
    n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
    n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
    n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
    n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
    n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
    n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
    n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
    n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
    n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
    n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
    n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
    n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
    n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
    n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
    n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
    n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
    n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
    n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
    n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
    n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
    n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
    n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
    n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
    n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
    n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
    n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
    n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
    n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
    n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
    n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
    n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
    n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
    n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
    n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
    n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
    n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
    n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
    n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
    n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
    n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
    n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
    n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
    n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
    n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
    n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
    n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
    n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
    n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
    n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
    n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
    n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
    n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
    n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
    n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
    n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
    n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
    n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
    n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
    n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
    n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
    n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
    n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
    n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
    n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
    n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
    n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
    n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
    n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
    n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
    n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
    n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
    n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
    n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
    n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
    n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
    n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
    n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
    n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
    n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
    n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
    n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
    n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
    n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
    n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
    n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
    n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
    n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
    n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
    n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
    n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
    n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
    n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
    n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
    n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
    n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
    n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
    n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
    n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
    n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
    n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
    n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
    n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
    n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
    n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
    n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
    n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
    n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
    n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
    n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
    n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
    n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
    n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
    n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
    n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
    n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
    n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
    n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
    n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
    n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
    n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
    n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
    n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
    n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
    n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
    n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
    n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
    n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
    n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
    n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
    n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
    n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
    n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
    n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
    n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
    n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
    n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
    n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
    n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
    n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
    n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
    n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
    n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
    n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
    n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
    n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
    n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
    n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
    n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
    n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
    n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
    n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
    n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
    n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
    n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
    n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
    n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
    n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
    n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
    n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
    n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
    n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
    n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
    n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
    n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
    n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
    n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
    n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
    n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
    n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
    n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
    n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
    n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
    n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
    n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
    n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
    n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
    n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
    n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
    n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
    n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
    n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
    n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
    n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
    n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
    n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
    n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
    n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
    n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
    n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
    n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
    n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
    n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
    n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
    n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
    n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
    n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
    n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
    n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
    n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
    n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
    n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
    n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
    n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
    n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
    n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
    n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
    n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
    n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
    n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
    n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
    n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
    n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
    n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
    n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
    n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
    n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
    n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
    n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
    n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
    n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
    n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
    n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
    n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
    n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
    n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
    n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
    n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
    n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
    n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
    n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
    n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
    n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
    n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
    n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
    n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
    n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
    n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
    n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
    n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
    n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
    n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
    n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
    n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
    n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
    n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
    n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
    n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
    n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
    n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
    n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
    n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
    n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
    n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
    n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
    n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
    n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
    n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
    n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
    n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
    n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
    n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
    n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
    n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
    n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
    n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
    n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
    n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
    n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
    n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
    n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
    n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
    n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
    n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
    n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
    n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
    n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
    n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369,
    n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379,
    n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
    n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
    n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409,
    n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
    n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429,
    n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439,
    n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449,
    n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
    n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469,
    n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479,
    n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489,
    n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499,
    n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509,
    n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519,
    n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
    n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539,
    n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549,
    n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
    n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
    n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
    n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
    n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
    n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
    n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
    n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
    n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
    n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
    n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
    n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
    n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
    n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
    n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
    n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
    n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
    n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
    n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
    n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
    n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
    n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
    n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
    n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
    n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
    n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
    n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
    n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
    n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
    n9840, n9841;
  assign n101 = ~g38 & g39;
  assign n102 = g38 & ~g39;
  assign n103 = ~n101 & ~n102;
  assign n104 = ~g37 & g38;
  assign n105 = g37 & ~g38;
  assign n106 = ~n104 & ~n105;
  assign n107 = n103 & ~n106;
  assign n108 = g2 & g3;
  assign n109 = g19 & ~g2;
  assign n110 = ~n108 & ~n109;
  assign n111 = ~g37 & n110;
  assign n112 = g37 & ~n110;
  assign n113 = ~n111 & ~n112;
  assign n114 = n107 & n113;
  assign n115 = g37 & ~n103;
  assign n116 = ~n114 & ~n115;
  assign n117 = ~g36 & g37;
  assign n118 = g36 & ~g37;
  assign n119 = ~n117 & ~n118;
  assign n120 = g35 & g36;
  assign n121 = ~g35 & ~g36;
  assign n122 = ~n120 & ~n121;
  assign n123 = n119 & n122;
  assign n124 = g2 & g5;
  assign n125 = ~g2 & g21;
  assign n126 = ~n124 & ~n125;
  assign n127 = ~g35 & ~n126;
  assign n128 = g35 & n126;
  assign n129 = ~n127 & ~n128;
  assign n130 = n123 & ~n129;
  assign n131 = g2 & g4;
  assign n132 = ~g2 & g20;
  assign n133 = ~n131 & ~n132;
  assign n134 = ~g35 & n133;
  assign n135 = g35 & ~n133;
  assign n136 = ~n134 & ~n135;
  assign n137 = ~n119 & n136;
  assign n138 = ~n130 & ~n137;
  assign n139 = g2 & ~g6;
  assign n140 = ~g2 & ~g22;
  assign n141 = ~n139 & ~n140;
  assign n142 = g35 & n141;
  assign n143 = ~n116 & n142;
  assign n144 = n116 & ~n142;
  assign n145 = ~n143 & ~n144;
  assign n146 = ~n138 & ~n145;
  assign n147 = n116 & n142;
  assign n148 = ~n146 & ~n147;
  assign n149 = ~n116 & n148;
  assign n150 = n116 & ~n148;
  assign n151 = ~n149 & ~n150;
  assign n152 = n123 & n136;
  assign n153 = ~g35 & n110;
  assign n154 = g35 & ~n110;
  assign n155 = ~n153 & ~n154;
  assign n156 = ~n119 & n155;
  assign n157 = ~n152 & ~n156;
  assign n158 = g35 & ~n126;
  assign n159 = n103 & ~n107;
  assign n160 = g37 & ~n159;
  assign n161 = n158 & n160;
  assign n162 = ~n158 & ~n160;
  assign n163 = ~n161 & ~n162;
  assign n164 = ~n157 & n163;
  assign n165 = n157 & ~n163;
  assign n166 = ~n164 & ~n165;
  assign n167 = ~n151 & n166;
  assign n168 = n151 & ~n166;
  assign n169 = ~n167 & ~n168;
  assign n170 = ~g39 & g40;
  assign n171 = g39 & ~g40;
  assign n172 = ~n170 & ~n171;
  assign n173 = ~g40 & g41;
  assign n174 = g40 & ~g41;
  assign n175 = ~n173 & ~n174;
  assign n176 = ~n172 & n175;
  assign n177 = g39 & n110;
  assign n178 = ~g39 & ~n110;
  assign n179 = ~n177 & ~n178;
  assign n180 = n176 & ~n179;
  assign n181 = g39 & ~n175;
  assign n182 = ~n180 & ~n181;
  assign n183 = ~g35 & n141;
  assign n184 = g35 & ~n141;
  assign n185 = ~n183 & ~n184;
  assign n186 = n123 & ~n185;
  assign n187 = ~n119 & ~n129;
  assign n188 = ~n186 & ~n187;
  assign n189 = ~n182 & ~n188;
  assign n190 = n182 & n188;
  assign n191 = ~n189 & ~n190;
  assign n192 = g2 & g8;
  assign n193 = ~g2 & g24;
  assign n194 = ~n192 & ~n193;
  assign n195 = g35 & ~n194;
  assign n196 = g2 & g7;
  assign n197 = ~g2 & g23;
  assign n198 = ~n196 & ~n197;
  assign n199 = g35 & ~n198;
  assign n200 = ~g35 & n198;
  assign n201 = ~n199 & ~n200;
  assign n202 = n123 & n201;
  assign n203 = ~n119 & ~n185;
  assign n204 = ~n202 & ~n203;
  assign n205 = n195 & ~n204;
  assign n206 = ~g37 & ~n126;
  assign n207 = g37 & n126;
  assign n208 = ~n206 & ~n207;
  assign n209 = n107 & ~n208;
  assign n210 = ~g37 & ~n133;
  assign n211 = g37 & n133;
  assign n212 = ~n210 & ~n211;
  assign n213 = ~n103 & ~n212;
  assign n214 = ~n209 & ~n213;
  assign n215 = ~n195 & ~n204;
  assign n216 = n195 & n204;
  assign n217 = ~n215 & ~n216;
  assign n218 = ~n214 & ~n217;
  assign n219 = ~n205 & ~n218;
  assign n220 = n191 & ~n219;
  assign n221 = ~n189 & ~n220;
  assign n222 = ~n103 & n113;
  assign n223 = n107 & ~n212;
  assign n224 = ~n222 & ~n223;
  assign n225 = n175 & ~n176;
  assign n226 = g39 & ~n225;
  assign n227 = ~n199 & ~n226;
  assign n228 = n199 & n226;
  assign n229 = ~n227 & ~n228;
  assign n230 = ~n224 & ~n229;
  assign n231 = n199 & ~n226;
  assign n232 = ~n230 & ~n231;
  assign n233 = n138 & ~n145;
  assign n234 = ~n138 & n145;
  assign n235 = ~n233 & ~n234;
  assign n236 = ~n232 & n235;
  assign n237 = n232 & ~n235;
  assign n238 = ~n236 & ~n237;
  assign n239 = ~n221 & ~n238;
  assign n240 = ~n232 & ~n235;
  assign n241 = ~n239 & ~n240;
  assign n242 = ~n169 & ~n241;
  assign n243 = n169 & n241;
  assign n244 = ~n242 & ~n243;
  assign n245 = ~n221 & n238;
  assign n246 = n221 & ~n238;
  assign n247 = ~n245 & ~n246;
  assign n248 = n224 & ~n229;
  assign n249 = ~n224 & n229;
  assign n250 = ~n248 & ~n249;
  assign n251 = ~n191 & ~n219;
  assign n252 = n191 & n219;
  assign n253 = ~n251 & ~n252;
  assign n254 = n250 & ~n253;
  assign n255 = ~n250 & n253;
  assign n256 = ~n254 & ~n255;
  assign n257 = n214 & ~n217;
  assign n258 = ~n214 & n217;
  assign n259 = ~n257 & ~n258;
  assign n260 = ~g42 & g43;
  assign n261 = g42 & ~g43;
  assign n262 = ~n260 & ~n261;
  assign n263 = ~g41 & g42;
  assign n264 = g41 & ~g42;
  assign n265 = ~n263 & ~n264;
  assign n266 = n262 & ~n265;
  assign n267 = n262 & ~n266;
  assign n268 = g41 & ~n267;
  assign n269 = ~n119 & n201;
  assign n270 = ~g35 & ~n194;
  assign n271 = g35 & n194;
  assign n272 = ~n270 & ~n271;
  assign n273 = n123 & ~n272;
  assign n274 = ~n269 & ~n273;
  assign n275 = ~n268 & ~n274;
  assign n276 = g39 & n133;
  assign n277 = ~g39 & ~n133;
  assign n278 = ~n276 & ~n277;
  assign n279 = n176 & ~n278;
  assign n280 = ~n175 & ~n179;
  assign n281 = ~n279 & ~n280;
  assign n282 = ~n268 & n274;
  assign n283 = n268 & ~n274;
  assign n284 = ~n282 & ~n283;
  assign n285 = ~n281 & ~n284;
  assign n286 = ~n275 & ~n285;
  assign n287 = n182 & n286;
  assign n288 = ~n182 & ~n286;
  assign n289 = ~n287 & ~n288;
  assign n290 = ~n259 & ~n289;
  assign n291 = n182 & ~n286;
  assign n292 = ~n290 & ~n291;
  assign n293 = ~n256 & ~n292;
  assign n294 = ~n250 & ~n253;
  assign n295 = ~n293 & ~n294;
  assign n296 = n247 & n295;
  assign n297 = n256 & ~n292;
  assign n298 = ~n256 & n292;
  assign n299 = ~n297 & ~n298;
  assign n300 = g41 & n110;
  assign n301 = ~g41 & ~n110;
  assign n302 = ~n300 & ~n301;
  assign n303 = n266 & ~n302;
  assign n304 = g41 & ~n262;
  assign n305 = ~n303 & ~n304;
  assign n306 = ~g10 & g2;
  assign n307 = ~g2 & ~g26;
  assign n308 = ~n306 & ~n307;
  assign n309 = g35 & n308;
  assign n310 = ~n305 & n309;
  assign n311 = ~n119 & ~n272;
  assign n312 = g2 & ~g9;
  assign n313 = ~g2 & ~g25;
  assign n314 = ~n312 & ~n313;
  assign n315 = ~g35 & ~n314;
  assign n316 = g35 & n314;
  assign n317 = ~n315 & ~n316;
  assign n318 = n123 & n317;
  assign n319 = ~n311 & ~n318;
  assign n320 = n305 & ~n309;
  assign n321 = ~n310 & ~n320;
  assign n322 = ~n319 & n321;
  assign n323 = ~n310 & ~n322;
  assign n324 = ~n281 & n284;
  assign n325 = n281 & ~n284;
  assign n326 = ~n324 & ~n325;
  assign n327 = ~n323 & ~n326;
  assign n328 = ~g37 & ~n141;
  assign n329 = g37 & n141;
  assign n330 = ~n328 & ~n329;
  assign n331 = n107 & n330;
  assign n332 = ~n103 & ~n208;
  assign n333 = ~n331 & ~n332;
  assign n334 = n316 & n333;
  assign n335 = ~n316 & ~n333;
  assign n336 = ~n334 & ~n335;
  assign n337 = g39 & n126;
  assign n338 = ~g39 & ~n126;
  assign n339 = ~n337 & ~n338;
  assign n340 = n176 & ~n339;
  assign n341 = ~n175 & ~n278;
  assign n342 = ~n340 & ~n341;
  assign n343 = ~n336 & ~n342;
  assign n344 = n336 & n342;
  assign n345 = ~n343 & ~n344;
  assign n346 = n323 & n326;
  assign n347 = ~n327 & ~n346;
  assign n348 = n345 & n347;
  assign n349 = ~n327 & ~n348;
  assign n350 = ~n259 & n289;
  assign n351 = n259 & ~n289;
  assign n352 = ~n350 & ~n351;
  assign n353 = n316 & ~n333;
  assign n354 = ~n343 & ~n353;
  assign n355 = ~n352 & n354;
  assign n356 = n352 & ~n354;
  assign n357 = ~n355 & ~n356;
  assign n358 = ~n349 & ~n357;
  assign n359 = ~n352 & ~n354;
  assign n360 = ~n358 & ~n359;
  assign n361 = n299 & n360;
  assign n362 = ~g41 & ~n133;
  assign n363 = g41 & n133;
  assign n364 = ~n362 & ~n363;
  assign n365 = n266 & ~n364;
  assign n366 = ~n262 & ~n302;
  assign n367 = ~n365 & ~n366;
  assign n368 = ~g44 & g45;
  assign n369 = g44 & ~g45;
  assign n370 = ~n368 & ~n369;
  assign n371 = ~g43 & ~g44;
  assign n372 = g43 & g44;
  assign n373 = ~n371 & ~n372;
  assign n374 = n370 & n373;
  assign n375 = n370 & ~n374;
  assign n376 = g43 & ~n375;
  assign n377 = g37 & n198;
  assign n378 = ~g37 & ~n198;
  assign n379 = ~n377 & ~n378;
  assign n380 = ~n103 & ~n379;
  assign n381 = ~g37 & ~n194;
  assign n382 = g37 & n194;
  assign n383 = ~n381 & ~n382;
  assign n384 = n107 & ~n383;
  assign n385 = ~n380 & ~n384;
  assign n386 = n376 & ~n385;
  assign n387 = ~n376 & n385;
  assign n388 = ~n386 & ~n387;
  assign n389 = ~n367 & ~n388;
  assign n390 = ~n376 & ~n385;
  assign n391 = ~n389 & ~n390;
  assign n392 = n319 & n321;
  assign n393 = ~n319 & ~n321;
  assign n394 = ~n392 & ~n393;
  assign n395 = ~n391 & ~n394;
  assign n396 = ~n119 & n317;
  assign n397 = ~g35 & n308;
  assign n398 = g35 & ~n308;
  assign n399 = ~n397 & ~n398;
  assign n400 = n123 & ~n399;
  assign n401 = ~n396 & ~n400;
  assign n402 = g11 & g2;
  assign n403 = ~g2 & g27;
  assign n404 = ~n402 & ~n403;
  assign n405 = g35 & ~n404;
  assign n406 = ~n175 & ~n339;
  assign n407 = g39 & ~n141;
  assign n408 = ~g39 & n141;
  assign n409 = ~n407 & ~n408;
  assign n410 = n176 & ~n409;
  assign n411 = ~n406 & ~n410;
  assign n412 = ~n405 & ~n411;
  assign n413 = n405 & n411;
  assign n414 = ~n412 & ~n413;
  assign n415 = ~n401 & ~n414;
  assign n416 = n405 & ~n411;
  assign n417 = ~n415 & ~n416;
  assign n418 = ~n103 & n330;
  assign n419 = n107 & ~n379;
  assign n420 = ~n418 & ~n419;
  assign n421 = n342 & ~n420;
  assign n422 = ~n342 & n420;
  assign n423 = ~n421 & ~n422;
  assign n424 = n417 & n423;
  assign n425 = ~n417 & ~n423;
  assign n426 = ~n424 & ~n425;
  assign n427 = n391 & n394;
  assign n428 = ~n395 & ~n427;
  assign n429 = ~n426 & n428;
  assign n430 = ~n395 & ~n429;
  assign n431 = ~n417 & n423;
  assign n432 = ~n421 & ~n431;
  assign n433 = n345 & ~n347;
  assign n434 = ~n345 & n347;
  assign n435 = ~n433 & ~n434;
  assign n436 = n432 & ~n435;
  assign n437 = ~n432 & n435;
  assign n438 = ~n436 & ~n437;
  assign n439 = ~n430 & ~n438;
  assign n440 = ~n432 & ~n435;
  assign n441 = ~n439 & ~n440;
  assign n442 = ~n349 & n357;
  assign n443 = n349 & ~n357;
  assign n444 = ~n442 & ~n443;
  assign n445 = n441 & n444;
  assign n446 = n401 & ~n414;
  assign n447 = ~n401 & n414;
  assign n448 = ~n446 & ~n447;
  assign n449 = g41 & n126;
  assign n450 = ~g41 & ~n126;
  assign n451 = ~n449 & ~n450;
  assign n452 = n266 & ~n451;
  assign n453 = ~n262 & ~n364;
  assign n454 = ~n452 & ~n453;
  assign n455 = g43 & n110;
  assign n456 = ~g43 & ~n110;
  assign n457 = ~n455 & ~n456;
  assign n458 = n374 & ~n457;
  assign n459 = g43 & ~n370;
  assign n460 = ~n458 & ~n459;
  assign n461 = ~g35 & n404;
  assign n462 = ~n405 & ~n461;
  assign n463 = n123 & n462;
  assign n464 = ~n119 & ~n399;
  assign n465 = ~n463 & ~n464;
  assign n466 = ~n460 & ~n465;
  assign n467 = g37 & ~n314;
  assign n468 = ~g37 & n314;
  assign n469 = ~n467 & ~n468;
  assign n470 = n107 & ~n469;
  assign n471 = ~n103 & ~n383;
  assign n472 = ~n470 & ~n471;
  assign n473 = n460 & n465;
  assign n474 = ~n472 & ~n473;
  assign n475 = ~n466 & ~n474;
  assign n476 = n454 & ~n475;
  assign n477 = ~n454 & n475;
  assign n478 = ~n476 & ~n477;
  assign n479 = ~n448 & ~n478;
  assign n480 = ~n454 & ~n475;
  assign n481 = ~n479 & ~n480;
  assign n482 = n426 & n428;
  assign n483 = ~n426 & ~n428;
  assign n484 = ~n482 & ~n483;
  assign n485 = ~n481 & ~n484;
  assign n486 = n448 & ~n478;
  assign n487 = ~n448 & n478;
  assign n488 = ~n486 & ~n487;
  assign n489 = g12 & g2;
  assign n490 = ~g2 & g28;
  assign n491 = ~n489 & ~n490;
  assign n492 = g35 & ~n491;
  assign n493 = ~n454 & n492;
  assign n494 = n454 & ~n492;
  assign n495 = ~n493 & ~n494;
  assign n496 = g39 & n198;
  assign n497 = ~g39 & ~n198;
  assign n498 = ~n496 & ~n497;
  assign n499 = n176 & ~n498;
  assign n500 = ~n175 & ~n409;
  assign n501 = ~n499 & ~n500;
  assign n502 = ~n495 & ~n501;
  assign n503 = n454 & n492;
  assign n504 = ~n502 & ~n503;
  assign n505 = n367 & ~n388;
  assign n506 = ~n367 & n388;
  assign n507 = ~n505 & ~n506;
  assign n508 = ~n504 & n507;
  assign n509 = n504 & ~n507;
  assign n510 = ~n508 & ~n509;
  assign n511 = ~n488 & ~n510;
  assign n512 = ~n504 & ~n507;
  assign n513 = ~n511 & ~n512;
  assign n514 = ~n481 & n484;
  assign n515 = n481 & ~n484;
  assign n516 = ~n514 & ~n515;
  assign n517 = ~n513 & ~n516;
  assign n518 = ~n485 & ~n517;
  assign n519 = n430 & ~n438;
  assign n520 = ~n430 & n438;
  assign n521 = ~n519 & ~n520;
  assign n522 = ~n518 & ~n521;
  assign n523 = n518 & n521;
  assign n524 = n513 & ~n516;
  assign n525 = ~n513 & n516;
  assign n526 = ~n524 & ~n525;
  assign n527 = ~g46 & g47;
  assign n528 = g46 & ~g47;
  assign n529 = ~n527 & ~n528;
  assign n530 = ~g45 & ~g46;
  assign n531 = g45 & g46;
  assign n532 = ~n530 & ~n531;
  assign n533 = n529 & n532;
  assign n534 = g45 & n110;
  assign n535 = ~g45 & ~n110;
  assign n536 = ~n534 & ~n535;
  assign n537 = n533 & ~n536;
  assign n538 = g45 & ~n529;
  assign n539 = ~n537 & ~n538;
  assign n540 = g13 & g2;
  assign n541 = ~g2 & g29;
  assign n542 = ~n540 & ~n541;
  assign n543 = g35 & ~n542;
  assign n544 = ~n539 & n543;
  assign n545 = n539 & ~n543;
  assign n546 = ~n544 & ~n545;
  assign n547 = ~g37 & n404;
  assign n548 = g37 & ~n404;
  assign n549 = ~n547 & ~n548;
  assign n550 = n107 & n549;
  assign n551 = ~g37 & n308;
  assign n552 = g37 & ~n308;
  assign n553 = ~n551 & ~n552;
  assign n554 = ~n103 & ~n553;
  assign n555 = ~n550 & ~n554;
  assign n556 = ~g43 & ~n126;
  assign n557 = g43 & n126;
  assign n558 = ~n556 & ~n557;
  assign n559 = n374 & ~n558;
  assign n560 = ~g43 & ~n133;
  assign n561 = g43 & n133;
  assign n562 = ~n560 & ~n561;
  assign n563 = ~n370 & ~n562;
  assign n564 = ~n559 & ~n563;
  assign n565 = ~n555 & ~n564;
  assign n566 = n555 & n564;
  assign n567 = ~g39 & n314;
  assign n568 = g39 & ~n314;
  assign n569 = ~n567 & ~n568;
  assign n570 = n176 & ~n569;
  assign n571 = ~g39 & ~n194;
  assign n572 = g39 & n194;
  assign n573 = ~n571 & ~n572;
  assign n574 = ~n175 & ~n573;
  assign n575 = ~n570 & ~n574;
  assign n576 = ~n566 & ~n575;
  assign n577 = ~n565 & ~n576;
  assign n578 = n546 & ~n577;
  assign n579 = ~n544 & ~n578;
  assign n580 = n495 & n501;
  assign n581 = ~n502 & ~n580;
  assign n582 = n579 & n581;
  assign n583 = ~n579 & ~n581;
  assign n584 = ~n582 & ~n583;
  assign n585 = g41 & ~n198;
  assign n586 = ~g41 & n198;
  assign n587 = ~n585 & ~n586;
  assign n588 = n266 & n587;
  assign n589 = ~g41 & ~n141;
  assign n590 = g41 & n141;
  assign n591 = ~n589 & ~n590;
  assign n592 = ~n262 & n591;
  assign n593 = ~n588 & ~n592;
  assign n594 = g14 & g2;
  assign n595 = ~g2 & g30;
  assign n596 = ~n594 & ~n595;
  assign n597 = g35 & ~n596;
  assign n598 = g35 & n491;
  assign n599 = ~g35 & ~n491;
  assign n600 = ~n598 & ~n599;
  assign n601 = ~n119 & ~n600;
  assign n602 = g35 & n542;
  assign n603 = ~g35 & ~n542;
  assign n604 = ~n602 & ~n603;
  assign n605 = n123 & ~n604;
  assign n606 = ~n601 & ~n605;
  assign n607 = n597 & n606;
  assign n608 = ~n597 & ~n606;
  assign n609 = ~n607 & ~n608;
  assign n610 = ~n593 & ~n609;
  assign n611 = n597 & ~n606;
  assign n612 = ~n610 & ~n611;
  assign n613 = ~n175 & ~n498;
  assign n614 = n176 & ~n573;
  assign n615 = ~n613 & ~n614;
  assign n616 = n529 & ~n533;
  assign n617 = g45 & ~n616;
  assign n618 = ~n370 & ~n457;
  assign n619 = n374 & ~n562;
  assign n620 = ~n618 & ~n619;
  assign n621 = n617 & ~n620;
  assign n622 = ~n617 & n620;
  assign n623 = ~n621 & ~n622;
  assign n624 = n615 & ~n623;
  assign n625 = ~n615 & n623;
  assign n626 = ~n624 & ~n625;
  assign n627 = n612 & ~n626;
  assign n628 = ~n612 & n626;
  assign n629 = ~n627 & ~n628;
  assign n630 = ~n262 & ~n451;
  assign n631 = n266 & n591;
  assign n632 = ~n630 & ~n631;
  assign n633 = ~n103 & ~n469;
  assign n634 = n107 & ~n553;
  assign n635 = ~n633 & ~n634;
  assign n636 = ~n632 & ~n635;
  assign n637 = n632 & n635;
  assign n638 = ~n636 & ~n637;
  assign n639 = n123 & ~n600;
  assign n640 = ~n119 & n462;
  assign n641 = ~n639 & ~n640;
  assign n642 = ~n638 & ~n641;
  assign n643 = n638 & n641;
  assign n644 = ~n642 & ~n643;
  assign n645 = ~n629 & ~n644;
  assign n646 = ~n612 & ~n626;
  assign n647 = ~n645 & ~n646;
  assign n648 = ~n584 & ~n647;
  assign n649 = ~n579 & n581;
  assign n650 = ~n648 & ~n649;
  assign n651 = ~n460 & n472;
  assign n652 = n460 & ~n472;
  assign n653 = ~n651 & ~n652;
  assign n654 = ~n465 & n653;
  assign n655 = n465 & ~n653;
  assign n656 = ~n654 & ~n655;
  assign n657 = ~n615 & ~n623;
  assign n658 = ~n617 & ~n620;
  assign n659 = ~n657 & ~n658;
  assign n660 = n638 & ~n641;
  assign n661 = ~n636 & ~n660;
  assign n662 = n659 & ~n661;
  assign n663 = ~n659 & n661;
  assign n664 = ~n662 & ~n663;
  assign n665 = ~n656 & ~n664;
  assign n666 = ~n659 & ~n661;
  assign n667 = ~n665 & ~n666;
  assign n668 = ~n488 & n510;
  assign n669 = n488 & ~n510;
  assign n670 = ~n668 & ~n669;
  assign n671 = ~n667 & n670;
  assign n672 = n667 & ~n670;
  assign n673 = ~n671 & ~n672;
  assign n674 = ~n650 & ~n673;
  assign n675 = ~n667 & ~n670;
  assign n676 = ~n674 & ~n675;
  assign n677 = ~n526 & ~n676;
  assign n678 = ~n523 & n677;
  assign n679 = ~n522 & ~n678;
  assign n680 = ~n445 & ~n679;
  assign n681 = ~n441 & ~n444;
  assign n682 = ~n680 & ~n681;
  assign n683 = ~n361 & ~n682;
  assign n684 = ~n299 & ~n360;
  assign n685 = ~n683 & ~n684;
  assign n686 = ~n296 & ~n685;
  assign n687 = ~n247 & ~n295;
  assign n688 = n526 & n676;
  assign n689 = ~n523 & ~n688;
  assign n690 = ~n445 & n689;
  assign n691 = n650 & ~n673;
  assign n692 = ~n650 & n673;
  assign n693 = ~n691 & ~n692;
  assign n694 = n194 & n198;
  assign n695 = ~n194 & ~n198;
  assign n696 = ~n194 & n314;
  assign n697 = n194 & ~n314;
  assign n698 = ~n696 & ~n697;
  assign n699 = ~n695 & ~n698;
  assign n700 = ~n694 & n699;
  assign n701 = g42 & ~n198;
  assign n702 = ~g42 & n198;
  assign n703 = ~n701 & ~n702;
  assign n704 = n700 & n703;
  assign n705 = n587 & n698;
  assign n706 = ~n704 & ~n705;
  assign n707 = g47 & ~n110;
  assign n708 = ~n308 & n404;
  assign n709 = n308 & ~n404;
  assign n710 = ~n708 & ~n709;
  assign n711 = ~n569 & n710;
  assign n712 = n308 & n314;
  assign n713 = ~n308 & ~n314;
  assign n714 = ~n712 & ~n713;
  assign n715 = ~n710 & n714;
  assign n716 = ~g40 & ~n314;
  assign n717 = g40 & n314;
  assign n718 = ~n716 & ~n717;
  assign n719 = n715 & n718;
  assign n720 = ~n711 & ~n719;
  assign n721 = n707 & n720;
  assign n722 = ~n707 & ~n720;
  assign n723 = ~n721 & ~n722;
  assign n724 = n706 & ~n723;
  assign n725 = ~n706 & n723;
  assign n726 = ~n724 & ~n725;
  assign n727 = ~n126 & n141;
  assign n728 = ~n141 & n198;
  assign n729 = n141 & ~n198;
  assign n730 = ~n728 & ~n729;
  assign n731 = n126 & ~n141;
  assign n732 = ~n730 & ~n731;
  assign n733 = ~n727 & n732;
  assign n734 = g44 & ~n126;
  assign n735 = ~g44 & n126;
  assign n736 = ~n734 & ~n735;
  assign n737 = n733 & n736;
  assign n738 = ~n558 & n730;
  assign n739 = ~n737 & ~n738;
  assign n740 = n491 & n542;
  assign n741 = ~n491 & ~n542;
  assign n742 = ~n740 & ~n741;
  assign n743 = n549 & n742;
  assign n744 = n404 & n491;
  assign n745 = ~n404 & ~n491;
  assign n746 = ~n744 & ~n745;
  assign n747 = ~n742 & n746;
  assign n748 = ~g38 & n404;
  assign n749 = g38 & ~n404;
  assign n750 = ~n748 & ~n749;
  assign n751 = n747 & n750;
  assign n752 = ~n743 & ~n751;
  assign n753 = ~n739 & n752;
  assign n754 = n739 & ~n752;
  assign n755 = ~n753 & ~n754;
  assign n756 = ~n126 & n133;
  assign n757 = n126 & ~n133;
  assign n758 = ~n756 & ~n757;
  assign n759 = n110 & n133;
  assign n760 = ~n110 & ~n133;
  assign n761 = ~n759 & ~n760;
  assign n762 = n758 & n761;
  assign n763 = g46 & ~n110;
  assign n764 = ~g46 & n110;
  assign n765 = ~n763 & ~n764;
  assign n766 = n762 & n765;
  assign n767 = ~n536 & ~n758;
  assign n768 = ~n766 & ~n767;
  assign n769 = ~n755 & n768;
  assign n770 = n755 & ~n768;
  assign n771 = ~n769 & ~n770;
  assign n772 = ~g15 & g2;
  assign n773 = ~g2 & ~g31;
  assign n774 = ~n772 & ~n773;
  assign n775 = ~n596 & ~n774;
  assign n776 = n596 & n774;
  assign n777 = ~n775 & ~n776;
  assign n778 = n542 & ~n596;
  assign n779 = ~n542 & n596;
  assign n780 = ~n778 & ~n779;
  assign n781 = n777 & ~n780;
  assign n782 = ~g36 & n542;
  assign n783 = g36 & ~n542;
  assign n784 = ~n782 & ~n783;
  assign n785 = n781 & n784;
  assign n786 = ~n604 & ~n777;
  assign n787 = ~n785 & ~n786;
  assign n788 = n774 & n787;
  assign n789 = ~n774 & ~n787;
  assign n790 = ~n788 & ~n789;
  assign n791 = n771 & ~n790;
  assign n792 = ~n771 & n790;
  assign n793 = ~n791 & ~n792;
  assign n794 = ~n726 & ~n793;
  assign n795 = ~n771 & ~n790;
  assign n796 = ~n794 & ~n795;
  assign n797 = g39 & ~n404;
  assign n798 = ~g39 & n404;
  assign n799 = ~n797 & ~n798;
  assign n800 = n747 & n799;
  assign n801 = n742 & n750;
  assign n802 = ~n800 & ~n801;
  assign n803 = ~g45 & ~n126;
  assign n804 = g45 & n126;
  assign n805 = ~n803 & ~n804;
  assign n806 = n733 & ~n805;
  assign n807 = n730 & n736;
  assign n808 = ~n806 & ~n807;
  assign n809 = ~n802 & ~n808;
  assign n810 = g47 & n110;
  assign n811 = ~g47 & ~n110;
  assign n812 = ~n810 & ~n811;
  assign n813 = n762 & ~n812;
  assign n814 = ~n758 & n765;
  assign n815 = ~n813 & ~n814;
  assign n816 = n802 & n808;
  assign n817 = ~n809 & ~n816;
  assign n818 = ~n815 & n817;
  assign n819 = ~n809 & ~n818;
  assign n820 = g16 & g2;
  assign n821 = ~g2 & g32;
  assign n822 = ~n820 & ~n821;
  assign n823 = n774 & n822;
  assign n824 = g35 & ~n774;
  assign n825 = ~g35 & n774;
  assign n826 = ~n824 & ~n825;
  assign n827 = n823 & ~n826;
  assign n828 = n774 & ~n822;
  assign n829 = ~n827 & ~n828;
  assign n830 = ~n777 & n784;
  assign n831 = ~g37 & n542;
  assign n832 = g37 & ~n542;
  assign n833 = ~n831 & ~n832;
  assign n834 = n781 & n833;
  assign n835 = ~n830 & ~n834;
  assign n836 = ~n829 & ~n835;
  assign n837 = g41 & ~n314;
  assign n838 = ~g41 & n314;
  assign n839 = ~n837 & ~n838;
  assign n840 = n715 & ~n839;
  assign n841 = n710 & n718;
  assign n842 = ~n840 & ~n841;
  assign n843 = g48 & ~n110;
  assign n844 = ~n842 & n843;
  assign n845 = ~g43 & ~n198;
  assign n846 = g43 & n198;
  assign n847 = ~n845 & ~n846;
  assign n848 = n700 & ~n847;
  assign n849 = n698 & n703;
  assign n850 = ~n848 & ~n849;
  assign n851 = n842 & ~n843;
  assign n852 = ~n844 & ~n851;
  assign n853 = ~n850 & n852;
  assign n854 = ~n844 & ~n853;
  assign n855 = n836 & n854;
  assign n856 = ~n836 & ~n854;
  assign n857 = ~n855 & ~n856;
  assign n858 = ~n819 & ~n857;
  assign n859 = n836 & ~n854;
  assign n860 = ~n858 & ~n859;
  assign n861 = ~n706 & ~n723;
  assign n862 = n707 & ~n720;
  assign n863 = ~n861 & ~n862;
  assign n864 = ~n604 & n781;
  assign n865 = ~n542 & ~n777;
  assign n866 = ~n864 & ~n865;
  assign n867 = ~n788 & n866;
  assign n868 = n788 & ~n866;
  assign n869 = ~n867 & ~n868;
  assign n870 = ~n863 & ~n869;
  assign n871 = n863 & n869;
  assign n872 = ~n870 & ~n871;
  assign n873 = ~n860 & n872;
  assign n874 = n860 & ~n872;
  assign n875 = ~n873 & ~n874;
  assign n876 = ~n796 & ~n875;
  assign n877 = ~n860 & ~n872;
  assign n878 = ~n876 & ~n877;
  assign n879 = ~g38 & ~n314;
  assign n880 = g38 & n314;
  assign n881 = ~n879 & ~n880;
  assign n882 = n710 & n881;
  assign n883 = ~n569 & n715;
  assign n884 = ~n882 & ~n883;
  assign n885 = ~n536 & n762;
  assign n886 = g44 & ~n110;
  assign n887 = ~g44 & n110;
  assign n888 = ~n886 & ~n887;
  assign n889 = ~n758 & n888;
  assign n890 = ~n885 & ~n889;
  assign n891 = n884 & ~n890;
  assign n892 = ~n884 & n890;
  assign n893 = ~n891 & ~n892;
  assign n894 = n763 & n893;
  assign n895 = ~n763 & ~n893;
  assign n896 = ~n894 & ~n895;
  assign n897 = ~n755 & ~n768;
  assign n898 = ~n739 & ~n752;
  assign n899 = ~n897 & ~n898;
  assign n900 = n896 & ~n899;
  assign n901 = ~n896 & n899;
  assign n902 = ~n900 & ~n901;
  assign n903 = ~n558 & n733;
  assign n904 = g42 & ~n126;
  assign n905 = ~g42 & n126;
  assign n906 = ~n904 & ~n905;
  assign n907 = n730 & n906;
  assign n908 = ~n903 & ~n907;
  assign n909 = n549 & n747;
  assign n910 = g36 & ~n404;
  assign n911 = ~g36 & n404;
  assign n912 = ~n910 & ~n911;
  assign n913 = n742 & n912;
  assign n914 = ~n909 & ~n913;
  assign n915 = n587 & n700;
  assign n916 = g40 & ~n198;
  assign n917 = ~g40 & n198;
  assign n918 = ~n916 & ~n917;
  assign n919 = n698 & n918;
  assign n920 = ~n915 & ~n919;
  assign n921 = n914 & ~n920;
  assign n922 = ~n914 & n920;
  assign n923 = ~n921 & ~n922;
  assign n924 = n908 & ~n923;
  assign n925 = ~n908 & n923;
  assign n926 = ~n924 & ~n925;
  assign n927 = ~n902 & ~n926;
  assign n928 = ~n896 & ~n899;
  assign n929 = ~n927 & ~n928;
  assign n930 = ~n863 & n869;
  assign n931 = ~n867 & ~n930;
  assign n932 = g45 & ~n110;
  assign n933 = ~n866 & n932;
  assign n934 = n866 & ~n932;
  assign n935 = ~n933 & ~n934;
  assign n936 = ~n908 & ~n923;
  assign n937 = ~n914 & ~n920;
  assign n938 = ~n936 & ~n937;
  assign n939 = n935 & n938;
  assign n940 = ~n935 & ~n938;
  assign n941 = ~n939 & ~n940;
  assign n942 = ~n931 & n941;
  assign n943 = n931 & ~n941;
  assign n944 = ~n942 & ~n943;
  assign n945 = ~n929 & n944;
  assign n946 = n929 & ~n944;
  assign n947 = ~n945 & ~n946;
  assign n948 = ~n457 & ~n758;
  assign n949 = n762 & n888;
  assign n950 = ~n948 & ~n949;
  assign n951 = ~n451 & n730;
  assign n952 = n733 & n906;
  assign n953 = ~n951 & ~n952;
  assign n954 = ~n469 & n710;
  assign n955 = n715 & n881;
  assign n956 = ~n954 & ~n955;
  assign n957 = ~n953 & n956;
  assign n958 = n953 & ~n956;
  assign n959 = ~n957 & ~n958;
  assign n960 = ~n950 & n959;
  assign n961 = n950 & ~n959;
  assign n962 = ~n960 & ~n961;
  assign n963 = n763 & ~n893;
  assign n964 = ~n884 & ~n890;
  assign n965 = ~n963 & ~n964;
  assign n966 = n962 & ~n965;
  assign n967 = ~n962 & n965;
  assign n968 = ~n966 & ~n967;
  assign n969 = n700 & n918;
  assign n970 = ~n498 & n698;
  assign n971 = ~n969 & ~n970;
  assign n972 = n777 & ~n781;
  assign n973 = ~n542 & ~n972;
  assign n974 = n747 & n912;
  assign n975 = n462 & n742;
  assign n976 = ~n974 & ~n975;
  assign n977 = ~n973 & n976;
  assign n978 = n973 & ~n976;
  assign n979 = ~n977 & ~n978;
  assign n980 = n971 & ~n979;
  assign n981 = ~n971 & n979;
  assign n982 = ~n980 & ~n981;
  assign n983 = n968 & ~n982;
  assign n984 = ~n968 & n982;
  assign n985 = ~n983 & ~n984;
  assign n986 = n947 & ~n985;
  assign n987 = ~n947 & n985;
  assign n988 = ~n986 & ~n987;
  assign n989 = ~n878 & ~n988;
  assign n990 = ~n947 & ~n985;
  assign n991 = ~n989 & ~n990;
  assign n992 = ~n929 & ~n944;
  assign n993 = ~n931 & ~n941;
  assign n994 = ~n992 & ~n993;
  assign n995 = ~n469 & n715;
  assign n996 = g36 & n314;
  assign n997 = ~g36 & ~n314;
  assign n998 = ~n996 & ~n997;
  assign n999 = n710 & n998;
  assign n1000 = ~n995 & ~n999;
  assign n1001 = ~n498 & n700;
  assign n1002 = g38 & ~n198;
  assign n1003 = ~g38 & n198;
  assign n1004 = ~n1002 & ~n1003;
  assign n1005 = n698 & n1004;
  assign n1006 = ~n1001 & ~n1005;
  assign n1007 = n886 & n1006;
  assign n1008 = ~n886 & ~n1006;
  assign n1009 = ~n1007 & ~n1008;
  assign n1010 = n1000 & n1009;
  assign n1011 = ~n1000 & ~n1009;
  assign n1012 = ~n1010 & ~n1011;
  assign n1013 = n935 & ~n938;
  assign n1014 = ~n933 & ~n1013;
  assign n1015 = ~n1012 & n1014;
  assign n1016 = n1012 & ~n1014;
  assign n1017 = ~n1015 & ~n1016;
  assign n1018 = ~n968 & ~n982;
  assign n1019 = ~n962 & ~n965;
  assign n1020 = ~n1018 & ~n1019;
  assign n1021 = n1017 & ~n1020;
  assign n1022 = ~n1017 & n1020;
  assign n1023 = ~n1021 & ~n1022;
  assign n1024 = n462 & n747;
  assign n1025 = ~n404 & n742;
  assign n1026 = ~n1024 & ~n1025;
  assign n1027 = ~n457 & n762;
  assign n1028 = ~g42 & n110;
  assign n1029 = g42 & ~n110;
  assign n1030 = ~n1028 & ~n1029;
  assign n1031 = ~n758 & n1030;
  assign n1032 = ~n1027 & ~n1031;
  assign n1033 = ~n451 & n733;
  assign n1034 = g40 & ~n126;
  assign n1035 = ~g40 & n126;
  assign n1036 = ~n1034 & ~n1035;
  assign n1037 = n730 & n1036;
  assign n1038 = ~n1033 & ~n1037;
  assign n1039 = n1032 & ~n1038;
  assign n1040 = ~n1032 & n1038;
  assign n1041 = ~n1039 & ~n1040;
  assign n1042 = n1026 & ~n1041;
  assign n1043 = ~n1026 & n1041;
  assign n1044 = ~n1042 & ~n1043;
  assign n1045 = ~n950 & ~n959;
  assign n1046 = ~n953 & ~n956;
  assign n1047 = ~n1045 & ~n1046;
  assign n1048 = ~n971 & ~n979;
  assign n1049 = ~n973 & ~n976;
  assign n1050 = ~n1048 & ~n1049;
  assign n1051 = n1047 & ~n1050;
  assign n1052 = ~n1047 & n1050;
  assign n1053 = ~n1051 & ~n1052;
  assign n1054 = ~n1044 & n1053;
  assign n1055 = n1044 & ~n1053;
  assign n1056 = ~n1054 & ~n1055;
  assign n1057 = n1023 & ~n1056;
  assign n1058 = ~n1023 & n1056;
  assign n1059 = ~n1057 & ~n1058;
  assign n1060 = ~n994 & n1059;
  assign n1061 = n994 & ~n1059;
  assign n1062 = ~n1060 & ~n1061;
  assign n1063 = n991 & n1062;
  assign n1064 = n850 & n852;
  assign n1065 = ~n850 & ~n852;
  assign n1066 = ~n1064 & ~n1065;
  assign n1067 = n730 & ~n805;
  assign n1068 = g46 & ~n126;
  assign n1069 = ~g46 & n126;
  assign n1070 = ~n1068 & ~n1069;
  assign n1071 = n733 & n1070;
  assign n1072 = ~n1067 & ~n1071;
  assign n1073 = g44 & ~n198;
  assign n1074 = ~g44 & n198;
  assign n1075 = ~n1073 & ~n1074;
  assign n1076 = n700 & n1075;
  assign n1077 = n698 & ~n847;
  assign n1078 = ~n1076 & ~n1077;
  assign n1079 = ~g40 & n404;
  assign n1080 = g40 & ~n404;
  assign n1081 = ~n1079 & ~n1080;
  assign n1082 = n747 & n1081;
  assign n1083 = n742 & n799;
  assign n1084 = ~n1082 & ~n1083;
  assign n1085 = n1078 & ~n1084;
  assign n1086 = ~n1078 & n1084;
  assign n1087 = ~n1085 & ~n1086;
  assign n1088 = ~n1072 & ~n1087;
  assign n1089 = ~n1078 & ~n1084;
  assign n1090 = ~n1088 & ~n1089;
  assign n1091 = n815 & n817;
  assign n1092 = ~n815 & ~n817;
  assign n1093 = ~n1091 & ~n1092;
  assign n1094 = n1090 & ~n1093;
  assign n1095 = ~n1090 & n1093;
  assign n1096 = ~n1094 & ~n1095;
  assign n1097 = ~n1066 & ~n1096;
  assign n1098 = ~n1090 & ~n1093;
  assign n1099 = ~n1097 & ~n1098;
  assign n1100 = n829 & ~n835;
  assign n1101 = ~n829 & n835;
  assign n1102 = ~n1100 & ~n1101;
  assign n1103 = ~g42 & ~n314;
  assign n1104 = g42 & n314;
  assign n1105 = ~n1103 & ~n1104;
  assign n1106 = n715 & n1105;
  assign n1107 = n710 & ~n839;
  assign n1108 = ~n1106 & ~n1107;
  assign n1109 = g49 & ~n110;
  assign n1110 = ~g38 & n542;
  assign n1111 = g38 & ~n542;
  assign n1112 = ~n1110 & ~n1111;
  assign n1113 = n781 & n1112;
  assign n1114 = ~n777 & n833;
  assign n1115 = ~n1113 & ~n1114;
  assign n1116 = ~n1109 & ~n1115;
  assign n1117 = n1109 & n1115;
  assign n1118 = ~n1116 & ~n1117;
  assign n1119 = ~n1108 & ~n1118;
  assign n1120 = n1109 & ~n1115;
  assign n1121 = ~n1119 & ~n1120;
  assign n1122 = ~n1102 & ~n1121;
  assign n1123 = ~n819 & n857;
  assign n1124 = n819 & ~n857;
  assign n1125 = ~n1123 & ~n1124;
  assign n1126 = ~n1122 & ~n1125;
  assign n1127 = n1122 & n1125;
  assign n1128 = ~n1126 & ~n1127;
  assign n1129 = ~n1099 & ~n1128;
  assign n1130 = n1122 & ~n1125;
  assign n1131 = ~n1129 & ~n1130;
  assign n1132 = n902 & ~n926;
  assign n1133 = ~n902 & n926;
  assign n1134 = ~n1132 & ~n1133;
  assign n1135 = n1131 & ~n1134;
  assign n1136 = ~n1131 & n1134;
  assign n1137 = ~n1135 & ~n1136;
  assign n1138 = ~n796 & n875;
  assign n1139 = n796 & ~n875;
  assign n1140 = ~n1138 & ~n1139;
  assign n1141 = n1137 & ~n1140;
  assign n1142 = ~n1137 & n1140;
  assign n1143 = ~n1141 & ~n1142;
  assign n1144 = ~n726 & n793;
  assign n1145 = n726 & ~n793;
  assign n1146 = ~n1144 & ~n1145;
  assign n1147 = ~g36 & ~n774;
  assign n1148 = g36 & n774;
  assign n1149 = ~n1147 & ~n1148;
  assign n1150 = n823 & n1149;
  assign n1151 = ~n822 & ~n826;
  assign n1152 = ~n1150 & ~n1151;
  assign n1153 = ~g48 & n110;
  assign n1154 = ~n843 & ~n1153;
  assign n1155 = n762 & n1154;
  assign n1156 = ~n758 & ~n812;
  assign n1157 = ~n1155 & ~n1156;
  assign n1158 = ~n1152 & ~n1157;
  assign n1159 = ~g39 & ~n542;
  assign n1160 = g39 & n542;
  assign n1161 = ~n1159 & ~n1160;
  assign n1162 = n781 & ~n1161;
  assign n1163 = ~n777 & n1112;
  assign n1164 = ~n1162 & ~n1163;
  assign n1165 = ~n822 & n1149;
  assign n1166 = g37 & n774;
  assign n1167 = ~g37 & ~n774;
  assign n1168 = ~n1166 & ~n1167;
  assign n1169 = n823 & n1168;
  assign n1170 = ~n1165 & ~n1169;
  assign n1171 = g50 & ~n110;
  assign n1172 = ~n1170 & ~n1171;
  assign n1173 = n1170 & n1171;
  assign n1174 = ~n1172 & ~n1173;
  assign n1175 = ~n1164 & ~n1174;
  assign n1176 = ~n1170 & n1171;
  assign n1177 = ~n1175 & ~n1176;
  assign n1178 = n1152 & ~n1157;
  assign n1179 = ~n1152 & n1157;
  assign n1180 = ~n1178 & ~n1179;
  assign n1181 = ~n1177 & ~n1180;
  assign n1182 = ~n1158 & ~n1181;
  assign n1183 = n1102 & n1121;
  assign n1184 = ~n1122 & ~n1183;
  assign n1185 = ~n1182 & ~n1184;
  assign n1186 = n1182 & n1184;
  assign n1187 = ~n1185 & ~n1186;
  assign n1188 = ~n1108 & n1118;
  assign n1189 = n1108 & ~n1118;
  assign n1190 = ~n1188 & ~n1189;
  assign n1191 = g41 & n404;
  assign n1192 = ~g41 & ~n404;
  assign n1193 = ~n1191 & ~n1192;
  assign n1194 = n747 & ~n1193;
  assign n1195 = n742 & n1081;
  assign n1196 = ~n1194 & ~n1195;
  assign n1197 = g45 & ~n198;
  assign n1198 = ~g45 & n198;
  assign n1199 = ~n1197 & ~n1198;
  assign n1200 = n700 & n1199;
  assign n1201 = n698 & n1075;
  assign n1202 = ~n1200 & ~n1201;
  assign n1203 = g43 & ~n314;
  assign n1204 = ~g43 & n314;
  assign n1205 = ~n1203 & ~n1204;
  assign n1206 = n715 & ~n1205;
  assign n1207 = n710 & n1105;
  assign n1208 = ~n1206 & ~n1207;
  assign n1209 = n1202 & ~n1208;
  assign n1210 = ~n1202 & n1208;
  assign n1211 = ~n1209 & ~n1210;
  assign n1212 = ~n1196 & ~n1211;
  assign n1213 = ~n1202 & ~n1208;
  assign n1214 = ~n1212 & ~n1213;
  assign n1215 = ~n1072 & n1087;
  assign n1216 = n1072 & ~n1087;
  assign n1217 = ~n1215 & ~n1216;
  assign n1218 = ~n1214 & n1217;
  assign n1219 = n1214 & ~n1217;
  assign n1220 = ~n1218 & ~n1219;
  assign n1221 = ~n1190 & ~n1220;
  assign n1222 = ~n1214 & ~n1217;
  assign n1223 = ~n1221 & ~n1222;
  assign n1224 = ~n1187 & ~n1223;
  assign n1225 = ~n1182 & n1184;
  assign n1226 = ~n1224 & ~n1225;
  assign n1227 = n1146 & ~n1226;
  assign n1228 = ~n1146 & n1226;
  assign n1229 = ~n1227 & ~n1228;
  assign n1230 = ~n1099 & n1128;
  assign n1231 = n1099 & ~n1128;
  assign n1232 = ~n1230 & ~n1231;
  assign n1233 = ~n1229 & ~n1232;
  assign n1234 = ~n1146 & ~n1226;
  assign n1235 = ~n1233 & ~n1234;
  assign n1236 = n1143 & n1235;
  assign n1237 = n1229 & ~n1232;
  assign n1238 = ~n1229 & n1232;
  assign n1239 = ~n1237 & ~n1238;
  assign n1240 = n1177 & ~n1180;
  assign n1241 = ~n1177 & n1180;
  assign n1242 = ~n1240 & ~n1241;
  assign n1243 = ~n758 & n1154;
  assign n1244 = ~g49 & ~n110;
  assign n1245 = g49 & n110;
  assign n1246 = ~n1244 & ~n1245;
  assign n1247 = n762 & ~n1246;
  assign n1248 = ~n1243 & ~n1247;
  assign n1249 = ~g47 & ~n126;
  assign n1250 = g47 & n126;
  assign n1251 = ~n1249 & ~n1250;
  assign n1252 = n733 & ~n1251;
  assign n1253 = n730 & n1070;
  assign n1254 = ~n1252 & ~n1253;
  assign n1255 = ~n1248 & ~n1254;
  assign n1256 = ~g50 & n126;
  assign n1257 = ~n133 & ~n1256;
  assign n1258 = g50 & ~n126;
  assign n1259 = ~n1257 & ~n1258;
  assign n1260 = ~n110 & n1259;
  assign n1261 = ~g38 & ~n774;
  assign n1262 = g38 & n774;
  assign n1263 = ~n1261 & ~n1262;
  assign n1264 = n823 & n1263;
  assign n1265 = ~n822 & n1168;
  assign n1266 = ~n1264 & ~n1265;
  assign n1267 = n1260 & ~n1266;
  assign n1268 = ~n1248 & n1254;
  assign n1269 = n1248 & ~n1254;
  assign n1270 = ~n1268 & ~n1269;
  assign n1271 = n1267 & ~n1270;
  assign n1272 = ~n1255 & ~n1271;
  assign n1273 = ~n1242 & n1272;
  assign n1274 = n1242 & ~n1272;
  assign n1275 = ~n1273 & ~n1274;
  assign n1276 = n1164 & ~n1174;
  assign n1277 = ~n1164 & n1174;
  assign n1278 = ~n1276 & ~n1277;
  assign n1279 = ~n758 & ~n1246;
  assign n1280 = ~g50 & n110;
  assign n1281 = ~n1171 & ~n1280;
  assign n1282 = n762 & n1281;
  assign n1283 = ~n1279 & ~n1282;
  assign n1284 = n742 & ~n1193;
  assign n1285 = g42 & ~n404;
  assign n1286 = ~g42 & n404;
  assign n1287 = ~n1285 & ~n1286;
  assign n1288 = n747 & n1287;
  assign n1289 = ~n1284 & ~n1288;
  assign n1290 = g48 & ~n126;
  assign n1291 = ~g48 & n126;
  assign n1292 = ~n1290 & ~n1291;
  assign n1293 = n733 & n1292;
  assign n1294 = n730 & ~n1251;
  assign n1295 = ~n1293 & ~n1294;
  assign n1296 = n1289 & ~n1295;
  assign n1297 = ~n1289 & n1295;
  assign n1298 = ~n1296 & ~n1297;
  assign n1299 = ~n1283 & ~n1298;
  assign n1300 = ~n1289 & ~n1295;
  assign n1301 = ~n1299 & ~n1300;
  assign n1302 = n698 & n1199;
  assign n1303 = ~g46 & n198;
  assign n1304 = g46 & ~n198;
  assign n1305 = ~n1303 & ~n1304;
  assign n1306 = n700 & n1305;
  assign n1307 = ~n1302 & ~n1306;
  assign n1308 = ~n777 & ~n1161;
  assign n1309 = ~g40 & n542;
  assign n1310 = g40 & ~n542;
  assign n1311 = ~n1309 & ~n1310;
  assign n1312 = n781 & n1311;
  assign n1313 = ~n1308 & ~n1312;
  assign n1314 = ~g44 & ~n314;
  assign n1315 = g44 & n314;
  assign n1316 = ~n1314 & ~n1315;
  assign n1317 = n715 & n1316;
  assign n1318 = n710 & ~n1205;
  assign n1319 = ~n1317 & ~n1318;
  assign n1320 = n1313 & ~n1319;
  assign n1321 = ~n1313 & n1319;
  assign n1322 = ~n1320 & ~n1321;
  assign n1323 = ~n1307 & ~n1322;
  assign n1324 = ~n1313 & ~n1319;
  assign n1325 = ~n1323 & ~n1324;
  assign n1326 = n1301 & ~n1325;
  assign n1327 = ~n1301 & n1325;
  assign n1328 = ~n1326 & ~n1327;
  assign n1329 = ~n1278 & ~n1328;
  assign n1330 = ~n1301 & ~n1325;
  assign n1331 = ~n1329 & ~n1330;
  assign n1332 = ~n1275 & ~n1331;
  assign n1333 = ~n1242 & ~n1272;
  assign n1334 = ~n1332 & ~n1333;
  assign n1335 = ~n1187 & n1223;
  assign n1336 = n1187 & ~n1223;
  assign n1337 = ~n1335 & ~n1336;
  assign n1338 = ~n1066 & n1096;
  assign n1339 = n1066 & ~n1096;
  assign n1340 = ~n1338 & ~n1339;
  assign n1341 = n1337 & ~n1340;
  assign n1342 = ~n1337 & n1340;
  assign n1343 = ~n1341 & ~n1342;
  assign n1344 = ~n1334 & ~n1343;
  assign n1345 = ~n1337 & ~n1340;
  assign n1346 = ~n1344 & ~n1345;
  assign n1347 = ~n1239 & ~n1346;
  assign n1348 = ~n1236 & n1347;
  assign n1349 = ~n1143 & ~n1235;
  assign n1350 = ~n1348 & ~n1349;
  assign n1351 = ~n1137 & ~n1140;
  assign n1352 = ~n1131 & ~n1134;
  assign n1353 = ~n1351 & ~n1352;
  assign n1354 = ~n878 & n988;
  assign n1355 = n878 & ~n988;
  assign n1356 = ~n1354 & ~n1355;
  assign n1357 = n1353 & n1356;
  assign n1358 = ~n1350 & ~n1357;
  assign n1359 = ~n1353 & ~n1356;
  assign n1360 = ~n1358 & ~n1359;
  assign n1361 = ~n1063 & ~n1360;
  assign n1362 = ~n1334 & n1343;
  assign n1363 = n1334 & ~n1343;
  assign n1364 = ~n1362 & ~n1363;
  assign n1365 = ~n1275 & n1331;
  assign n1366 = n1275 & ~n1331;
  assign n1367 = ~n1365 & ~n1366;
  assign n1368 = g45 & ~n314;
  assign n1369 = ~g45 & n314;
  assign n1370 = ~n1368 & ~n1369;
  assign n1371 = n715 & ~n1370;
  assign n1372 = n710 & n1316;
  assign n1373 = ~n1371 & ~n1372;
  assign n1374 = g50 & ~n758;
  assign n1375 = g41 & n542;
  assign n1376 = ~g41 & ~n542;
  assign n1377 = ~n1375 & ~n1376;
  assign n1378 = n781 & ~n1377;
  assign n1379 = ~n777 & n1311;
  assign n1380 = ~n1378 & ~n1379;
  assign n1381 = ~n1374 & ~n1380;
  assign n1382 = n1374 & n1380;
  assign n1383 = ~n1381 & ~n1382;
  assign n1384 = ~n1373 & ~n1383;
  assign n1385 = n1374 & ~n1380;
  assign n1386 = ~n1384 & ~n1385;
  assign n1387 = ~n1260 & ~n1266;
  assign n1388 = n1260 & n1266;
  assign n1389 = ~n1387 & ~n1388;
  assign n1390 = n1386 & ~n1389;
  assign n1391 = ~n1386 & n1389;
  assign n1392 = ~n1390 & ~n1391;
  assign n1393 = g49 & ~n126;
  assign n1394 = ~g49 & n126;
  assign n1395 = ~n1393 & ~n1394;
  assign n1396 = n733 & n1395;
  assign n1397 = n730 & n1292;
  assign n1398 = ~n1396 & ~n1397;
  assign n1399 = ~g39 & ~n774;
  assign n1400 = g39 & n774;
  assign n1401 = ~n1399 & ~n1400;
  assign n1402 = n823 & n1401;
  assign n1403 = ~n822 & n1263;
  assign n1404 = ~n1402 & ~n1403;
  assign n1405 = ~g47 & ~n198;
  assign n1406 = g47 & n198;
  assign n1407 = ~n1405 & ~n1406;
  assign n1408 = n700 & ~n1407;
  assign n1409 = n698 & n1305;
  assign n1410 = ~n1408 & ~n1409;
  assign n1411 = ~n1404 & n1410;
  assign n1412 = n1404 & ~n1410;
  assign n1413 = ~n1411 & ~n1412;
  assign n1414 = ~n1398 & ~n1413;
  assign n1415 = ~n1404 & ~n1410;
  assign n1416 = ~n1414 & ~n1415;
  assign n1417 = ~n1392 & ~n1416;
  assign n1418 = ~n1386 & ~n1389;
  assign n1419 = ~n1417 & ~n1418;
  assign n1420 = n1196 & ~n1211;
  assign n1421 = ~n1196 & n1211;
  assign n1422 = ~n1420 & ~n1421;
  assign n1423 = ~n1267 & ~n1270;
  assign n1424 = n1267 & n1270;
  assign n1425 = ~n1423 & ~n1424;
  assign n1426 = ~n1422 & n1425;
  assign n1427 = n1422 & ~n1425;
  assign n1428 = ~n1426 & ~n1427;
  assign n1429 = ~n1419 & ~n1428;
  assign n1430 = ~n1422 & ~n1425;
  assign n1431 = ~n1429 & ~n1430;
  assign n1432 = n1190 & ~n1220;
  assign n1433 = ~n1190 & n1220;
  assign n1434 = ~n1432 & ~n1433;
  assign n1435 = n1431 & ~n1434;
  assign n1436 = ~n1431 & n1434;
  assign n1437 = ~n1435 & ~n1436;
  assign n1438 = ~n1367 & ~n1437;
  assign n1439 = ~n1431 & ~n1434;
  assign n1440 = ~n1438 & ~n1439;
  assign n1441 = n1364 & n1440;
  assign n1442 = ~n1364 & ~n1440;
  assign n1443 = g50 & ~n728;
  assign n1444 = ~n126 & ~n1443;
  assign n1445 = ~n729 & n1444;
  assign n1446 = ~g42 & n542;
  assign n1447 = g42 & ~n542;
  assign n1448 = ~n1446 & ~n1447;
  assign n1449 = n781 & n1448;
  assign n1450 = ~n777 & ~n1377;
  assign n1451 = ~n1449 & ~n1450;
  assign n1452 = n1445 & ~n1451;
  assign n1453 = n742 & n1287;
  assign n1454 = g43 & ~n404;
  assign n1455 = ~g43 & n404;
  assign n1456 = ~n1454 & ~n1455;
  assign n1457 = n747 & n1456;
  assign n1458 = ~n1453 & ~n1457;
  assign n1459 = ~n1452 & ~n1458;
  assign n1460 = n1452 & n1458;
  assign n1461 = ~n1459 & ~n1460;
  assign n1462 = g40 & n774;
  assign n1463 = ~g40 & ~n774;
  assign n1464 = ~n1462 & ~n1463;
  assign n1465 = n823 & n1464;
  assign n1466 = ~n822 & n1401;
  assign n1467 = ~n1465 & ~n1466;
  assign n1468 = g48 & ~n198;
  assign n1469 = ~g48 & n198;
  assign n1470 = ~n1468 & ~n1469;
  assign n1471 = n700 & n1470;
  assign n1472 = n698 & ~n1407;
  assign n1473 = ~n1471 & ~n1472;
  assign n1474 = g46 & n314;
  assign n1475 = ~g46 & ~n314;
  assign n1476 = ~n1474 & ~n1475;
  assign n1477 = n715 & n1476;
  assign n1478 = n710 & ~n1370;
  assign n1479 = ~n1477 & ~n1478;
  assign n1480 = ~n1473 & n1479;
  assign n1481 = n1473 & ~n1479;
  assign n1482 = ~n1480 & ~n1481;
  assign n1483 = ~n1467 & ~n1482;
  assign n1484 = ~n1473 & ~n1479;
  assign n1485 = ~n1483 & ~n1484;
  assign n1486 = ~n1461 & ~n1485;
  assign n1487 = n1452 & ~n1458;
  assign n1488 = ~n1486 & ~n1487;
  assign n1489 = ~n1307 & n1322;
  assign n1490 = n1307 & ~n1322;
  assign n1491 = ~n1489 & ~n1490;
  assign n1492 = ~n1283 & n1298;
  assign n1493 = n1283 & ~n1298;
  assign n1494 = ~n1492 & ~n1493;
  assign n1495 = ~n1491 & n1494;
  assign n1496 = n1491 & ~n1494;
  assign n1497 = ~n1495 & ~n1496;
  assign n1498 = ~n1488 & ~n1497;
  assign n1499 = ~n1491 & ~n1494;
  assign n1500 = ~n1498 & ~n1499;
  assign n1501 = ~n1419 & n1428;
  assign n1502 = n1419 & ~n1428;
  assign n1503 = ~n1501 & ~n1502;
  assign n1504 = n1278 & ~n1328;
  assign n1505 = ~n1278 & n1328;
  assign n1506 = ~n1504 & ~n1505;
  assign n1507 = n1503 & ~n1506;
  assign n1508 = ~n1503 & n1506;
  assign n1509 = ~n1507 & ~n1508;
  assign n1510 = n1500 & ~n1509;
  assign n1511 = ~n1500 & n1509;
  assign n1512 = ~n1510 & ~n1511;
  assign n1513 = n1488 & ~n1497;
  assign n1514 = ~n1488 & n1497;
  assign n1515 = ~n1513 & ~n1514;
  assign n1516 = n1392 & ~n1416;
  assign n1517 = ~n1392 & n1416;
  assign n1518 = ~n1516 & ~n1517;
  assign n1519 = g44 & ~n404;
  assign n1520 = ~g44 & n404;
  assign n1521 = ~n1519 & ~n1520;
  assign n1522 = n747 & n1521;
  assign n1523 = n742 & n1456;
  assign n1524 = ~n1522 & ~n1523;
  assign n1525 = ~n1256 & ~n1258;
  assign n1526 = n733 & n1525;
  assign n1527 = n730 & n1395;
  assign n1528 = ~n1526 & ~n1527;
  assign n1529 = ~n1524 & ~n1528;
  assign n1530 = n1445 & n1451;
  assign n1531 = ~n1445 & ~n1451;
  assign n1532 = ~n1530 & ~n1531;
  assign n1533 = ~n1524 & n1528;
  assign n1534 = n1524 & ~n1528;
  assign n1535 = ~n1533 & ~n1534;
  assign n1536 = ~n1532 & ~n1535;
  assign n1537 = ~n1529 & ~n1536;
  assign n1538 = n1373 & ~n1383;
  assign n1539 = ~n1373 & n1383;
  assign n1540 = ~n1538 & ~n1539;
  assign n1541 = ~n1398 & n1413;
  assign n1542 = n1398 & ~n1413;
  assign n1543 = ~n1541 & ~n1542;
  assign n1544 = ~n1540 & n1543;
  assign n1545 = n1540 & ~n1543;
  assign n1546 = ~n1544 & ~n1545;
  assign n1547 = ~n1537 & ~n1546;
  assign n1548 = ~n1540 & ~n1543;
  assign n1549 = ~n1547 & ~n1548;
  assign n1550 = n1518 & ~n1549;
  assign n1551 = ~n1518 & n1549;
  assign n1552 = ~n1550 & ~n1551;
  assign n1553 = ~n1515 & ~n1552;
  assign n1554 = ~n1518 & ~n1549;
  assign n1555 = ~n1553 & ~n1554;
  assign n1556 = n1512 & n1555;
  assign n1557 = ~g45 & ~n404;
  assign n1558 = g45 & n404;
  assign n1559 = ~n1557 & ~n1558;
  assign n1560 = n742 & ~n1559;
  assign n1561 = g46 & ~n404;
  assign n1562 = ~g46 & n404;
  assign n1563 = ~n1561 & ~n1562;
  assign n1564 = n747 & n1563;
  assign n1565 = ~n1560 & ~n1564;
  assign n1566 = g50 & ~n697;
  assign n1567 = ~n198 & ~n1566;
  assign n1568 = ~n696 & n1567;
  assign n1569 = g44 & ~n542;
  assign n1570 = ~g44 & n542;
  assign n1571 = ~n1569 & ~n1570;
  assign n1572 = n781 & n1571;
  assign n1573 = g43 & n542;
  assign n1574 = ~g43 & ~n542;
  assign n1575 = ~n1573 & ~n1574;
  assign n1576 = ~n777 & ~n1575;
  assign n1577 = ~n1572 & ~n1576;
  assign n1578 = ~n1568 & ~n1577;
  assign n1579 = n1568 & n1577;
  assign n1580 = ~n1578 & ~n1579;
  assign n1581 = n1565 & ~n1580;
  assign n1582 = ~n1565 & n1580;
  assign n1583 = ~n1581 & ~n1582;
  assign n1584 = g50 & n698;
  assign n1585 = g42 & ~n774;
  assign n1586 = ~g42 & n774;
  assign n1587 = ~n1585 & ~n1586;
  assign n1588 = ~n822 & ~n1587;
  assign n1589 = ~g43 & n774;
  assign n1590 = g43 & ~n774;
  assign n1591 = ~n1589 & ~n1590;
  assign n1592 = n823 & ~n1591;
  assign n1593 = ~n1588 & ~n1592;
  assign n1594 = n1584 & n1593;
  assign n1595 = ~n1584 & ~n1593;
  assign n1596 = ~n1594 & ~n1595;
  assign n1597 = ~g48 & n314;
  assign n1598 = g48 & ~n314;
  assign n1599 = ~n1597 & ~n1598;
  assign n1600 = n710 & ~n1599;
  assign n1601 = ~g49 & ~n314;
  assign n1602 = g49 & n314;
  assign n1603 = ~n1601 & ~n1602;
  assign n1604 = n715 & n1603;
  assign n1605 = ~n1600 & ~n1604;
  assign n1606 = ~n1596 & ~n1605;
  assign n1607 = n1584 & ~n1593;
  assign n1608 = ~n1606 & ~n1607;
  assign n1609 = n1583 & ~n1608;
  assign n1610 = ~n1583 & n1608;
  assign n1611 = ~n1609 & ~n1610;
  assign n1612 = n823 & ~n1587;
  assign n1613 = g41 & ~n774;
  assign n1614 = ~g41 & n774;
  assign n1615 = ~n1613 & ~n1614;
  assign n1616 = ~n822 & ~n1615;
  assign n1617 = ~n1612 & ~n1616;
  assign n1618 = n715 & ~n1599;
  assign n1619 = g47 & ~n314;
  assign n1620 = ~g47 & n314;
  assign n1621 = ~n1619 & ~n1620;
  assign n1622 = n710 & ~n1621;
  assign n1623 = ~n1618 & ~n1622;
  assign n1624 = g49 & n198;
  assign n1625 = ~g49 & ~n198;
  assign n1626 = ~n1624 & ~n1625;
  assign n1627 = n698 & ~n1626;
  assign n1628 = ~g50 & n198;
  assign n1629 = g50 & ~n198;
  assign n1630 = ~n1628 & ~n1629;
  assign n1631 = n700 & n1630;
  assign n1632 = ~n1627 & ~n1631;
  assign n1633 = n1623 & ~n1632;
  assign n1634 = ~n1623 & n1632;
  assign n1635 = ~n1633 & ~n1634;
  assign n1636 = ~n1617 & n1635;
  assign n1637 = n1617 & ~n1635;
  assign n1638 = ~n1636 & ~n1637;
  assign n1639 = ~g50 & n404;
  assign n1640 = n308 & ~n1639;
  assign n1641 = g50 & ~n404;
  assign n1642 = n314 & ~n1641;
  assign n1643 = ~n1640 & n1642;
  assign n1644 = ~g44 & ~n774;
  assign n1645 = g44 & n774;
  assign n1646 = ~n1644 & ~n1645;
  assign n1647 = n823 & n1646;
  assign n1648 = ~n822 & ~n1591;
  assign n1649 = ~n1647 & ~n1648;
  assign n1650 = n1643 & ~n1649;
  assign n1651 = g45 & n542;
  assign n1652 = ~g45 & ~n542;
  assign n1653 = ~n1651 & ~n1652;
  assign n1654 = n781 & ~n1653;
  assign n1655 = ~n777 & n1571;
  assign n1656 = ~n1654 & ~n1655;
  assign n1657 = g47 & n404;
  assign n1658 = ~g47 & ~n404;
  assign n1659 = ~n1657 & ~n1658;
  assign n1660 = n747 & ~n1659;
  assign n1661 = n742 & n1563;
  assign n1662 = ~n1660 & ~n1661;
  assign n1663 = ~n1656 & n1662;
  assign n1664 = n1656 & ~n1662;
  assign n1665 = ~n1663 & ~n1664;
  assign n1666 = n1650 & ~n1665;
  assign n1667 = ~n1656 & ~n1662;
  assign n1668 = ~n1666 & ~n1667;
  assign n1669 = ~n1638 & n1668;
  assign n1670 = n1638 & ~n1668;
  assign n1671 = ~n1669 & ~n1670;
  assign n1672 = ~n1611 & ~n1671;
  assign n1673 = ~n1638 & ~n1668;
  assign n1674 = ~n1672 & ~n1673;
  assign n1675 = ~n1623 & ~n1632;
  assign n1676 = ~n1617 & ~n1635;
  assign n1677 = ~n1675 & ~n1676;
  assign n1678 = n1568 & ~n1577;
  assign n1679 = n1677 & n1678;
  assign n1680 = ~n1677 & ~n1678;
  assign n1681 = ~n1679 & ~n1680;
  assign n1682 = n781 & ~n1575;
  assign n1683 = ~n777 & n1448;
  assign n1684 = ~n1682 & ~n1683;
  assign n1685 = g50 & n730;
  assign n1686 = ~n1684 & n1685;
  assign n1687 = n1684 & ~n1685;
  assign n1688 = ~n1686 & ~n1687;
  assign n1689 = n715 & ~n1621;
  assign n1690 = n710 & n1476;
  assign n1691 = ~n1689 & ~n1690;
  assign n1692 = ~n1688 & ~n1691;
  assign n1693 = n1688 & n1691;
  assign n1694 = ~n1692 & ~n1693;
  assign n1695 = n1681 & n1694;
  assign n1696 = ~n1681 & ~n1694;
  assign n1697 = ~n1695 & ~n1696;
  assign n1698 = ~n1583 & ~n1608;
  assign n1699 = ~n1565 & ~n1580;
  assign n1700 = ~n1698 & ~n1699;
  assign n1701 = n823 & ~n1615;
  assign n1702 = ~n822 & n1464;
  assign n1703 = ~n1701 & ~n1702;
  assign n1704 = n700 & ~n1626;
  assign n1705 = n698 & n1470;
  assign n1706 = ~n1704 & ~n1705;
  assign n1707 = n1703 & ~n1706;
  assign n1708 = ~n1703 & n1706;
  assign n1709 = ~n1707 & ~n1708;
  assign n1710 = n747 & ~n1559;
  assign n1711 = n742 & n1521;
  assign n1712 = ~n1710 & ~n1711;
  assign n1713 = n1709 & ~n1712;
  assign n1714 = ~n1709 & n1712;
  assign n1715 = ~n1713 & ~n1714;
  assign n1716 = ~n1700 & n1715;
  assign n1717 = n1700 & ~n1715;
  assign n1718 = ~n1716 & ~n1717;
  assign n1719 = ~n1697 & ~n1718;
  assign n1720 = n1697 & n1718;
  assign n1721 = ~n1719 & ~n1720;
  assign n1722 = ~n1674 & ~n1721;
  assign n1723 = ~n1674 & n1721;
  assign n1724 = n1674 & ~n1721;
  assign n1725 = ~n1723 & ~n1724;
  assign n1726 = n742 & ~n1659;
  assign n1727 = g48 & ~n404;
  assign n1728 = ~g48 & n404;
  assign n1729 = ~n1727 & ~n1728;
  assign n1730 = n747 & n1729;
  assign n1731 = ~n1726 & ~n1730;
  assign n1732 = g46 & n542;
  assign n1733 = ~g46 & ~n542;
  assign n1734 = ~n1732 & ~n1733;
  assign n1735 = n781 & ~n1734;
  assign n1736 = ~n777 & ~n1653;
  assign n1737 = ~n1735 & ~n1736;
  assign n1738 = n710 & n1603;
  assign n1739 = ~g50 & ~n314;
  assign n1740 = g50 & n314;
  assign n1741 = ~n1739 & ~n1740;
  assign n1742 = n715 & n1741;
  assign n1743 = ~n1738 & ~n1742;
  assign n1744 = n1737 & ~n1743;
  assign n1745 = ~n1737 & n1743;
  assign n1746 = ~n1744 & ~n1745;
  assign n1747 = ~n1731 & ~n1746;
  assign n1748 = ~n1737 & ~n1743;
  assign n1749 = ~n1747 & ~n1748;
  assign n1750 = n1596 & ~n1605;
  assign n1751 = ~n1596 & n1605;
  assign n1752 = ~n1750 & ~n1751;
  assign n1753 = n1749 & ~n1752;
  assign n1754 = ~n1749 & n1752;
  assign n1755 = ~n1753 & ~n1754;
  assign n1756 = n1650 & n1665;
  assign n1757 = ~n1650 & ~n1665;
  assign n1758 = ~n1756 & ~n1757;
  assign n1759 = ~n1755 & ~n1758;
  assign n1760 = ~n1749 & ~n1752;
  assign n1761 = ~n1759 & ~n1760;
  assign n1762 = ~n1611 & n1671;
  assign n1763 = n1611 & ~n1671;
  assign n1764 = ~n1762 & ~n1763;
  assign n1765 = ~n1761 & n1764;
  assign n1766 = n1761 & ~n1764;
  assign n1767 = ~n1765 & ~n1766;
  assign n1768 = ~g47 & n542;
  assign n1769 = g47 & ~n542;
  assign n1770 = ~n1768 & ~n1769;
  assign n1771 = n781 & n1770;
  assign n1772 = ~n777 & ~n1734;
  assign n1773 = ~n1771 & ~n1772;
  assign n1774 = ~g45 & n774;
  assign n1775 = g45 & ~n774;
  assign n1776 = ~n1774 & ~n1775;
  assign n1777 = n823 & ~n1776;
  assign n1778 = ~n822 & n1646;
  assign n1779 = ~n1777 & ~n1778;
  assign n1780 = g50 & n710;
  assign n1781 = n1779 & n1780;
  assign n1782 = ~n1779 & ~n1780;
  assign n1783 = ~n1781 & ~n1782;
  assign n1784 = ~n1773 & ~n1783;
  assign n1785 = ~n1779 & n1780;
  assign n1786 = ~n1784 & ~n1785;
  assign n1787 = ~n1643 & ~n1649;
  assign n1788 = n1643 & n1649;
  assign n1789 = ~n1787 & ~n1788;
  assign n1790 = ~n1786 & ~n1789;
  assign n1791 = n1786 & n1789;
  assign n1792 = ~n1790 & ~n1791;
  assign n1793 = ~n1731 & n1746;
  assign n1794 = n1731 & ~n1746;
  assign n1795 = ~n1793 & ~n1794;
  assign n1796 = n1792 & ~n1795;
  assign n1797 = ~n1790 & ~n1796;
  assign n1798 = ~n1755 & n1758;
  assign n1799 = n1755 & ~n1758;
  assign n1800 = ~n1798 & ~n1799;
  assign n1801 = n1797 & n1800;
  assign n1802 = ~g50 & n542;
  assign n1803 = ~n491 & ~n1802;
  assign n1804 = g50 & ~n542;
  assign n1805 = ~n404 & ~n1804;
  assign n1806 = ~n1803 & n1805;
  assign n1807 = ~n822 & ~n1776;
  assign n1808 = ~g46 & ~n774;
  assign n1809 = g46 & n774;
  assign n1810 = ~n1808 & ~n1809;
  assign n1811 = n823 & n1810;
  assign n1812 = ~n1807 & ~n1811;
  assign n1813 = n1806 & ~n1812;
  assign n1814 = g49 & ~n404;
  assign n1815 = ~g49 & n404;
  assign n1816 = ~n1814 & ~n1815;
  assign n1817 = n747 & n1816;
  assign n1818 = n742 & n1729;
  assign n1819 = ~n1817 & ~n1818;
  assign n1820 = ~n1813 & ~n1819;
  assign n1821 = n1813 & n1819;
  assign n1822 = ~n1820 & ~n1821;
  assign n1823 = ~n1773 & n1783;
  assign n1824 = n1773 & ~n1783;
  assign n1825 = ~n1823 & ~n1824;
  assign n1826 = ~n1822 & ~n1825;
  assign n1827 = n1813 & ~n1819;
  assign n1828 = ~n1826 & ~n1827;
  assign n1829 = n1792 & n1795;
  assign n1830 = ~n1792 & ~n1795;
  assign n1831 = ~n1829 & ~n1830;
  assign n1832 = n1828 & n1831;
  assign n1833 = ~n1806 & ~n1812;
  assign n1834 = n1806 & n1812;
  assign n1835 = ~n1833 & ~n1834;
  assign n1836 = g48 & ~n542;
  assign n1837 = ~g48 & n542;
  assign n1838 = ~n1836 & ~n1837;
  assign n1839 = n781 & n1838;
  assign n1840 = ~n777 & n1770;
  assign n1841 = ~n1839 & ~n1840;
  assign n1842 = n742 & n1816;
  assign n1843 = ~n1639 & ~n1641;
  assign n1844 = n747 & n1843;
  assign n1845 = ~n1842 & ~n1844;
  assign n1846 = ~n1841 & n1845;
  assign n1847 = n1841 & ~n1845;
  assign n1848 = ~n1846 & ~n1847;
  assign n1849 = ~n1835 & ~n1848;
  assign n1850 = ~n1841 & ~n1845;
  assign n1851 = ~n1849 & ~n1850;
  assign n1852 = n1822 & ~n1825;
  assign n1853 = ~n1822 & n1825;
  assign n1854 = ~n1852 & ~n1853;
  assign n1855 = n1851 & n1854;
  assign n1856 = ~n822 & n1810;
  assign n1857 = g47 & ~n774;
  assign n1858 = ~g47 & n774;
  assign n1859 = ~n1857 & ~n1858;
  assign n1860 = n823 & ~n1859;
  assign n1861 = ~n1856 & ~n1860;
  assign n1862 = g50 & n742;
  assign n1863 = ~g49 & ~n542;
  assign n1864 = g49 & n542;
  assign n1865 = ~n1863 & ~n1864;
  assign n1866 = n781 & ~n1865;
  assign n1867 = ~n777 & n1838;
  assign n1868 = ~n1866 & ~n1867;
  assign n1869 = n1862 & n1868;
  assign n1870 = ~n1862 & ~n1868;
  assign n1871 = ~n1869 & ~n1870;
  assign n1872 = ~n1861 & ~n1871;
  assign n1873 = n1862 & ~n1868;
  assign n1874 = ~n1872 & ~n1873;
  assign n1875 = ~n1835 & n1848;
  assign n1876 = n1835 & ~n1848;
  assign n1877 = ~n1875 & ~n1876;
  assign n1878 = n1874 & n1877;
  assign n1879 = ~g50 & ~n774;
  assign n1880 = ~n596 & ~n1879;
  assign n1881 = g50 & n774;
  assign n1882 = ~n542 & ~n1881;
  assign n1883 = ~n1880 & n1882;
  assign n1884 = g48 & n774;
  assign n1885 = ~g48 & ~n774;
  assign n1886 = ~n1884 & ~n1885;
  assign n1887 = n823 & n1886;
  assign n1888 = ~n822 & ~n1859;
  assign n1889 = ~n1887 & ~n1888;
  assign n1890 = n1883 & ~n1889;
  assign n1891 = n1861 & ~n1871;
  assign n1892 = ~n1861 & n1871;
  assign n1893 = ~n1891 & ~n1892;
  assign n1894 = ~n1890 & n1893;
  assign n1895 = g50 & ~n822;
  assign n1896 = n774 & ~n1895;
  assign n1897 = ~g50 & n823;
  assign n1898 = ~g49 & n774;
  assign n1899 = g49 & ~n774;
  assign n1900 = ~n1898 & ~n1899;
  assign n1901 = ~n822 & ~n1900;
  assign n1902 = ~n1897 & ~n1901;
  assign n1903 = n1896 & ~n1902;
  assign n1904 = g50 & ~n777;
  assign n1905 = ~n822 & n1886;
  assign n1906 = n823 & ~n1900;
  assign n1907 = ~n1905 & ~n1906;
  assign n1908 = ~n1904 & n1907;
  assign n1909 = n1903 & ~n1908;
  assign n1910 = n1904 & ~n1907;
  assign n1911 = ~n1909 & ~n1910;
  assign n1912 = n781 & ~n1802;
  assign n1913 = ~n1804 & n1912;
  assign n1914 = ~n777 & ~n1865;
  assign n1915 = ~n1913 & ~n1914;
  assign n1916 = ~n1883 & n1889;
  assign n1917 = ~n1890 & ~n1916;
  assign n1918 = n1915 & ~n1917;
  assign n1919 = ~n1911 & ~n1918;
  assign n1920 = ~n1915 & n1917;
  assign n1921 = ~n1919 & ~n1920;
  assign n1922 = ~n1894 & ~n1921;
  assign n1923 = n1890 & ~n1893;
  assign n1924 = ~n1922 & ~n1923;
  assign n1925 = ~n1878 & ~n1924;
  assign n1926 = ~n1874 & ~n1877;
  assign n1927 = ~n1925 & ~n1926;
  assign n1928 = ~n1855 & ~n1927;
  assign n1929 = ~n1851 & ~n1854;
  assign n1930 = ~n1928 & ~n1929;
  assign n1931 = ~n1832 & ~n1930;
  assign n1932 = ~n1828 & ~n1831;
  assign n1933 = ~n1931 & ~n1932;
  assign n1934 = ~n1801 & ~n1933;
  assign n1935 = ~n1797 & ~n1800;
  assign n1936 = ~n1934 & ~n1935;
  assign n1937 = ~n1767 & ~n1936;
  assign n1938 = ~n1761 & ~n1764;
  assign n1939 = ~n1937 & ~n1938;
  assign n1940 = ~n1725 & ~n1939;
  assign n1941 = ~n1722 & ~n1940;
  assign n1942 = ~n1532 & n1535;
  assign n1943 = n1532 & ~n1535;
  assign n1944 = ~n1942 & ~n1943;
  assign n1945 = ~n1467 & n1482;
  assign n1946 = n1467 & ~n1482;
  assign n1947 = ~n1945 & ~n1946;
  assign n1948 = ~n1709 & ~n1712;
  assign n1949 = ~n1703 & ~n1706;
  assign n1950 = ~n1948 & ~n1949;
  assign n1951 = n1688 & ~n1691;
  assign n1952 = ~n1686 & ~n1951;
  assign n1953 = ~n1950 & n1952;
  assign n1954 = n1950 & ~n1952;
  assign n1955 = ~n1953 & ~n1954;
  assign n1956 = ~n1947 & n1955;
  assign n1957 = n1947 & ~n1955;
  assign n1958 = ~n1956 & ~n1957;
  assign n1959 = n1944 & ~n1958;
  assign n1960 = ~n1944 & n1958;
  assign n1961 = ~n1959 & ~n1960;
  assign n1962 = ~n1677 & n1678;
  assign n1963 = ~n1696 & ~n1962;
  assign n1964 = ~n1961 & n1963;
  assign n1965 = n1961 & ~n1963;
  assign n1966 = ~n1964 & ~n1965;
  assign n1967 = n1697 & ~n1718;
  assign n1968 = ~n1700 & ~n1715;
  assign n1969 = ~n1967 & ~n1968;
  assign n1970 = n1966 & ~n1969;
  assign n1971 = ~n1966 & n1969;
  assign n1972 = ~n1970 & ~n1971;
  assign n1973 = ~n1941 & ~n1972;
  assign n1974 = ~n1966 & ~n1969;
  assign n1975 = ~n1973 & ~n1974;
  assign n1976 = ~n1961 & ~n1963;
  assign n1977 = ~n1944 & ~n1958;
  assign n1978 = ~n1976 & ~n1977;
  assign n1979 = ~n1537 & n1546;
  assign n1980 = n1537 & ~n1546;
  assign n1981 = ~n1979 & ~n1980;
  assign n1982 = ~n1947 & ~n1955;
  assign n1983 = ~n1950 & ~n1952;
  assign n1984 = ~n1982 & ~n1983;
  assign n1985 = ~n1461 & n1485;
  assign n1986 = n1461 & ~n1485;
  assign n1987 = ~n1985 & ~n1986;
  assign n1988 = ~n1984 & n1987;
  assign n1989 = n1984 & ~n1987;
  assign n1990 = ~n1988 & ~n1989;
  assign n1991 = ~n1981 & n1990;
  assign n1992 = n1981 & ~n1990;
  assign n1993 = ~n1991 & ~n1992;
  assign n1994 = ~n1978 & n1993;
  assign n1995 = n1978 & ~n1993;
  assign n1996 = ~n1994 & ~n1995;
  assign n1997 = ~n1975 & ~n1996;
  assign n1998 = ~n1978 & ~n1993;
  assign n1999 = ~n1997 & ~n1998;
  assign n2000 = ~n1981 & ~n1990;
  assign n2001 = ~n1984 & ~n1987;
  assign n2002 = ~n2000 & ~n2001;
  assign n2003 = n1515 & ~n1552;
  assign n2004 = ~n1515 & n1552;
  assign n2005 = ~n2003 & ~n2004;
  assign n2006 = ~n2002 & n2005;
  assign n2007 = n2002 & ~n2005;
  assign n2008 = ~n2006 & ~n2007;
  assign n2009 = ~n1999 & ~n2008;
  assign n2010 = ~n2002 & ~n2005;
  assign n2011 = ~n2009 & ~n2010;
  assign n2012 = ~n1556 & ~n2011;
  assign n2013 = ~n1512 & ~n1555;
  assign n2014 = ~n2012 & ~n2013;
  assign n2015 = ~n1367 & n1437;
  assign n2016 = n1367 & ~n1437;
  assign n2017 = ~n2015 & ~n2016;
  assign n2018 = ~n1500 & ~n1509;
  assign n2019 = ~n1503 & ~n1506;
  assign n2020 = ~n2018 & ~n2019;
  assign n2021 = ~n2017 & ~n2020;
  assign n2022 = n2014 & ~n2021;
  assign n2023 = n2017 & n2020;
  assign n2024 = ~n2022 & ~n2023;
  assign n2025 = ~n1442 & ~n2024;
  assign n2026 = ~n1063 & ~n2025;
  assign n2027 = ~n1441 & n2026;
  assign n2028 = n1239 & n1346;
  assign n2029 = ~n1236 & ~n2028;
  assign n2030 = ~n1357 & n2029;
  assign n2031 = n2027 & n2030;
  assign n2032 = ~n991 & ~n1062;
  assign n2033 = ~n2031 & ~n2032;
  assign n2034 = ~n1361 & n2033;
  assign n2035 = n656 & n664;
  assign n2036 = ~n665 & ~n2035;
  assign n2037 = ~n546 & ~n577;
  assign n2038 = n546 & n577;
  assign n2039 = ~n2037 & ~n2038;
  assign n2040 = ~n262 & n587;
  assign n2041 = g41 & n194;
  assign n2042 = ~g41 & ~n194;
  assign n2043 = ~n2041 & ~n2042;
  assign n2044 = n266 & ~n2043;
  assign n2045 = ~n2040 & ~n2044;
  assign n2046 = ~g47 & g48;
  assign n2047 = g47 & ~g48;
  assign n2048 = ~n2046 & ~n2047;
  assign n2049 = ~g48 & g49;
  assign n2050 = g48 & ~g49;
  assign n2051 = ~n2049 & ~n2050;
  assign n2052 = n2048 & n2051;
  assign n2053 = g47 & ~n2052;
  assign n2054 = ~n529 & ~n536;
  assign n2055 = g45 & ~n133;
  assign n2056 = ~g45 & n133;
  assign n2057 = ~n2055 & ~n2056;
  assign n2058 = n533 & n2057;
  assign n2059 = ~n2054 & ~n2058;
  assign n2060 = n2053 & ~n2059;
  assign n2061 = ~n2053 & n2059;
  assign n2062 = ~n2060 & ~n2061;
  assign n2063 = ~n2045 & ~n2062;
  assign n2064 = ~n2053 & ~n2059;
  assign n2065 = ~n2063 & ~n2064;
  assign n2066 = ~n539 & ~n2065;
  assign n2067 = n539 & n2065;
  assign n2068 = ~n2066 & ~n2067;
  assign n2069 = ~n370 & ~n558;
  assign n2070 = g43 & ~n141;
  assign n2071 = ~g43 & n141;
  assign n2072 = ~n2070 & ~n2071;
  assign n2073 = n374 & ~n2072;
  assign n2074 = ~n2069 & ~n2073;
  assign n2075 = g35 & n774;
  assign n2076 = ~n175 & ~n569;
  assign n2077 = ~g39 & n308;
  assign n2078 = g39 & ~n308;
  assign n2079 = ~n2077 & ~n2078;
  assign n2080 = n176 & ~n2079;
  assign n2081 = ~n2076 & ~n2080;
  assign n2082 = ~n2075 & ~n2081;
  assign n2083 = n2075 & n2081;
  assign n2084 = ~n2082 & ~n2083;
  assign n2085 = ~n2074 & ~n2084;
  assign n2086 = n2075 & ~n2081;
  assign n2087 = ~n2085 & ~n2086;
  assign n2088 = ~n2068 & ~n2087;
  assign n2089 = n539 & ~n2065;
  assign n2090 = ~n2088 & ~n2089;
  assign n2091 = ~n2039 & ~n2090;
  assign n2092 = n593 & ~n609;
  assign n2093 = ~n593 & n609;
  assign n2094 = ~n2092 & ~n2093;
  assign n2095 = ~n2048 & n2051;
  assign n2096 = ~n812 & n2095;
  assign n2097 = g47 & ~n2051;
  assign n2098 = ~n2096 & ~n2097;
  assign n2099 = ~g35 & ~n596;
  assign n2100 = g35 & n596;
  assign n2101 = ~n2099 & ~n2100;
  assign n2102 = n123 & ~n2101;
  assign n2103 = ~n119 & ~n604;
  assign n2104 = ~n2102 & ~n2103;
  assign n2105 = ~n2098 & ~n2104;
  assign n2106 = n2098 & n2104;
  assign n2107 = g37 & ~n491;
  assign n2108 = ~g37 & n491;
  assign n2109 = ~n2107 & ~n2108;
  assign n2110 = n107 & n2109;
  assign n2111 = ~n103 & n549;
  assign n2112 = ~n2110 & ~n2111;
  assign n2113 = ~n2106 & ~n2112;
  assign n2114 = ~n2105 & ~n2113;
  assign n2115 = ~n2094 & ~n2114;
  assign n2116 = ~n565 & ~n566;
  assign n2117 = n575 & n2116;
  assign n2118 = ~n575 & ~n2116;
  assign n2119 = ~n2117 & ~n2118;
  assign n2120 = n2094 & n2114;
  assign n2121 = ~n2115 & ~n2120;
  assign n2122 = ~n2119 & n2121;
  assign n2123 = ~n2115 & ~n2122;
  assign n2124 = n2039 & n2090;
  assign n2125 = ~n2091 & ~n2124;
  assign n2126 = ~n2123 & n2125;
  assign n2127 = ~n2091 & ~n2126;
  assign n2128 = n2036 & n2127;
  assign n2129 = ~n2036 & ~n2127;
  assign n2130 = ~n2128 & ~n2129;
  assign n2131 = n584 & ~n647;
  assign n2132 = ~n584 & n647;
  assign n2133 = ~n2131 & ~n2132;
  assign n2134 = n2130 & ~n2133;
  assign n2135 = ~n2130 & n2133;
  assign n2136 = ~n2134 & ~n2135;
  assign n2137 = n629 & ~n644;
  assign n2138 = ~n629 & n644;
  assign n2139 = ~n2137 & ~n2138;
  assign n2140 = n2123 & n2125;
  assign n2141 = ~n2123 & ~n2125;
  assign n2142 = ~n2140 & ~n2141;
  assign n2143 = n2139 & ~n2142;
  assign n2144 = ~n2139 & n2142;
  assign n2145 = ~n2143 & ~n2144;
  assign n2146 = n2119 & n2121;
  assign n2147 = ~n2119 & ~n2121;
  assign n2148 = ~n2146 & ~n2147;
  assign n2149 = ~n2068 & n2087;
  assign n2150 = n2068 & ~n2087;
  assign n2151 = ~n2149 & ~n2150;
  assign n2152 = g35 & ~n822;
  assign n2153 = n533 & ~n805;
  assign n2154 = ~n529 & n2057;
  assign n2155 = ~n2153 & ~n2154;
  assign n2156 = n2152 & ~n2155;
  assign n2157 = ~n2152 & n2155;
  assign n2158 = n266 & ~n839;
  assign n2159 = ~n262 & ~n2043;
  assign n2160 = ~n2158 & ~n2159;
  assign n2161 = ~n2157 & ~n2160;
  assign n2162 = ~n2156 & ~n2161;
  assign n2163 = n2045 & n2062;
  assign n2164 = ~n2063 & ~n2163;
  assign n2165 = ~n2162 & n2164;
  assign n2166 = n176 & n799;
  assign n2167 = ~n175 & ~n2079;
  assign n2168 = ~n2166 & ~n2167;
  assign n2169 = ~n103 & n2109;
  assign n2170 = n107 & n833;
  assign n2171 = ~n2169 & ~n2170;
  assign n2172 = ~n2168 & ~n2171;
  assign n2173 = n374 & ~n847;
  assign n2174 = ~n370 & ~n2072;
  assign n2175 = ~n2173 & ~n2174;
  assign n2176 = n2168 & n2171;
  assign n2177 = ~n2172 & ~n2176;
  assign n2178 = ~n2175 & n2177;
  assign n2179 = ~n2172 & ~n2178;
  assign n2180 = n2162 & ~n2164;
  assign n2181 = ~n2165 & ~n2180;
  assign n2182 = ~n2179 & n2181;
  assign n2183 = ~n2165 & ~n2182;
  assign n2184 = n2151 & ~n2183;
  assign n2185 = ~n2151 & n2183;
  assign n2186 = ~n2184 & ~n2185;
  assign n2187 = ~n2148 & ~n2186;
  assign n2188 = ~n2151 & ~n2183;
  assign n2189 = ~n2187 & ~n2188;
  assign n2190 = ~n2145 & ~n2189;
  assign n2191 = ~n2139 & ~n2142;
  assign n2192 = ~n2190 & ~n2191;
  assign n2193 = ~n2136 & ~n2192;
  assign n2194 = ~n2148 & n2186;
  assign n2195 = n2148 & ~n2186;
  assign n2196 = ~n2194 & ~n2195;
  assign n2197 = n2104 & ~n2112;
  assign n2198 = ~n2104 & n2112;
  assign n2199 = ~n2197 & ~n2198;
  assign n2200 = n2098 & n2199;
  assign n2201 = ~n2098 & ~n2199;
  assign n2202 = ~n2200 & ~n2201;
  assign n2203 = ~n370 & ~n847;
  assign n2204 = g43 & n194;
  assign n2205 = ~g43 & ~n194;
  assign n2206 = ~n2204 & ~n2205;
  assign n2207 = n374 & ~n2206;
  assign n2208 = ~n2203 & ~n2207;
  assign n2209 = ~n119 & ~n2101;
  assign n2210 = n123 & ~n826;
  assign n2211 = ~n2209 & ~n2210;
  assign n2212 = n2098 & n2211;
  assign n2213 = ~n2098 & ~n2211;
  assign n2214 = ~n2212 & ~n2213;
  assign n2215 = ~n2208 & ~n2214;
  assign n2216 = n2098 & ~n2211;
  assign n2217 = ~n2215 & ~n2216;
  assign n2218 = n2074 & ~n2084;
  assign n2219 = ~n2074 & n2084;
  assign n2220 = ~n2218 & ~n2219;
  assign n2221 = n2217 & ~n2220;
  assign n2222 = ~n2217 & n2220;
  assign n2223 = ~n2221 & ~n2222;
  assign n2224 = n2202 & ~n2223;
  assign n2225 = ~n2217 & ~n2220;
  assign n2226 = ~n2224 & ~n2225;
  assign n2227 = ~n2152 & ~n2155;
  assign n2228 = n2152 & n2155;
  assign n2229 = ~n2227 & ~n2228;
  assign n2230 = ~n2160 & n2229;
  assign n2231 = n2160 & ~n2229;
  assign n2232 = ~n2230 & ~n2231;
  assign n2233 = n2208 & ~n2214;
  assign n2234 = ~n2208 & n2214;
  assign n2235 = ~n2233 & ~n2234;
  assign n2236 = ~n2232 & ~n2235;
  assign n2237 = n2232 & n2235;
  assign n2238 = ~n2236 & ~n2237;
  assign n2239 = n266 & ~n1193;
  assign n2240 = ~g41 & n308;
  assign n2241 = g41 & ~n308;
  assign n2242 = ~n2240 & ~n2241;
  assign n2243 = ~n262 & ~n2242;
  assign n2244 = ~n2239 & ~n2243;
  assign n2245 = n374 & ~n1205;
  assign n2246 = ~n370 & ~n2206;
  assign n2247 = ~n2245 & ~n2246;
  assign n2248 = n2244 & ~n2247;
  assign n2249 = ~n2244 & n2247;
  assign n2250 = ~n2248 & ~n2249;
  assign n2251 = g35 & n822;
  assign n2252 = ~g35 & ~n822;
  assign n2253 = ~n2251 & ~n2252;
  assign n2254 = ~n119 & ~n2253;
  assign n2255 = g17 & g2;
  assign n2256 = ~g2 & g33;
  assign n2257 = ~n2255 & ~n2256;
  assign n2258 = ~g35 & n2257;
  assign n2259 = g35 & ~n2257;
  assign n2260 = ~n2258 & ~n2259;
  assign n2261 = n123 & n2260;
  assign n2262 = ~n2254 & ~n2261;
  assign n2263 = ~n2250 & ~n2262;
  assign n2264 = ~n2244 & ~n2247;
  assign n2265 = ~n2263 & ~n2264;
  assign n2266 = n107 & n1168;
  assign n2267 = ~g37 & n596;
  assign n2268 = g37 & ~n596;
  assign n2269 = ~n2267 & ~n2268;
  assign n2270 = ~n103 & n2269;
  assign n2271 = ~n2266 & ~n2270;
  assign n2272 = n533 & n1199;
  assign n2273 = ~g45 & n141;
  assign n2274 = g45 & ~n141;
  assign n2275 = ~n2273 & ~n2274;
  assign n2276 = ~n529 & ~n2275;
  assign n2277 = ~n2272 & ~n2276;
  assign n2278 = ~n2271 & ~n2277;
  assign n2279 = n176 & ~n1161;
  assign n2280 = g39 & n491;
  assign n2281 = ~g39 & ~n491;
  assign n2282 = ~n2280 & ~n2281;
  assign n2283 = ~n175 & ~n2282;
  assign n2284 = ~n2279 & ~n2283;
  assign n2285 = n2271 & n2277;
  assign n2286 = ~n2278 & ~n2285;
  assign n2287 = ~n2284 & n2286;
  assign n2288 = ~n2278 & ~n2287;
  assign n2289 = ~n1251 & n2095;
  assign n2290 = ~g47 & ~n133;
  assign n2291 = g47 & n133;
  assign n2292 = ~n2290 & ~n2291;
  assign n2293 = ~n2051 & ~n2292;
  assign n2294 = ~n2289 & ~n2293;
  assign n2295 = g49 & ~g50;
  assign n2296 = ~n1246 & n2295;
  assign n2297 = g49 & g50;
  assign n2298 = ~n2296 & ~n2297;
  assign n2299 = ~g2 & g34;
  assign n2300 = ~g18 & g34;
  assign n2301 = g2 & ~n2300;
  assign n2302 = ~n2299 & ~n2301;
  assign n2303 = g35 & ~n2302;
  assign n2304 = ~n2298 & ~n2303;
  assign n2305 = n2298 & n2303;
  assign n2306 = ~n2304 & ~n2305;
  assign n2307 = ~n2294 & ~n2306;
  assign n2308 = ~n2298 & n2303;
  assign n2309 = ~n2307 & ~n2308;
  assign n2310 = ~n2288 & n2309;
  assign n2311 = n2288 & ~n2309;
  assign n2312 = ~n2310 & ~n2311;
  assign n2313 = ~n2265 & ~n2312;
  assign n2314 = ~n2288 & ~n2309;
  assign n2315 = ~n2313 & ~n2314;
  assign n2316 = n2238 & ~n2315;
  assign n2317 = ~n2236 & ~n2316;
  assign n2318 = ~n262 & ~n839;
  assign n2319 = n266 & ~n2242;
  assign n2320 = ~n2318 & ~n2319;
  assign n2321 = ~n529 & ~n805;
  assign n2322 = n533 & ~n2275;
  assign n2323 = ~n2321 & ~n2322;
  assign n2324 = ~n2320 & ~n2323;
  assign n2325 = n2320 & n2323;
  assign n2326 = n2095 & ~n2292;
  assign n2327 = ~n812 & ~n2051;
  assign n2328 = ~n2326 & ~n2327;
  assign n2329 = ~n2325 & ~n2328;
  assign n2330 = ~n2324 & ~n2329;
  assign n2331 = g49 & ~n2259;
  assign n2332 = ~n119 & ~n826;
  assign n2333 = n123 & ~n2253;
  assign n2334 = ~n2332 & ~n2333;
  assign n2335 = ~n2331 & ~n2334;
  assign n2336 = ~g49 & n2259;
  assign n2337 = ~n2335 & ~n2336;
  assign n2338 = ~n2330 & ~n2337;
  assign n2339 = n2330 & n2337;
  assign n2340 = ~n2338 & ~n2339;
  assign n2341 = ~n2175 & ~n2177;
  assign n2342 = n2175 & n2177;
  assign n2343 = ~n2341 & ~n2342;
  assign n2344 = n2340 & ~n2343;
  assign n2345 = ~n2338 & ~n2344;
  assign n2346 = ~n2179 & ~n2181;
  assign n2347 = n2179 & n2181;
  assign n2348 = ~n2346 & ~n2347;
  assign n2349 = n2345 & ~n2348;
  assign n2350 = ~n2345 & n2348;
  assign n2351 = ~n2349 & ~n2350;
  assign n2352 = ~n2317 & ~n2351;
  assign n2353 = ~n2345 & ~n2348;
  assign n2354 = ~n2352 & ~n2353;
  assign n2355 = ~n2226 & n2354;
  assign n2356 = n2226 & ~n2354;
  assign n2357 = ~n2355 & ~n2356;
  assign n2358 = n2196 & ~n2357;
  assign n2359 = ~n2196 & n2357;
  assign n2360 = ~n2358 & ~n2359;
  assign n2361 = ~n2202 & ~n2223;
  assign n2362 = n2202 & n2223;
  assign n2363 = ~n2361 & ~n2362;
  assign n2364 = ~g45 & ~n194;
  assign n2365 = g45 & n194;
  assign n2366 = ~n2364 & ~n2365;
  assign n2367 = n533 & ~n2366;
  assign n2368 = ~n529 & n1199;
  assign n2369 = ~n2367 & ~n2368;
  assign n2370 = g39 & n596;
  assign n2371 = ~g39 & ~n596;
  assign n2372 = ~n2370 & ~n2371;
  assign n2373 = n176 & ~n2372;
  assign n2374 = ~n175 & ~n1161;
  assign n2375 = ~n2373 & ~n2374;
  assign n2376 = ~n262 & ~n1193;
  assign n2377 = ~g41 & n491;
  assign n2378 = g41 & ~n491;
  assign n2379 = ~n2377 & ~n2378;
  assign n2380 = n266 & n2379;
  assign n2381 = ~n2376 & ~n2380;
  assign n2382 = n2375 & ~n2381;
  assign n2383 = ~n2375 & n2381;
  assign n2384 = ~n2382 & ~n2383;
  assign n2385 = ~n2369 & ~n2384;
  assign n2386 = ~n2375 & ~n2381;
  assign n2387 = ~n2385 & ~n2386;
  assign n2388 = g50 & ~n1246;
  assign n2389 = ~g49 & n133;
  assign n2390 = g49 & ~n133;
  assign n2391 = ~n2389 & ~n2390;
  assign n2392 = n2295 & n2391;
  assign n2393 = ~n2388 & ~n2392;
  assign n2394 = ~g36 & ~g37;
  assign n2395 = ~n2302 & ~n2394;
  assign n2396 = g36 & g37;
  assign n2397 = g35 & ~n2396;
  assign n2398 = ~n2395 & n2397;
  assign n2399 = ~n2393 & n2398;
  assign n2400 = ~g43 & ~n308;
  assign n2401 = g43 & n308;
  assign n2402 = ~n2400 & ~n2401;
  assign n2403 = n374 & n2402;
  assign n2404 = ~n370 & ~n1205;
  assign n2405 = ~n2403 & ~n2404;
  assign n2406 = g35 & n2302;
  assign n2407 = ~g35 & ~n2302;
  assign n2408 = ~n2406 & ~n2407;
  assign n2409 = n123 & ~n2408;
  assign n2410 = ~n119 & n2260;
  assign n2411 = ~n2409 & ~n2410;
  assign n2412 = ~n2405 & ~n2411;
  assign n2413 = n2405 & n2411;
  assign n2414 = ~n1251 & ~n2051;
  assign n2415 = ~g47 & n141;
  assign n2416 = g47 & ~n141;
  assign n2417 = ~n2415 & ~n2416;
  assign n2418 = n2095 & ~n2417;
  assign n2419 = ~n2414 & ~n2418;
  assign n2420 = ~n2413 & ~n2419;
  assign n2421 = ~n2412 & ~n2420;
  assign n2422 = n2399 & n2421;
  assign n2423 = ~n2399 & ~n2421;
  assign n2424 = ~n2422 & ~n2423;
  assign n2425 = ~n2387 & ~n2424;
  assign n2426 = n2399 & ~n2421;
  assign n2427 = ~n2425 & ~n2426;
  assign n2428 = ~n2331 & ~n2336;
  assign n2429 = n2334 & ~n2428;
  assign n2430 = ~n2334 & n2428;
  assign n2431 = ~n2429 & ~n2430;
  assign n2432 = ~n2320 & n2328;
  assign n2433 = n2320 & ~n2328;
  assign n2434 = ~n2432 & ~n2433;
  assign n2435 = ~n2323 & ~n2434;
  assign n2436 = n2323 & n2434;
  assign n2437 = ~n2435 & ~n2436;
  assign n2438 = ~n2431 & n2437;
  assign n2439 = n2431 & ~n2437;
  assign n2440 = ~n2438 & ~n2439;
  assign n2441 = ~n2427 & ~n2440;
  assign n2442 = n2431 & n2437;
  assign n2443 = ~n2441 & ~n2442;
  assign n2444 = n176 & ~n2282;
  assign n2445 = ~n175 & n799;
  assign n2446 = ~n2444 & ~n2445;
  assign n2447 = ~n103 & n833;
  assign n2448 = n107 & n2269;
  assign n2449 = ~n2447 & ~n2448;
  assign n2450 = n2446 & ~n2449;
  assign n2451 = ~n2446 & n2449;
  assign n2452 = ~n2450 & ~n2451;
  assign n2453 = n2208 & ~n2452;
  assign n2454 = ~n2446 & ~n2449;
  assign n2455 = ~n2453 & ~n2454;
  assign n2456 = ~n2340 & ~n2343;
  assign n2457 = n2340 & n2343;
  assign n2458 = ~n2456 & ~n2457;
  assign n2459 = n2455 & ~n2458;
  assign n2460 = ~n2455 & n2458;
  assign n2461 = ~n2459 & ~n2460;
  assign n2462 = ~n2443 & ~n2461;
  assign n2463 = ~n2455 & ~n2458;
  assign n2464 = ~n2462 & ~n2463;
  assign n2465 = ~n2363 & ~n2464;
  assign n2466 = ~n2317 & n2351;
  assign n2467 = n2317 & ~n2351;
  assign n2468 = ~n2466 & ~n2467;
  assign n2469 = n2363 & n2464;
  assign n2470 = ~n2465 & ~n2469;
  assign n2471 = ~n2468 & n2470;
  assign n2472 = ~n2465 & ~n2471;
  assign n2473 = ~n2360 & ~n2472;
  assign n2474 = n2145 & ~n2189;
  assign n2475 = ~n2145 & n2189;
  assign n2476 = ~n2474 & ~n2475;
  assign n2477 = ~n2196 & ~n2357;
  assign n2478 = ~n2226 & ~n2354;
  assign n2479 = ~n2477 & ~n2478;
  assign n2480 = n2476 & n2479;
  assign n2481 = n2473 & ~n2480;
  assign n2482 = ~n2476 & ~n2479;
  assign n2483 = ~n2481 & ~n2482;
  assign n2484 = n2136 & n2192;
  assign n2485 = ~n2483 & ~n2484;
  assign n2486 = ~n2443 & n2461;
  assign n2487 = n2443 & ~n2461;
  assign n2488 = ~n2486 & ~n2487;
  assign n2489 = ~n2238 & n2315;
  assign n2490 = ~n2316 & ~n2489;
  assign n2491 = ~n2208 & n2452;
  assign n2492 = ~n2453 & ~n2491;
  assign n2493 = n2250 & n2262;
  assign n2494 = ~n2263 & ~n2493;
  assign n2495 = n2284 & ~n2286;
  assign n2496 = ~n2287 & ~n2495;
  assign n2497 = n2294 & ~n2306;
  assign n2498 = ~n2294 & n2306;
  assign n2499 = ~n2497 & ~n2498;
  assign n2500 = ~n2496 & n2499;
  assign n2501 = n2494 & ~n2500;
  assign n2502 = n2496 & ~n2499;
  assign n2503 = ~n2501 & ~n2502;
  assign n2504 = n2492 & ~n2503;
  assign n2505 = n2265 & n2312;
  assign n2506 = ~n2313 & ~n2505;
  assign n2507 = ~n2492 & n2503;
  assign n2508 = ~n2504 & ~n2507;
  assign n2509 = n2506 & n2508;
  assign n2510 = ~n2504 & ~n2509;
  assign n2511 = n2490 & n2510;
  assign n2512 = ~n2490 & ~n2510;
  assign n2513 = ~n2511 & ~n2512;
  assign n2514 = ~n2488 & ~n2513;
  assign n2515 = n2490 & ~n2510;
  assign n2516 = ~n2514 & ~n2515;
  assign n2517 = ~n2468 & ~n2470;
  assign n2518 = n2468 & n2470;
  assign n2519 = ~n2517 & ~n2518;
  assign n2520 = n2516 & n2519;
  assign n2521 = n2427 & n2440;
  assign n2522 = ~n2441 & ~n2521;
  assign n2523 = n2506 & ~n2508;
  assign n2524 = ~n2506 & n2508;
  assign n2525 = ~n2523 & ~n2524;
  assign n2526 = n2522 & ~n2525;
  assign n2527 = ~n2412 & ~n2413;
  assign n2528 = ~n2419 & n2527;
  assign n2529 = n2419 & ~n2527;
  assign n2530 = ~n2528 & ~n2529;
  assign n2531 = n266 & ~n1377;
  assign n2532 = ~n262 & n2379;
  assign n2533 = ~n2531 & ~n2532;
  assign n2534 = n374 & n1456;
  assign n2535 = ~n370 & n2402;
  assign n2536 = ~n2534 & ~n2535;
  assign n2537 = ~n2533 & ~n2536;
  assign n2538 = n2533 & n2536;
  assign n2539 = ~n529 & ~n2366;
  assign n2540 = n533 & ~n1370;
  assign n2541 = ~n2539 & ~n2540;
  assign n2542 = ~n2538 & ~n2541;
  assign n2543 = ~n2537 & ~n2542;
  assign n2544 = n2369 & ~n2384;
  assign n2545 = ~n2369 & n2384;
  assign n2546 = ~n2544 & ~n2545;
  assign n2547 = ~n2543 & n2546;
  assign n2548 = n2543 & ~n2546;
  assign n2549 = ~n2547 & ~n2548;
  assign n2550 = n2530 & ~n2549;
  assign n2551 = ~n2543 & ~n2546;
  assign n2552 = ~n2550 & ~n2551;
  assign n2553 = ~n1407 & n2095;
  assign n2554 = ~n2051 & ~n2417;
  assign n2555 = ~n2553 & ~n2554;
  assign n2556 = ~n119 & ~n2302;
  assign n2557 = n1395 & n2295;
  assign n2558 = g50 & n2391;
  assign n2559 = ~n2557 & ~n2558;
  assign n2560 = n2556 & n2559;
  assign n2561 = ~n2556 & ~n2559;
  assign n2562 = ~n2560 & ~n2561;
  assign n2563 = ~n2555 & ~n2562;
  assign n2564 = n2556 & ~n2559;
  assign n2565 = ~n2563 & ~n2564;
  assign n2566 = n2393 & n2398;
  assign n2567 = ~n2393 & ~n2398;
  assign n2568 = ~n2566 & ~n2567;
  assign n2569 = ~n103 & n1168;
  assign n2570 = g37 & n822;
  assign n2571 = ~g37 & ~n822;
  assign n2572 = ~n2570 & ~n2571;
  assign n2573 = n107 & ~n2572;
  assign n2574 = ~n2569 & ~n2573;
  assign n2575 = n2568 & ~n2574;
  assign n2576 = ~n2568 & n2574;
  assign n2577 = ~n2575 & ~n2576;
  assign n2578 = ~n2565 & ~n2577;
  assign n2579 = ~n2568 & ~n2574;
  assign n2580 = ~n2578 & ~n2579;
  assign n2581 = n2387 & ~n2424;
  assign n2582 = ~n2387 & n2424;
  assign n2583 = ~n2581 & ~n2582;
  assign n2584 = n2580 & ~n2583;
  assign n2585 = ~n2580 & n2583;
  assign n2586 = ~n2584 & ~n2585;
  assign n2587 = ~n2552 & ~n2586;
  assign n2588 = ~n2580 & ~n2583;
  assign n2589 = ~n2587 & ~n2588;
  assign n2590 = ~n2522 & n2525;
  assign n2591 = ~n2526 & ~n2590;
  assign n2592 = ~n2589 & n2591;
  assign n2593 = ~n2526 & ~n2592;
  assign n2594 = n2488 & ~n2513;
  assign n2595 = ~n2488 & n2513;
  assign n2596 = ~n2594 & ~n2595;
  assign n2597 = ~n2593 & ~n2596;
  assign n2598 = ~n2520 & n2597;
  assign n2599 = n2555 & n2562;
  assign n2600 = ~n2563 & ~n2599;
  assign n2601 = ~n175 & n1401;
  assign n2602 = g39 & n822;
  assign n2603 = ~g39 & ~n822;
  assign n2604 = ~n2602 & ~n2603;
  assign n2605 = n176 & ~n2604;
  assign n2606 = ~n2601 & ~n2605;
  assign n2607 = ~n529 & ~n1370;
  assign n2608 = g45 & ~n308;
  assign n2609 = ~g45 & n308;
  assign n2610 = ~n2608 & ~n2609;
  assign n2611 = n533 & ~n2610;
  assign n2612 = ~n2607 & ~n2611;
  assign n2613 = n2606 & n2612;
  assign n2614 = ~n2606 & ~n2612;
  assign n2615 = g37 & n2302;
  assign n2616 = ~g37 & ~n2302;
  assign n2617 = ~n2615 & ~n2616;
  assign n2618 = n107 & ~n2617;
  assign n2619 = g37 & ~n2257;
  assign n2620 = ~g37 & n2257;
  assign n2621 = ~n2619 & ~n2620;
  assign n2622 = ~n103 & n2621;
  assign n2623 = ~n2618 & ~n2622;
  assign n2624 = ~n2614 & n2623;
  assign n2625 = ~n2613 & ~n2624;
  assign n2626 = ~n2600 & n2625;
  assign n2627 = n2600 & ~n2625;
  assign n2628 = ~n2626 & ~n2627;
  assign n2629 = ~n370 & n1456;
  assign n2630 = ~g43 & n491;
  assign n2631 = g43 & ~n491;
  assign n2632 = ~n2630 & ~n2631;
  assign n2633 = n374 & n2632;
  assign n2634 = ~n2629 & ~n2633;
  assign n2635 = ~n262 & ~n1377;
  assign n2636 = ~g41 & n596;
  assign n2637 = g41 & ~n596;
  assign n2638 = ~n2636 & ~n2637;
  assign n2639 = n266 & n2638;
  assign n2640 = ~n2635 & ~n2639;
  assign n2641 = n2634 & ~n2640;
  assign n2642 = ~n2634 & n2640;
  assign n2643 = ~n2641 & ~n2642;
  assign n2644 = ~n1407 & ~n2051;
  assign n2645 = g47 & n194;
  assign n2646 = ~g47 & ~n194;
  assign n2647 = ~n2645 & ~n2646;
  assign n2648 = n2095 & ~n2647;
  assign n2649 = ~n2644 & ~n2648;
  assign n2650 = ~n2643 & ~n2649;
  assign n2651 = ~n2634 & ~n2640;
  assign n2652 = ~n2650 & ~n2651;
  assign n2653 = ~n2628 & ~n2652;
  assign n2654 = n2600 & n2625;
  assign n2655 = ~n2653 & ~n2654;
  assign n2656 = ~n2565 & n2577;
  assign n2657 = n2565 & ~n2577;
  assign n2658 = ~n2656 & ~n2657;
  assign n2659 = g38 & g39;
  assign n2660 = n2302 & ~n2659;
  assign n2661 = ~g38 & ~g39;
  assign n2662 = ~n2660 & ~n2661;
  assign n2663 = g37 & ~n2662;
  assign n2664 = g50 & n1395;
  assign n2665 = ~g49 & n141;
  assign n2666 = g49 & ~n141;
  assign n2667 = ~n2665 & ~n2666;
  assign n2668 = n2295 & ~n2667;
  assign n2669 = ~n2664 & ~n2668;
  assign n2670 = n2663 & ~n2669;
  assign n2671 = n107 & n2621;
  assign n2672 = ~n103 & ~n2572;
  assign n2673 = ~n2671 & ~n2672;
  assign n2674 = n176 & n1401;
  assign n2675 = ~n175 & ~n2372;
  assign n2676 = ~n2674 & ~n2675;
  assign n2677 = n2673 & ~n2676;
  assign n2678 = ~n2673 & n2676;
  assign n2679 = ~n2677 & ~n2678;
  assign n2680 = n2670 & ~n2679;
  assign n2681 = ~n2673 & ~n2676;
  assign n2682 = ~n2680 & ~n2681;
  assign n2683 = ~n2658 & n2682;
  assign n2684 = n2658 & ~n2682;
  assign n2685 = ~n2683 & ~n2684;
  assign n2686 = n2655 & ~n2685;
  assign n2687 = ~n2655 & n2685;
  assign n2688 = ~n2686 & ~n2687;
  assign n2689 = ~n2530 & n2549;
  assign n2690 = ~n2550 & ~n2689;
  assign n2691 = n374 & ~n1575;
  assign n2692 = ~n370 & n2632;
  assign n2693 = ~n2691 & ~n2692;
  assign n2694 = ~n103 & ~n2302;
  assign n2695 = ~n2693 & n2694;
  assign n2696 = ~n2051 & ~n2647;
  assign n2697 = ~n1621 & n2095;
  assign n2698 = ~n2696 & ~n2697;
  assign n2699 = n2693 & ~n2694;
  assign n2700 = ~n2695 & ~n2699;
  assign n2701 = ~n2698 & n2700;
  assign n2702 = ~n2695 & ~n2701;
  assign n2703 = n2663 & n2669;
  assign n2704 = ~n2663 & ~n2669;
  assign n2705 = ~n2703 & ~n2704;
  assign n2706 = ~n2702 & ~n2705;
  assign n2707 = ~n1626 & n2295;
  assign n2708 = g50 & ~n2667;
  assign n2709 = ~n2707 & ~n2708;
  assign n2710 = ~n262 & n2638;
  assign n2711 = n266 & ~n1615;
  assign n2712 = ~n2710 & ~n2711;
  assign n2713 = n2709 & ~n2712;
  assign n2714 = ~n2709 & n2712;
  assign n2715 = ~n2713 & ~n2714;
  assign n2716 = g39 & n2257;
  assign n2717 = ~g39 & ~n2257;
  assign n2718 = ~n2716 & ~n2717;
  assign n2719 = n176 & ~n2718;
  assign n2720 = ~n175 & ~n2604;
  assign n2721 = ~n2719 & ~n2720;
  assign n2722 = ~n2715 & ~n2721;
  assign n2723 = ~n2709 & ~n2712;
  assign n2724 = ~n2722 & ~n2723;
  assign n2725 = n2702 & n2705;
  assign n2726 = ~n2706 & ~n2725;
  assign n2727 = ~n2724 & n2726;
  assign n2728 = ~n2706 & ~n2727;
  assign n2729 = ~n2670 & n2679;
  assign n2730 = ~n2680 & ~n2729;
  assign n2731 = n2538 & ~n2541;
  assign n2732 = ~n2533 & ~n2541;
  assign n2733 = ~n2536 & n2732;
  assign n2734 = ~n2731 & ~n2733;
  assign n2735 = n2533 & ~n2536;
  assign n2736 = ~n2533 & n2536;
  assign n2737 = ~n2735 & ~n2736;
  assign n2738 = n2541 & ~n2737;
  assign n2739 = n2734 & ~n2738;
  assign n2740 = n2730 & n2739;
  assign n2741 = ~n2730 & ~n2739;
  assign n2742 = ~n2740 & ~n2741;
  assign n2743 = ~n2728 & ~n2742;
  assign n2744 = n2730 & ~n2739;
  assign n2745 = ~n2743 & ~n2744;
  assign n2746 = ~n2690 & ~n2745;
  assign n2747 = n2690 & n2745;
  assign n2748 = ~n2746 & ~n2747;
  assign n2749 = ~n2688 & n2748;
  assign n2750 = n2688 & ~n2748;
  assign n2751 = ~n2749 & ~n2750;
  assign n2752 = n2628 & ~n2652;
  assign n2753 = ~n2628 & n2652;
  assign n2754 = ~n2752 & ~n2753;
  assign n2755 = ~g40 & ~g41;
  assign n2756 = ~n2302 & ~n2755;
  assign n2757 = n226 & ~n2756;
  assign n2758 = g47 & ~n308;
  assign n2759 = ~g47 & n308;
  assign n2760 = ~n2758 & ~n2759;
  assign n2761 = n2095 & ~n2760;
  assign n2762 = ~n1621 & ~n2051;
  assign n2763 = ~n2761 & ~n2762;
  assign n2764 = n2757 & ~n2763;
  assign n2765 = ~n529 & ~n2610;
  assign n2766 = n533 & ~n1559;
  assign n2767 = ~n2765 & ~n2766;
  assign n2768 = ~n2764 & ~n2767;
  assign n2769 = n2757 & n2767;
  assign n2770 = ~n2763 & n2769;
  assign n2771 = ~n2768 & ~n2770;
  assign n2772 = g50 & ~n1626;
  assign n2773 = g49 & ~n194;
  assign n2774 = ~g49 & n194;
  assign n2775 = ~n2773 & ~n2774;
  assign n2776 = n2295 & n2775;
  assign n2777 = ~n2772 & ~n2776;
  assign n2778 = ~n262 & ~n1615;
  assign n2779 = ~g41 & n822;
  assign n2780 = g41 & ~n822;
  assign n2781 = ~n2779 & ~n2780;
  assign n2782 = n266 & n2781;
  assign n2783 = ~n2778 & ~n2782;
  assign n2784 = ~n2777 & ~n2783;
  assign n2785 = ~n370 & ~n1575;
  assign n2786 = ~g43 & n596;
  assign n2787 = g43 & ~n596;
  assign n2788 = ~n2786 & ~n2787;
  assign n2789 = n374 & n2788;
  assign n2790 = ~n2785 & ~n2789;
  assign n2791 = ~n2777 & n2783;
  assign n2792 = n2777 & ~n2783;
  assign n2793 = ~n2791 & ~n2792;
  assign n2794 = ~n2790 & ~n2793;
  assign n2795 = ~n2784 & ~n2794;
  assign n2796 = ~n2771 & ~n2795;
  assign n2797 = n2764 & ~n2767;
  assign n2798 = ~n2796 & ~n2797;
  assign n2799 = n2643 & ~n2649;
  assign n2800 = ~n2643 & n2649;
  assign n2801 = ~n2799 & ~n2800;
  assign n2802 = n2612 & n2623;
  assign n2803 = ~n2612 & ~n2623;
  assign n2804 = ~n2802 & ~n2803;
  assign n2805 = ~n2606 & n2804;
  assign n2806 = n2606 & ~n2804;
  assign n2807 = ~n2805 & ~n2806;
  assign n2808 = ~n2801 & ~n2807;
  assign n2809 = n2801 & n2807;
  assign n2810 = ~n2808 & ~n2809;
  assign n2811 = ~n2798 & ~n2810;
  assign n2812 = ~n2801 & n2807;
  assign n2813 = ~n2811 & ~n2812;
  assign n2814 = ~n2754 & ~n2813;
  assign n2815 = n2728 & ~n2742;
  assign n2816 = ~n2728 & n2742;
  assign n2817 = ~n2815 & ~n2816;
  assign n2818 = n2754 & n2813;
  assign n2819 = ~n2814 & ~n2818;
  assign n2820 = ~n2817 & n2819;
  assign n2821 = ~n2814 & ~n2820;
  assign n2822 = ~n2751 & ~n2821;
  assign n2823 = n2751 & n2821;
  assign n2824 = n2798 & n2810;
  assign n2825 = ~n2811 & ~n2824;
  assign n2826 = n2724 & ~n2726;
  assign n2827 = ~n2727 & ~n2826;
  assign n2828 = n2715 & ~n2721;
  assign n2829 = ~n2715 & n2721;
  assign n2830 = ~n2828 & ~n2829;
  assign n2831 = n2698 & ~n2700;
  assign n2832 = ~n2701 & ~n2831;
  assign n2833 = g45 & n491;
  assign n2834 = ~g45 & ~n491;
  assign n2835 = ~n2833 & ~n2834;
  assign n2836 = n533 & ~n2835;
  assign n2837 = ~n529 & ~n1559;
  assign n2838 = ~n2836 & ~n2837;
  assign n2839 = ~n2757 & ~n2763;
  assign n2840 = n2757 & n2763;
  assign n2841 = ~n2839 & ~n2840;
  assign n2842 = ~n2838 & ~n2841;
  assign n2843 = n2838 & n2841;
  assign n2844 = ~n175 & ~n2718;
  assign n2845 = ~g39 & n2302;
  assign n2846 = n176 & ~n2845;
  assign n2847 = g39 & ~n2302;
  assign n2848 = n2846 & ~n2847;
  assign n2849 = ~n2844 & ~n2848;
  assign n2850 = ~n2843 & ~n2849;
  assign n2851 = ~n2842 & ~n2850;
  assign n2852 = ~n2832 & ~n2851;
  assign n2853 = n2832 & n2851;
  assign n2854 = ~n2852 & ~n2853;
  assign n2855 = ~n2830 & ~n2854;
  assign n2856 = n2832 & ~n2851;
  assign n2857 = ~n2855 & ~n2856;
  assign n2858 = n2827 & n2857;
  assign n2859 = ~n2827 & ~n2857;
  assign n2860 = ~n2858 & ~n2859;
  assign n2861 = n2825 & ~n2860;
  assign n2862 = ~n2825 & n2860;
  assign n2863 = ~n2861 & ~n2862;
  assign n2864 = n2771 & n2795;
  assign n2865 = ~n2796 & ~n2864;
  assign n2866 = g41 & n2257;
  assign n2867 = ~g41 & ~n2257;
  assign n2868 = ~n2866 & ~n2867;
  assign n2869 = n266 & ~n2868;
  assign n2870 = ~n262 & n2781;
  assign n2871 = ~n2869 & ~n2870;
  assign n2872 = n1603 & n2295;
  assign n2873 = g50 & n2775;
  assign n2874 = ~n2872 & ~n2873;
  assign n2875 = ~n2871 & ~n2874;
  assign n2876 = n2871 & n2874;
  assign n2877 = ~n529 & ~n2835;
  assign n2878 = n533 & ~n1653;
  assign n2879 = ~n2877 & ~n2878;
  assign n2880 = ~n2876 & ~n2879;
  assign n2881 = ~n2875 & ~n2880;
  assign n2882 = ~n175 & ~n2302;
  assign n2883 = ~n1659 & n2095;
  assign n2884 = ~n2051 & ~n2760;
  assign n2885 = ~n2883 & ~n2884;
  assign n2886 = n2882 & ~n2885;
  assign n2887 = n374 & ~n1591;
  assign n2888 = ~n370 & n2788;
  assign n2889 = ~n2887 & ~n2888;
  assign n2890 = ~n2882 & n2885;
  assign n2891 = ~n2886 & ~n2890;
  assign n2892 = ~n2889 & n2891;
  assign n2893 = ~n2886 & ~n2892;
  assign n2894 = n2881 & ~n2893;
  assign n2895 = ~n2881 & n2893;
  assign n2896 = ~n2894 & ~n2895;
  assign n2897 = ~n2790 & n2793;
  assign n2898 = n2790 & ~n2793;
  assign n2899 = ~n2897 & ~n2898;
  assign n2900 = ~n2896 & ~n2899;
  assign n2901 = ~n2881 & ~n2893;
  assign n2902 = ~n2900 & ~n2901;
  assign n2903 = n2865 & ~n2902;
  assign n2904 = ~n2830 & n2854;
  assign n2905 = n2830 & ~n2854;
  assign n2906 = ~n2904 & ~n2905;
  assign n2907 = ~n2865 & ~n2902;
  assign n2908 = n2865 & n2902;
  assign n2909 = ~n2907 & ~n2908;
  assign n2910 = ~n2906 & ~n2909;
  assign n2911 = ~n2903 & ~n2910;
  assign n2912 = ~n2863 & n2911;
  assign n2913 = ~n2817 & ~n2819;
  assign n2914 = n2817 & n2819;
  assign n2915 = ~n2913 & ~n2914;
  assign n2916 = n2827 & ~n2857;
  assign n2917 = ~n2861 & ~n2916;
  assign n2918 = n2915 & n2917;
  assign n2919 = n2896 & n2899;
  assign n2920 = ~n2900 & ~n2919;
  assign n2921 = n2838 & ~n2849;
  assign n2922 = ~n2838 & n2849;
  assign n2923 = ~n2921 & ~n2922;
  assign n2924 = ~n2841 & n2923;
  assign n2925 = n2841 & ~n2923;
  assign n2926 = ~n2924 & ~n2925;
  assign n2927 = n2889 & ~n2891;
  assign n2928 = ~n2892 & ~n2927;
  assign n2929 = g42 & g43;
  assign n2930 = n2302 & ~n2929;
  assign n2931 = ~g42 & ~g43;
  assign n2932 = ~n2930 & ~n2931;
  assign n2933 = g41 & ~n2932;
  assign n2934 = g47 & ~n491;
  assign n2935 = ~g47 & n491;
  assign n2936 = ~n2934 & ~n2935;
  assign n2937 = n2095 & n2936;
  assign n2938 = ~n1659 & ~n2051;
  assign n2939 = ~n2937 & ~n2938;
  assign n2940 = n2933 & ~n2939;
  assign n2941 = n2928 & n2940;
  assign n2942 = ~n370 & ~n1591;
  assign n2943 = ~g43 & n822;
  assign n2944 = g43 & ~n822;
  assign n2945 = ~n2943 & ~n2944;
  assign n2946 = n374 & n2945;
  assign n2947 = ~n2942 & ~n2946;
  assign n2948 = g50 & n1603;
  assign n2949 = ~g49 & n308;
  assign n2950 = g49 & ~n308;
  assign n2951 = ~n2949 & ~n2950;
  assign n2952 = n2295 & ~n2951;
  assign n2953 = ~n2948 & ~n2952;
  assign n2954 = g41 & n2302;
  assign n2955 = ~g41 & ~n2302;
  assign n2956 = ~n2954 & ~n2955;
  assign n2957 = n266 & ~n2956;
  assign n2958 = ~n262 & ~n2868;
  assign n2959 = ~n2957 & ~n2958;
  assign n2960 = ~n2953 & n2959;
  assign n2961 = n2953 & ~n2959;
  assign n2962 = ~n2960 & ~n2961;
  assign n2963 = ~n2947 & ~n2962;
  assign n2964 = ~n2953 & ~n2959;
  assign n2965 = ~n2963 & ~n2964;
  assign n2966 = ~n2928 & ~n2940;
  assign n2967 = ~n2941 & ~n2966;
  assign n2968 = ~n2965 & n2967;
  assign n2969 = ~n2941 & ~n2968;
  assign n2970 = ~n2926 & n2969;
  assign n2971 = n2926 & ~n2969;
  assign n2972 = ~n2970 & ~n2971;
  assign n2973 = n2920 & ~n2972;
  assign n2974 = ~n2926 & ~n2969;
  assign n2975 = ~n2973 & ~n2974;
  assign n2976 = n2906 & n2909;
  assign n2977 = ~n2910 & ~n2976;
  assign n2978 = n2975 & ~n2977;
  assign n2979 = ~n2918 & ~n2978;
  assign n2980 = ~n2912 & n2979;
  assign n2981 = n2871 & ~n2874;
  assign n2982 = ~n2871 & n2874;
  assign n2983 = ~n2981 & ~n2982;
  assign n2984 = n2879 & ~n2983;
  assign n2985 = ~n2879 & n2983;
  assign n2986 = ~n2984 & ~n2985;
  assign n2987 = ~n262 & ~n2302;
  assign n2988 = ~n370 & n2945;
  assign n2989 = ~g43 & ~n2257;
  assign n2990 = g43 & n2257;
  assign n2991 = ~n2989 & ~n2990;
  assign n2992 = n374 & ~n2991;
  assign n2993 = ~n2988 & ~n2992;
  assign n2994 = n2987 & ~n2993;
  assign n2995 = ~n2987 & n2993;
  assign n2996 = n1816 & n2295;
  assign n2997 = g50 & ~n2951;
  assign n2998 = ~n2996 & ~n2997;
  assign n2999 = ~n2995 & ~n2998;
  assign n3000 = ~n2994 & ~n2999;
  assign n3001 = ~g45 & n596;
  assign n3002 = g45 & ~n596;
  assign n3003 = ~n3001 & ~n3002;
  assign n3004 = n533 & n3003;
  assign n3005 = ~n529 & ~n1653;
  assign n3006 = ~n3004 & ~n3005;
  assign n3007 = ~n2933 & ~n2939;
  assign n3008 = n2933 & n2939;
  assign n3009 = ~n3007 & ~n3008;
  assign n3010 = ~n3006 & n3009;
  assign n3011 = n3006 & ~n3009;
  assign n3012 = ~n3010 & ~n3011;
  assign n3013 = ~n3000 & ~n3012;
  assign n3014 = ~n3006 & ~n3009;
  assign n3015 = ~n3013 & ~n3014;
  assign n3016 = ~n2986 & n3015;
  assign n3017 = n2986 & ~n3015;
  assign n3018 = ~n3016 & ~n3017;
  assign n3019 = n2965 & n2967;
  assign n3020 = ~n2965 & ~n2967;
  assign n3021 = ~n3019 & ~n3020;
  assign n3022 = ~n3018 & ~n3021;
  assign n3023 = ~n2986 & ~n3015;
  assign n3024 = ~n3022 & ~n3023;
  assign n3025 = ~n2920 & ~n2972;
  assign n3026 = n2920 & n2972;
  assign n3027 = ~n3025 & ~n3026;
  assign n3028 = n3024 & n3027;
  assign n3029 = n3018 & ~n3021;
  assign n3030 = ~n3018 & n3021;
  assign n3031 = ~n3029 & ~n3030;
  assign n3032 = n3000 & n3012;
  assign n3033 = ~n3013 & ~n3032;
  assign n3034 = n1770 & n2095;
  assign n3035 = ~n2051 & n2936;
  assign n3036 = ~n3034 & ~n3035;
  assign n3037 = n533 & ~n1776;
  assign n3038 = ~n529 & n3003;
  assign n3039 = ~n3037 & ~n3038;
  assign n3040 = ~n3036 & ~n3039;
  assign n3041 = g44 & g45;
  assign n3042 = ~g44 & ~g45;
  assign n3043 = ~n2302 & ~n3042;
  assign n3044 = g43 & ~n3043;
  assign n3045 = ~n3041 & n3044;
  assign n3046 = g50 & n1816;
  assign n3047 = ~g49 & n491;
  assign n3048 = g49 & ~n491;
  assign n3049 = ~n3047 & ~n3048;
  assign n3050 = n2295 & n3049;
  assign n3051 = ~n3046 & ~n3050;
  assign n3052 = n3045 & ~n3051;
  assign n3053 = n3036 & n3039;
  assign n3054 = ~n3040 & ~n3053;
  assign n3055 = n3052 & n3054;
  assign n3056 = ~n3040 & ~n3055;
  assign n3057 = n2947 & ~n2962;
  assign n3058 = ~n2947 & n2962;
  assign n3059 = ~n3057 & ~n3058;
  assign n3060 = ~n3056 & n3059;
  assign n3061 = n3056 & ~n3059;
  assign n3062 = ~n3060 & ~n3061;
  assign n3063 = n3033 & ~n3062;
  assign n3064 = ~n3056 & ~n3059;
  assign n3065 = ~n3063 & ~n3064;
  assign n3066 = n3031 & n3065;
  assign n3067 = n3052 & ~n3054;
  assign n3068 = ~n3052 & n3054;
  assign n3069 = ~n3067 & ~n3068;
  assign n3070 = g47 & n596;
  assign n3071 = ~g47 & ~n596;
  assign n3072 = ~n3070 & ~n3071;
  assign n3073 = n2095 & ~n3072;
  assign n3074 = n1770 & ~n2051;
  assign n3075 = ~n3073 & ~n3074;
  assign n3076 = ~n529 & ~n1776;
  assign n3077 = ~g45 & ~n822;
  assign n3078 = g45 & n822;
  assign n3079 = ~n3077 & ~n3078;
  assign n3080 = n533 & ~n3079;
  assign n3081 = ~n3076 & ~n3080;
  assign n3082 = g43 & ~n2302;
  assign n3083 = ~g43 & n2302;
  assign n3084 = ~n3082 & ~n3083;
  assign n3085 = n374 & n3084;
  assign n3086 = ~n370 & ~n2991;
  assign n3087 = ~n3085 & ~n3086;
  assign n3088 = ~n3081 & n3087;
  assign n3089 = n3081 & ~n3087;
  assign n3090 = ~n3088 & ~n3089;
  assign n3091 = ~n3075 & ~n3090;
  assign n3092 = ~n3081 & ~n3087;
  assign n3093 = ~n3091 & ~n3092;
  assign n3094 = n2987 & ~n2998;
  assign n3095 = ~n2987 & n2998;
  assign n3096 = ~n3094 & ~n3095;
  assign n3097 = ~n2993 & n3096;
  assign n3098 = n2993 & ~n3096;
  assign n3099 = ~n3097 & ~n3098;
  assign n3100 = n3093 & n3099;
  assign n3101 = ~n3093 & ~n3099;
  assign n3102 = ~n3100 & ~n3101;
  assign n3103 = ~n3069 & ~n3102;
  assign n3104 = ~n3093 & n3099;
  assign n3105 = ~n3103 & ~n3104;
  assign n3106 = n3033 & n3062;
  assign n3107 = ~n3033 & ~n3062;
  assign n3108 = ~n3106 & ~n3107;
  assign n3109 = ~n3105 & ~n3108;
  assign n3110 = ~n2051 & ~n3072;
  assign n3111 = ~n1859 & n2095;
  assign n3112 = ~n3110 & ~n3111;
  assign n3113 = ~n370 & ~n2302;
  assign n3114 = g50 & n3049;
  assign n3115 = ~n1865 & n2295;
  assign n3116 = ~n3114 & ~n3115;
  assign n3117 = n3113 & n3116;
  assign n3118 = ~n3113 & ~n3116;
  assign n3119 = ~n3117 & ~n3118;
  assign n3120 = ~n3112 & ~n3119;
  assign n3121 = n3113 & ~n3116;
  assign n3122 = ~n3120 & ~n3121;
  assign n3123 = n3045 & n3051;
  assign n3124 = ~n3045 & ~n3051;
  assign n3125 = ~n3123 & ~n3124;
  assign n3126 = ~n3122 & ~n3125;
  assign n3127 = ~n3075 & n3090;
  assign n3128 = n3075 & ~n3090;
  assign n3129 = ~n3127 & ~n3128;
  assign n3130 = n3122 & n3125;
  assign n3131 = ~n3126 & ~n3130;
  assign n3132 = ~n3129 & n3131;
  assign n3133 = ~n3126 & ~n3132;
  assign n3134 = n3069 & ~n3102;
  assign n3135 = ~n3069 & n3102;
  assign n3136 = ~n3134 & ~n3135;
  assign n3137 = ~n3133 & ~n3136;
  assign n3138 = ~n3109 & ~n3137;
  assign n3139 = n3105 & n3108;
  assign n3140 = ~n3138 & ~n3139;
  assign n3141 = ~n3066 & n3140;
  assign n3142 = ~n3031 & ~n3065;
  assign n3143 = ~n3024 & ~n3027;
  assign n3144 = ~n3142 & ~n3143;
  assign n3145 = ~n3141 & n3144;
  assign n3146 = ~n3028 & ~n3145;
  assign n3147 = ~g45 & ~n2257;
  assign n3148 = g45 & n2257;
  assign n3149 = ~n3147 & ~n3148;
  assign n3150 = n533 & ~n3149;
  assign n3151 = ~n529 & ~n3079;
  assign n3152 = ~n3150 & ~n3151;
  assign n3153 = g46 & g47;
  assign n3154 = ~g46 & ~g47;
  assign n3155 = ~n2302 & ~n3154;
  assign n3156 = g45 & ~n3155;
  assign n3157 = ~n3153 & n3156;
  assign n3158 = g50 & ~n1865;
  assign n3159 = ~g49 & n596;
  assign n3160 = g49 & ~n596;
  assign n3161 = ~n3159 & ~n3160;
  assign n3162 = n2295 & n3161;
  assign n3163 = ~n3158 & ~n3162;
  assign n3164 = n3157 & ~n3163;
  assign n3165 = ~n3152 & ~n3164;
  assign n3166 = n3152 & n3164;
  assign n3167 = ~n3165 & ~n3166;
  assign n3168 = n3112 & ~n3119;
  assign n3169 = ~n3112 & n3119;
  assign n3170 = ~n3168 & ~n3169;
  assign n3171 = ~n3167 & ~n3170;
  assign n3172 = ~n3152 & n3164;
  assign n3173 = ~n3171 & ~n3172;
  assign n3174 = ~n3129 & ~n3131;
  assign n3175 = n3129 & n3131;
  assign n3176 = ~n3174 & ~n3175;
  assign n3177 = n3173 & n3176;
  assign n3178 = g45 & n2302;
  assign n3179 = ~g45 & ~n2302;
  assign n3180 = ~n3178 & ~n3179;
  assign n3181 = n533 & ~n3180;
  assign n3182 = ~n529 & ~n3149;
  assign n3183 = ~n3181 & ~n3182;
  assign n3184 = g47 & n822;
  assign n3185 = ~g47 & ~n822;
  assign n3186 = ~n3184 & ~n3185;
  assign n3187 = n2095 & ~n3186;
  assign n3188 = ~n1859 & ~n2051;
  assign n3189 = ~n3187 & ~n3188;
  assign n3190 = ~n3183 & ~n3189;
  assign n3191 = ~n3157 & ~n3163;
  assign n3192 = n3157 & n3163;
  assign n3193 = ~n3191 & ~n3192;
  assign n3194 = n3183 & n3189;
  assign n3195 = ~n3190 & ~n3194;
  assign n3196 = ~n3193 & n3195;
  assign n3197 = ~n3190 & ~n3196;
  assign n3198 = ~n3167 & n3170;
  assign n3199 = n3167 & ~n3170;
  assign n3200 = ~n3198 & ~n3199;
  assign n3201 = n3197 & n3200;
  assign n3202 = g47 & n2257;
  assign n3203 = ~g47 & ~n2257;
  assign n3204 = ~n3202 & ~n3203;
  assign n3205 = n2095 & ~n3204;
  assign n3206 = ~n2051 & ~n3186;
  assign n3207 = ~n3205 & ~n3206;
  assign n3208 = ~n1900 & n2295;
  assign n3209 = g50 & n3161;
  assign n3210 = ~n3208 & ~n3209;
  assign n3211 = ~n529 & ~n2302;
  assign n3212 = n3210 & n3211;
  assign n3213 = ~n3210 & ~n3211;
  assign n3214 = ~n3212 & ~n3213;
  assign n3215 = ~n3207 & ~n3214;
  assign n3216 = ~n3210 & n3211;
  assign n3217 = ~n3215 & ~n3216;
  assign n3218 = ~n3193 & ~n3195;
  assign n3219 = n3193 & n3195;
  assign n3220 = ~n3218 & ~n3219;
  assign n3221 = n3217 & n3220;
  assign n3222 = g48 & g49;
  assign n3223 = n2302 & ~n3222;
  assign n3224 = ~g48 & ~g49;
  assign n3225 = ~n3223 & ~n3224;
  assign n3226 = g47 & ~n3225;
  assign n3227 = g50 & ~n1900;
  assign n3228 = ~g49 & ~n822;
  assign n3229 = g49 & n822;
  assign n3230 = ~n3228 & ~n3229;
  assign n3231 = n2295 & ~n3230;
  assign n3232 = ~n3227 & ~n3231;
  assign n3233 = n3226 & ~n3232;
  assign n3234 = n3207 & ~n3214;
  assign n3235 = ~n3207 & n3214;
  assign n3236 = ~n3234 & ~n3235;
  assign n3237 = n3233 & ~n3236;
  assign n3238 = ~n3233 & n3236;
  assign n3239 = ~n2051 & ~n2302;
  assign n3240 = g49 & n2257;
  assign n3241 = ~g49 & ~n2257;
  assign n3242 = ~n3240 & ~n3241;
  assign n3243 = ~n2295 & n3242;
  assign n3244 = g49 & n2302;
  assign n3245 = ~n3243 & n3244;
  assign n3246 = ~n3239 & ~n3245;
  assign n3247 = n2295 & ~n3242;
  assign n3248 = g50 & ~n3230;
  assign n3249 = ~n3247 & ~n3248;
  assign n3250 = ~n3246 & ~n3249;
  assign n3251 = g47 & n2302;
  assign n3252 = ~g47 & ~n2302;
  assign n3253 = ~n3251 & ~n3252;
  assign n3254 = n2095 & ~n3253;
  assign n3255 = ~n2051 & ~n3204;
  assign n3256 = ~n3254 & ~n3255;
  assign n3257 = n3226 & n3232;
  assign n3258 = ~n3226 & ~n3232;
  assign n3259 = ~n3257 & ~n3258;
  assign n3260 = n3256 & n3259;
  assign n3261 = n3250 & ~n3260;
  assign n3262 = ~n3256 & ~n3259;
  assign n3263 = ~n3261 & ~n3262;
  assign n3264 = ~n3238 & ~n3263;
  assign n3265 = ~n3237 & ~n3264;
  assign n3266 = ~n3221 & ~n3265;
  assign n3267 = ~n3217 & ~n3220;
  assign n3268 = ~n3266 & ~n3267;
  assign n3269 = ~n3201 & ~n3268;
  assign n3270 = ~n3197 & ~n3200;
  assign n3271 = ~n3269 & ~n3270;
  assign n3272 = ~n3177 & ~n3271;
  assign n3273 = ~n3173 & ~n3176;
  assign n3274 = ~n3272 & ~n3273;
  assign n3275 = n3133 & n3136;
  assign n3276 = ~n3139 & ~n3275;
  assign n3277 = ~n3274 & n3276;
  assign n3278 = ~n3028 & ~n3066;
  assign n3279 = n3277 & n3278;
  assign n3280 = ~n3146 & ~n3279;
  assign n3281 = n2980 & ~n3280;
  assign n3282 = ~n2823 & n3281;
  assign n3283 = ~n2915 & ~n2917;
  assign n3284 = ~n2975 & n2977;
  assign n3285 = ~n2912 & n3284;
  assign n3286 = n2863 & ~n2911;
  assign n3287 = ~n3285 & ~n3286;
  assign n3288 = ~n2918 & ~n3287;
  assign n3289 = ~n3283 & ~n3288;
  assign n3290 = ~n2823 & ~n3289;
  assign n3291 = ~n3282 & ~n3290;
  assign n3292 = ~n2822 & n3291;
  assign n3293 = n2593 & n2596;
  assign n3294 = ~n2520 & ~n3293;
  assign n3295 = n2552 & ~n2586;
  assign n3296 = ~n2552 & n2586;
  assign n3297 = ~n3295 & ~n3296;
  assign n3298 = ~n2494 & ~n2499;
  assign n3299 = ~n2496 & n3298;
  assign n3300 = ~n2494 & n2499;
  assign n3301 = n2496 & n3300;
  assign n3302 = n2494 & ~n2499;
  assign n3303 = n2496 & n3302;
  assign n3304 = n2494 & n2499;
  assign n3305 = ~n2496 & n3304;
  assign n3306 = ~n3303 & ~n3305;
  assign n3307 = ~n3301 & n3306;
  assign n3308 = ~n3299 & n3307;
  assign n3309 = ~n2655 & ~n2685;
  assign n3310 = ~n2658 & ~n2682;
  assign n3311 = ~n3309 & ~n3310;
  assign n3312 = ~n3308 & n3311;
  assign n3313 = n3308 & ~n3311;
  assign n3314 = ~n3312 & ~n3313;
  assign n3315 = ~n3297 & ~n3314;
  assign n3316 = ~n3308 & ~n3311;
  assign n3317 = ~n3315 & ~n3316;
  assign n3318 = ~n2589 & ~n2591;
  assign n3319 = n2589 & n2591;
  assign n3320 = ~n3318 & ~n3319;
  assign n3321 = n3317 & n3320;
  assign n3322 = ~n2688 & ~n2748;
  assign n3323 = n2690 & ~n2745;
  assign n3324 = ~n3322 & ~n3323;
  assign n3325 = n3297 & ~n3314;
  assign n3326 = ~n3297 & n3314;
  assign n3327 = ~n3325 & ~n3326;
  assign n3328 = n3324 & n3327;
  assign n3329 = ~n3321 & ~n3328;
  assign n3330 = n3294 & n3329;
  assign n3331 = ~n3292 & n3330;
  assign n3332 = ~n3324 & ~n3327;
  assign n3333 = ~n3321 & n3332;
  assign n3334 = ~n3317 & ~n3320;
  assign n3335 = ~n3333 & ~n3334;
  assign n3336 = n3294 & ~n3335;
  assign n3337 = ~n2516 & ~n2519;
  assign n3338 = ~n3336 & ~n3337;
  assign n3339 = ~n3331 & n3338;
  assign n3340 = ~n2598 & n3339;
  assign n3341 = n2360 & n2472;
  assign n3342 = ~n2480 & ~n2484;
  assign n3343 = ~n3341 & n3342;
  assign n3344 = ~n3340 & n3343;
  assign n3345 = ~n2485 & ~n3344;
  assign n3346 = ~n2193 & n3345;
  assign n3347 = ~n2193 & n2483;
  assign n3348 = n1000 & ~n1009;
  assign n3349 = n886 & ~n1006;
  assign n3350 = ~n3348 & ~n3349;
  assign n3351 = n715 & n998;
  assign n3352 = n317 & n710;
  assign n3353 = ~n3351 & ~n3352;
  assign n3354 = ~n742 & ~n747;
  assign n3355 = ~n404 & ~n3354;
  assign n3356 = ~n3353 & n3355;
  assign n3357 = n3353 & ~n3355;
  assign n3358 = ~n3356 & ~n3357;
  assign n3359 = n733 & n1036;
  assign n3360 = ~n339 & n730;
  assign n3361 = ~n3359 & ~n3360;
  assign n3362 = ~n3358 & n3361;
  assign n3363 = n3358 & ~n3361;
  assign n3364 = ~n3362 & ~n3363;
  assign n3365 = n3350 & ~n3364;
  assign n3366 = ~n3350 & n3364;
  assign n3367 = ~n3365 & ~n3366;
  assign n3368 = ~n379 & n698;
  assign n3369 = n700 & n1004;
  assign n3370 = ~n3368 & ~n3369;
  assign n3371 = n762 & n1030;
  assign n3372 = ~n302 & ~n758;
  assign n3373 = ~n3371 & ~n3372;
  assign n3374 = ~n3370 & n3373;
  assign n3375 = n3370 & ~n3373;
  assign n3376 = ~n3374 & ~n3375;
  assign n3377 = g43 & ~n110;
  assign n3378 = ~n3376 & ~n3377;
  assign n3379 = n3376 & n3377;
  assign n3380 = ~n3378 & ~n3379;
  assign n3381 = ~n1026 & ~n1041;
  assign n3382 = ~n1032 & ~n1038;
  assign n3383 = ~n3381 & ~n3382;
  assign n3384 = ~n1000 & ~n3383;
  assign n3385 = n1000 & n3383;
  assign n3386 = ~n3384 & ~n3385;
  assign n3387 = n3380 & n3386;
  assign n3388 = ~n3380 & ~n3386;
  assign n3389 = ~n3387 & ~n3388;
  assign n3390 = n3367 & ~n3389;
  assign n3391 = ~n3367 & n3389;
  assign n3392 = ~n3390 & ~n3391;
  assign n3393 = ~n1044 & ~n1053;
  assign n3394 = ~n1047 & ~n1050;
  assign n3395 = ~n3393 & ~n3394;
  assign n3396 = ~n3392 & n3395;
  assign n3397 = n3392 & ~n3395;
  assign n3398 = ~n3396 & ~n3397;
  assign n3399 = ~n1017 & ~n1020;
  assign n3400 = ~n1012 & ~n1014;
  assign n3401 = ~n3399 & ~n3400;
  assign n3402 = n3398 & ~n3401;
  assign n3403 = ~n3398 & n3401;
  assign n3404 = ~n3402 & ~n3403;
  assign n3405 = ~n994 & ~n1059;
  assign n3406 = ~n1023 & ~n1056;
  assign n3407 = ~n3405 & ~n3406;
  assign n3408 = ~n3404 & ~n3407;
  assign n3409 = n3404 & n3407;
  assign n3410 = ~n3408 & ~n3409;
  assign n3411 = n3347 & n3410;
  assign n3412 = n3346 & n3411;
  assign n3413 = n2034 & n3412;
  assign n3414 = ~n3347 & ~n3410;
  assign n3415 = n3346 & n3414;
  assign n3416 = ~n2034 & n3415;
  assign n3417 = ~n3346 & n3411;
  assign n3418 = ~n2034 & n3417;
  assign n3419 = ~n3346 & n3414;
  assign n3420 = n2034 & n3419;
  assign n3421 = n2034 & n3417;
  assign n3422 = ~n3420 & ~n3421;
  assign n3423 = ~n3418 & n3422;
  assign n3424 = ~n3416 & n3423;
  assign n3425 = ~n3347 & n3410;
  assign n3426 = ~n3346 & n3425;
  assign n3427 = ~n2034 & n3426;
  assign n3428 = n3346 & n3425;
  assign n3429 = n2034 & n3428;
  assign n3430 = n3347 & ~n3410;
  assign n3431 = n3346 & n3430;
  assign n3432 = ~n2034 & n3431;
  assign n3433 = ~n3429 & ~n3432;
  assign n3434 = ~n3427 & n3433;
  assign n3435 = n3424 & n3434;
  assign n3436 = ~n3413 & n3435;
  assign n3437 = n693 & n3436;
  assign n3438 = n3331 & n3343;
  assign n3439 = ~n3437 & n3438;
  assign n3440 = ~n2484 & ~n3437;
  assign n3441 = ~n3347 & n3440;
  assign n3442 = ~n2480 & ~n3341;
  assign n3443 = ~n2520 & n3440;
  assign n3444 = ~n3293 & ~n3335;
  assign n3445 = ~n2597 & ~n3337;
  assign n3446 = ~n3444 & n3445;
  assign n3447 = n3443 & ~n3446;
  assign n3448 = n3442 & n3447;
  assign n3449 = n2484 & ~n3410;
  assign n3450 = n2034 & n3449;
  assign n3451 = ~n2193 & ~n2484;
  assign n3452 = ~n3346 & n3451;
  assign n3453 = ~n3410 & n3452;
  assign n3454 = n2483 & n3453;
  assign n3455 = n2034 & n3454;
  assign n3456 = n2193 & ~n3410;
  assign n3457 = n2483 & n3456;
  assign n3458 = ~n2034 & n3457;
  assign n3459 = ~n2034 & n3428;
  assign n3460 = n2193 & n3410;
  assign n3461 = n2483 & n3460;
  assign n3462 = n2034 & n3461;
  assign n3463 = ~n3459 & ~n3462;
  assign n3464 = ~n3458 & n3463;
  assign n3465 = ~n3455 & n3464;
  assign n3466 = n3410 & n3452;
  assign n3467 = ~n2483 & n3466;
  assign n3468 = n2034 & n3467;
  assign n3469 = ~n2034 & n3454;
  assign n3470 = n3346 & n3451;
  assign n3471 = n3410 & n3470;
  assign n3472 = ~n2034 & n3471;
  assign n3473 = ~n2483 & n3453;
  assign n3474 = ~n2034 & n3473;
  assign n3475 = ~n3472 & ~n3474;
  assign n3476 = ~n3469 & n3475;
  assign n3477 = ~n3468 & n3476;
  assign n3478 = ~n3410 & n3470;
  assign n3479 = n2034 & n3478;
  assign n3480 = n2484 & n3410;
  assign n3481 = n2483 & n3480;
  assign n3482 = ~n2034 & n3481;
  assign n3483 = ~n3479 & ~n3482;
  assign n3484 = n3477 & n3483;
  assign n3485 = n3465 & n3484;
  assign n3486 = ~n3450 & n3485;
  assign n3487 = ~n693 & ~n3486;
  assign n3488 = ~n3448 & ~n3487;
  assign n3489 = ~n3441 & n3488;
  assign n3490 = ~n3439 & n3489;
  assign n3491 = ~n296 & ~n3490;
  assign n3492 = ~n361 & n3491;
  assign n3493 = n690 & n3492;
  assign n3494 = ~n687 & ~n3493;
  assign n3495 = ~n686 & n3494;
  assign n3496 = n244 & ~n3495;
  assign n3497 = g1 & ~n3496;
  assign n3498 = ~n244 & n3495;
  assign n3499 = n3497 & ~n3498;
  assign n3500 = g35 & g56;
  assign n3501 = ~g35 & ~g56;
  assign n3502 = ~n3500 & ~n3501;
  assign n3503 = n123 & n3502;
  assign n3504 = ~g35 & g55;
  assign n3505 = g35 & ~g55;
  assign n3506 = ~n3504 & ~n3505;
  assign n3507 = ~n119 & ~n3506;
  assign n3508 = ~n3503 & ~n3507;
  assign n3509 = n268 & ~n3508;
  assign n3510 = ~n268 & n3508;
  assign n3511 = ~n3509 & ~n3510;
  assign n3512 = g39 & g52;
  assign n3513 = ~g39 & ~g52;
  assign n3514 = ~n3512 & ~n3513;
  assign n3515 = n176 & n3514;
  assign n3516 = g39 & g51;
  assign n3517 = ~g39 & ~g51;
  assign n3518 = ~n3516 & ~n3517;
  assign n3519 = ~n175 & n3518;
  assign n3520 = ~n3515 & ~n3519;
  assign n3521 = ~n3511 & ~n3520;
  assign n3522 = ~n268 & ~n3508;
  assign n3523 = ~n3521 & ~n3522;
  assign n3524 = n176 & n3518;
  assign n3525 = ~n181 & ~n3524;
  assign n3526 = ~g37 & ~g53;
  assign n3527 = g37 & g53;
  assign n3528 = ~n3526 & ~n3527;
  assign n3529 = n107 & n3528;
  assign n3530 = ~g37 & ~g52;
  assign n3531 = g37 & g52;
  assign n3532 = ~n3530 & ~n3531;
  assign n3533 = ~n103 & n3532;
  assign n3534 = ~n3529 & ~n3533;
  assign n3535 = n123 & ~n3506;
  assign n3536 = ~g35 & ~g54;
  assign n3537 = g35 & g54;
  assign n3538 = ~n3536 & ~n3537;
  assign n3539 = ~n119 & n3538;
  assign n3540 = ~n3535 & ~n3539;
  assign n3541 = n3500 & ~n3540;
  assign n3542 = ~n3500 & n3540;
  assign n3543 = ~n3541 & ~n3542;
  assign n3544 = ~n3534 & ~n3543;
  assign n3545 = n3534 & n3543;
  assign n3546 = ~n3544 & ~n3545;
  assign n3547 = n3525 & n3546;
  assign n3548 = ~n3525 & ~n3546;
  assign n3549 = ~n3547 & ~n3548;
  assign n3550 = ~n3523 & ~n3549;
  assign n3551 = n3525 & ~n3546;
  assign n3552 = ~n3550 & ~n3551;
  assign n3553 = n123 & n3538;
  assign n3554 = ~g35 & ~g53;
  assign n3555 = g35 & g53;
  assign n3556 = ~n3554 & ~n3555;
  assign n3557 = ~n119 & n3556;
  assign n3558 = ~n3553 & ~n3557;
  assign n3559 = ~n3525 & ~n3558;
  assign n3560 = n3525 & n3558;
  assign n3561 = ~n3559 & ~n3560;
  assign n3562 = ~n3534 & n3543;
  assign n3563 = ~n3541 & ~n3562;
  assign n3564 = n3561 & n3563;
  assign n3565 = ~n3561 & ~n3563;
  assign n3566 = ~n3564 & ~n3565;
  assign n3567 = g35 & g55;
  assign n3568 = n107 & n3532;
  assign n3569 = ~g37 & ~g51;
  assign n3570 = g37 & g51;
  assign n3571 = ~n3569 & ~n3570;
  assign n3572 = ~n103 & n3571;
  assign n3573 = ~n3568 & ~n3572;
  assign n3574 = ~n3567 & ~n3573;
  assign n3575 = n3567 & n3573;
  assign n3576 = ~n3574 & ~n3575;
  assign n3577 = n226 & ~n3576;
  assign n3578 = ~n226 & n3576;
  assign n3579 = ~n3577 & ~n3578;
  assign n3580 = n3566 & ~n3579;
  assign n3581 = ~n3566 & n3579;
  assign n3582 = ~n3580 & ~n3581;
  assign n3583 = n3552 & ~n3582;
  assign n3584 = ~n3552 & n3582;
  assign n3585 = ~n3583 & ~n3584;
  assign n3586 = g35 & g58;
  assign n3587 = ~g35 & g57;
  assign n3588 = g35 & ~g57;
  assign n3589 = ~n3587 & ~n3588;
  assign n3590 = n123 & ~n3589;
  assign n3591 = ~n119 & n3502;
  assign n3592 = ~n3590 & ~n3591;
  assign n3593 = n3586 & ~n3592;
  assign n3594 = g41 & g51;
  assign n3595 = ~g41 & ~g51;
  assign n3596 = ~n3594 & ~n3595;
  assign n3597 = n266 & n3596;
  assign n3598 = ~n304 & ~n3597;
  assign n3599 = ~n3586 & ~n3592;
  assign n3600 = n3586 & n3592;
  assign n3601 = ~n3599 & ~n3600;
  assign n3602 = ~n3598 & ~n3601;
  assign n3603 = ~n3593 & ~n3602;
  assign n3604 = ~g39 & g53;
  assign n3605 = g39 & ~g53;
  assign n3606 = ~n3604 & ~n3605;
  assign n3607 = n176 & ~n3606;
  assign n3608 = ~n175 & n3514;
  assign n3609 = ~n3607 & ~n3608;
  assign n3610 = g35 & g57;
  assign n3611 = g37 & g54;
  assign n3612 = ~g37 & ~g54;
  assign n3613 = ~n3611 & ~n3612;
  assign n3614 = n107 & n3613;
  assign n3615 = ~n103 & n3528;
  assign n3616 = ~n3614 & ~n3615;
  assign n3617 = ~n3610 & ~n3616;
  assign n3618 = n3610 & n3616;
  assign n3619 = ~n3617 & ~n3618;
  assign n3620 = ~n3609 & ~n3619;
  assign n3621 = n3609 & n3619;
  assign n3622 = ~n3620 & ~n3621;
  assign n3623 = ~n3603 & n3622;
  assign n3624 = n3511 & ~n3520;
  assign n3625 = ~n3511 & n3520;
  assign n3626 = ~n3624 & ~n3625;
  assign n3627 = n3603 & ~n3622;
  assign n3628 = ~n3623 & ~n3627;
  assign n3629 = ~n3626 & n3628;
  assign n3630 = ~n3623 & ~n3629;
  assign n3631 = n3523 & n3549;
  assign n3632 = ~n3550 & ~n3631;
  assign n3633 = n3610 & ~n3616;
  assign n3634 = ~n3620 & ~n3633;
  assign n3635 = ~n3632 & ~n3634;
  assign n3636 = n3632 & n3634;
  assign n3637 = ~n3635 & ~n3636;
  assign n3638 = ~n3630 & ~n3637;
  assign n3639 = n3632 & ~n3634;
  assign n3640 = ~n3638 & ~n3639;
  assign n3641 = n3585 & n3640;
  assign n3642 = n3561 & ~n3563;
  assign n3643 = ~n3559 & ~n3642;
  assign n3644 = n123 & n3556;
  assign n3645 = ~g35 & ~g52;
  assign n3646 = g35 & g52;
  assign n3647 = ~n3645 & ~n3646;
  assign n3648 = ~n119 & n3647;
  assign n3649 = ~n3644 & ~n3648;
  assign n3650 = n3537 & n3649;
  assign n3651 = ~n3537 & ~n3649;
  assign n3652 = ~n3650 & ~n3651;
  assign n3653 = n107 & n3571;
  assign n3654 = ~n115 & ~n3653;
  assign n3655 = n3652 & n3654;
  assign n3656 = ~n3652 & ~n3654;
  assign n3657 = ~n3655 & ~n3656;
  assign n3658 = ~n226 & ~n3576;
  assign n3659 = n3567 & ~n3573;
  assign n3660 = ~n3658 & ~n3659;
  assign n3661 = ~n3657 & n3660;
  assign n3662 = n3657 & ~n3660;
  assign n3663 = ~n3661 & ~n3662;
  assign n3664 = ~n3643 & n3663;
  assign n3665 = n3643 & ~n3663;
  assign n3666 = ~n3664 & ~n3665;
  assign n3667 = ~n3552 & ~n3582;
  assign n3668 = ~n3566 & ~n3579;
  assign n3669 = ~n3667 & ~n3668;
  assign n3670 = n3666 & n3669;
  assign n3671 = ~n370 & n373;
  assign n3672 = ~g43 & g57;
  assign n3673 = g43 & ~g57;
  assign n3674 = ~n3672 & ~n3673;
  assign n3675 = n3671 & ~n3674;
  assign n3676 = g43 & g56;
  assign n3677 = ~g43 & ~g56;
  assign n3678 = ~n3676 & ~n3677;
  assign n3679 = n370 & n3678;
  assign n3680 = ~n3675 & ~n3679;
  assign n3681 = ~g35 & g65;
  assign n3682 = g35 & ~g65;
  assign n3683 = ~n3681 & ~n3682;
  assign n3684 = n123 & ~n3683;
  assign n3685 = ~g35 & g64;
  assign n3686 = g35 & ~g64;
  assign n3687 = ~n3685 & ~n3686;
  assign n3688 = ~n119 & ~n3687;
  assign n3689 = ~n3684 & ~n3688;
  assign n3690 = ~n3680 & ~n3689;
  assign n3691 = ~g41 & g59;
  assign n3692 = g41 & ~g59;
  assign n3693 = ~n3691 & ~n3692;
  assign n3694 = n266 & ~n3693;
  assign n3695 = ~g41 & g58;
  assign n3696 = g41 & ~g58;
  assign n3697 = ~n3695 & ~n3696;
  assign n3698 = ~n262 & ~n3697;
  assign n3699 = ~n3694 & ~n3698;
  assign n3700 = n3680 & n3689;
  assign n3701 = ~n3690 & ~n3700;
  assign n3702 = ~n3699 & n3701;
  assign n3703 = ~n3690 & ~n3702;
  assign n3704 = g35 & g66;
  assign n3705 = ~g49 & g51;
  assign n3706 = g49 & ~g51;
  assign n3707 = ~n3705 & ~n3706;
  assign n3708 = n2295 & ~n3707;
  assign n3709 = ~n2297 & ~n3708;
  assign n3710 = ~n3704 & ~n3709;
  assign n3711 = n3704 & n3709;
  assign n3712 = ~n3710 & ~n3711;
  assign n3713 = ~g47 & g53;
  assign n3714 = g47 & ~g53;
  assign n3715 = ~n3713 & ~n3714;
  assign n3716 = n2095 & ~n3715;
  assign n3717 = ~g47 & g52;
  assign n3718 = g47 & ~g52;
  assign n3719 = ~n3717 & ~n3718;
  assign n3720 = ~n2051 & ~n3719;
  assign n3721 = ~n3716 & ~n3720;
  assign n3722 = ~n3712 & ~n3721;
  assign n3723 = n3704 & ~n3709;
  assign n3724 = ~n3722 & ~n3723;
  assign n3725 = ~n3703 & ~n3724;
  assign n3726 = ~g45 & g54;
  assign n3727 = g45 & ~g54;
  assign n3728 = ~n3726 & ~n3727;
  assign n3729 = ~n529 & ~n3728;
  assign n3730 = ~n529 & ~n530;
  assign n3731 = ~n531 & n3730;
  assign n3732 = ~g45 & g55;
  assign n3733 = g45 & ~g55;
  assign n3734 = ~n3732 & ~n3733;
  assign n3735 = n3731 & ~n3734;
  assign n3736 = ~n3729 & ~n3735;
  assign n3737 = ~g37 & g63;
  assign n3738 = g37 & ~g63;
  assign n3739 = ~n3737 & ~n3738;
  assign n3740 = n107 & ~n3739;
  assign n3741 = ~g37 & g62;
  assign n3742 = g37 & ~g62;
  assign n3743 = ~n3741 & ~n3742;
  assign n3744 = ~n103 & ~n3743;
  assign n3745 = ~n3740 & ~n3744;
  assign n3746 = ~g39 & g61;
  assign n3747 = g39 & ~g61;
  assign n3748 = ~n3746 & ~n3747;
  assign n3749 = n176 & ~n3748;
  assign n3750 = ~g39 & g60;
  assign n3751 = g39 & ~g60;
  assign n3752 = ~n3750 & ~n3751;
  assign n3753 = ~n175 & ~n3752;
  assign n3754 = ~n3749 & ~n3753;
  assign n3755 = ~n3745 & n3754;
  assign n3756 = n3745 & ~n3754;
  assign n3757 = ~n3755 & ~n3756;
  assign n3758 = ~n3736 & ~n3757;
  assign n3759 = ~n3745 & ~n3754;
  assign n3760 = ~n3758 & ~n3759;
  assign n3761 = n3703 & n3724;
  assign n3762 = ~n3725 & ~n3761;
  assign n3763 = ~n3760 & n3762;
  assign n3764 = ~n3725 & ~n3763;
  assign n3765 = ~g45 & g53;
  assign n3766 = g45 & ~g53;
  assign n3767 = ~n3765 & ~n3766;
  assign n3768 = n3731 & ~n3767;
  assign n3769 = ~g45 & g52;
  assign n3770 = g45 & ~g52;
  assign n3771 = ~n3769 & ~n3770;
  assign n3772 = n529 & ~n3771;
  assign n3773 = ~n3768 & ~n3772;
  assign n3774 = ~g41 & g57;
  assign n3775 = g41 & ~g57;
  assign n3776 = ~n3774 & ~n3775;
  assign n3777 = n266 & ~n3776;
  assign n3778 = ~g41 & g56;
  assign n3779 = g41 & ~g56;
  assign n3780 = ~n3778 & ~n3779;
  assign n3781 = ~n262 & ~n3780;
  assign n3782 = ~n3777 & ~n3781;
  assign n3783 = g35 & g64;
  assign n3784 = n3782 & n3783;
  assign n3785 = ~n3782 & ~n3783;
  assign n3786 = ~n3784 & ~n3785;
  assign n3787 = ~n3773 & n3786;
  assign n3788 = n3773 & ~n3786;
  assign n3789 = ~n3787 & ~n3788;
  assign n3790 = ~g47 & g51;
  assign n3791 = g47 & ~g51;
  assign n3792 = ~n3790 & ~n3791;
  assign n3793 = n2095 & ~n3792;
  assign n3794 = ~n2097 & ~n3793;
  assign n3795 = ~g43 & g55;
  assign n3796 = g43 & ~g55;
  assign n3797 = ~n3795 & ~n3796;
  assign n3798 = n370 & ~n3797;
  assign n3799 = n3671 & n3678;
  assign n3800 = ~n3798 & ~n3799;
  assign n3801 = ~g35 & g63;
  assign n3802 = g35 & ~g63;
  assign n3803 = ~n3801 & ~n3802;
  assign n3804 = n123 & ~n3803;
  assign n3805 = ~g35 & g62;
  assign n3806 = g35 & ~g62;
  assign n3807 = ~n3805 & ~n3806;
  assign n3808 = ~n119 & ~n3807;
  assign n3809 = ~n3804 & ~n3808;
  assign n3810 = ~n3800 & ~n3809;
  assign n3811 = n3800 & n3809;
  assign n3812 = ~n3810 & ~n3811;
  assign n3813 = n3794 & ~n3812;
  assign n3814 = ~n3794 & n3812;
  assign n3815 = ~n3813 & ~n3814;
  assign n3816 = n3789 & ~n3815;
  assign n3817 = ~n3789 & n3815;
  assign n3818 = ~n3816 & ~n3817;
  assign n3819 = ~n3764 & ~n3818;
  assign n3820 = ~n3789 & ~n3815;
  assign n3821 = ~n3819 & ~n3820;
  assign n3822 = ~g37 & g61;
  assign n3823 = g37 & ~g61;
  assign n3824 = ~n3822 & ~n3823;
  assign n3825 = n107 & ~n3824;
  assign n3826 = ~g37 & g60;
  assign n3827 = g37 & ~g60;
  assign n3828 = ~n3826 & ~n3827;
  assign n3829 = ~n103 & ~n3828;
  assign n3830 = ~n3825 & ~n3829;
  assign n3831 = ~g39 & g59;
  assign n3832 = g39 & ~g59;
  assign n3833 = ~n3831 & ~n3832;
  assign n3834 = n176 & ~n3833;
  assign n3835 = ~g39 & g58;
  assign n3836 = g39 & ~g58;
  assign n3837 = ~n3835 & ~n3836;
  assign n3838 = ~n175 & ~n3837;
  assign n3839 = ~n3834 & ~n3838;
  assign n3840 = g43 & g54;
  assign n3841 = ~g43 & ~g54;
  assign n3842 = ~n3840 & ~n3841;
  assign n3843 = n370 & n3842;
  assign n3844 = n3671 & ~n3797;
  assign n3845 = ~n3843 & ~n3844;
  assign n3846 = ~n3839 & ~n3845;
  assign n3847 = n3839 & n3845;
  assign n3848 = ~n3846 & ~n3847;
  assign n3849 = ~n3830 & n3848;
  assign n3850 = n3830 & ~n3848;
  assign n3851 = ~n3849 & ~n3850;
  assign n3852 = n123 & ~n3687;
  assign n3853 = ~n119 & ~n3803;
  assign n3854 = ~n3852 & ~n3853;
  assign n3855 = g35 & g65;
  assign n3856 = g49 & n3855;
  assign n3857 = ~g49 & ~n3855;
  assign n3858 = ~n3856 & ~n3857;
  assign n3859 = ~n3854 & ~n3858;
  assign n3860 = ~g49 & n3855;
  assign n3861 = ~n3859 & ~n3860;
  assign n3862 = n266 & ~n3697;
  assign n3863 = ~n262 & ~n3776;
  assign n3864 = ~n3862 & ~n3863;
  assign n3865 = n2095 & ~n3719;
  assign n3866 = ~n2051 & ~n3792;
  assign n3867 = ~n3865 & ~n3866;
  assign n3868 = ~n3864 & ~n3867;
  assign n3869 = ~n3728 & n3731;
  assign n3870 = n529 & ~n3767;
  assign n3871 = ~n3869 & ~n3870;
  assign n3872 = n3864 & n3867;
  assign n3873 = ~n3871 & ~n3872;
  assign n3874 = ~n3868 & ~n3873;
  assign n3875 = ~n3861 & n3874;
  assign n3876 = n3861 & ~n3874;
  assign n3877 = ~n3875 & ~n3876;
  assign n3878 = n3851 & ~n3877;
  assign n3879 = ~n3861 & ~n3874;
  assign n3880 = ~n3878 & ~n3879;
  assign n3881 = n3731 & ~n3771;
  assign n3882 = g45 & g51;
  assign n3883 = ~g45 & ~g51;
  assign n3884 = ~n3882 & ~n3883;
  assign n3885 = n529 & n3884;
  assign n3886 = ~n3881 & ~n3885;
  assign n3887 = n266 & ~n3780;
  assign n3888 = ~g41 & g55;
  assign n3889 = g41 & ~g55;
  assign n3890 = ~n3888 & ~n3889;
  assign n3891 = ~n262 & ~n3890;
  assign n3892 = ~n3887 & ~n3891;
  assign n3893 = ~n2053 & n3892;
  assign n3894 = n2053 & ~n3892;
  assign n3895 = ~n3893 & ~n3894;
  assign n3896 = ~n3886 & n3895;
  assign n3897 = n3886 & ~n3895;
  assign n3898 = ~n3896 & ~n3897;
  assign n3899 = ~n3773 & ~n3786;
  assign n3900 = ~n3782 & n3783;
  assign n3901 = ~n3899 & ~n3900;
  assign n3902 = ~n3830 & ~n3847;
  assign n3903 = ~n3846 & ~n3902;
  assign n3904 = ~n3901 & n3903;
  assign n3905 = n3901 & ~n3903;
  assign n3906 = ~n3904 & ~n3905;
  assign n3907 = ~n3898 & n3906;
  assign n3908 = n3898 & ~n3906;
  assign n3909 = ~n3907 & ~n3908;
  assign n3910 = n3880 & n3909;
  assign n3911 = ~n3880 & ~n3909;
  assign n3912 = ~n3910 & ~n3911;
  assign n3913 = n3821 & n3912;
  assign n3914 = ~n3821 & ~n3912;
  assign n3915 = ~n3913 & ~n3914;
  assign n3916 = n123 & ~n3807;
  assign n3917 = ~g35 & g61;
  assign n3918 = g35 & ~g61;
  assign n3919 = ~n3917 & ~n3918;
  assign n3920 = ~n119 & ~n3919;
  assign n3921 = ~n3916 & ~n3920;
  assign n3922 = n107 & ~n3828;
  assign n3923 = ~g37 & g59;
  assign n3924 = g37 & ~g59;
  assign n3925 = ~n3923 & ~n3924;
  assign n3926 = ~n103 & ~n3925;
  assign n3927 = ~n3922 & ~n3926;
  assign n3928 = n3921 & ~n3927;
  assign n3929 = ~n3921 & n3927;
  assign n3930 = ~n3928 & ~n3929;
  assign n3931 = n3794 & ~n3930;
  assign n3932 = ~n3794 & n3930;
  assign n3933 = ~n3931 & ~n3932;
  assign n3934 = n3794 & n3812;
  assign n3935 = ~n3810 & ~n3934;
  assign n3936 = n176 & ~n3837;
  assign n3937 = ~g39 & g57;
  assign n3938 = g39 & ~g57;
  assign n3939 = ~n3937 & ~n3938;
  assign n3940 = ~n175 & ~n3939;
  assign n3941 = ~n3936 & ~n3940;
  assign n3942 = g35 & g63;
  assign n3943 = ~g43 & g53;
  assign n3944 = g43 & ~g53;
  assign n3945 = ~n3943 & ~n3944;
  assign n3946 = n370 & ~n3945;
  assign n3947 = n3671 & n3842;
  assign n3948 = ~n3946 & ~n3947;
  assign n3949 = n3942 & ~n3948;
  assign n3950 = ~n3942 & n3948;
  assign n3951 = ~n3949 & ~n3950;
  assign n3952 = ~n3941 & ~n3951;
  assign n3953 = n3941 & n3951;
  assign n3954 = ~n3952 & ~n3953;
  assign n3955 = n3935 & ~n3954;
  assign n3956 = ~n3935 & n3954;
  assign n3957 = ~n3955 & ~n3956;
  assign n3958 = n3933 & n3957;
  assign n3959 = ~n3933 & ~n3957;
  assign n3960 = ~n3958 & ~n3959;
  assign n3961 = ~n3851 & ~n3877;
  assign n3962 = n3851 & n3877;
  assign n3963 = ~n3961 & ~n3962;
  assign n3964 = n107 & ~n3743;
  assign n3965 = ~n103 & ~n3824;
  assign n3966 = ~n3964 & ~n3965;
  assign n3967 = n3800 & ~n3966;
  assign n3968 = n176 & ~n3752;
  assign n3969 = ~n175 & ~n3833;
  assign n3970 = ~n3968 & ~n3969;
  assign n3971 = ~n3800 & n3966;
  assign n3972 = ~n3967 & ~n3971;
  assign n3973 = ~n3970 & n3972;
  assign n3974 = ~n3967 & ~n3973;
  assign n3975 = ~n3963 & ~n3974;
  assign n3976 = ~g39 & g62;
  assign n3977 = g39 & ~g62;
  assign n3978 = ~n3976 & ~n3977;
  assign n3979 = n176 & ~n3978;
  assign n3980 = ~n175 & ~n3748;
  assign n3981 = ~n3979 & ~n3980;
  assign n3982 = ~g45 & g56;
  assign n3983 = g45 & ~g56;
  assign n3984 = ~n3982 & ~n3983;
  assign n3985 = n3731 & ~n3984;
  assign n3986 = n529 & ~n3734;
  assign n3987 = ~n3985 & ~n3986;
  assign n3988 = ~n3981 & ~n3987;
  assign n3989 = ~g41 & g60;
  assign n3990 = g41 & ~g60;
  assign n3991 = ~n3989 & ~n3990;
  assign n3992 = n266 & ~n3991;
  assign n3993 = ~n262 & ~n3693;
  assign n3994 = ~n3992 & ~n3993;
  assign n3995 = n3981 & n3987;
  assign n3996 = ~n3988 & ~n3995;
  assign n3997 = ~n3994 & n3996;
  assign n3998 = ~n3988 & ~n3997;
  assign n3999 = ~g66 & ~n2396;
  assign n4000 = ~n2394 & ~n3999;
  assign n4001 = g35 & ~n4000;
  assign n4002 = ~g49 & g52;
  assign n4003 = g49 & ~g52;
  assign n4004 = ~n4002 & ~n4003;
  assign n4005 = n2295 & ~n4004;
  assign n4006 = g50 & ~n3707;
  assign n4007 = ~n4005 & ~n4006;
  assign n4008 = n4001 & ~n4007;
  assign n4009 = ~n119 & ~n3683;
  assign n4010 = ~g35 & ~g66;
  assign n4011 = ~n3704 & ~n4010;
  assign n4012 = n123 & n4011;
  assign n4013 = ~n4009 & ~n4012;
  assign n4014 = ~g47 & g54;
  assign n4015 = g47 & ~g54;
  assign n4016 = ~n4014 & ~n4015;
  assign n4017 = n2095 & ~n4016;
  assign n4018 = ~n2051 & ~n3715;
  assign n4019 = ~n4017 & ~n4018;
  assign n4020 = ~n4013 & ~n4019;
  assign n4021 = n4013 & n4019;
  assign n4022 = n370 & ~n3674;
  assign n4023 = ~g43 & g58;
  assign n4024 = g43 & ~g58;
  assign n4025 = ~n4023 & ~n4024;
  assign n4026 = n3671 & ~n4025;
  assign n4027 = ~n4022 & ~n4026;
  assign n4028 = ~n4021 & ~n4027;
  assign n4029 = ~n4020 & ~n4028;
  assign n4030 = ~n4008 & ~n4029;
  assign n4031 = n4008 & n4029;
  assign n4032 = ~n4030 & ~n4031;
  assign n4033 = ~n3998 & ~n4032;
  assign n4034 = n4008 & ~n4029;
  assign n4035 = ~n4033 & ~n4034;
  assign n4036 = n3854 & ~n3858;
  assign n4037 = ~n3854 & n3858;
  assign n4038 = ~n4036 & ~n4037;
  assign n4039 = n3864 & ~n3871;
  assign n4040 = ~n3864 & n3871;
  assign n4041 = ~n4039 & ~n4040;
  assign n4042 = ~n3867 & n4041;
  assign n4043 = n3867 & ~n4041;
  assign n4044 = ~n4042 & ~n4043;
  assign n4045 = n4038 & ~n4044;
  assign n4046 = ~n4038 & n4044;
  assign n4047 = ~n4045 & ~n4046;
  assign n4048 = ~n4035 & ~n4047;
  assign n4049 = ~n4038 & ~n4044;
  assign n4050 = ~n4048 & ~n4049;
  assign n4051 = n3963 & n3974;
  assign n4052 = ~n3975 & ~n4051;
  assign n4053 = ~n4050 & n4052;
  assign n4054 = ~n3975 & ~n4053;
  assign n4055 = ~n3960 & ~n4054;
  assign n4056 = n3960 & n4054;
  assign n4057 = ~n4055 & ~n4056;
  assign n4058 = ~n3915 & ~n4057;
  assign n4059 = n3960 & ~n4054;
  assign n4060 = ~n4058 & ~n4059;
  assign n4061 = n266 & ~n3890;
  assign n4062 = g41 & g54;
  assign n4063 = ~g41 & ~g54;
  assign n4064 = ~n4062 & ~n4063;
  assign n4065 = ~n262 & n4064;
  assign n4066 = ~n4061 & ~n4065;
  assign n4067 = n123 & ~n3919;
  assign n4068 = ~g35 & g60;
  assign n4069 = g35 & ~g60;
  assign n4070 = ~n4068 & ~n4069;
  assign n4071 = ~n119 & ~n4070;
  assign n4072 = ~n4067 & ~n4071;
  assign n4073 = g35 & g62;
  assign n4074 = n4072 & n4073;
  assign n4075 = ~n4072 & ~n4073;
  assign n4076 = ~n4074 & ~n4075;
  assign n4077 = ~n4066 & n4076;
  assign n4078 = n4066 & ~n4076;
  assign n4079 = ~n4077 & ~n4078;
  assign n4080 = ~n3794 & ~n3921;
  assign n4081 = n3794 & n3921;
  assign n4082 = ~n3927 & ~n4081;
  assign n4083 = ~n4080 & ~n4082;
  assign n4084 = n176 & ~n3939;
  assign n4085 = g39 & g56;
  assign n4086 = ~g39 & ~g56;
  assign n4087 = ~n4085 & ~n4086;
  assign n4088 = ~n175 & n4087;
  assign n4089 = ~n4084 & ~n4088;
  assign n4090 = ~g43 & g52;
  assign n4091 = g43 & ~g52;
  assign n4092 = ~n4090 & ~n4091;
  assign n4093 = n370 & ~n4092;
  assign n4094 = n3671 & ~n3945;
  assign n4095 = ~n4093 & ~n4094;
  assign n4096 = n107 & ~n3925;
  assign n4097 = ~g37 & g58;
  assign n4098 = g37 & ~g58;
  assign n4099 = ~n4097 & ~n4098;
  assign n4100 = ~n103 & ~n4099;
  assign n4101 = ~n4096 & ~n4100;
  assign n4102 = n4095 & ~n4101;
  assign n4103 = ~n4095 & n4101;
  assign n4104 = ~n4102 & ~n4103;
  assign n4105 = ~n4089 & n4104;
  assign n4106 = n4089 & ~n4104;
  assign n4107 = ~n4105 & ~n4106;
  assign n4108 = ~n4083 & n4107;
  assign n4109 = n4083 & ~n4107;
  assign n4110 = ~n4108 & ~n4109;
  assign n4111 = ~n4079 & ~n4110;
  assign n4112 = n4079 & n4110;
  assign n4113 = ~n4111 & ~n4112;
  assign n4114 = ~n3886 & ~n3895;
  assign n4115 = ~n2053 & ~n3892;
  assign n4116 = ~n4114 & ~n4115;
  assign n4117 = n3731 & n3884;
  assign n4118 = g45 & n529;
  assign n4119 = ~n4117 & ~n4118;
  assign n4120 = ~n3941 & n3951;
  assign n4121 = ~n3949 & ~n4120;
  assign n4122 = n4119 & n4121;
  assign n4123 = ~n4119 & ~n4121;
  assign n4124 = ~n4122 & ~n4123;
  assign n4125 = n4116 & ~n4124;
  assign n4126 = ~n4116 & n4124;
  assign n4127 = ~n4125 & ~n4126;
  assign n4128 = ~n3898 & ~n3906;
  assign n4129 = ~n3901 & ~n3903;
  assign n4130 = ~n4128 & ~n4129;
  assign n4131 = n4127 & ~n4130;
  assign n4132 = ~n4127 & n4130;
  assign n4133 = ~n4131 & ~n4132;
  assign n4134 = ~n4113 & ~n4133;
  assign n4135 = n4113 & n4133;
  assign n4136 = ~n4134 & ~n4135;
  assign n4137 = ~n3935 & ~n3954;
  assign n4138 = ~n3959 & ~n4137;
  assign n4139 = ~n3821 & n3912;
  assign n4140 = ~n3911 & ~n4139;
  assign n4141 = ~n4138 & n4140;
  assign n4142 = n4138 & ~n4140;
  assign n4143 = ~n4141 & ~n4142;
  assign n4144 = ~n4136 & n4143;
  assign n4145 = n4136 & ~n4143;
  assign n4146 = ~n4144 & ~n4145;
  assign n4147 = n4060 & n4146;
  assign n4148 = ~g41 & g53;
  assign n4149 = g41 & ~g53;
  assign n4150 = ~n4148 & ~n4149;
  assign n4151 = n266 & ~n4150;
  assign n4152 = g41 & ~g52;
  assign n4153 = ~g41 & g52;
  assign n4154 = ~n4152 & ~n4153;
  assign n4155 = ~n262 & ~n4154;
  assign n4156 = ~n4151 & ~n4155;
  assign n4157 = g35 & g60;
  assign n4158 = ~g39 & g55;
  assign n4159 = g39 & ~g55;
  assign n4160 = ~n4158 & ~n4159;
  assign n4161 = n176 & ~n4160;
  assign n4162 = g39 & g54;
  assign n4163 = ~g39 & ~g54;
  assign n4164 = ~n4162 & ~n4163;
  assign n4165 = ~n175 & n4164;
  assign n4166 = ~n4161 & ~n4165;
  assign n4167 = ~n4157 & ~n4166;
  assign n4168 = n4157 & n4166;
  assign n4169 = ~n4167 & ~n4168;
  assign n4170 = ~n4156 & ~n4169;
  assign n4171 = n4156 & n4169;
  assign n4172 = ~n4170 & ~n4171;
  assign n4173 = g35 & g61;
  assign n4174 = ~n4119 & n4173;
  assign n4175 = n4119 & ~n4173;
  assign n4176 = ~n4089 & ~n4104;
  assign n4177 = ~n4095 & ~n4101;
  assign n4178 = ~n4176 & ~n4177;
  assign n4179 = ~n4175 & ~n4178;
  assign n4180 = ~n4174 & ~n4179;
  assign n4181 = n4172 & ~n4180;
  assign n4182 = ~n4172 & n4180;
  assign n4183 = ~n4181 & ~n4182;
  assign n4184 = n107 & ~n4099;
  assign n4185 = ~g37 & g57;
  assign n4186 = g37 & ~g57;
  assign n4187 = ~n4185 & ~n4186;
  assign n4188 = ~n103 & ~n4187;
  assign n4189 = ~n4184 & ~n4188;
  assign n4190 = n123 & ~n4070;
  assign n4191 = ~g35 & g59;
  assign n4192 = g35 & ~g59;
  assign n4193 = ~n4191 & ~n4192;
  assign n4194 = ~n119 & ~n4193;
  assign n4195 = ~n4190 & ~n4194;
  assign n4196 = ~n4189 & ~n4195;
  assign n4197 = n4189 & n4195;
  assign n4198 = ~n4196 & ~n4197;
  assign n4199 = n266 & n4064;
  assign n4200 = ~n262 & ~n4150;
  assign n4201 = ~n4199 & ~n4200;
  assign n4202 = ~n4198 & ~n4201;
  assign n4203 = n4198 & n4201;
  assign n4204 = ~n4202 & ~n4203;
  assign n4205 = ~n4066 & ~n4076;
  assign n4206 = ~n4072 & n4073;
  assign n4207 = ~n4205 & ~n4206;
  assign n4208 = g43 & g51;
  assign n4209 = ~g43 & ~g51;
  assign n4210 = ~n4208 & ~n4209;
  assign n4211 = n370 & n4210;
  assign n4212 = n3671 & ~n4092;
  assign n4213 = ~n4211 & ~n4212;
  assign n4214 = ~n538 & n4213;
  assign n4215 = n538 & ~n4213;
  assign n4216 = ~n4214 & ~n4215;
  assign n4217 = n176 & n4087;
  assign n4218 = ~n175 & ~n4160;
  assign n4219 = ~n4217 & ~n4218;
  assign n4220 = n4216 & ~n4219;
  assign n4221 = ~n4216 & n4219;
  assign n4222 = ~n4220 & ~n4221;
  assign n4223 = n4207 & ~n4222;
  assign n4224 = ~n4207 & n4222;
  assign n4225 = ~n4223 & ~n4224;
  assign n4226 = ~n4204 & ~n4225;
  assign n4227 = ~n4207 & ~n4222;
  assign n4228 = ~n4226 & ~n4227;
  assign n4229 = ~n4183 & n4228;
  assign n4230 = n4183 & ~n4228;
  assign n4231 = ~n4229 & ~n4230;
  assign n4232 = ~n4083 & ~n4107;
  assign n4233 = ~n4111 & ~n4232;
  assign n4234 = ~n4116 & ~n4124;
  assign n4235 = n4119 & ~n4121;
  assign n4236 = ~n4234 & ~n4235;
  assign n4237 = ~n4119 & ~n4173;
  assign n4238 = n4119 & n4173;
  assign n4239 = ~n4237 & ~n4238;
  assign n4240 = n4178 & ~n4239;
  assign n4241 = ~n4178 & n4239;
  assign n4242 = ~n4240 & ~n4241;
  assign n4243 = ~n4236 & n4242;
  assign n4244 = n4236 & ~n4242;
  assign n4245 = ~n4243 & ~n4244;
  assign n4246 = ~n4233 & ~n4245;
  assign n4247 = ~n4236 & ~n4242;
  assign n4248 = ~n4246 & ~n4247;
  assign n4249 = ~n4216 & ~n4219;
  assign n4250 = ~n538 & ~n4213;
  assign n4251 = ~n4249 & ~n4250;
  assign n4252 = n123 & ~n4193;
  assign n4253 = ~g35 & g58;
  assign n4254 = g35 & ~g58;
  assign n4255 = ~n4253 & ~n4254;
  assign n4256 = ~n119 & ~n4255;
  assign n4257 = ~n4252 & ~n4256;
  assign n4258 = g43 & n370;
  assign n4259 = n3671 & n4210;
  assign n4260 = ~n4258 & ~n4259;
  assign n4261 = n107 & ~n4187;
  assign n4262 = ~g37 & g56;
  assign n4263 = g37 & ~g56;
  assign n4264 = ~n4262 & ~n4263;
  assign n4265 = ~n103 & ~n4264;
  assign n4266 = ~n4261 & ~n4265;
  assign n4267 = n4260 & ~n4266;
  assign n4268 = ~n4260 & n4266;
  assign n4269 = ~n4267 & ~n4268;
  assign n4270 = n4257 & ~n4269;
  assign n4271 = ~n4257 & n4269;
  assign n4272 = ~n4270 & ~n4271;
  assign n4273 = n4251 & ~n4272;
  assign n4274 = ~n4251 & n4272;
  assign n4275 = ~n4273 & ~n4274;
  assign n4276 = n4198 & ~n4201;
  assign n4277 = ~n4196 & ~n4276;
  assign n4278 = ~n4275 & n4277;
  assign n4279 = n4275 & ~n4277;
  assign n4280 = ~n4278 & ~n4279;
  assign n4281 = n4248 & ~n4280;
  assign n4282 = ~n4248 & n4280;
  assign n4283 = ~n4281 & ~n4282;
  assign n4284 = ~n4231 & n4283;
  assign n4285 = n4231 & ~n4283;
  assign n4286 = ~n4284 & ~n4285;
  assign n4287 = n4204 & ~n4225;
  assign n4288 = ~n4204 & n4225;
  assign n4289 = ~n4287 & ~n4288;
  assign n4290 = n4233 & ~n4245;
  assign n4291 = ~n4233 & n4245;
  assign n4292 = ~n4290 & ~n4291;
  assign n4293 = ~n4289 & ~n4292;
  assign n4294 = n4113 & ~n4133;
  assign n4295 = ~n4127 & ~n4130;
  assign n4296 = ~n4294 & ~n4295;
  assign n4297 = n4289 & n4292;
  assign n4298 = ~n4293 & ~n4297;
  assign n4299 = ~n4296 & n4298;
  assign n4300 = ~n4293 & ~n4299;
  assign n4301 = n4286 & n4300;
  assign n4302 = ~n4296 & ~n4298;
  assign n4303 = n4296 & n4298;
  assign n4304 = ~n4302 & ~n4303;
  assign n4305 = ~n4136 & ~n4143;
  assign n4306 = ~n4138 & ~n4140;
  assign n4307 = ~n4305 & ~n4306;
  assign n4308 = n4304 & n4307;
  assign n4309 = ~n4301 & ~n4308;
  assign n4310 = ~n4147 & n4309;
  assign n4311 = ~g43 & g59;
  assign n4312 = g43 & ~g59;
  assign n4313 = ~n4311 & ~n4312;
  assign n4314 = n370 & ~n4313;
  assign n4315 = ~g43 & g60;
  assign n4316 = g43 & ~g60;
  assign n4317 = ~n4315 & ~n4316;
  assign n4318 = n3671 & ~n4317;
  assign n4319 = ~n4314 & ~n4318;
  assign n4320 = ~g41 & g62;
  assign n4321 = g41 & ~g62;
  assign n4322 = ~n4320 & ~n4321;
  assign n4323 = n266 & ~n4322;
  assign n4324 = ~g41 & g61;
  assign n4325 = g41 & ~g61;
  assign n4326 = ~n4324 & ~n4325;
  assign n4327 = ~n262 & ~n4326;
  assign n4328 = ~n4323 & ~n4327;
  assign n4329 = ~g47 & g56;
  assign n4330 = g47 & ~g56;
  assign n4331 = ~n4329 & ~n4330;
  assign n4332 = n2095 & ~n4331;
  assign n4333 = ~g47 & g55;
  assign n4334 = g47 & ~g55;
  assign n4335 = ~n4333 & ~n4334;
  assign n4336 = ~n2051 & ~n4335;
  assign n4337 = ~n4332 & ~n4336;
  assign n4338 = n4328 & ~n4337;
  assign n4339 = ~n4328 & n4337;
  assign n4340 = ~n4338 & ~n4339;
  assign n4341 = ~n4319 & ~n4340;
  assign n4342 = ~n4328 & ~n4337;
  assign n4343 = ~n4341 & ~n4342;
  assign n4344 = n2095 & ~n4335;
  assign n4345 = ~n2051 & ~n4016;
  assign n4346 = ~n4344 & ~n4345;
  assign n4347 = ~g49 & g53;
  assign n4348 = g49 & ~g53;
  assign n4349 = ~n4347 & ~n4348;
  assign n4350 = n2295 & ~n4349;
  assign n4351 = g50 & ~n4004;
  assign n4352 = ~n4350 & ~n4351;
  assign n4353 = g66 & ~n119;
  assign n4354 = ~n4352 & ~n4353;
  assign n4355 = n4352 & n4353;
  assign n4356 = ~n4354 & ~n4355;
  assign n4357 = ~n4346 & n4356;
  assign n4358 = n4346 & ~n4356;
  assign n4359 = ~n4357 & ~n4358;
  assign n4360 = ~g37 & g66;
  assign n4361 = g37 & ~g66;
  assign n4362 = ~n4360 & ~n4361;
  assign n4363 = n107 & ~n4362;
  assign n4364 = ~g37 & g65;
  assign n4365 = g37 & ~g65;
  assign n4366 = ~n4364 & ~n4365;
  assign n4367 = ~n103 & ~n4366;
  assign n4368 = ~n4363 & ~n4367;
  assign n4369 = ~g39 & g64;
  assign n4370 = g39 & ~g64;
  assign n4371 = ~n4369 & ~n4370;
  assign n4372 = n176 & ~n4371;
  assign n4373 = ~g39 & g63;
  assign n4374 = g39 & ~g63;
  assign n4375 = ~n4373 & ~n4374;
  assign n4376 = ~n175 & ~n4375;
  assign n4377 = ~n4372 & ~n4376;
  assign n4378 = ~n4368 & ~n4377;
  assign n4379 = g45 & ~g58;
  assign n4380 = ~g45 & g58;
  assign n4381 = ~n4379 & ~n4380;
  assign n4382 = n3731 & ~n4381;
  assign n4383 = ~g45 & g57;
  assign n4384 = g45 & ~g57;
  assign n4385 = ~n4383 & ~n4384;
  assign n4386 = ~n529 & ~n4385;
  assign n4387 = ~n4382 & ~n4386;
  assign n4388 = n4368 & n4377;
  assign n4389 = ~n4378 & ~n4388;
  assign n4390 = ~n4387 & n4389;
  assign n4391 = ~n4378 & ~n4390;
  assign n4392 = n4359 & ~n4391;
  assign n4393 = ~n4359 & n4391;
  assign n4394 = ~n4392 & ~n4393;
  assign n4395 = ~n4343 & ~n4394;
  assign n4396 = ~n4359 & ~n4391;
  assign n4397 = ~n4395 & ~n4396;
  assign n4398 = ~g37 & g64;
  assign n4399 = g37 & ~g64;
  assign n4400 = ~n4398 & ~n4399;
  assign n4401 = n107 & ~n4400;
  assign n4402 = ~n103 & ~n3739;
  assign n4403 = ~n4401 & ~n4402;
  assign n4404 = ~n4001 & n4007;
  assign n4405 = ~n4008 & ~n4404;
  assign n4406 = ~n4403 & ~n4405;
  assign n4407 = n4403 & n4405;
  assign n4408 = ~n4406 & ~n4407;
  assign n4409 = ~n4352 & n4353;
  assign n4410 = ~n4346 & ~n4356;
  assign n4411 = ~n4409 & ~n4410;
  assign n4412 = ~n4408 & ~n4411;
  assign n4413 = n4408 & n4411;
  assign n4414 = ~n4412 & ~n4413;
  assign n4415 = n176 & ~n4375;
  assign n4416 = ~n175 & ~n3978;
  assign n4417 = ~n4415 & ~n4416;
  assign n4418 = ~g66 & ~n2659;
  assign n4419 = ~n2661 & ~n4418;
  assign n4420 = g37 & ~n4419;
  assign n4421 = ~g49 & g54;
  assign n4422 = g49 & ~g54;
  assign n4423 = ~n4421 & ~n4422;
  assign n4424 = n2295 & ~n4423;
  assign n4425 = g50 & ~n4349;
  assign n4426 = ~n4424 & ~n4425;
  assign n4427 = n4420 & ~n4426;
  assign n4428 = ~n4417 & n4427;
  assign n4429 = n107 & ~n4366;
  assign n4430 = ~n103 & ~n4400;
  assign n4431 = ~n4429 & ~n4430;
  assign n4432 = n4417 & ~n4427;
  assign n4433 = ~n4428 & ~n4432;
  assign n4434 = ~n4431 & n4433;
  assign n4435 = ~n4428 & ~n4434;
  assign n4436 = n4414 & n4435;
  assign n4437 = ~n4414 & ~n4435;
  assign n4438 = ~n4436 & ~n4437;
  assign n4439 = ~n4397 & ~n4438;
  assign n4440 = n4397 & n4438;
  assign n4441 = ~n4439 & ~n4440;
  assign n4442 = n4420 & n4426;
  assign n4443 = ~n4420 & ~n4426;
  assign n4444 = ~n4442 & ~n4443;
  assign n4445 = ~g47 & g57;
  assign n4446 = g47 & ~g57;
  assign n4447 = ~n4445 & ~n4446;
  assign n4448 = n2095 & ~n4447;
  assign n4449 = ~n2051 & ~n4331;
  assign n4450 = ~n4448 & ~n4449;
  assign n4451 = g66 & ~n103;
  assign n4452 = ~g43 & g61;
  assign n4453 = g43 & ~g61;
  assign n4454 = ~n4452 & ~n4453;
  assign n4455 = n3671 & ~n4454;
  assign n4456 = n370 & ~n4317;
  assign n4457 = ~n4455 & ~n4456;
  assign n4458 = ~n4451 & ~n4457;
  assign n4459 = n4451 & n4457;
  assign n4460 = ~n4458 & ~n4459;
  assign n4461 = ~n4450 & ~n4460;
  assign n4462 = n4451 & ~n4457;
  assign n4463 = ~n4461 & ~n4462;
  assign n4464 = ~n4444 & ~n4463;
  assign n4465 = ~g39 & g65;
  assign n4466 = g39 & ~g65;
  assign n4467 = ~n4465 & ~n4466;
  assign n4468 = n176 & ~n4467;
  assign n4469 = ~n175 & ~n4371;
  assign n4470 = ~n4468 & ~n4469;
  assign n4471 = ~g41 & g63;
  assign n4472 = g41 & ~g63;
  assign n4473 = ~n4471 & ~n4472;
  assign n4474 = n266 & ~n4473;
  assign n4475 = ~n262 & ~n4322;
  assign n4476 = ~n4474 & ~n4475;
  assign n4477 = ~g49 & g55;
  assign n4478 = g49 & ~g55;
  assign n4479 = ~n4477 & ~n4478;
  assign n4480 = n2295 & ~n4479;
  assign n4481 = g50 & ~n4423;
  assign n4482 = ~n4480 & ~n4481;
  assign n4483 = n4476 & ~n4482;
  assign n4484 = ~n4476 & n4482;
  assign n4485 = ~n4483 & ~n4484;
  assign n4486 = ~n4470 & ~n4485;
  assign n4487 = ~n4476 & ~n4482;
  assign n4488 = ~n4486 & ~n4487;
  assign n4489 = n4444 & n4463;
  assign n4490 = ~n4464 & ~n4489;
  assign n4491 = ~n4488 & n4490;
  assign n4492 = ~n4464 & ~n4491;
  assign n4493 = n4431 & ~n4433;
  assign n4494 = ~n4434 & ~n4493;
  assign n4495 = n3731 & ~n4385;
  assign n4496 = ~n529 & ~n3984;
  assign n4497 = ~n4495 & ~n4496;
  assign n4498 = n370 & ~n4025;
  assign n4499 = n3671 & ~n4313;
  assign n4500 = ~n4498 & ~n4499;
  assign n4501 = n266 & ~n4326;
  assign n4502 = ~n262 & ~n3991;
  assign n4503 = ~n4501 & ~n4502;
  assign n4504 = n4500 & ~n4503;
  assign n4505 = ~n4500 & n4503;
  assign n4506 = ~n4504 & ~n4505;
  assign n4507 = n4497 & ~n4506;
  assign n4508 = ~n4497 & n4506;
  assign n4509 = ~n4507 & ~n4508;
  assign n4510 = ~n4494 & ~n4509;
  assign n4511 = n4494 & n4509;
  assign n4512 = ~n4510 & ~n4511;
  assign n4513 = ~n4492 & ~n4512;
  assign n4514 = n4494 & ~n4509;
  assign n4515 = ~n4513 & ~n4514;
  assign n4516 = n3994 & n3996;
  assign n4517 = ~n3994 & ~n3996;
  assign n4518 = ~n4516 & ~n4517;
  assign n4519 = n4013 & ~n4019;
  assign n4520 = ~n4013 & n4019;
  assign n4521 = ~n4519 & ~n4520;
  assign n4522 = n4027 & n4521;
  assign n4523 = ~n4027 & ~n4521;
  assign n4524 = ~n4522 & ~n4523;
  assign n4525 = n4500 & n4503;
  assign n4526 = ~n4497 & ~n4525;
  assign n4527 = ~n4500 & ~n4503;
  assign n4528 = ~n4526 & ~n4527;
  assign n4529 = ~n4524 & ~n4528;
  assign n4530 = n4524 & n4528;
  assign n4531 = ~n4529 & ~n4530;
  assign n4532 = ~n4518 & n4531;
  assign n4533 = n4518 & ~n4531;
  assign n4534 = ~n4532 & ~n4533;
  assign n4535 = ~n4515 & n4534;
  assign n4536 = n4515 & ~n4534;
  assign n4537 = ~n4535 & ~n4536;
  assign n4538 = ~n4441 & ~n4537;
  assign n4539 = n4441 & n4537;
  assign n4540 = ~n4538 & ~n4539;
  assign n4541 = n4492 & ~n4512;
  assign n4542 = ~n4492 & n4512;
  assign n4543 = ~n4541 & ~n4542;
  assign n4544 = ~n4343 & n4394;
  assign n4545 = n4343 & ~n4394;
  assign n4546 = ~n4544 & ~n4545;
  assign n4547 = ~g45 & g59;
  assign n4548 = g45 & ~g59;
  assign n4549 = ~n4547 & ~n4548;
  assign n4550 = n3731 & ~n4549;
  assign n4551 = ~n529 & ~n4381;
  assign n4552 = ~n4550 & ~n4551;
  assign n4553 = g66 & ~n2755;
  assign n4554 = n226 & ~n4553;
  assign n4555 = ~g47 & g58;
  assign n4556 = g47 & ~g58;
  assign n4557 = ~n4555 & ~n4556;
  assign n4558 = n2095 & ~n4557;
  assign n4559 = ~n2051 & ~n4447;
  assign n4560 = ~n4558 & ~n4559;
  assign n4561 = n4554 & ~n4560;
  assign n4562 = n4552 & n4561;
  assign n4563 = ~n4552 & ~n4561;
  assign n4564 = ~n4562 & ~n4563;
  assign n4565 = n370 & ~n4454;
  assign n4566 = ~g43 & g62;
  assign n4567 = g43 & ~g62;
  assign n4568 = ~n4566 & ~n4567;
  assign n4569 = n3671 & ~n4568;
  assign n4570 = ~n4565 & ~n4569;
  assign n4571 = ~g49 & g56;
  assign n4572 = g49 & ~g56;
  assign n4573 = ~n4571 & ~n4572;
  assign n4574 = n2295 & ~n4573;
  assign n4575 = g50 & ~n4479;
  assign n4576 = ~n4574 & ~n4575;
  assign n4577 = ~g41 & g64;
  assign n4578 = g41 & ~g64;
  assign n4579 = ~n4577 & ~n4578;
  assign n4580 = n266 & ~n4579;
  assign n4581 = ~n262 & ~n4473;
  assign n4582 = ~n4580 & ~n4581;
  assign n4583 = n4576 & ~n4582;
  assign n4584 = ~n4576 & n4582;
  assign n4585 = ~n4583 & ~n4584;
  assign n4586 = ~n4570 & ~n4585;
  assign n4587 = ~n4576 & ~n4582;
  assign n4588 = ~n4586 & ~n4587;
  assign n4589 = ~n4564 & ~n4588;
  assign n4590 = ~n4552 & n4561;
  assign n4591 = ~n4589 & ~n4590;
  assign n4592 = n4319 & ~n4340;
  assign n4593 = ~n4319 & n4340;
  assign n4594 = ~n4592 & ~n4593;
  assign n4595 = n4387 & n4389;
  assign n4596 = ~n4387 & ~n4389;
  assign n4597 = ~n4595 & ~n4596;
  assign n4598 = n4594 & ~n4597;
  assign n4599 = ~n4594 & n4597;
  assign n4600 = ~n4598 & ~n4599;
  assign n4601 = ~n4591 & ~n4600;
  assign n4602 = ~n4594 & ~n4597;
  assign n4603 = ~n4601 & ~n4602;
  assign n4604 = ~n4546 & n4603;
  assign n4605 = n4546 & ~n4603;
  assign n4606 = ~n4604 & ~n4605;
  assign n4607 = ~n4543 & ~n4606;
  assign n4608 = ~n4546 & ~n4603;
  assign n4609 = ~n4607 & ~n4608;
  assign n4610 = ~n4540 & ~n4609;
  assign n4611 = n4543 & ~n4606;
  assign n4612 = ~n4543 & n4606;
  assign n4613 = ~n4611 & ~n4612;
  assign n4614 = n4591 & n4600;
  assign n4615 = ~n4601 & ~n4614;
  assign n4616 = n4488 & n4490;
  assign n4617 = ~n4488 & ~n4490;
  assign n4618 = ~n4616 & ~n4617;
  assign n4619 = n4470 & n4485;
  assign n4620 = ~n4486 & ~n4619;
  assign n4621 = n4450 & n4460;
  assign n4622 = ~n4461 & ~n4621;
  assign n4623 = ~n175 & ~n4467;
  assign n4624 = g39 & g66;
  assign n4625 = ~g39 & ~g66;
  assign n4626 = n176 & ~n4625;
  assign n4627 = ~n4624 & n4626;
  assign n4628 = ~n4623 & ~n4627;
  assign n4629 = ~g45 & g60;
  assign n4630 = g45 & ~g60;
  assign n4631 = ~n4629 & ~n4630;
  assign n4632 = n3731 & ~n4631;
  assign n4633 = ~n529 & ~n4549;
  assign n4634 = ~n4632 & ~n4633;
  assign n4635 = ~n4628 & ~n4634;
  assign n4636 = ~n4554 & ~n4560;
  assign n4637 = n4554 & n4560;
  assign n4638 = ~n4636 & ~n4637;
  assign n4639 = n4628 & ~n4634;
  assign n4640 = ~n4628 & n4634;
  assign n4641 = ~n4639 & ~n4640;
  assign n4642 = ~n4638 & ~n4641;
  assign n4643 = ~n4635 & ~n4642;
  assign n4644 = n4622 & n4643;
  assign n4645 = ~n4622 & ~n4643;
  assign n4646 = ~n4644 & ~n4645;
  assign n4647 = n4620 & ~n4646;
  assign n4648 = n4622 & ~n4643;
  assign n4649 = ~n4647 & ~n4648;
  assign n4650 = ~n4618 & n4649;
  assign n4651 = n4618 & ~n4649;
  assign n4652 = ~n4650 & ~n4651;
  assign n4653 = n4615 & ~n4652;
  assign n4654 = ~n4618 & ~n4649;
  assign n4655 = ~n4653 & ~n4654;
  assign n4656 = n4613 & n4655;
  assign n4657 = ~n4564 & n4588;
  assign n4658 = n4564 & ~n4588;
  assign n4659 = ~n4657 & ~n4658;
  assign n4660 = n4570 & ~n4585;
  assign n4661 = ~n4570 & n4585;
  assign n4662 = ~n4660 & ~n4661;
  assign n4663 = ~n529 & ~n4631;
  assign n4664 = ~g45 & g61;
  assign n4665 = g45 & ~g61;
  assign n4666 = ~n4664 & ~n4665;
  assign n4667 = n3731 & ~n4666;
  assign n4668 = ~n4663 & ~n4667;
  assign n4669 = ~g49 & g57;
  assign n4670 = g49 & ~g57;
  assign n4671 = ~n4669 & ~n4670;
  assign n4672 = n2295 & ~n4671;
  assign n4673 = g50 & ~n4573;
  assign n4674 = ~n4672 & ~n4673;
  assign n4675 = ~g41 & g65;
  assign n4676 = g41 & ~g65;
  assign n4677 = ~n4675 & ~n4676;
  assign n4678 = n266 & ~n4677;
  assign n4679 = ~n262 & ~n4579;
  assign n4680 = ~n4678 & ~n4679;
  assign n4681 = ~n4674 & n4680;
  assign n4682 = n4674 & ~n4680;
  assign n4683 = ~n4681 & ~n4682;
  assign n4684 = ~n4668 & ~n4683;
  assign n4685 = ~n4674 & ~n4680;
  assign n4686 = ~n4684 & ~n4685;
  assign n4687 = g66 & ~n175;
  assign n4688 = ~g47 & g59;
  assign n4689 = g47 & ~g59;
  assign n4690 = ~n4688 & ~n4689;
  assign n4691 = n2095 & ~n4690;
  assign n4692 = ~n2051 & ~n4557;
  assign n4693 = ~n4691 & ~n4692;
  assign n4694 = n4687 & ~n4693;
  assign n4695 = ~n4687 & n4693;
  assign n4696 = n370 & ~n4568;
  assign n4697 = ~g43 & g63;
  assign n4698 = g43 & ~g63;
  assign n4699 = ~n4697 & ~n4698;
  assign n4700 = n3671 & ~n4699;
  assign n4701 = ~n4696 & ~n4700;
  assign n4702 = ~n4695 & ~n4701;
  assign n4703 = ~n4694 & ~n4702;
  assign n4704 = n4686 & ~n4703;
  assign n4705 = ~n4686 & n4703;
  assign n4706 = ~n4704 & ~n4705;
  assign n4707 = ~n4662 & ~n4706;
  assign n4708 = ~n4686 & ~n4703;
  assign n4709 = ~n4707 & ~n4708;
  assign n4710 = n4659 & n4709;
  assign n4711 = ~n4659 & ~n4709;
  assign n4712 = ~n4710 & ~n4711;
  assign n4713 = n4620 & n4646;
  assign n4714 = ~n4620 & ~n4646;
  assign n4715 = ~n4713 & ~n4714;
  assign n4716 = n4712 & n4715;
  assign n4717 = ~n4712 & ~n4715;
  assign n4718 = ~n4716 & ~n4717;
  assign n4719 = n4662 & ~n4706;
  assign n4720 = ~n4662 & n4706;
  assign n4721 = ~n4719 & ~n4720;
  assign n4722 = ~n4638 & n4641;
  assign n4723 = n4638 & ~n4641;
  assign n4724 = ~n4722 & ~n4723;
  assign n4725 = ~n4721 & ~n4724;
  assign n4726 = ~g66 & n266;
  assign n4727 = ~n262 & ~n4677;
  assign n4728 = ~n4726 & ~n4727;
  assign n4729 = ~g49 & g58;
  assign n4730 = g49 & ~g58;
  assign n4731 = ~n4729 & ~n4730;
  assign n4732 = n2295 & ~n4731;
  assign n4733 = g50 & ~n4671;
  assign n4734 = ~n4732 & ~n4733;
  assign n4735 = n370 & ~n4699;
  assign n4736 = ~g43 & g64;
  assign n4737 = g43 & ~g64;
  assign n4738 = ~n4736 & ~n4737;
  assign n4739 = n3671 & ~n4738;
  assign n4740 = ~n4735 & ~n4739;
  assign n4741 = ~n4734 & n4740;
  assign n4742 = n4734 & ~n4740;
  assign n4743 = ~n4741 & ~n4742;
  assign n4744 = ~n4728 & ~n4743;
  assign n4745 = ~n4734 & ~n4740;
  assign n4746 = ~n4744 & ~n4745;
  assign n4747 = ~g66 & ~n2929;
  assign n4748 = ~n2931 & ~n4747;
  assign n4749 = g41 & ~n4748;
  assign n4750 = ~g47 & g60;
  assign n4751 = g47 & ~g60;
  assign n4752 = ~n4750 & ~n4751;
  assign n4753 = n2095 & ~n4752;
  assign n4754 = ~n2051 & ~n4690;
  assign n4755 = ~n4753 & ~n4754;
  assign n4756 = n4749 & ~n4755;
  assign n4757 = ~n4694 & ~n4695;
  assign n4758 = ~n4701 & n4757;
  assign n4759 = n4701 & ~n4757;
  assign n4760 = ~n4758 & ~n4759;
  assign n4761 = ~n4756 & n4760;
  assign n4762 = n4756 & ~n4760;
  assign n4763 = ~n4761 & ~n4762;
  assign n4764 = ~n4746 & ~n4763;
  assign n4765 = n4756 & n4760;
  assign n4766 = ~n4764 & ~n4765;
  assign n4767 = n4721 & n4724;
  assign n4768 = ~n4725 & ~n4767;
  assign n4769 = ~n4766 & n4768;
  assign n4770 = ~n4725 & ~n4769;
  assign n4771 = ~n4718 & ~n4770;
  assign n4772 = n4712 & ~n4715;
  assign n4773 = ~n4711 & ~n4772;
  assign n4774 = ~n4615 & ~n4652;
  assign n4775 = n4615 & n4652;
  assign n4776 = ~n4774 & ~n4775;
  assign n4777 = n4773 & n4776;
  assign n4778 = n4771 & ~n4777;
  assign n4779 = ~n4773 & ~n4776;
  assign n4780 = ~n4778 & ~n4779;
  assign n4781 = ~n4656 & ~n4780;
  assign n4782 = ~n4613 & ~n4655;
  assign n4783 = ~n4781 & ~n4782;
  assign n4784 = n4540 & n4609;
  assign n4785 = ~n4783 & ~n4784;
  assign n4786 = ~n4746 & n4763;
  assign n4787 = n4746 & ~n4763;
  assign n4788 = ~n4786 & ~n4787;
  assign n4789 = n4668 & n4683;
  assign n4790 = ~n4684 & ~n4789;
  assign n4791 = n370 & ~n4738;
  assign n4792 = ~g43 & g65;
  assign n4793 = g43 & ~g65;
  assign n4794 = ~n4792 & ~n4793;
  assign n4795 = n3671 & ~n4794;
  assign n4796 = ~n4791 & ~n4795;
  assign n4797 = g66 & ~n262;
  assign n4798 = ~g49 & g59;
  assign n4799 = g49 & ~g59;
  assign n4800 = ~n4798 & ~n4799;
  assign n4801 = n2295 & ~n4800;
  assign n4802 = g50 & ~n4731;
  assign n4803 = ~n4801 & ~n4802;
  assign n4804 = n4797 & n4803;
  assign n4805 = ~n4797 & ~n4803;
  assign n4806 = ~n4804 & ~n4805;
  assign n4807 = ~n4796 & ~n4806;
  assign n4808 = n4797 & ~n4803;
  assign n4809 = ~n4807 & ~n4808;
  assign n4810 = ~g45 & g62;
  assign n4811 = g45 & ~g62;
  assign n4812 = ~n4810 & ~n4811;
  assign n4813 = n3731 & ~n4812;
  assign n4814 = ~n529 & ~n4666;
  assign n4815 = ~n4813 & ~n4814;
  assign n4816 = n4749 & n4755;
  assign n4817 = ~n4749 & ~n4755;
  assign n4818 = ~n4816 & ~n4817;
  assign n4819 = ~n4815 & n4818;
  assign n4820 = n4815 & ~n4818;
  assign n4821 = ~n4819 & ~n4820;
  assign n4822 = ~n4809 & ~n4821;
  assign n4823 = ~n4815 & ~n4818;
  assign n4824 = ~n4822 & ~n4823;
  assign n4825 = ~n4790 & ~n4824;
  assign n4826 = n4790 & n4824;
  assign n4827 = ~n4825 & ~n4826;
  assign n4828 = ~n4788 & ~n4827;
  assign n4829 = n4790 & ~n4824;
  assign n4830 = ~n4828 & ~n4829;
  assign n4831 = n4766 & ~n4768;
  assign n4832 = ~n4769 & ~n4831;
  assign n4833 = n4830 & ~n4832;
  assign n4834 = ~n4830 & n4832;
  assign n4835 = ~g47 & g62;
  assign n4836 = g47 & ~g62;
  assign n4837 = ~n4835 & ~n4836;
  assign n4838 = n2095 & ~n4837;
  assign n4839 = ~g47 & g61;
  assign n4840 = g47 & ~g61;
  assign n4841 = ~n4839 & ~n4840;
  assign n4842 = ~n2051 & ~n4841;
  assign n4843 = ~n4838 & ~n4842;
  assign n4844 = ~g45 & g64;
  assign n4845 = g45 & ~g64;
  assign n4846 = ~n4844 & ~n4845;
  assign n4847 = n3731 & ~n4846;
  assign n4848 = ~g45 & ~g63;
  assign n4849 = g45 & g63;
  assign n4850 = ~n4848 & ~n4849;
  assign n4851 = ~n529 & n4850;
  assign n4852 = ~n4847 & ~n4851;
  assign n4853 = ~n4843 & ~n4852;
  assign n4854 = n370 & ~n4794;
  assign n4855 = g43 & g66;
  assign n4856 = ~g43 & ~g66;
  assign n4857 = n3671 & ~n4856;
  assign n4858 = ~n4855 & n4857;
  assign n4859 = ~n4854 & ~n4858;
  assign n4860 = n4843 & n4852;
  assign n4861 = ~n4853 & ~n4860;
  assign n4862 = ~n4859 & n4861;
  assign n4863 = ~n4853 & ~n4862;
  assign n4864 = n4796 & ~n4806;
  assign n4865 = ~n4796 & n4806;
  assign n4866 = ~n4864 & ~n4865;
  assign n4867 = ~n4863 & ~n4866;
  assign n4868 = ~g49 & g60;
  assign n4869 = g49 & ~g60;
  assign n4870 = ~n4868 & ~n4869;
  assign n4871 = n2295 & ~n4870;
  assign n4872 = g50 & ~n4800;
  assign n4873 = ~n4871 & ~n4872;
  assign n4874 = g66 & ~n3042;
  assign n4875 = n376 & ~n4874;
  assign n4876 = ~n4873 & n4875;
  assign n4877 = n2095 & ~n4841;
  assign n4878 = ~n2051 & ~n4752;
  assign n4879 = ~n4877 & ~n4878;
  assign n4880 = ~n4876 & ~n4879;
  assign n4881 = n4876 & n4879;
  assign n4882 = ~n4880 & ~n4881;
  assign n4883 = n3731 & n4850;
  assign n4884 = ~n529 & ~n4812;
  assign n4885 = ~n4883 & ~n4884;
  assign n4886 = ~n4882 & ~n4885;
  assign n4887 = n4882 & n4885;
  assign n4888 = ~n4886 & ~n4887;
  assign n4889 = n4863 & n4866;
  assign n4890 = ~n4867 & ~n4889;
  assign n4891 = n4888 & n4890;
  assign n4892 = ~n4867 & ~n4891;
  assign n4893 = n4809 & n4821;
  assign n4894 = ~n4822 & ~n4893;
  assign n4895 = n4876 & ~n4879;
  assign n4896 = ~n4886 & ~n4895;
  assign n4897 = ~n4728 & n4743;
  assign n4898 = n4728 & ~n4743;
  assign n4899 = ~n4897 & ~n4898;
  assign n4900 = n4896 & ~n4899;
  assign n4901 = ~n4896 & n4899;
  assign n4902 = ~n4900 & ~n4901;
  assign n4903 = ~n4894 & ~n4902;
  assign n4904 = n4894 & n4902;
  assign n4905 = ~n4903 & ~n4904;
  assign n4906 = ~n4892 & ~n4905;
  assign n4907 = n4859 & n4861;
  assign n4908 = ~n4859 & ~n4861;
  assign n4909 = ~n4907 & ~n4908;
  assign n4910 = ~n4873 & ~n4875;
  assign n4911 = n4873 & n4875;
  assign n4912 = ~n4910 & ~n4911;
  assign n4913 = g66 & n370;
  assign n4914 = ~g49 & g61;
  assign n4915 = g49 & ~g61;
  assign n4916 = ~n4914 & ~n4915;
  assign n4917 = n2295 & ~n4916;
  assign n4918 = g50 & ~n4870;
  assign n4919 = ~n4917 & ~n4918;
  assign n4920 = n4913 & ~n4919;
  assign n4921 = ~g47 & g63;
  assign n4922 = g47 & ~g63;
  assign n4923 = ~n4921 & ~n4922;
  assign n4924 = n2095 & ~n4923;
  assign n4925 = ~n2051 & ~n4837;
  assign n4926 = ~n4924 & ~n4925;
  assign n4927 = ~n4913 & n4919;
  assign n4928 = ~n4920 & ~n4927;
  assign n4929 = ~n4926 & n4928;
  assign n4930 = ~n4920 & ~n4929;
  assign n4931 = n4912 & ~n4930;
  assign n4932 = ~n4912 & n4930;
  assign n4933 = ~n4931 & ~n4932;
  assign n4934 = ~n4909 & ~n4933;
  assign n4935 = ~n4912 & ~n4930;
  assign n4936 = ~n4934 & ~n4935;
  assign n4937 = n4888 & ~n4890;
  assign n4938 = ~n4888 & n4890;
  assign n4939 = ~n4937 & ~n4938;
  assign n4940 = ~n4936 & ~n4939;
  assign n4941 = ~n4906 & ~n4940;
  assign n4942 = n4892 & n4905;
  assign n4943 = ~n4941 & ~n4942;
  assign n4944 = ~n4788 & n4827;
  assign n4945 = n4788 & ~n4827;
  assign n4946 = ~n4944 & ~n4945;
  assign n4947 = n4894 & ~n4902;
  assign n4948 = ~n4896 & ~n4899;
  assign n4949 = ~n4947 & ~n4948;
  assign n4950 = n4946 & n4949;
  assign n4951 = n4943 & ~n4950;
  assign n4952 = ~n4946 & ~n4949;
  assign n4953 = ~n4951 & ~n4952;
  assign n4954 = ~n4834 & n4953;
  assign n4955 = ~n4833 & ~n4954;
  assign n4956 = g66 & ~n3154;
  assign n4957 = n617 & ~n4956;
  assign n4958 = ~g49 & g62;
  assign n4959 = g49 & ~g62;
  assign n4960 = ~n4958 & ~n4959;
  assign n4961 = n2295 & ~n4960;
  assign n4962 = g50 & ~n4916;
  assign n4963 = ~n4961 & ~n4962;
  assign n4964 = n4957 & ~n4963;
  assign n4965 = ~n529 & ~n4846;
  assign n4966 = ~g45 & g65;
  assign n4967 = g45 & ~g65;
  assign n4968 = ~n4966 & ~n4967;
  assign n4969 = n3731 & ~n4968;
  assign n4970 = ~n4965 & ~n4969;
  assign n4971 = ~n4964 & ~n4970;
  assign n4972 = n4926 & ~n4928;
  assign n4973 = ~n4929 & ~n4972;
  assign n4974 = n4964 & ~n4970;
  assign n4975 = ~n4964 & n4970;
  assign n4976 = ~n4974 & ~n4975;
  assign n4977 = n4973 & ~n4976;
  assign n4978 = ~n4971 & ~n4977;
  assign n4979 = n4909 & ~n4933;
  assign n4980 = ~n4909 & n4933;
  assign n4981 = ~n4979 & ~n4980;
  assign n4982 = n4978 & n4981;
  assign n4983 = ~n529 & ~n4968;
  assign n4984 = ~g45 & g66;
  assign n4985 = g45 & ~g66;
  assign n4986 = ~n4984 & ~n4985;
  assign n4987 = n3731 & ~n4986;
  assign n4988 = ~n4983 & ~n4987;
  assign n4989 = ~g47 & g64;
  assign n4990 = g47 & ~g64;
  assign n4991 = ~n4989 & ~n4990;
  assign n4992 = n2095 & ~n4991;
  assign n4993 = ~n2051 & ~n4923;
  assign n4994 = ~n4992 & ~n4993;
  assign n4995 = ~n4988 & ~n4994;
  assign n4996 = ~n4957 & ~n4963;
  assign n4997 = n4957 & n4963;
  assign n4998 = ~n4996 & ~n4997;
  assign n4999 = n4988 & n4994;
  assign n5000 = ~n4995 & ~n4999;
  assign n5001 = ~n4998 & n5000;
  assign n5002 = ~n4995 & ~n5001;
  assign n5003 = ~n4973 & ~n4976;
  assign n5004 = n4973 & n4976;
  assign n5005 = ~n5003 & ~n5004;
  assign n5006 = n5002 & ~n5005;
  assign n5007 = ~g66 & ~n3222;
  assign n5008 = ~n3224 & ~n5007;
  assign n5009 = g47 & ~n5008;
  assign n5010 = ~g49 & g64;
  assign n5011 = g49 & ~g64;
  assign n5012 = ~n5010 & ~n5011;
  assign n5013 = n2295 & ~n5012;
  assign n5014 = ~g49 & g63;
  assign n5015 = g49 & ~g63;
  assign n5016 = ~n5014 & ~n5015;
  assign n5017 = g50 & ~n5016;
  assign n5018 = ~n5013 & ~n5017;
  assign n5019 = n5009 & ~n5018;
  assign n5020 = ~g47 & g65;
  assign n5021 = g47 & ~g65;
  assign n5022 = ~n5020 & ~n5021;
  assign n5023 = n2095 & ~n5022;
  assign n5024 = ~n2051 & ~n4991;
  assign n5025 = ~n5023 & ~n5024;
  assign n5026 = g66 & ~n529;
  assign n5027 = n2295 & ~n5016;
  assign n5028 = g50 & ~n4960;
  assign n5029 = ~n5027 & ~n5028;
  assign n5030 = n5026 & n5029;
  assign n5031 = ~n5026 & ~n5029;
  assign n5032 = ~n5030 & ~n5031;
  assign n5033 = n5025 & ~n5032;
  assign n5034 = ~n5025 & n5032;
  assign n5035 = ~n5033 & ~n5034;
  assign n5036 = ~n5019 & n5035;
  assign n5037 = g49 & g66;
  assign n5038 = g66 & ~n2051;
  assign n5039 = ~g49 & g65;
  assign n5040 = g49 & ~g65;
  assign n5041 = ~n5039 & ~n5040;
  assign n5042 = n2295 & ~n5041;
  assign n5043 = g50 & ~n5012;
  assign n5044 = ~n5042 & ~n5043;
  assign n5045 = ~n5038 & n5044;
  assign n5046 = ~n2295 & n5041;
  assign n5047 = ~n5045 & ~n5046;
  assign n5048 = n5037 & n5047;
  assign n5049 = n5038 & ~n5044;
  assign n5050 = ~n5048 & ~n5049;
  assign n5051 = ~n5009 & ~n5018;
  assign n5052 = n5009 & n5018;
  assign n5053 = ~n5051 & ~n5052;
  assign n5054 = ~g66 & n2095;
  assign n5055 = ~n2051 & ~n5022;
  assign n5056 = ~n5054 & ~n5055;
  assign n5057 = n5053 & n5056;
  assign n5058 = ~n5050 & ~n5057;
  assign n5059 = ~n5053 & ~n5056;
  assign n5060 = ~n5058 & ~n5059;
  assign n5061 = ~n5036 & ~n5060;
  assign n5062 = n5019 & ~n5035;
  assign n5063 = ~n5061 & ~n5062;
  assign n5064 = ~n5025 & ~n5032;
  assign n5065 = n5026 & ~n5029;
  assign n5066 = ~n5064 & ~n5065;
  assign n5067 = ~n4998 & ~n5000;
  assign n5068 = n4998 & n5000;
  assign n5069 = ~n5067 & ~n5068;
  assign n5070 = n5066 & ~n5069;
  assign n5071 = ~n5066 & n5069;
  assign n5072 = ~n5070 & ~n5071;
  assign n5073 = ~n5063 & ~n5072;
  assign n5074 = ~n5066 & ~n5069;
  assign n5075 = ~n5073 & ~n5074;
  assign n5076 = ~n5006 & ~n5075;
  assign n5077 = ~n5002 & n5005;
  assign n5078 = ~n5076 & ~n5077;
  assign n5079 = ~n4982 & ~n5078;
  assign n5080 = ~n4978 & ~n4981;
  assign n5081 = ~n5079 & ~n5080;
  assign n5082 = ~n4950 & ~n5081;
  assign n5083 = n4936 & n4939;
  assign n5084 = ~n4942 & ~n5083;
  assign n5085 = n5082 & n5084;
  assign n5086 = ~n4833 & n5085;
  assign n5087 = ~n4955 & ~n5086;
  assign n5088 = n4718 & n4770;
  assign n5089 = ~n4777 & ~n5088;
  assign n5090 = ~n4656 & n5089;
  assign n5091 = ~n4784 & n5090;
  assign n5092 = ~n5087 & n5091;
  assign n5093 = ~n4785 & ~n5092;
  assign n5094 = ~n4610 & n5093;
  assign n5095 = ~n4183 & ~n4228;
  assign n5096 = ~n4172 & ~n4180;
  assign n5097 = ~n5095 & ~n5096;
  assign n5098 = n4156 & ~n4169;
  assign n5099 = n4157 & ~n4166;
  assign n5100 = ~n5098 & ~n5099;
  assign n5101 = n266 & ~n4154;
  assign n5102 = ~n262 & n3596;
  assign n5103 = ~n5101 & ~n5102;
  assign n5104 = ~n370 & ~n3671;
  assign n5105 = g43 & ~n5104;
  assign n5106 = n107 & ~n4264;
  assign n5107 = ~g37 & ~g55;
  assign n5108 = g37 & g55;
  assign n5109 = ~n5107 & ~n5108;
  assign n5110 = ~n103 & n5109;
  assign n5111 = ~n5106 & ~n5110;
  assign n5112 = n5105 & ~n5111;
  assign n5113 = ~n5105 & n5111;
  assign n5114 = ~n5112 & ~n5113;
  assign n5115 = n5103 & ~n5114;
  assign n5116 = ~n5103 & n5114;
  assign n5117 = ~n5115 & ~n5116;
  assign n5118 = ~n5100 & n5117;
  assign n5119 = n5100 & ~n5117;
  assign n5120 = ~n5118 & ~n5119;
  assign n5121 = n123 & ~n4255;
  assign n5122 = ~n119 & ~n3589;
  assign n5123 = ~n5121 & ~n5122;
  assign n5124 = g35 & g59;
  assign n5125 = n176 & n4164;
  assign n5126 = ~n175 & ~n3606;
  assign n5127 = ~n5125 & ~n5126;
  assign n5128 = ~n5124 & ~n5127;
  assign n5129 = n5124 & n5127;
  assign n5130 = ~n5128 & ~n5129;
  assign n5131 = n5123 & ~n5130;
  assign n5132 = ~n5123 & n5130;
  assign n5133 = ~n5131 & ~n5132;
  assign n5134 = ~n4257 & ~n4260;
  assign n5135 = n4257 & n4260;
  assign n5136 = ~n4266 & ~n5135;
  assign n5137 = ~n5134 & ~n5136;
  assign n5138 = ~n4156 & n5137;
  assign n5139 = n4156 & ~n5137;
  assign n5140 = ~n5138 & ~n5139;
  assign n5141 = n5133 & ~n5140;
  assign n5142 = ~n5133 & n5140;
  assign n5143 = ~n5141 & ~n5142;
  assign n5144 = ~n5120 & n5143;
  assign n5145 = n5120 & ~n5143;
  assign n5146 = ~n5144 & ~n5145;
  assign n5147 = ~n4275 & ~n4277;
  assign n5148 = ~n4251 & ~n4272;
  assign n5149 = ~n5147 & ~n5148;
  assign n5150 = ~n5146 & n5149;
  assign n5151 = n5146 & ~n5149;
  assign n5152 = ~n5150 & ~n5151;
  assign n5153 = n5097 & ~n5152;
  assign n5154 = ~n5097 & n5152;
  assign n5155 = ~n5153 & ~n5154;
  assign n5156 = ~n4231 & ~n4283;
  assign n5157 = ~n4248 & ~n4280;
  assign n5158 = ~n5156 & ~n5157;
  assign n5159 = n5155 & n5158;
  assign n5160 = n4050 & n4052;
  assign n5161 = ~n4050 & ~n4052;
  assign n5162 = ~n5160 & ~n5161;
  assign n5163 = ~n3764 & n3818;
  assign n5164 = n3764 & ~n3818;
  assign n5165 = ~n5163 & ~n5164;
  assign n5166 = n3970 & ~n3972;
  assign n5167 = ~n3973 & ~n5166;
  assign n5168 = n3736 & ~n3757;
  assign n5169 = ~n3736 & n3757;
  assign n5170 = ~n5168 & ~n5169;
  assign n5171 = n3712 & ~n3721;
  assign n5172 = ~n3712 & n3721;
  assign n5173 = ~n5171 & ~n5172;
  assign n5174 = ~n3699 & ~n3701;
  assign n5175 = n3699 & n3701;
  assign n5176 = ~n5174 & ~n5175;
  assign n5177 = n5173 & n5176;
  assign n5178 = ~n5170 & ~n5177;
  assign n5179 = ~n5173 & ~n5176;
  assign n5180 = ~n5178 & ~n5179;
  assign n5181 = n5167 & ~n5180;
  assign n5182 = n3760 & ~n3762;
  assign n5183 = ~n3763 & ~n5182;
  assign n5184 = ~n5167 & n5180;
  assign n5185 = ~n5181 & ~n5184;
  assign n5186 = n5183 & n5185;
  assign n5187 = ~n5181 & ~n5186;
  assign n5188 = n5165 & ~n5187;
  assign n5189 = ~n5165 & n5187;
  assign n5190 = ~n5188 & ~n5189;
  assign n5191 = ~n5162 & ~n5190;
  assign n5192 = ~n5165 & ~n5187;
  assign n5193 = ~n5191 & ~n5192;
  assign n5194 = n3915 & ~n4057;
  assign n5195 = ~n3915 & n4057;
  assign n5196 = ~n5194 & ~n5195;
  assign n5197 = n5193 & n5196;
  assign n5198 = ~n4035 & n4047;
  assign n5199 = n4035 & ~n4047;
  assign n5200 = ~n5198 & ~n5199;
  assign n5201 = n5183 & ~n5185;
  assign n5202 = ~n5183 & n5185;
  assign n5203 = ~n5201 & ~n5202;
  assign n5204 = ~n5200 & ~n5203;
  assign n5205 = ~n4518 & ~n4531;
  assign n5206 = n4524 & ~n4528;
  assign n5207 = ~n5205 & ~n5206;
  assign n5208 = ~n4403 & n4405;
  assign n5209 = ~n4412 & ~n5208;
  assign n5210 = n3998 & ~n4032;
  assign n5211 = ~n3998 & n4032;
  assign n5212 = ~n5210 & ~n5211;
  assign n5213 = n5209 & ~n5212;
  assign n5214 = ~n5209 & n5212;
  assign n5215 = ~n5213 & ~n5214;
  assign n5216 = ~n5207 & ~n5215;
  assign n5217 = ~n5209 & ~n5212;
  assign n5218 = ~n5216 & ~n5217;
  assign n5219 = n5200 & n5203;
  assign n5220 = ~n5204 & ~n5219;
  assign n5221 = ~n5218 & n5220;
  assign n5222 = ~n5204 & ~n5221;
  assign n5223 = n5162 & ~n5190;
  assign n5224 = ~n5162 & n5190;
  assign n5225 = ~n5223 & ~n5224;
  assign n5226 = n5222 & n5225;
  assign n5227 = ~n5197 & ~n5226;
  assign n5228 = n5207 & ~n5215;
  assign n5229 = ~n5207 & n5215;
  assign n5230 = ~n5228 & ~n5229;
  assign n5231 = ~n5170 & n5179;
  assign n5232 = ~n5170 & n5173;
  assign n5233 = n5176 & n5232;
  assign n5234 = ~n5231 & ~n5233;
  assign n5235 = ~n5177 & ~n5179;
  assign n5236 = n5170 & n5235;
  assign n5237 = n5234 & ~n5236;
  assign n5238 = n4414 & ~n4435;
  assign n5239 = ~n4439 & ~n5238;
  assign n5240 = ~n5237 & n5239;
  assign n5241 = n5237 & ~n5239;
  assign n5242 = ~n5240 & ~n5241;
  assign n5243 = ~n5230 & ~n5242;
  assign n5244 = ~n5237 & ~n5239;
  assign n5245 = ~n5243 & ~n5244;
  assign n5246 = ~n5218 & ~n5220;
  assign n5247 = n5218 & n5220;
  assign n5248 = ~n5246 & ~n5247;
  assign n5249 = n5245 & n5248;
  assign n5250 = n4441 & ~n4537;
  assign n5251 = ~n4515 & ~n4534;
  assign n5252 = ~n5250 & ~n5251;
  assign n5253 = ~n5230 & n5242;
  assign n5254 = n5230 & ~n5242;
  assign n5255 = ~n5253 & ~n5254;
  assign n5256 = n5252 & n5255;
  assign n5257 = ~n5249 & ~n5256;
  assign n5258 = n5227 & n5257;
  assign n5259 = ~n5159 & n5258;
  assign n5260 = ~n5094 & n5259;
  assign n5261 = n4310 & n5260;
  assign n5262 = ~n4301 & ~n5197;
  assign n5263 = ~n5159 & n5262;
  assign n5264 = ~n5193 & ~n5196;
  assign n5265 = ~n5222 & ~n5225;
  assign n5266 = ~n5264 & ~n5265;
  assign n5267 = ~n5252 & ~n5255;
  assign n5268 = ~n5249 & n5267;
  assign n5269 = ~n5245 & ~n5248;
  assign n5270 = ~n5268 & ~n5269;
  assign n5271 = ~n5226 & ~n5270;
  assign n5272 = n5266 & ~n5271;
  assign n5273 = ~n4147 & ~n4308;
  assign n5274 = ~n5272 & n5273;
  assign n5275 = n5263 & n5274;
  assign n5276 = ~n4304 & ~n4307;
  assign n5277 = ~n4060 & ~n4146;
  assign n5278 = ~n4308 & n5277;
  assign n5279 = ~n5276 & ~n5278;
  assign n5280 = ~n4286 & ~n4300;
  assign n5281 = n5279 & ~n5280;
  assign n5282 = ~n4301 & ~n5159;
  assign n5283 = ~n5281 & n5282;
  assign n5284 = ~n5155 & ~n5158;
  assign n5285 = ~n5283 & ~n5284;
  assign n5286 = ~n5275 & n5285;
  assign n5287 = ~n5261 & n5286;
  assign n5288 = n3630 & ~n3637;
  assign n5289 = ~n3630 & n3637;
  assign n5290 = ~n5288 & ~n5289;
  assign n5291 = ~n5123 & ~n5130;
  assign n5292 = n5124 & ~n5127;
  assign n5293 = ~n5291 & ~n5292;
  assign n5294 = ~n103 & n3613;
  assign n5295 = n107 & n5109;
  assign n5296 = ~n5294 & ~n5295;
  assign n5297 = n3609 & n5296;
  assign n5298 = ~n3609 & ~n5296;
  assign n5299 = ~n5297 & ~n5298;
  assign n5300 = ~n5293 & ~n5299;
  assign n5301 = n3609 & ~n5296;
  assign n5302 = ~n5300 & ~n5301;
  assign n5303 = ~n3626 & ~n3628;
  assign n5304 = n3626 & n3628;
  assign n5305 = ~n5303 & ~n5304;
  assign n5306 = ~n5302 & ~n5305;
  assign n5307 = ~n5302 & n5305;
  assign n5308 = n5302 & ~n5305;
  assign n5309 = ~n5307 & ~n5308;
  assign n5310 = ~n5103 & ~n5114;
  assign n5311 = ~n5105 & ~n5111;
  assign n5312 = ~n5310 & ~n5311;
  assign n5313 = n3598 & ~n3601;
  assign n5314 = ~n3598 & n3601;
  assign n5315 = ~n5313 & ~n5314;
  assign n5316 = n5312 & ~n5315;
  assign n5317 = ~n5312 & n5315;
  assign n5318 = ~n5316 & ~n5317;
  assign n5319 = n5293 & ~n5299;
  assign n5320 = ~n5293 & n5299;
  assign n5321 = ~n5319 & ~n5320;
  assign n5322 = ~n5318 & ~n5321;
  assign n5323 = ~n5312 & ~n5315;
  assign n5324 = ~n5322 & ~n5323;
  assign n5325 = ~n5309 & ~n5324;
  assign n5326 = ~n5306 & ~n5325;
  assign n5327 = n5290 & n5326;
  assign n5328 = n5309 & ~n5324;
  assign n5329 = ~n5309 & n5324;
  assign n5330 = ~n5328 & ~n5329;
  assign n5331 = ~n5318 & n5321;
  assign n5332 = n5318 & ~n5321;
  assign n5333 = ~n5331 & ~n5332;
  assign n5334 = ~n5133 & ~n5140;
  assign n5335 = ~n4156 & ~n5137;
  assign n5336 = ~n5334 & ~n5335;
  assign n5337 = n5333 & ~n5336;
  assign n5338 = ~n5333 & n5336;
  assign n5339 = ~n5337 & ~n5338;
  assign n5340 = ~n5100 & ~n5117;
  assign n5341 = ~n5120 & ~n5143;
  assign n5342 = ~n5340 & ~n5341;
  assign n5343 = ~n5339 & ~n5342;
  assign n5344 = ~n5333 & ~n5336;
  assign n5345 = ~n5343 & ~n5344;
  assign n5346 = n5330 & n5345;
  assign n5347 = ~n5339 & n5342;
  assign n5348 = n5339 & ~n5342;
  assign n5349 = ~n5347 & ~n5348;
  assign n5350 = ~n5097 & ~n5152;
  assign n5351 = ~n5146 & ~n5149;
  assign n5352 = ~n5350 & ~n5351;
  assign n5353 = n5349 & n5352;
  assign n5354 = ~n5346 & ~n5353;
  assign n5355 = ~n5327 & n5354;
  assign n5356 = ~n5287 & n5355;
  assign n5357 = ~n3670 & n5356;
  assign n5358 = ~n3641 & n5357;
  assign n5359 = ~n5349 & ~n5352;
  assign n5360 = ~n5346 & n5359;
  assign n5361 = ~n5330 & ~n5345;
  assign n5362 = ~n5360 & ~n5361;
  assign n5363 = ~n5327 & ~n5362;
  assign n5364 = ~n5290 & ~n5326;
  assign n5365 = ~n5363 & ~n5364;
  assign n5366 = ~n3641 & ~n5365;
  assign n5367 = ~n3585 & ~n3640;
  assign n5368 = ~n5366 & ~n5367;
  assign n5369 = ~n3670 & ~n5368;
  assign n5370 = ~n3666 & ~n3669;
  assign n5371 = ~n5369 & ~n5370;
  assign n5372 = ~n5358 & n5371;
  assign n5373 = ~n3652 & n3654;
  assign n5374 = n3537 & ~n3649;
  assign n5375 = ~n5373 & ~n5374;
  assign n5376 = ~n3654 & n5375;
  assign n5377 = n3654 & ~n5375;
  assign n5378 = ~n5376 & ~n5377;
  assign n5379 = n123 & n3647;
  assign n5380 = ~g35 & ~g51;
  assign n5381 = g35 & g51;
  assign n5382 = ~n5380 & ~n5381;
  assign n5383 = ~n119 & n5382;
  assign n5384 = ~n5379 & ~n5383;
  assign n5385 = n160 & n3555;
  assign n5386 = ~n160 & ~n3555;
  assign n5387 = ~n5385 & ~n5386;
  assign n5388 = n5384 & ~n5387;
  assign n5389 = ~n5384 & n5387;
  assign n5390 = ~n5388 & ~n5389;
  assign n5391 = ~n5378 & n5390;
  assign n5392 = n5378 & ~n5390;
  assign n5393 = ~n5391 & ~n5392;
  assign n5394 = ~n3643 & ~n3663;
  assign n5395 = ~n3657 & ~n3660;
  assign n5396 = ~n5394 & ~n5395;
  assign n5397 = ~n5393 & ~n5396;
  assign n5398 = n5393 & n5396;
  assign n5399 = ~n5397 & ~n5398;
  assign n5400 = n5372 & n5399;
  assign n5401 = ~n5372 & ~n5399;
  assign n5402 = ~n5400 & ~n5401;
  assign n5403 = ~g1 & ~n5402;
  assign n5404 = ~n3499 & ~n5403;
  assign n5405 = ~n157 & ~n163;
  assign n5406 = n158 & ~n160;
  assign n5407 = ~n5405 & ~n5406;
  assign n5408 = n123 & n155;
  assign n5409 = g35 & ~n119;
  assign n5410 = ~n5408 & ~n5409;
  assign n5411 = ~n135 & ~n5410;
  assign n5412 = n135 & n5410;
  assign n5413 = ~n5411 & ~n5412;
  assign n5414 = n5407 & n5413;
  assign n5415 = ~n5407 & ~n5413;
  assign n5416 = ~n5414 & ~n5415;
  assign n5417 = ~n151 & ~n166;
  assign n5418 = ~n116 & ~n148;
  assign n5419 = ~n5417 & ~n5418;
  assign n5420 = ~n5416 & ~n5419;
  assign n5421 = n5416 & n5419;
  assign n5422 = ~n5420 & ~n5421;
  assign n5423 = ~n243 & ~n3495;
  assign n5424 = ~n242 & ~n5423;
  assign n5425 = n5422 & ~n5424;
  assign n5426 = g1 & ~n5425;
  assign n5427 = ~n5422 & n5424;
  assign n5428 = n5426 & ~n5427;
  assign n5429 = n123 & n5382;
  assign n5430 = ~n5409 & ~n5429;
  assign n5431 = ~n3646 & n5430;
  assign n5432 = n3646 & ~n5430;
  assign n5433 = ~n5431 & ~n5432;
  assign n5434 = ~n5384 & ~n5387;
  assign n5435 = ~n160 & n3555;
  assign n5436 = ~n5434 & ~n5435;
  assign n5437 = ~n5433 & n5436;
  assign n5438 = n5433 & ~n5436;
  assign n5439 = ~n5437 & ~n5438;
  assign n5440 = ~n5378 & ~n5390;
  assign n5441 = ~n3654 & ~n5375;
  assign n5442 = ~n5440 & ~n5441;
  assign n5443 = ~n5439 & ~n5442;
  assign n5444 = n5439 & n5442;
  assign n5445 = ~n5443 & ~n5444;
  assign n5446 = ~n5372 & ~n5398;
  assign n5447 = ~n5397 & ~n5446;
  assign n5448 = ~n5445 & ~n5447;
  assign n5449 = n5445 & n5447;
  assign n5450 = ~n5448 & ~n5449;
  assign n5451 = ~g1 & ~n5450;
  assign n5452 = ~n5428 & ~n5451;
  assign n5453 = n5404 & ~n5452;
  assign n5454 = n690 & ~n3490;
  assign n5455 = ~n361 & n5454;
  assign n5456 = n685 & ~n5455;
  assign n5457 = ~n296 & ~n687;
  assign n5458 = ~n5456 & n5457;
  assign n5459 = n5456 & ~n5457;
  assign n5460 = ~n5458 & ~n5459;
  assign n5461 = g1 & n5460;
  assign n5462 = ~n3670 & ~n5370;
  assign n5463 = ~n3641 & n5356;
  assign n5464 = ~n5462 & ~n5463;
  assign n5465 = n5368 & n5464;
  assign n5466 = n5368 & ~n5463;
  assign n5467 = n5462 & ~n5466;
  assign n5468 = ~g1 & ~n5467;
  assign n5469 = ~n5465 & n5468;
  assign n5470 = ~n5461 & ~n5469;
  assign n5471 = n5404 & ~n5470;
  assign n5472 = ~n5453 & n5471;
  assign n5473 = ~n5404 & n5452;
  assign n5474 = ~n5404 & n5470;
  assign n5475 = ~n5453 & ~n5474;
  assign n5476 = n682 & ~n5454;
  assign n5477 = ~n361 & ~n684;
  assign n5478 = ~n5476 & n5477;
  assign n5479 = n5476 & ~n5477;
  assign n5480 = ~n5478 & ~n5479;
  assign n5481 = g1 & n5480;
  assign n5482 = ~n3641 & ~n5367;
  assign n5483 = n5365 & n5482;
  assign n5484 = ~n5356 & n5365;
  assign n5485 = ~n5483 & n5484;
  assign n5486 = ~n5356 & n5483;
  assign n5487 = n5482 & ~n5486;
  assign n5488 = ~g1 & ~n5487;
  assign n5489 = ~n5485 & n5488;
  assign n5490 = ~n5481 & ~n5489;
  assign n5491 = ~n5470 & n5490;
  assign n5492 = n689 & ~n3490;
  assign n5493 = ~n445 & ~n681;
  assign n5494 = g1 & n5493;
  assign n5495 = ~n5492 & n5494;
  assign n5496 = n679 & n5495;
  assign n5497 = ~n5327 & ~n5364;
  assign n5498 = ~n5287 & n5354;
  assign n5499 = ~n5497 & ~n5498;
  assign n5500 = n5362 & n5499;
  assign n5501 = n5362 & ~n5498;
  assign n5502 = n5497 & ~n5501;
  assign n5503 = ~g1 & ~n5502;
  assign n5504 = ~n5500 & n5503;
  assign n5505 = n679 & ~n5492;
  assign n5506 = g1 & ~n5493;
  assign n5507 = ~n5505 & n5506;
  assign n5508 = ~n5504 & ~n5507;
  assign n5509 = ~n5496 & n5508;
  assign n5510 = n5490 & ~n5509;
  assign n5511 = ~n5491 & n5510;
  assign n5512 = n5470 & ~n5490;
  assign n5513 = ~n5511 & ~n5512;
  assign n5514 = n5475 & ~n5513;
  assign n5515 = ~n5473 & ~n5514;
  assign n5516 = ~n5472 & n5515;
  assign n5517 = ~n688 & ~n3490;
  assign n5518 = ~n677 & ~n5517;
  assign n5519 = ~n522 & ~n523;
  assign n5520 = g1 & ~n5519;
  assign n5521 = ~n5518 & n5520;
  assign n5522 = ~n5287 & ~n5353;
  assign n5523 = ~n5359 & ~n5522;
  assign n5524 = ~n5346 & ~n5361;
  assign n5525 = ~g1 & ~n5524;
  assign n5526 = ~n5523 & n5525;
  assign n5527 = ~n5521 & ~n5526;
  assign n5528 = ~g1 & n5523;
  assign n5529 = n5524 & n5528;
  assign n5530 = g1 & ~n5517;
  assign n5531 = n5519 & n5530;
  assign n5532 = ~n677 & n5531;
  assign n5533 = ~n5529 & ~n5532;
  assign n5534 = n5527 & n5533;
  assign n5535 = n5509 & ~n5534;
  assign n5536 = ~n5353 & ~n5359;
  assign n5537 = ~n5287 & n5536;
  assign n5538 = n5287 & ~n5536;
  assign n5539 = ~n5537 & ~n5538;
  assign n5540 = ~g1 & n5539;
  assign n5541 = ~n677 & ~n688;
  assign n5542 = n3490 & ~n5541;
  assign n5543 = ~n3490 & n5541;
  assign n5544 = g1 & ~n5543;
  assign n5545 = ~n5542 & n5544;
  assign n5546 = ~n5540 & ~n5545;
  assign n5547 = ~n5534 & n5546;
  assign n5548 = ~n5509 & n5534;
  assign n5549 = ~n5547 & ~n5548;
  assign n5550 = ~n3340 & n3442;
  assign n5551 = n2483 & ~n5550;
  assign n5552 = ~n3451 & ~n5551;
  assign n5553 = ~n3470 & ~n5552;
  assign n5554 = g1 & ~n5553;
  assign n5555 = ~n5094 & n5258;
  assign n5556 = ~n5265 & ~n5271;
  assign n5557 = ~n5197 & ~n5556;
  assign n5558 = ~n5264 & ~n5557;
  assign n5559 = ~n5555 & n5558;
  assign n5560 = n5273 & ~n5559;
  assign n5561 = n5279 & ~n5560;
  assign n5562 = ~n4301 & ~n5280;
  assign n5563 = ~n5561 & n5562;
  assign n5564 = n5561 & ~n5562;
  assign n5565 = ~g1 & ~n5564;
  assign n5566 = ~n5563 & n5565;
  assign n5567 = ~n5554 & ~n5566;
  assign n5568 = ~n3437 & ~n3487;
  assign n5569 = ~n3346 & n5568;
  assign n5570 = n3346 & ~n5568;
  assign n5571 = ~n5569 & ~n5570;
  assign n5572 = g1 & n5571;
  assign n5573 = ~n4301 & ~n5279;
  assign n5574 = ~n5280 & ~n5573;
  assign n5575 = ~n5159 & ~n5284;
  assign n5576 = n4310 & ~n5559;
  assign n5577 = ~n5575 & ~n5576;
  assign n5578 = n5574 & n5577;
  assign n5579 = n5574 & ~n5576;
  assign n5580 = n5575 & ~n5579;
  assign n5581 = ~g1 & ~n5580;
  assign n5582 = ~n5578 & n5581;
  assign n5583 = ~n5572 & ~n5582;
  assign n5584 = n5567 & n5583;
  assign n5585 = n5546 & ~n5584;
  assign n5586 = n5549 & n5585;
  assign n5587 = n5527 & ~n5546;
  assign n5588 = ~n5532 & n5587;
  assign n5589 = ~n5529 & n5588;
  assign n5590 = ~n5548 & n5589;
  assign n5591 = ~n5586 & ~n5590;
  assign n5592 = ~n5546 & n5583;
  assign n5593 = n5567 & ~n5583;
  assign n5594 = ~n5592 & ~n5593;
  assign n5595 = ~n3340 & ~n3341;
  assign n5596 = ~n2473 & ~n5595;
  assign n5597 = ~n2480 & ~n2482;
  assign n5598 = n5596 & ~n5597;
  assign n5599 = ~n5596 & n5597;
  assign n5600 = ~n5598 & ~n5599;
  assign n5601 = g1 & n5600;
  assign n5602 = ~n4308 & ~n5276;
  assign n5603 = ~n4147 & ~n5559;
  assign n5604 = ~n5277 & ~n5603;
  assign n5605 = ~n5602 & ~n5604;
  assign n5606 = n5602 & n5604;
  assign n5607 = ~n5605 & ~n5606;
  assign n5608 = ~g1 & ~n5607;
  assign n5609 = ~n5601 & ~n5608;
  assign n5610 = ~n2597 & ~n3293;
  assign n5611 = ~n3292 & n3329;
  assign n5612 = n3335 & ~n5611;
  assign n5613 = ~n5610 & n5612;
  assign n5614 = n5610 & ~n5612;
  assign n5615 = g1 & ~n5614;
  assign n5616 = ~n5613 & n5615;
  assign n5617 = ~n5226 & ~n5265;
  assign n5618 = ~n5094 & n5257;
  assign n5619 = n5270 & ~n5618;
  assign n5620 = ~n5617 & ~n5619;
  assign n5621 = n5617 & n5619;
  assign n5622 = ~n5620 & ~n5621;
  assign n5623 = ~g1 & ~n5622;
  assign n5624 = ~g83 & ~n5623;
  assign n5625 = ~n5616 & n5624;
  assign n5626 = ~n2473 & ~n3341;
  assign n5627 = ~n3340 & n5626;
  assign n5628 = n3340 & ~n5626;
  assign n5629 = ~n5627 & ~n5628;
  assign n5630 = g1 & n5629;
  assign n5631 = ~n4147 & ~n5277;
  assign n5632 = n5559 & n5631;
  assign n5633 = ~n5559 & ~n5631;
  assign n5634 = ~n5632 & ~n5633;
  assign n5635 = ~g1 & ~n5634;
  assign n5636 = ~n5630 & ~n5635;
  assign n5637 = ~n3293 & ~n5612;
  assign n5638 = ~n2597 & ~n5637;
  assign n5639 = ~n2520 & ~n3337;
  assign n5640 = g1 & ~n5639;
  assign n5641 = ~n5638 & n5640;
  assign n5642 = ~n5226 & ~n5619;
  assign n5643 = ~n5265 & ~n5642;
  assign n5644 = ~n5197 & ~n5264;
  assign n5645 = ~g1 & ~n5644;
  assign n5646 = ~n5643 & n5645;
  assign n5647 = ~n5641 & ~n5646;
  assign n5648 = ~n2520 & n3445;
  assign n5649 = g1 & n5648;
  assign n5650 = ~n5637 & n5649;
  assign n5651 = ~g1 & n5266;
  assign n5652 = ~n5197 & n5651;
  assign n5653 = ~n5642 & n5652;
  assign n5654 = ~n5650 & ~n5653;
  assign n5655 = n5647 & n5654;
  assign n5656 = n5636 & n5655;
  assign n5657 = n5625 & n5656;
  assign n5658 = n5609 & n5657;
  assign n5659 = n5567 & ~n5658;
  assign n5660 = n5549 & n5659;
  assign n5661 = n5594 & n5660;
  assign n5662 = n5591 & ~n5661;
  assign n5663 = ~n5535 & n5662;
  assign n5664 = n5516 & n5663;
  assign n5665 = ~n2397 & ~n5381;
  assign n5666 = n2397 & n5381;
  assign n5667 = ~n5665 & ~n5666;
  assign n5668 = ~n3646 & ~n5667;
  assign n5669 = n3646 & n5667;
  assign n5670 = ~n5668 & ~n5669;
  assign n5671 = ~n5433 & ~n5436;
  assign n5672 = ~n3646 & ~n5430;
  assign n5673 = ~n5671 & ~n5672;
  assign n5674 = ~n5670 & n5673;
  assign n5675 = n5670 & ~n5673;
  assign n5676 = ~n5674 & ~n5675;
  assign n5677 = ~n5444 & ~n5447;
  assign n5678 = ~n5443 & ~n5677;
  assign n5679 = n5676 & n5678;
  assign n5680 = ~n5676 & ~n5678;
  assign n5681 = ~n5679 & ~n5680;
  assign n5682 = ~g1 & n5681;
  assign n5683 = n135 & ~n154;
  assign n5684 = ~n135 & n154;
  assign n5685 = ~n5683 & ~n5684;
  assign n5686 = ~n2397 & ~n5685;
  assign n5687 = n2397 & n5685;
  assign n5688 = ~n5686 & ~n5687;
  assign n5689 = ~n5407 & n5413;
  assign n5690 = ~n5411 & ~n5689;
  assign n5691 = n5688 & n5690;
  assign n5692 = ~n5688 & ~n5690;
  assign n5693 = ~n5691 & ~n5692;
  assign n5694 = ~n5421 & ~n5424;
  assign n5695 = ~n5420 & ~n5694;
  assign n5696 = g1 & n5695;
  assign n5697 = ~n5693 & n5696;
  assign n5698 = g1 & n5693;
  assign n5699 = ~n5695 & n5698;
  assign n5700 = ~n5697 & ~n5699;
  assign n5701 = ~n5682 & n5700;
  assign n5702 = n5452 & n5701;
  assign n5703 = ~n5490 & n5509;
  assign n5704 = ~n5491 & ~n5703;
  assign n5705 = n5625 & ~n5655;
  assign n5706 = ~n5636 & n5655;
  assign n5707 = ~n5705 & ~n5706;
  assign n5708 = ~n5609 & n5636;
  assign n5709 = ~n5567 & n5609;
  assign n5710 = ~n5708 & ~n5709;
  assign n5711 = n5707 & n5710;
  assign n5712 = ~n3292 & ~n3328;
  assign n5713 = ~n3332 & ~n5712;
  assign n5714 = ~n3321 & ~n3334;
  assign n5715 = n5713 & n5714;
  assign n5716 = g1 & n5715;
  assign n5717 = g1 & ~n5713;
  assign n5718 = ~n5714 & n5717;
  assign n5719 = ~n5094 & ~n5256;
  assign n5720 = ~n5267 & ~n5719;
  assign n5721 = ~n5249 & ~n5269;
  assign n5722 = n5720 & ~n5721;
  assign n5723 = ~n5720 & n5721;
  assign n5724 = ~n5722 & ~n5723;
  assign n5725 = ~g1 & n5724;
  assign n5726 = ~g84 & ~n5725;
  assign n5727 = ~n5718 & n5726;
  assign n5728 = ~n5716 & n5727;
  assign n5729 = ~n5616 & ~n5623;
  assign n5730 = g83 & ~n5729;
  assign n5731 = ~n5625 & ~n5730;
  assign n5732 = ~n5728 & ~n5731;
  assign n5733 = ~n5716 & ~n5725;
  assign n5734 = ~n5718 & n5733;
  assign n5735 = g84 & ~n5734;
  assign n5736 = ~n5728 & ~n5735;
  assign n5737 = ~n3328 & ~n3332;
  assign n5738 = n3292 & ~n5737;
  assign n5739 = g1 & ~n5738;
  assign n5740 = ~n3292 & n5737;
  assign n5741 = n5739 & ~n5740;
  assign n5742 = ~n5256 & ~n5267;
  assign n5743 = n5094 & ~n5742;
  assign n5744 = ~n5094 & n5742;
  assign n5745 = ~g1 & ~n5744;
  assign n5746 = ~n5743 & n5745;
  assign n5747 = ~n5741 & ~n5746;
  assign n5748 = ~g85 & n5747;
  assign n5749 = ~n5736 & ~n5748;
  assign n5750 = ~n5732 & ~n5749;
  assign n5751 = ~n2822 & ~n2823;
  assign n5752 = ~n2912 & ~n2978;
  assign n5753 = ~n3280 & n5752;
  assign n5754 = n3287 & ~n5753;
  assign n5755 = ~n2918 & ~n5754;
  assign n5756 = ~n3283 & ~n5755;
  assign n5757 = g1 & ~n5756;
  assign n5758 = ~n5751 & n5757;
  assign n5759 = ~n4610 & ~n4784;
  assign n5760 = ~n5087 & n5089;
  assign n5761 = n4780 & ~n5760;
  assign n5762 = ~n4656 & ~n5761;
  assign n5763 = ~n4782 & ~n5762;
  assign n5764 = ~g1 & n5763;
  assign n5765 = n5759 & n5764;
  assign n5766 = n5751 & n5756;
  assign n5767 = g1 & n5766;
  assign n5768 = ~g1 & ~n5763;
  assign n5769 = ~n5759 & n5768;
  assign n5770 = ~n5767 & ~n5769;
  assign n5771 = ~g86 & n5770;
  assign n5772 = ~n5765 & n5771;
  assign n5773 = ~n5758 & n5772;
  assign n5774 = g85 & ~n5747;
  assign n5775 = ~n5748 & ~n5774;
  assign n5776 = n5773 & n5775;
  assign n5777 = n5736 & n5748;
  assign n5778 = ~n5773 & ~n5775;
  assign n5779 = ~n5758 & ~n5765;
  assign n5780 = n5770 & n5779;
  assign n5781 = g86 & ~n5780;
  assign n5782 = ~n5773 & ~n5781;
  assign n5783 = ~n2918 & ~n3283;
  assign n5784 = n5754 & n5783;
  assign n5785 = g1 & ~n5784;
  assign n5786 = ~n4656 & ~n4782;
  assign n5787 = n5761 & n5786;
  assign n5788 = ~g1 & ~n5787;
  assign n5789 = ~n5785 & ~n5788;
  assign n5790 = ~n5754 & ~n5783;
  assign n5791 = g1 & ~n5790;
  assign n5792 = ~n5761 & ~n5786;
  assign n5793 = ~g1 & ~n5792;
  assign n5794 = ~n5791 & ~n5793;
  assign n5795 = ~g87 & ~n5794;
  assign n5796 = ~n5789 & n5795;
  assign n5797 = ~n5782 & ~n5796;
  assign n5798 = ~n5778 & ~n5797;
  assign n5799 = ~n5777 & ~n5798;
  assign n5800 = ~n5776 & n5799;
  assign n5801 = n5750 & ~n5800;
  assign n5802 = n5728 & n5731;
  assign n5803 = ~n5801 & ~n5802;
  assign n5804 = n5782 & n5796;
  assign n5805 = ~n5776 & ~n5804;
  assign n5806 = ~n5087 & ~n5088;
  assign n5807 = ~n4771 & ~n5806;
  assign n5808 = ~n4777 & ~n4779;
  assign n5809 = ~n5807 & ~n5808;
  assign n5810 = ~g1 & n5809;
  assign n5811 = ~n2978 & ~n3280;
  assign n5812 = ~n3284 & ~n5811;
  assign n5813 = ~n2912 & ~n3286;
  assign n5814 = g1 & ~n5813;
  assign n5815 = ~n5812 & n5814;
  assign n5816 = ~n5810 & ~n5815;
  assign n5817 = n5812 & n5813;
  assign n5818 = g1 & n5817;
  assign n5819 = n5807 & n5808;
  assign n5820 = ~g1 & n5819;
  assign n5821 = ~n5818 & ~n5820;
  assign n5822 = n5816 & n5821;
  assign n5823 = ~g88 & n5822;
  assign n5824 = ~n5789 & ~n5794;
  assign n5825 = g87 & ~n5824;
  assign n5826 = ~n5796 & ~n5825;
  assign n5827 = ~n5823 & ~n5826;
  assign n5828 = ~n4771 & ~n5088;
  assign n5829 = ~n5087 & ~n5828;
  assign n5830 = n5087 & n5828;
  assign n5831 = ~n5829 & ~n5830;
  assign n5832 = ~g1 & ~n5831;
  assign n5833 = ~n2978 & ~n3284;
  assign n5834 = ~n3280 & n5833;
  assign n5835 = n3280 & ~n5833;
  assign n5836 = g1 & ~n5835;
  assign n5837 = ~n5834 & n5836;
  assign n5838 = ~n5832 & ~n5837;
  assign n5839 = ~g89 & n5838;
  assign n5840 = g88 & ~n5822;
  assign n5841 = n5839 & ~n5840;
  assign n5842 = ~n5823 & n5841;
  assign n5843 = ~n5796 & n5823;
  assign n5844 = ~n5825 & n5843;
  assign n5845 = ~n3028 & ~n3143;
  assign n5846 = ~n3140 & ~n3277;
  assign n5847 = ~n3066 & ~n5846;
  assign n5848 = ~n3142 & ~n5847;
  assign n5849 = g1 & n5848;
  assign n5850 = n5845 & n5849;
  assign n5851 = ~n5081 & n5084;
  assign n5852 = ~n4943 & ~n5851;
  assign n5853 = ~n4950 & ~n5852;
  assign n5854 = ~n4952 & ~n5853;
  assign n5855 = ~n4833 & ~n4834;
  assign n5856 = n5854 & n5855;
  assign n5857 = ~g1 & n5856;
  assign n5858 = ~n5854 & ~n5855;
  assign n5859 = ~g1 & n5858;
  assign n5860 = g1 & ~n5845;
  assign n5861 = ~n5848 & n5860;
  assign n5862 = ~n5859 & ~n5861;
  assign n5863 = ~n5857 & n5862;
  assign n5864 = ~n5850 & n5863;
  assign n5865 = g90 & ~n5864;
  assign n5866 = ~n5850 & ~n5859;
  assign n5867 = ~n5857 & ~n5861;
  assign n5868 = ~g90 & n5867;
  assign n5869 = n5866 & n5868;
  assign n5870 = ~n5865 & ~n5869;
  assign n5871 = ~n3066 & ~n3142;
  assign n5872 = n5846 & n5871;
  assign n5873 = ~n5846 & ~n5871;
  assign n5874 = ~n5872 & ~n5873;
  assign n5875 = g1 & ~n5874;
  assign n5876 = ~n4950 & ~n4952;
  assign n5877 = ~n5852 & n5876;
  assign n5878 = ~g1 & ~n5877;
  assign n5879 = n5852 & ~n5876;
  assign n5880 = n5878 & ~n5879;
  assign n5881 = ~n5875 & ~n5880;
  assign n5882 = ~g91 & n5881;
  assign n5883 = ~n5870 & ~n5882;
  assign n5884 = g89 & ~n5838;
  assign n5885 = ~n5839 & n5869;
  assign n5886 = ~n5884 & n5885;
  assign n5887 = n5883 & ~n5886;
  assign n5888 = ~n5839 & ~n5884;
  assign n5889 = ~n5869 & ~n5888;
  assign n5890 = ~n5887 & ~n5889;
  assign n5891 = ~n5844 & ~n5890;
  assign n5892 = ~n5842 & n5891;
  assign n5893 = ~n5823 & ~n5840;
  assign n5894 = ~n5839 & ~n5893;
  assign n5895 = ~n5844 & n5894;
  assign n5896 = ~n5892 & ~n5895;
  assign n5897 = ~n5827 & n5896;
  assign n5898 = ~n3109 & ~n3139;
  assign n5899 = ~n3274 & ~n3275;
  assign n5900 = ~n3137 & ~n5899;
  assign n5901 = ~n5898 & n5900;
  assign n5902 = n5898 & ~n5900;
  assign n5903 = g1 & ~n5902;
  assign n5904 = ~n5901 & n5903;
  assign n5905 = ~n4906 & ~n4942;
  assign n5906 = ~n5081 & ~n5083;
  assign n5907 = ~n4940 & ~n5906;
  assign n5908 = ~n5905 & ~n5907;
  assign n5909 = n5905 & n5907;
  assign n5910 = ~n5908 & ~n5909;
  assign n5911 = ~g1 & ~n5910;
  assign n5912 = ~n5904 & ~n5911;
  assign n5913 = ~g92 & n5912;
  assign n5914 = g91 & ~n5881;
  assign n5915 = ~n5882 & ~n5914;
  assign n5916 = ~n5913 & ~n5915;
  assign n5917 = n5913 & n5915;
  assign n5918 = ~n3137 & ~n3275;
  assign n5919 = ~n3274 & ~n5918;
  assign n5920 = n3274 & n5918;
  assign n5921 = ~n5919 & ~n5920;
  assign n5922 = g1 & ~n5921;
  assign n5923 = ~n4940 & ~n5083;
  assign n5924 = n5081 & ~n5923;
  assign n5925 = ~n5081 & n5923;
  assign n5926 = ~g1 & ~n5925;
  assign n5927 = ~n5924 & n5926;
  assign n5928 = ~n5922 & ~n5927;
  assign n5929 = ~g93 & n5928;
  assign n5930 = g92 & n5912;
  assign n5931 = ~g92 & ~n5912;
  assign n5932 = ~n5930 & ~n5931;
  assign n5933 = ~n5929 & n5932;
  assign n5934 = ~n5917 & n5933;
  assign n5935 = n5929 & ~n5932;
  assign n5936 = g93 & ~n5928;
  assign n5937 = ~n5929 & ~n5936;
  assign n5938 = ~n4982 & ~n5080;
  assign n5939 = ~n5078 & ~n5938;
  assign n5940 = n5078 & n5938;
  assign n5941 = ~n5939 & ~n5940;
  assign n5942 = ~g1 & ~n5941;
  assign n5943 = ~n3177 & ~n3273;
  assign n5944 = ~n3271 & n5943;
  assign n5945 = n3271 & ~n5943;
  assign n5946 = ~n5944 & ~n5945;
  assign n5947 = g1 & n5946;
  assign n5948 = ~n5942 & ~n5947;
  assign n5949 = ~n5937 & ~n5948;
  assign n5950 = g94 & n5948;
  assign n5951 = ~n5937 & n5950;
  assign n5952 = ~n5949 & ~n5951;
  assign n5953 = ~n5917 & ~n5952;
  assign n5954 = ~n5935 & n5953;
  assign n5955 = ~n5006 & ~n5077;
  assign n5956 = ~n5075 & ~n5955;
  assign n5957 = n5075 & n5955;
  assign n5958 = ~n5956 & ~n5957;
  assign n5959 = ~g1 & ~n5958;
  assign n5960 = ~n3201 & ~n3270;
  assign n5961 = ~n3268 & n5960;
  assign n5962 = n3268 & ~n5960;
  assign n5963 = ~n5961 & ~n5962;
  assign n5964 = g1 & n5963;
  assign n5965 = ~n5959 & ~n5964;
  assign n5966 = ~g95 & n5965;
  assign n5967 = n3217 & ~n3220;
  assign n5968 = ~n3217 & n3220;
  assign n5969 = ~n5967 & ~n5968;
  assign n5970 = ~n3265 & ~n5969;
  assign n5971 = n3265 & n5969;
  assign n5972 = g1 & ~n5971;
  assign n5973 = ~n5970 & n5972;
  assign n5974 = ~n5063 & n5072;
  assign n5975 = n5063 & ~n5072;
  assign n5976 = ~n5974 & ~n5975;
  assign n5977 = ~g1 & ~n5976;
  assign n5978 = ~n5973 & ~n5977;
  assign n5979 = ~g96 & n5978;
  assign n5980 = ~n5036 & ~n5062;
  assign n5981 = n5060 & ~n5980;
  assign n5982 = ~n5061 & ~n5981;
  assign n5983 = ~g1 & n5982;
  assign n5984 = ~n3237 & ~n3238;
  assign n5985 = ~n3263 & n5984;
  assign n5986 = n3263 & ~n5984;
  assign n5987 = g1 & ~n5986;
  assign n5988 = ~n5985 & n5987;
  assign n5989 = ~n5983 & ~n5988;
  assign n5990 = g97 & ~n5989;
  assign n5991 = ~n5057 & ~n5059;
  assign n5992 = n5050 & n5991;
  assign n5993 = ~n5050 & ~n5991;
  assign n5994 = ~n5992 & ~n5993;
  assign n5995 = ~g1 & ~n5994;
  assign n5996 = ~n3260 & ~n3262;
  assign n5997 = n3250 & n5996;
  assign n5998 = ~n3250 & ~n5996;
  assign n5999 = ~n5997 & ~n5998;
  assign n6000 = g1 & n5999;
  assign n6001 = ~n5995 & ~n6000;
  assign n6002 = g98 & ~n6001;
  assign n6003 = ~g97 & ~n5989;
  assign n6004 = g97 & n5989;
  assign n6005 = ~n6003 & ~n6004;
  assign n6006 = n6002 & ~n6005;
  assign n6007 = ~n5990 & ~n6006;
  assign n6008 = ~n5979 & ~n6007;
  assign n6009 = g96 & ~n5978;
  assign n6010 = ~n6008 & ~n6009;
  assign n6011 = ~n5966 & ~n6010;
  assign n6012 = g95 & ~n5965;
  assign n6013 = ~n6011 & ~n6012;
  assign n6014 = ~g94 & ~n5948;
  assign n6015 = ~n6013 & ~n6014;
  assign n6016 = n5937 & n5948;
  assign n6017 = n6015 & ~n6016;
  assign n6018 = ~n5917 & n6017;
  assign n6019 = ~n5935 & n6018;
  assign n6020 = ~n5954 & ~n6019;
  assign n6021 = ~n5934 & n6020;
  assign n6022 = ~n5916 & n6021;
  assign n6023 = n5870 & n5882;
  assign n6024 = ~n5886 & ~n6023;
  assign n6025 = ~n6022 & n6024;
  assign n6026 = ~n5844 & n6025;
  assign n6027 = ~n5842 & n6026;
  assign n6028 = n5897 & ~n6027;
  assign n6029 = ~n5802 & ~n6028;
  assign n6030 = n5805 & n6029;
  assign n6031 = ~n5777 & n6030;
  assign n6032 = ~n5803 & ~n6031;
  assign n6033 = n5549 & ~n6032;
  assign n6034 = n5711 & n6033;
  assign n6035 = n5594 & n6034;
  assign n6036 = n5452 & ~n5701;
  assign n6037 = n5475 & ~n6036;
  assign n6038 = n6035 & n6037;
  assign n6039 = n5704 & n6038;
  assign n6040 = g0 & ~n6039;
  assign n6041 = n5702 & n6040;
  assign n6042 = n5664 & n6041;
  assign n6043 = ~g1 & n5402;
  assign n6044 = ~n5638 & n5639;
  assign n6045 = n2036 & ~n2127;
  assign n6046 = ~n2130 & ~n2133;
  assign n6047 = ~n6045 & ~n6046;
  assign n6048 = ~n693 & n6047;
  assign n6049 = n693 & ~n6047;
  assign n6050 = ~n6048 & ~n6049;
  assign n6051 = n3451 & ~n6050;
  assign n6052 = n5597 & n6051;
  assign n6053 = n5626 & n6052;
  assign n6054 = n6044 & n6053;
  assign n6055 = n5597 & n5626;
  assign n6056 = n3337 & n6055;
  assign n6057 = n2483 & ~n6056;
  assign n6058 = n6051 & ~n6057;
  assign n6059 = n2193 & ~n6050;
  assign n6060 = ~n6058 & ~n6059;
  assign n6061 = ~n6054 & n6060;
  assign n6062 = ~n693 & ~n6047;
  assign n6063 = n6061 & ~n6062;
  assign n6064 = n5541 & ~n6063;
  assign n6065 = ~n677 & ~n6064;
  assign n6066 = n5519 & ~n6065;
  assign n6067 = ~n522 & ~n6066;
  assign n6068 = n5493 & ~n6067;
  assign n6069 = ~n681 & ~n6068;
  assign n6070 = n5477 & ~n6069;
  assign n6071 = ~n684 & ~n6070;
  assign n6072 = n5457 & ~n6071;
  assign n6073 = ~n687 & ~n6072;
  assign n6074 = n244 & ~n6073;
  assign n6075 = ~n244 & n6073;
  assign n6076 = ~n6074 & ~n6075;
  assign n6077 = g1 & ~n6076;
  assign n6078 = ~n6043 & ~n6077;
  assign n6079 = ~n242 & ~n6074;
  assign n6080 = ~n5422 & ~n6079;
  assign n6081 = n5422 & n6079;
  assign n6082 = ~n6080 & ~n6081;
  assign n6083 = g1 & n6082;
  assign n6084 = ~g1 & n5450;
  assign n6085 = ~n6083 & ~n6084;
  assign n6086 = ~n6078 & n6085;
  assign n6087 = ~n5485 & ~n5487;
  assign n6088 = ~g1 & ~n6087;
  assign n6089 = ~n5477 & n6069;
  assign n6090 = ~n6070 & ~n6089;
  assign n6091 = g1 & ~n6090;
  assign n6092 = ~n6088 & ~n6091;
  assign n6093 = ~n5465 & ~n5467;
  assign n6094 = ~g1 & ~n6093;
  assign n6095 = n5457 & n6071;
  assign n6096 = ~n5457 & ~n6071;
  assign n6097 = ~n6095 & ~n6096;
  assign n6098 = g1 & n6097;
  assign n6099 = ~n6094 & ~n6098;
  assign n6100 = ~n6092 & ~n6099;
  assign n6101 = ~n5493 & n6067;
  assign n6102 = ~n6068 & ~n6101;
  assign n6103 = g1 & ~n6102;
  assign n6104 = ~n5500 & ~n5502;
  assign n6105 = ~g1 & ~n6104;
  assign n6106 = ~n6103 & ~n6105;
  assign n6107 = n6092 & n6106;
  assign n6108 = ~n6100 & ~n6107;
  assign n6109 = ~n6078 & ~n6108;
  assign n6110 = n6099 & n6107;
  assign n6111 = ~n6109 & ~n6110;
  assign n6112 = ~n5523 & ~n5524;
  assign n6113 = n5523 & n5524;
  assign n6114 = ~n6112 & ~n6113;
  assign n6115 = ~g1 & n6114;
  assign n6116 = ~n5519 & n6065;
  assign n6117 = ~n6066 & ~n6116;
  assign n6118 = g1 & ~n6117;
  assign n6119 = ~n6115 & ~n6118;
  assign n6120 = ~g1 & ~n5539;
  assign n6121 = ~n5541 & n6063;
  assign n6122 = ~n6064 & ~n6121;
  assign n6123 = g1 & ~n6122;
  assign n6124 = ~n6120 & ~n6123;
  assign n6125 = ~n5578 & ~n5580;
  assign n6126 = ~g1 & ~n6125;
  assign n6127 = ~n2193 & n6050;
  assign n6128 = ~n3452 & n6127;
  assign n6129 = n6061 & ~n6128;
  assign n6130 = g1 & ~n6129;
  assign n6131 = ~n6126 & ~n6130;
  assign n6132 = n6124 & n6131;
  assign n6133 = n6119 & n6132;
  assign n6134 = ~n6119 & ~n6124;
  assign n6135 = ~n6106 & n6134;
  assign n6136 = ~n6133 & ~n6135;
  assign n6137 = n5707 & ~n6032;
  assign n6138 = ~n5609 & ~n5636;
  assign n6139 = ~n5567 & n6138;
  assign n6140 = n6131 & ~n6139;
  assign n6141 = n6137 & ~n6140;
  assign n6142 = ~n6136 & n6141;
  assign n6143 = ~n6111 & n6142;
  assign n6144 = ~n6086 & n6143;
  assign n6145 = ~g1 & ~n5681;
  assign n6146 = n5422 & ~n6079;
  assign n6147 = ~n5420 & ~n6146;
  assign n6148 = ~n5693 & ~n6147;
  assign n6149 = n5693 & n6147;
  assign n6150 = ~n6148 & ~n6149;
  assign n6151 = g1 & ~n6150;
  assign n6152 = ~n6145 & ~n6151;
  assign n6153 = ~n6085 & n6152;
  assign n6154 = n6144 & ~n6153;
  assign n6155 = g0 & n5609;
  assign n6156 = n5625 & n6155;
  assign n6157 = n5656 & n6156;
  assign n6158 = n5567 & ~n6131;
  assign n6159 = n6157 & n6158;
  assign n6160 = n6135 & n6159;
  assign n6161 = ~n6085 & ~n6111;
  assign n6162 = n6160 & n6161;
  assign n6163 = ~n6152 & n6162;
  assign n6164 = ~n6154 & n6163;
  assign n6165 = ~n6042 & n6164;
  assign n6166 = n6042 & ~n6164;
  assign n6167 = ~n6165 & ~n6166;
  assign n6168 = g72 & g83;
  assign n6169 = g71 & g84;
  assign n6170 = g69 & g86;
  assign n6171 = n6169 & ~n6170;
  assign n6172 = ~n6169 & n6170;
  assign n6173 = ~n6171 & ~n6172;
  assign n6174 = n6168 & ~n6173;
  assign n6175 = n6169 & n6170;
  assign n6176 = ~n6174 & ~n6175;
  assign n6177 = g71 & g83;
  assign n6178 = g69 & g85;
  assign n6179 = ~n6177 & n6178;
  assign n6180 = n6177 & ~n6178;
  assign n6181 = ~n6179 & ~n6180;
  assign n6182 = n6176 & ~n6181;
  assign n6183 = ~n6176 & n6181;
  assign n6184 = ~n6182 & ~n6183;
  assign n6185 = g70 & g84;
  assign n6186 = g68 & g86;
  assign n6187 = g67 & g87;
  assign n6188 = n6186 & ~n6187;
  assign n6189 = ~n6186 & n6187;
  assign n6190 = ~n6188 & ~n6189;
  assign n6191 = ~n6185 & ~n6190;
  assign n6192 = n6185 & n6190;
  assign n6193 = ~n6191 & ~n6192;
  assign n6194 = g70 & g85;
  assign n6195 = g68 & g87;
  assign n6196 = g67 & g88;
  assign n6197 = n6195 & ~n6196;
  assign n6198 = ~n6195 & n6196;
  assign n6199 = ~n6197 & ~n6198;
  assign n6200 = n6194 & ~n6199;
  assign n6201 = n6195 & n6196;
  assign n6202 = ~n6200 & ~n6201;
  assign n6203 = n6193 & ~n6202;
  assign n6204 = ~n6193 & n6202;
  assign n6205 = ~n6203 & ~n6204;
  assign n6206 = ~n6184 & ~n6205;
  assign n6207 = ~n6193 & ~n6202;
  assign n6208 = ~n6206 & ~n6207;
  assign n6209 = ~n6176 & ~n6181;
  assign n6210 = n6177 & n6178;
  assign n6211 = ~n6209 & ~n6210;
  assign n6212 = g70 & g83;
  assign n6213 = g68 & g85;
  assign n6214 = g67 & g86;
  assign n6215 = n6213 & ~n6214;
  assign n6216 = ~n6213 & n6214;
  assign n6217 = ~n6215 & ~n6216;
  assign n6218 = ~n6212 & ~n6217;
  assign n6219 = n6212 & n6217;
  assign n6220 = ~n6218 & ~n6219;
  assign n6221 = n6185 & ~n6190;
  assign n6222 = n6186 & n6187;
  assign n6223 = ~n6221 & ~n6222;
  assign n6224 = g69 & g84;
  assign n6225 = n6223 & n6224;
  assign n6226 = ~n6223 & ~n6224;
  assign n6227 = ~n6225 & ~n6226;
  assign n6228 = n6220 & ~n6227;
  assign n6229 = ~n6220 & n6227;
  assign n6230 = ~n6228 & ~n6229;
  assign n6231 = ~n6211 & n6230;
  assign n6232 = n6211 & ~n6230;
  assign n6233 = ~n6231 & ~n6232;
  assign n6234 = n6208 & ~n6233;
  assign n6235 = ~n6208 & n6233;
  assign n6236 = ~n6234 & ~n6235;
  assign n6237 = ~n6194 & ~n6199;
  assign n6238 = n6194 & n6199;
  assign n6239 = ~n6237 & ~n6238;
  assign n6240 = g72 & g84;
  assign n6241 = g71 & g85;
  assign n6242 = g69 & g87;
  assign n6243 = n6241 & ~n6242;
  assign n6244 = ~n6241 & n6242;
  assign n6245 = ~n6243 & ~n6244;
  assign n6246 = n6240 & ~n6245;
  assign n6247 = n6241 & n6242;
  assign n6248 = ~n6246 & ~n6247;
  assign n6249 = g70 & g86;
  assign n6250 = g68 & g88;
  assign n6251 = g67 & g89;
  assign n6252 = n6250 & ~n6251;
  assign n6253 = ~n6250 & n6251;
  assign n6254 = ~n6252 & ~n6253;
  assign n6255 = n6249 & ~n6254;
  assign n6256 = n6250 & n6251;
  assign n6257 = ~n6255 & ~n6256;
  assign n6258 = n6248 & ~n6257;
  assign n6259 = ~n6248 & n6257;
  assign n6260 = ~n6258 & ~n6259;
  assign n6261 = n6239 & ~n6260;
  assign n6262 = ~n6239 & n6260;
  assign n6263 = ~n6261 & ~n6262;
  assign n6264 = n6168 & n6173;
  assign n6265 = ~n6168 & ~n6173;
  assign n6266 = ~n6264 & ~n6265;
  assign n6267 = g69 & g88;
  assign n6268 = g74 & g83;
  assign n6269 = g71 & g86;
  assign n6270 = n6268 & ~n6269;
  assign n6271 = ~n6268 & n6269;
  assign n6272 = ~n6270 & ~n6271;
  assign n6273 = n6267 & ~n6272;
  assign n6274 = n6268 & n6269;
  assign n6275 = ~n6273 & ~n6274;
  assign n6276 = g73 & g83;
  assign n6277 = g70 & g87;
  assign n6278 = g68 & g89;
  assign n6279 = g67 & g90;
  assign n6280 = n6278 & ~n6279;
  assign n6281 = ~n6278 & n6279;
  assign n6282 = ~n6280 & ~n6281;
  assign n6283 = n6277 & ~n6282;
  assign n6284 = n6278 & n6279;
  assign n6285 = ~n6283 & ~n6284;
  assign n6286 = ~n6276 & ~n6285;
  assign n6287 = n6276 & n6285;
  assign n6288 = ~n6286 & ~n6287;
  assign n6289 = ~n6275 & ~n6288;
  assign n6290 = n6276 & ~n6285;
  assign n6291 = ~n6289 & ~n6290;
  assign n6292 = ~n6266 & n6291;
  assign n6293 = n6266 & ~n6291;
  assign n6294 = ~n6292 & ~n6293;
  assign n6295 = ~n6263 & ~n6294;
  assign n6296 = ~n6266 & ~n6291;
  assign n6297 = ~n6295 & ~n6296;
  assign n6298 = n6184 & ~n6205;
  assign n6299 = ~n6184 & n6205;
  assign n6300 = ~n6298 & ~n6299;
  assign n6301 = ~n6239 & ~n6260;
  assign n6302 = ~n6248 & ~n6257;
  assign n6303 = ~n6301 & ~n6302;
  assign n6304 = ~n6300 & n6303;
  assign n6305 = n6300 & ~n6303;
  assign n6306 = ~n6304 & ~n6305;
  assign n6307 = ~n6297 & ~n6306;
  assign n6308 = ~n6300 & ~n6303;
  assign n6309 = ~n6307 & ~n6308;
  assign n6310 = n6236 & n6309;
  assign n6311 = n6297 & ~n6306;
  assign n6312 = ~n6297 & n6306;
  assign n6313 = ~n6311 & ~n6312;
  assign n6314 = g72 & g87;
  assign n6315 = g76 & g83;
  assign n6316 = g69 & g90;
  assign n6317 = n6315 & ~n6316;
  assign n6318 = ~n6315 & n6316;
  assign n6319 = ~n6317 & ~n6318;
  assign n6320 = n6314 & ~n6319;
  assign n6321 = n6315 & n6316;
  assign n6322 = ~n6320 & ~n6321;
  assign n6323 = g71 & g88;
  assign n6324 = g75 & g84;
  assign n6325 = g74 & g85;
  assign n6326 = n6324 & ~n6325;
  assign n6327 = ~n6324 & n6325;
  assign n6328 = ~n6326 & ~n6327;
  assign n6329 = n6323 & ~n6328;
  assign n6330 = n6324 & n6325;
  assign n6331 = ~n6329 & ~n6330;
  assign n6332 = g70 & g89;
  assign n6333 = g67 & g92;
  assign n6334 = g68 & g91;
  assign n6335 = ~n6333 & n6334;
  assign n6336 = n6333 & ~n6334;
  assign n6337 = ~n6335 & ~n6336;
  assign n6338 = n6332 & ~n6337;
  assign n6339 = n6333 & n6334;
  assign n6340 = ~n6338 & ~n6339;
  assign n6341 = n6331 & ~n6340;
  assign n6342 = ~n6331 & n6340;
  assign n6343 = ~n6341 & ~n6342;
  assign n6344 = ~n6322 & ~n6343;
  assign n6345 = ~n6331 & ~n6340;
  assign n6346 = ~n6344 & ~n6345;
  assign n6347 = g73 & g85;
  assign n6348 = g69 & g89;
  assign n6349 = g72 & g86;
  assign n6350 = ~n6348 & n6349;
  assign n6351 = n6348 & ~n6349;
  assign n6352 = ~n6350 & ~n6351;
  assign n6353 = n6347 & ~n6352;
  assign n6354 = n6348 & n6349;
  assign n6355 = ~n6353 & ~n6354;
  assign n6356 = g72 & g85;
  assign n6357 = g73 & g84;
  assign n6358 = ~n6356 & n6357;
  assign n6359 = n6356 & ~n6357;
  assign n6360 = ~n6358 & ~n6359;
  assign n6361 = n6355 & ~n6360;
  assign n6362 = ~n6355 & n6360;
  assign n6363 = ~n6361 & ~n6362;
  assign n6364 = n6267 & n6272;
  assign n6365 = ~n6267 & ~n6272;
  assign n6366 = ~n6364 & ~n6365;
  assign n6367 = ~n6363 & n6366;
  assign n6368 = n6363 & ~n6366;
  assign n6369 = ~n6367 & ~n6368;
  assign n6370 = ~n6346 & ~n6369;
  assign n6371 = ~n6363 & ~n6366;
  assign n6372 = ~n6370 & ~n6371;
  assign n6373 = n6275 & ~n6288;
  assign n6374 = ~n6275 & n6288;
  assign n6375 = ~n6373 & ~n6374;
  assign n6376 = ~n6277 & ~n6282;
  assign n6377 = n6277 & n6282;
  assign n6378 = ~n6376 & ~n6377;
  assign n6379 = g71 & g87;
  assign n6380 = g75 & g83;
  assign n6381 = g74 & g84;
  assign n6382 = n6380 & ~n6381;
  assign n6383 = ~n6380 & n6381;
  assign n6384 = ~n6382 & ~n6383;
  assign n6385 = n6379 & ~n6384;
  assign n6386 = n6380 & n6381;
  assign n6387 = ~n6385 & ~n6386;
  assign n6388 = g70 & g88;
  assign n6389 = g68 & g90;
  assign n6390 = g67 & g91;
  assign n6391 = n6389 & ~n6390;
  assign n6392 = ~n6389 & n6390;
  assign n6393 = ~n6391 & ~n6392;
  assign n6394 = n6388 & ~n6393;
  assign n6395 = n6389 & n6390;
  assign n6396 = ~n6394 & ~n6395;
  assign n6397 = n6387 & ~n6396;
  assign n6398 = ~n6387 & n6396;
  assign n6399 = ~n6397 & ~n6398;
  assign n6400 = ~n6378 & ~n6399;
  assign n6401 = ~n6387 & ~n6396;
  assign n6402 = ~n6400 & ~n6401;
  assign n6403 = ~n6375 & n6402;
  assign n6404 = n6375 & ~n6402;
  assign n6405 = ~n6403 & ~n6404;
  assign n6406 = ~n6372 & ~n6405;
  assign n6407 = ~n6375 & ~n6402;
  assign n6408 = ~n6406 & ~n6407;
  assign n6409 = n6263 & ~n6294;
  assign n6410 = ~n6263 & n6294;
  assign n6411 = ~n6409 & ~n6410;
  assign n6412 = ~n6355 & ~n6360;
  assign n6413 = n6356 & n6357;
  assign n6414 = ~n6412 & ~n6413;
  assign n6415 = n6249 & n6254;
  assign n6416 = ~n6249 & ~n6254;
  assign n6417 = ~n6415 & ~n6416;
  assign n6418 = n6240 & n6245;
  assign n6419 = ~n6240 & ~n6245;
  assign n6420 = ~n6418 & ~n6419;
  assign n6421 = ~n6417 & n6420;
  assign n6422 = n6417 & ~n6420;
  assign n6423 = ~n6421 & ~n6422;
  assign n6424 = ~n6414 & ~n6423;
  assign n6425 = ~n6417 & ~n6420;
  assign n6426 = ~n6424 & ~n6425;
  assign n6427 = n6411 & ~n6426;
  assign n6428 = ~n6411 & n6426;
  assign n6429 = ~n6427 & ~n6428;
  assign n6430 = ~n6408 & ~n6429;
  assign n6431 = ~n6411 & ~n6426;
  assign n6432 = ~n6430 & ~n6431;
  assign n6433 = n6313 & n6432;
  assign n6434 = ~n6408 & n6429;
  assign n6435 = n6408 & ~n6429;
  assign n6436 = ~n6434 & ~n6435;
  assign n6437 = ~n6347 & n6352;
  assign n6438 = ~n6353 & ~n6437;
  assign n6439 = ~n6388 & ~n6393;
  assign n6440 = n6388 & n6393;
  assign n6441 = ~n6439 & ~n6440;
  assign n6442 = n6438 & ~n6441;
  assign n6443 = ~n6379 & ~n6384;
  assign n6444 = n6379 & n6384;
  assign n6445 = ~n6443 & ~n6444;
  assign n6446 = ~n6438 & ~n6441;
  assign n6447 = n6438 & n6441;
  assign n6448 = ~n6446 & ~n6447;
  assign n6449 = ~n6445 & ~n6448;
  assign n6450 = ~n6442 & ~n6449;
  assign n6451 = n6378 & ~n6399;
  assign n6452 = ~n6378 & n6399;
  assign n6453 = ~n6451 & ~n6452;
  assign n6454 = ~n6450 & n6453;
  assign n6455 = n6450 & ~n6453;
  assign n6456 = ~n6454 & ~n6455;
  assign n6457 = ~n6322 & n6343;
  assign n6458 = n6322 & ~n6343;
  assign n6459 = ~n6457 & ~n6458;
  assign n6460 = g73 & g86;
  assign n6461 = g70 & g90;
  assign n6462 = g67 & g93;
  assign n6463 = g68 & g92;
  assign n6464 = ~n6462 & n6463;
  assign n6465 = n6462 & ~n6463;
  assign n6466 = ~n6464 & ~n6465;
  assign n6467 = n6461 & ~n6466;
  assign n6468 = n6462 & n6463;
  assign n6469 = ~n6467 & ~n6468;
  assign n6470 = n6460 & ~n6469;
  assign n6471 = g75 & g85;
  assign n6472 = g74 & g86;
  assign n6473 = n6471 & n6472;
  assign n6474 = g71 & g89;
  assign n6475 = ~n6471 & ~n6472;
  assign n6476 = ~n6473 & ~n6475;
  assign n6477 = n6474 & n6476;
  assign n6478 = ~n6473 & ~n6477;
  assign n6479 = n6460 & n6469;
  assign n6480 = ~n6460 & ~n6469;
  assign n6481 = ~n6479 & ~n6480;
  assign n6482 = ~n6478 & ~n6481;
  assign n6483 = ~n6470 & ~n6482;
  assign n6484 = g69 & g91;
  assign n6485 = g77 & g83;
  assign n6486 = g76 & g84;
  assign n6487 = n6485 & ~n6486;
  assign n6488 = ~n6485 & n6486;
  assign n6489 = ~n6487 & ~n6488;
  assign n6490 = n6484 & ~n6489;
  assign n6491 = n6485 & n6486;
  assign n6492 = ~n6490 & ~n6491;
  assign n6493 = ~n6332 & n6337;
  assign n6494 = ~n6338 & ~n6493;
  assign n6495 = ~n6492 & n6494;
  assign n6496 = n6323 & n6328;
  assign n6497 = ~n6323 & ~n6328;
  assign n6498 = ~n6496 & ~n6497;
  assign n6499 = ~n6492 & ~n6494;
  assign n6500 = n6492 & n6494;
  assign n6501 = ~n6499 & ~n6500;
  assign n6502 = ~n6498 & ~n6501;
  assign n6503 = ~n6495 & ~n6502;
  assign n6504 = n6483 & ~n6503;
  assign n6505 = ~n6483 & n6503;
  assign n6506 = ~n6504 & ~n6505;
  assign n6507 = ~n6459 & ~n6506;
  assign n6508 = ~n6483 & ~n6503;
  assign n6509 = ~n6507 & ~n6508;
  assign n6510 = ~n6456 & ~n6509;
  assign n6511 = ~n6450 & ~n6453;
  assign n6512 = ~n6510 & ~n6511;
  assign n6513 = ~n6372 & n6405;
  assign n6514 = n6372 & ~n6405;
  assign n6515 = ~n6513 & ~n6514;
  assign n6516 = n6414 & ~n6423;
  assign n6517 = ~n6414 & n6423;
  assign n6518 = ~n6516 & ~n6517;
  assign n6519 = n6515 & ~n6518;
  assign n6520 = ~n6515 & n6518;
  assign n6521 = ~n6519 & ~n6520;
  assign n6522 = ~n6512 & ~n6521;
  assign n6523 = ~n6515 & ~n6518;
  assign n6524 = ~n6522 & ~n6523;
  assign n6525 = n6436 & n6524;
  assign n6526 = ~n6433 & ~n6525;
  assign n6527 = ~n6310 & n6526;
  assign n6528 = g69 & g83;
  assign n6529 = g68 & g84;
  assign n6530 = g67 & g85;
  assign n6531 = n6529 & ~n6530;
  assign n6532 = ~n6529 & n6530;
  assign n6533 = ~n6531 & ~n6532;
  assign n6534 = n6528 & ~n6533;
  assign n6535 = n6529 & n6530;
  assign n6536 = ~n6534 & ~n6535;
  assign n6537 = g67 & g84;
  assign n6538 = g68 & g83;
  assign n6539 = ~n6537 & n6538;
  assign n6540 = n6537 & ~n6538;
  assign n6541 = ~n6539 & ~n6540;
  assign n6542 = n6536 & ~n6541;
  assign n6543 = ~n6536 & n6541;
  assign n6544 = ~n6542 & ~n6543;
  assign n6545 = ~n6528 & ~n6533;
  assign n6546 = n6528 & n6533;
  assign n6547 = ~n6545 & ~n6546;
  assign n6548 = n6212 & ~n6217;
  assign n6549 = n6213 & n6214;
  assign n6550 = ~n6548 & ~n6549;
  assign n6551 = n6547 & ~n6550;
  assign n6552 = ~n6547 & n6550;
  assign n6553 = ~n6551 & ~n6552;
  assign n6554 = ~n6220 & ~n6227;
  assign n6555 = ~n6223 & n6224;
  assign n6556 = ~n6554 & ~n6555;
  assign n6557 = ~n6553 & ~n6556;
  assign n6558 = ~n6547 & ~n6550;
  assign n6559 = ~n6557 & ~n6558;
  assign n6560 = n6544 & n6559;
  assign n6561 = n6553 & n6556;
  assign n6562 = ~n6557 & ~n6561;
  assign n6563 = ~n6208 & ~n6233;
  assign n6564 = ~n6211 & ~n6230;
  assign n6565 = ~n6563 & ~n6564;
  assign n6566 = ~n6562 & n6565;
  assign n6567 = ~n6560 & ~n6566;
  assign n6568 = g67 & g83;
  assign n6569 = ~n6536 & ~n6541;
  assign n6570 = n6537 & n6538;
  assign n6571 = ~n6569 & ~n6570;
  assign n6572 = ~n6568 & n6571;
  assign n6573 = n6567 & ~n6572;
  assign n6574 = ~n6512 & n6521;
  assign n6575 = n6512 & ~n6521;
  assign n6576 = ~n6574 & ~n6575;
  assign n6577 = ~n6498 & n6501;
  assign n6578 = n6498 & ~n6501;
  assign n6579 = ~n6577 & ~n6578;
  assign n6580 = n6478 & n6481;
  assign n6581 = ~n6482 & ~n6580;
  assign n6582 = n6461 & n6466;
  assign n6583 = ~n6461 & ~n6466;
  assign n6584 = ~n6582 & ~n6583;
  assign n6585 = ~n6484 & n6489;
  assign n6586 = ~n6490 & ~n6585;
  assign n6587 = ~n6474 & ~n6476;
  assign n6588 = ~n6477 & ~n6587;
  assign n6589 = n6586 & ~n6588;
  assign n6590 = ~n6586 & n6588;
  assign n6591 = ~n6589 & ~n6590;
  assign n6592 = ~n6584 & ~n6591;
  assign n6593 = n6586 & n6588;
  assign n6594 = ~n6592 & ~n6593;
  assign n6595 = n6581 & n6594;
  assign n6596 = ~n6581 & ~n6594;
  assign n6597 = ~n6595 & ~n6596;
  assign n6598 = ~n6579 & ~n6597;
  assign n6599 = n6581 & ~n6594;
  assign n6600 = ~n6598 & ~n6599;
  assign n6601 = g69 & g92;
  assign n6602 = g76 & g85;
  assign n6603 = g77 & g84;
  assign n6604 = n6602 & ~n6603;
  assign n6605 = ~n6602 & n6603;
  assign n6606 = ~n6604 & ~n6605;
  assign n6607 = n6601 & ~n6606;
  assign n6608 = n6602 & n6603;
  assign n6609 = ~n6607 & ~n6608;
  assign n6610 = g70 & g91;
  assign n6611 = g67 & g94;
  assign n6612 = g68 & g93;
  assign n6613 = ~n6611 & n6612;
  assign n6614 = n6611 & ~n6612;
  assign n6615 = ~n6613 & ~n6614;
  assign n6616 = n6610 & ~n6615;
  assign n6617 = n6611 & n6612;
  assign n6618 = ~n6616 & ~n6617;
  assign n6619 = g74 & g87;
  assign n6620 = g75 & g86;
  assign n6621 = n6619 & n6620;
  assign n6622 = g71 & g90;
  assign n6623 = ~n6619 & ~n6620;
  assign n6624 = ~n6621 & ~n6623;
  assign n6625 = n6622 & n6624;
  assign n6626 = ~n6621 & ~n6625;
  assign n6627 = n6618 & ~n6626;
  assign n6628 = ~n6618 & n6626;
  assign n6629 = ~n6627 & ~n6628;
  assign n6630 = ~n6609 & ~n6629;
  assign n6631 = ~n6618 & ~n6626;
  assign n6632 = ~n6630 & ~n6631;
  assign n6633 = n6314 & n6319;
  assign n6634 = ~n6314 & ~n6319;
  assign n6635 = ~n6633 & ~n6634;
  assign n6636 = ~n6632 & ~n6635;
  assign n6637 = g72 & g88;
  assign n6638 = g73 & g87;
  assign n6639 = ~n6637 & n6638;
  assign n6640 = n6637 & ~n6638;
  assign n6641 = ~n6639 & ~n6640;
  assign n6642 = g73 & g88;
  assign n6643 = g72 & g89;
  assign n6644 = g78 & g83;
  assign n6645 = n6643 & ~n6644;
  assign n6646 = ~n6643 & n6644;
  assign n6647 = ~n6645 & ~n6646;
  assign n6648 = n6642 & ~n6647;
  assign n6649 = n6643 & n6644;
  assign n6650 = ~n6648 & ~n6649;
  assign n6651 = ~n6641 & ~n6650;
  assign n6652 = n6637 & n6638;
  assign n6653 = ~n6651 & ~n6652;
  assign n6654 = n6632 & n6635;
  assign n6655 = ~n6636 & ~n6654;
  assign n6656 = ~n6653 & n6655;
  assign n6657 = ~n6636 & ~n6656;
  assign n6658 = ~n6445 & n6448;
  assign n6659 = n6445 & ~n6448;
  assign n6660 = ~n6658 & ~n6659;
  assign n6661 = n6657 & ~n6660;
  assign n6662 = ~n6657 & n6660;
  assign n6663 = ~n6661 & ~n6662;
  assign n6664 = ~n6600 & ~n6663;
  assign n6665 = ~n6657 & ~n6660;
  assign n6666 = ~n6664 & ~n6665;
  assign n6667 = n6346 & ~n6369;
  assign n6668 = ~n6346 & n6369;
  assign n6669 = ~n6667 & ~n6668;
  assign n6670 = ~n6456 & n6509;
  assign n6671 = n6456 & ~n6509;
  assign n6672 = ~n6670 & ~n6671;
  assign n6673 = ~n6669 & n6672;
  assign n6674 = n6669 & ~n6672;
  assign n6675 = ~n6673 & ~n6674;
  assign n6676 = ~n6666 & ~n6675;
  assign n6677 = ~n6669 & ~n6672;
  assign n6678 = ~n6676 & ~n6677;
  assign n6679 = n6576 & n6678;
  assign n6680 = ~n6666 & n6675;
  assign n6681 = n6666 & ~n6675;
  assign n6682 = ~n6680 & ~n6681;
  assign n6683 = ~n6579 & n6597;
  assign n6684 = n6579 & ~n6597;
  assign n6685 = ~n6683 & ~n6684;
  assign n6686 = ~n6653 & ~n6655;
  assign n6687 = n6653 & n6655;
  assign n6688 = ~n6686 & ~n6687;
  assign n6689 = ~n6609 & n6629;
  assign n6690 = n6609 & ~n6629;
  assign n6691 = ~n6689 & ~n6690;
  assign n6692 = g75 & g87;
  assign n6693 = g74 & g88;
  assign n6694 = n6692 & n6693;
  assign n6695 = g71 & g91;
  assign n6696 = ~n6692 & ~n6693;
  assign n6697 = ~n6694 & ~n6696;
  assign n6698 = n6695 & n6697;
  assign n6699 = ~n6694 & ~n6698;
  assign n6700 = g70 & g92;
  assign n6701 = g67 & g95;
  assign n6702 = g68 & g94;
  assign n6703 = ~n6701 & n6702;
  assign n6704 = n6701 & ~n6702;
  assign n6705 = ~n6703 & ~n6704;
  assign n6706 = n6700 & ~n6705;
  assign n6707 = n6701 & n6702;
  assign n6708 = ~n6706 & ~n6707;
  assign n6709 = g79 & g83;
  assign n6710 = g72 & g90;
  assign n6711 = g78 & g84;
  assign n6712 = ~n6710 & n6711;
  assign n6713 = n6710 & ~n6711;
  assign n6714 = ~n6712 & ~n6713;
  assign n6715 = n6709 & ~n6714;
  assign n6716 = n6710 & n6711;
  assign n6717 = ~n6715 & ~n6716;
  assign n6718 = ~n6708 & n6717;
  assign n6719 = n6708 & ~n6717;
  assign n6720 = ~n6718 & ~n6719;
  assign n6721 = ~n6699 & ~n6720;
  assign n6722 = ~n6708 & ~n6717;
  assign n6723 = ~n6721 & ~n6722;
  assign n6724 = ~n6641 & n6650;
  assign n6725 = n6641 & ~n6650;
  assign n6726 = ~n6724 & ~n6725;
  assign n6727 = n6723 & ~n6726;
  assign n6728 = ~n6723 & n6726;
  assign n6729 = ~n6727 & ~n6728;
  assign n6730 = ~n6691 & ~n6729;
  assign n6731 = ~n6723 & ~n6726;
  assign n6732 = ~n6730 & ~n6731;
  assign n6733 = n6688 & ~n6732;
  assign n6734 = ~n6688 & n6732;
  assign n6735 = ~n6733 & ~n6734;
  assign n6736 = ~n6685 & ~n6735;
  assign n6737 = ~n6688 & ~n6732;
  assign n6738 = ~n6736 & ~n6737;
  assign n6739 = ~n6600 & n6663;
  assign n6740 = n6600 & ~n6663;
  assign n6741 = ~n6739 & ~n6740;
  assign n6742 = n6459 & ~n6506;
  assign n6743 = ~n6459 & n6506;
  assign n6744 = ~n6742 & ~n6743;
  assign n6745 = n6741 & ~n6744;
  assign n6746 = ~n6741 & n6744;
  assign n6747 = ~n6745 & ~n6746;
  assign n6748 = ~n6738 & ~n6747;
  assign n6749 = ~n6741 & ~n6744;
  assign n6750 = ~n6748 & ~n6749;
  assign n6751 = n6682 & n6750;
  assign n6752 = g70 & g95;
  assign n6753 = g82 & g83;
  assign n6754 = g74 & g91;
  assign n6755 = n6753 & ~n6754;
  assign n6756 = ~n6753 & n6754;
  assign n6757 = ~n6755 & ~n6756;
  assign n6758 = ~n6752 & ~n6757;
  assign n6759 = n6752 & n6757;
  assign n6760 = ~n6758 & ~n6759;
  assign n6761 = g80 & g85;
  assign n6762 = g72 & g93;
  assign n6763 = g79 & g86;
  assign n6764 = n6762 & ~n6763;
  assign n6765 = ~n6762 & n6763;
  assign n6766 = ~n6764 & ~n6765;
  assign n6767 = ~n6761 & ~n6766;
  assign n6768 = n6761 & n6766;
  assign n6769 = ~n6767 & ~n6768;
  assign n6770 = g81 & g84;
  assign n6771 = g69 & g96;
  assign n6772 = g73 & g92;
  assign n6773 = ~n6771 & ~n6772;
  assign n6774 = n6771 & n6772;
  assign n6775 = ~n6773 & ~n6774;
  assign n6776 = ~n6770 & n6775;
  assign n6777 = n6770 & ~n6775;
  assign n6778 = ~n6776 & ~n6777;
  assign n6779 = ~n6769 & n6778;
  assign n6780 = n6769 & ~n6778;
  assign n6781 = ~n6779 & ~n6780;
  assign n6782 = ~n6760 & ~n6781;
  assign n6783 = ~n6769 & ~n6778;
  assign n6784 = ~n6782 & ~n6783;
  assign n6785 = g69 & g98;
  assign n6786 = g5 & n6785;
  assign n6787 = g80 & g86;
  assign n6788 = g81 & g85;
  assign n6789 = ~n6787 & n6788;
  assign n6790 = n6787 & ~n6788;
  assign n6791 = ~n6789 & ~n6790;
  assign n6792 = n6786 & ~n6791;
  assign n6793 = n6787 & n6788;
  assign n6794 = ~n6792 & ~n6793;
  assign n6795 = g68 & g97;
  assign n6796 = g75 & g90;
  assign n6797 = g76 & g89;
  assign n6798 = ~n6796 & n6797;
  assign n6799 = n6796 & ~n6797;
  assign n6800 = ~n6798 & ~n6799;
  assign n6801 = n6795 & ~n6800;
  assign n6802 = ~n6795 & n6800;
  assign n6803 = ~n6801 & ~n6802;
  assign n6804 = g78 & g87;
  assign n6805 = g71 & g94;
  assign n6806 = g77 & g88;
  assign n6807 = ~n6805 & n6806;
  assign n6808 = n6805 & ~n6806;
  assign n6809 = ~n6807 & ~n6808;
  assign n6810 = n6804 & ~n6809;
  assign n6811 = ~n6804 & n6809;
  assign n6812 = ~n6810 & ~n6811;
  assign n6813 = ~n6803 & n6812;
  assign n6814 = n6803 & ~n6812;
  assign n6815 = ~n6813 & ~n6814;
  assign n6816 = ~n6794 & ~n6815;
  assign n6817 = n6803 & n6812;
  assign n6818 = ~n6816 & ~n6817;
  assign n6819 = ~n6784 & ~n6818;
  assign n6820 = g81 & g83;
  assign n6821 = g80 & g84;
  assign n6822 = g73 & g91;
  assign n6823 = ~n6821 & ~n6822;
  assign n6824 = n6821 & n6822;
  assign n6825 = ~n6823 & ~n6824;
  assign n6826 = n6820 & n6825;
  assign n6827 = ~n6820 & ~n6825;
  assign n6828 = ~n6826 & ~n6827;
  assign n6829 = g71 & g93;
  assign n6830 = g75 & g89;
  assign n6831 = g74 & g90;
  assign n6832 = ~n6830 & n6831;
  assign n6833 = n6830 & ~n6831;
  assign n6834 = ~n6832 & ~n6833;
  assign n6835 = ~n6829 & ~n6834;
  assign n6836 = n6829 & n6834;
  assign n6837 = ~n6835 & ~n6836;
  assign n6838 = g70 & g94;
  assign n6839 = g68 & g96;
  assign n6840 = g67 & g97;
  assign n6841 = ~n6839 & n6840;
  assign n6842 = n6839 & ~n6840;
  assign n6843 = ~n6841 & ~n6842;
  assign n6844 = ~n6838 & ~n6843;
  assign n6845 = n6838 & n6843;
  assign n6846 = ~n6844 & ~n6845;
  assign n6847 = ~n6837 & n6846;
  assign n6848 = n6837 & ~n6846;
  assign n6849 = ~n6847 & ~n6848;
  assign n6850 = n6828 & n6849;
  assign n6851 = ~n6828 & ~n6849;
  assign n6852 = ~n6850 & ~n6851;
  assign n6853 = n6784 & n6818;
  assign n6854 = ~n6819 & ~n6853;
  assign n6855 = ~n6852 & n6854;
  assign n6856 = ~n6819 & ~n6855;
  assign n6857 = g79 & g84;
  assign n6858 = g78 & g85;
  assign n6859 = g72 & g91;
  assign n6860 = n6858 & ~n6859;
  assign n6861 = ~n6858 & n6859;
  assign n6862 = ~n6860 & ~n6861;
  assign n6863 = n6857 & n6862;
  assign n6864 = ~n6857 & ~n6862;
  assign n6865 = ~n6863 & ~n6864;
  assign n6866 = g69 & g94;
  assign n6867 = g76 & g87;
  assign n6868 = g77 & g86;
  assign n6869 = ~n6867 & n6868;
  assign n6870 = n6867 & ~n6868;
  assign n6871 = ~n6869 & ~n6870;
  assign n6872 = ~n6866 & ~n6871;
  assign n6873 = n6866 & n6871;
  assign n6874 = ~n6872 & ~n6873;
  assign n6875 = n6865 & ~n6874;
  assign n6876 = ~n6865 & n6874;
  assign n6877 = ~n6875 & ~n6876;
  assign n6878 = ~n6824 & ~n6826;
  assign n6879 = g80 & g83;
  assign n6880 = g73 & g90;
  assign n6881 = n6879 & ~n6880;
  assign n6882 = ~n6879 & n6880;
  assign n6883 = ~n6881 & ~n6882;
  assign n6884 = ~n6878 & n6883;
  assign n6885 = n6878 & ~n6883;
  assign n6886 = ~n6884 & ~n6885;
  assign n6887 = ~n6877 & n6886;
  assign n6888 = n6877 & ~n6886;
  assign n6889 = ~n6887 & ~n6888;
  assign n6890 = n6828 & ~n6849;
  assign n6891 = ~n6837 & ~n6846;
  assign n6892 = ~n6890 & ~n6891;
  assign n6893 = n6838 & ~n6843;
  assign n6894 = n6839 & n6840;
  assign n6895 = ~n6893 & ~n6894;
  assign n6896 = g71 & g92;
  assign n6897 = g74 & g89;
  assign n6898 = g75 & g88;
  assign n6899 = ~n6897 & n6898;
  assign n6900 = n6897 & ~n6898;
  assign n6901 = ~n6899 & ~n6900;
  assign n6902 = ~n6896 & ~n6901;
  assign n6903 = n6896 & n6901;
  assign n6904 = ~n6902 & ~n6903;
  assign n6905 = ~n6895 & n6904;
  assign n6906 = n6895 & ~n6904;
  assign n6907 = ~n6905 & ~n6906;
  assign n6908 = g70 & g93;
  assign n6909 = g67 & g96;
  assign n6910 = g68 & g95;
  assign n6911 = n6909 & n6910;
  assign n6912 = ~n6909 & ~n6910;
  assign n6913 = ~n6911 & ~n6912;
  assign n6914 = n6908 & n6913;
  assign n6915 = ~n6908 & ~n6913;
  assign n6916 = ~n6914 & ~n6915;
  assign n6917 = ~n6907 & n6916;
  assign n6918 = n6907 & ~n6916;
  assign n6919 = ~n6917 & ~n6918;
  assign n6920 = n6892 & n6919;
  assign n6921 = ~n6892 & ~n6919;
  assign n6922 = ~n6920 & ~n6921;
  assign n6923 = ~n6889 & ~n6922;
  assign n6924 = n6889 & n6922;
  assign n6925 = ~n6923 & ~n6924;
  assign n6926 = ~n6856 & ~n6925;
  assign n6927 = n6856 & n6925;
  assign n6928 = ~n6926 & ~n6927;
  assign n6929 = n6752 & ~n6757;
  assign n6930 = n6753 & n6754;
  assign n6931 = ~n6929 & ~n6930;
  assign n6932 = g67 & g98;
  assign n6933 = g3 & n6932;
  assign n6934 = n6770 & n6775;
  assign n6935 = ~n6774 & ~n6934;
  assign n6936 = ~n6933 & ~n6935;
  assign n6937 = n6933 & n6935;
  assign n6938 = ~n6936 & ~n6937;
  assign n6939 = n6931 & ~n6938;
  assign n6940 = ~n6931 & n6938;
  assign n6941 = ~n6939 & ~n6940;
  assign n6942 = g68 & g98;
  assign n6943 = g4 & n6942;
  assign n6944 = ~g3 & n6932;
  assign n6945 = g3 & ~n6932;
  assign n6946 = ~n6944 & ~n6945;
  assign n6947 = n6943 & ~n6946;
  assign n6948 = g74 & g92;
  assign n6949 = g70 & g96;
  assign n6950 = n6948 & n6949;
  assign n6951 = g82 & g84;
  assign n6952 = ~n6948 & ~n6949;
  assign n6953 = ~n6950 & ~n6952;
  assign n6954 = n6951 & n6953;
  assign n6955 = ~n6950 & ~n6954;
  assign n6956 = ~n6943 & ~n6946;
  assign n6957 = n6943 & n6946;
  assign n6958 = ~n6956 & ~n6957;
  assign n6959 = ~n6955 & ~n6958;
  assign n6960 = ~n6947 & ~n6959;
  assign n6961 = n6805 & n6806;
  assign n6962 = ~n6810 & ~n6961;
  assign n6963 = n6796 & n6797;
  assign n6964 = ~n6801 & ~n6963;
  assign n6965 = n6962 & ~n6964;
  assign n6966 = ~n6962 & n6964;
  assign n6967 = ~n6965 & ~n6966;
  assign n6968 = n6761 & ~n6766;
  assign n6969 = n6762 & n6763;
  assign n6970 = ~n6968 & ~n6969;
  assign n6971 = ~n6967 & ~n6970;
  assign n6972 = n6967 & n6970;
  assign n6973 = ~n6971 & ~n6972;
  assign n6974 = n6960 & n6973;
  assign n6975 = ~n6960 & ~n6973;
  assign n6976 = ~n6974 & ~n6975;
  assign n6977 = ~n6941 & ~n6976;
  assign n6978 = ~n6960 & n6973;
  assign n6979 = ~n6977 & ~n6978;
  assign n6980 = g78 & g86;
  assign n6981 = g72 & g92;
  assign n6982 = n6980 & ~n6981;
  assign n6983 = ~n6980 & n6981;
  assign n6984 = ~n6982 & ~n6983;
  assign n6985 = g79 & g85;
  assign n6986 = ~n6984 & ~n6985;
  assign n6987 = n6984 & n6985;
  assign n6988 = ~n6986 & ~n6987;
  assign n6989 = g76 & g88;
  assign n6990 = g77 & g87;
  assign n6991 = ~n6989 & n6990;
  assign n6992 = n6989 & ~n6990;
  assign n6993 = ~n6991 & ~n6992;
  assign n6994 = g69 & g95;
  assign n6995 = ~n6993 & ~n6994;
  assign n6996 = n6993 & n6994;
  assign n6997 = ~n6995 & ~n6996;
  assign n6998 = n6988 & ~n6997;
  assign n6999 = ~n6988 & n6997;
  assign n7000 = ~n6998 & ~n6999;
  assign n7001 = g73 & g93;
  assign n7002 = g78 & g88;
  assign n7003 = g79 & g87;
  assign n7004 = ~n7002 & n7003;
  assign n7005 = n7002 & ~n7003;
  assign n7006 = ~n7004 & ~n7005;
  assign n7007 = n7001 & ~n7006;
  assign n7008 = n7002 & n7003;
  assign n7009 = ~n7007 & ~n7008;
  assign n7010 = g76 & g90;
  assign n7011 = g71 & g95;
  assign n7012 = g75 & g91;
  assign n7013 = ~n7011 & n7012;
  assign n7014 = n7011 & ~n7012;
  assign n7015 = ~n7013 & ~n7014;
  assign n7016 = n7010 & ~n7015;
  assign n7017 = n7011 & n7012;
  assign n7018 = ~n7016 & ~n7017;
  assign n7019 = g72 & g94;
  assign n7020 = g77 & g89;
  assign n7021 = g69 & g97;
  assign n7022 = ~n7020 & n7021;
  assign n7023 = n7020 & ~n7021;
  assign n7024 = ~n7022 & ~n7023;
  assign n7025 = n7019 & ~n7024;
  assign n7026 = n7020 & n7021;
  assign n7027 = ~n7025 & ~n7026;
  assign n7028 = n7018 & ~n7027;
  assign n7029 = ~n7018 & n7027;
  assign n7030 = ~n7028 & ~n7029;
  assign n7031 = ~n7009 & ~n7030;
  assign n7032 = ~n7018 & ~n7027;
  assign n7033 = ~n7031 & ~n7032;
  assign n7034 = ~n7000 & ~n7033;
  assign n7035 = ~n6988 & ~n6997;
  assign n7036 = ~n7034 & ~n7035;
  assign n7037 = n6829 & ~n6834;
  assign n7038 = n6830 & n6831;
  assign n7039 = ~n7037 & ~n7038;
  assign n7040 = ~n6993 & n6994;
  assign n7041 = n6989 & n6990;
  assign n7042 = ~n7040 & ~n7041;
  assign n7043 = ~n7039 & n7042;
  assign n7044 = n7039 & ~n7042;
  assign n7045 = ~n7043 & ~n7044;
  assign n7046 = ~n6984 & n6985;
  assign n7047 = n6980 & n6981;
  assign n7048 = ~n7046 & ~n7047;
  assign n7049 = n7045 & ~n7048;
  assign n7050 = ~n7045 & n7048;
  assign n7051 = ~n7049 & ~n7050;
  assign n7052 = ~n6931 & ~n6938;
  assign n7053 = n6933 & ~n6935;
  assign n7054 = ~n7052 & ~n7053;
  assign n7055 = ~n6962 & ~n6964;
  assign n7056 = ~n6971 & ~n7055;
  assign n7057 = n7054 & ~n7056;
  assign n7058 = ~n7054 & n7056;
  assign n7059 = ~n7057 & ~n7058;
  assign n7060 = ~n7051 & ~n7059;
  assign n7061 = n7051 & n7059;
  assign n7062 = ~n7060 & ~n7061;
  assign n7063 = n7036 & ~n7062;
  assign n7064 = ~n7036 & n7062;
  assign n7065 = ~n7063 & ~n7064;
  assign n7066 = n6979 & n7065;
  assign n7067 = ~n6979 & ~n7065;
  assign n7068 = ~n7066 & ~n7067;
  assign n7069 = ~n6928 & ~n7068;
  assign n7070 = ~n6856 & n6925;
  assign n7071 = ~n7069 & ~n7070;
  assign n7072 = n6857 & ~n6862;
  assign n7073 = n6858 & n6859;
  assign n7074 = ~n7072 & ~n7073;
  assign n7075 = g73 & g89;
  assign n7076 = n6866 & ~n6871;
  assign n7077 = n6867 & n6868;
  assign n7078 = ~n7076 & ~n7077;
  assign n7079 = n7075 & ~n7078;
  assign n7080 = ~n7075 & n7078;
  assign n7081 = ~n7079 & ~n7080;
  assign n7082 = n7074 & n7081;
  assign n7083 = ~n7074 & ~n7081;
  assign n7084 = ~n7082 & ~n7083;
  assign n7085 = ~n7039 & ~n7042;
  assign n7086 = ~n7045 & ~n7048;
  assign n7087 = ~n7085 & ~n7086;
  assign n7088 = ~n6878 & ~n6883;
  assign n7089 = n6879 & n6880;
  assign n7090 = ~n7088 & ~n7089;
  assign n7091 = n7087 & ~n7090;
  assign n7092 = ~n7087 & n7090;
  assign n7093 = ~n7091 & ~n7092;
  assign n7094 = ~n7084 & ~n7093;
  assign n7095 = n7084 & n7093;
  assign n7096 = ~n7094 & ~n7095;
  assign n7097 = ~n6877 & ~n6886;
  assign n7098 = ~n6865 & ~n6874;
  assign n7099 = ~n7097 & ~n7098;
  assign n7100 = ~n7054 & ~n7056;
  assign n7101 = ~n7060 & ~n7100;
  assign n7102 = ~n7099 & ~n7101;
  assign n7103 = n7099 & n7101;
  assign n7104 = ~n7102 & ~n7103;
  assign n7105 = ~n7096 & n7104;
  assign n7106 = n7096 & ~n7104;
  assign n7107 = ~n7105 & ~n7106;
  assign n7108 = ~n6979 & n7065;
  assign n7109 = ~n7064 & ~n7108;
  assign n7110 = ~n6892 & n6919;
  assign n7111 = ~n6923 & ~n7110;
  assign n7112 = ~n6695 & n6697;
  assign n7113 = n6695 & ~n6697;
  assign n7114 = ~n7112 & ~n7113;
  assign n7115 = g69 & g93;
  assign n7116 = g76 & g86;
  assign n7117 = g77 & g85;
  assign n7118 = ~n7116 & n7117;
  assign n7119 = n7116 & ~n7117;
  assign n7120 = ~n7118 & ~n7119;
  assign n7121 = ~n7115 & ~n7120;
  assign n7122 = n7115 & n7120;
  assign n7123 = ~n7121 & ~n7122;
  assign n7124 = ~n6700 & n6705;
  assign n7125 = ~n6706 & ~n7124;
  assign n7126 = ~n7123 & ~n7125;
  assign n7127 = n7123 & n7125;
  assign n7128 = ~n7126 & ~n7127;
  assign n7129 = ~n7114 & n7128;
  assign n7130 = n7114 & ~n7128;
  assign n7131 = ~n7129 & ~n7130;
  assign n7132 = ~n6895 & ~n6904;
  assign n7133 = ~n6917 & ~n7132;
  assign n7134 = n6709 & n6714;
  assign n7135 = ~n6709 & ~n6714;
  assign n7136 = ~n7134 & ~n7135;
  assign n7137 = n6896 & ~n6901;
  assign n7138 = n6897 & n6898;
  assign n7139 = ~n7137 & ~n7138;
  assign n7140 = ~n6911 & ~n6914;
  assign n7141 = n7139 & ~n7140;
  assign n7142 = ~n7139 & n7140;
  assign n7143 = ~n7141 & ~n7142;
  assign n7144 = ~n7136 & n7143;
  assign n7145 = n7136 & ~n7143;
  assign n7146 = ~n7144 & ~n7145;
  assign n7147 = n7133 & ~n7146;
  assign n7148 = ~n7133 & n7146;
  assign n7149 = ~n7147 & ~n7148;
  assign n7150 = n7131 & ~n7149;
  assign n7151 = ~n7131 & n7149;
  assign n7152 = ~n7150 & ~n7151;
  assign n7153 = ~n7111 & ~n7152;
  assign n7154 = n7111 & n7152;
  assign n7155 = ~n7153 & ~n7154;
  assign n7156 = n7109 & n7155;
  assign n7157 = ~n7109 & ~n7155;
  assign n7158 = ~n7156 & ~n7157;
  assign n7159 = ~n7107 & n7158;
  assign n7160 = n7107 & ~n7158;
  assign n7161 = ~n7159 & ~n7160;
  assign n7162 = ~n7071 & ~n7161;
  assign n7163 = ~n7107 & ~n7158;
  assign n7164 = ~n7162 & ~n7163;
  assign n7165 = ~n7109 & n7155;
  assign n7166 = ~n7153 & ~n7165;
  assign n7167 = ~n7074 & n7081;
  assign n7168 = ~n7079 & ~n7167;
  assign n7169 = n6610 & n6615;
  assign n7170 = ~n6610 & ~n6615;
  assign n7171 = ~n7169 & ~n7170;
  assign n7172 = ~n6622 & n6624;
  assign n7173 = n6622 & ~n6624;
  assign n7174 = ~n7172 & ~n7173;
  assign n7175 = ~n7171 & n7174;
  assign n7176 = n7171 & ~n7174;
  assign n7177 = ~n7175 & ~n7176;
  assign n7178 = ~n7168 & n7177;
  assign n7179 = n7168 & ~n7177;
  assign n7180 = ~n7178 & ~n7179;
  assign n7181 = ~n6642 & ~n6647;
  assign n7182 = n6642 & n6647;
  assign n7183 = ~n7181 & ~n7182;
  assign n7184 = ~n6601 & n6606;
  assign n7185 = ~n6607 & ~n7184;
  assign n7186 = n7115 & ~n7120;
  assign n7187 = n7116 & n7117;
  assign n7188 = ~n7186 & ~n7187;
  assign n7189 = n7185 & ~n7188;
  assign n7190 = ~n7185 & n7188;
  assign n7191 = ~n7189 & ~n7190;
  assign n7192 = n7183 & n7191;
  assign n7193 = ~n7183 & ~n7191;
  assign n7194 = ~n7192 & ~n7193;
  assign n7195 = n7180 & ~n7194;
  assign n7196 = ~n7180 & n7194;
  assign n7197 = ~n7195 & ~n7196;
  assign n7198 = ~n7087 & ~n7090;
  assign n7199 = ~n7094 & ~n7198;
  assign n7200 = n7197 & ~n7199;
  assign n7201 = ~n7197 & n7199;
  assign n7202 = ~n7200 & ~n7201;
  assign n7203 = n7096 & n7104;
  assign n7204 = ~n7102 & ~n7203;
  assign n7205 = ~n7136 & ~n7143;
  assign n7206 = ~n7139 & ~n7140;
  assign n7207 = ~n7205 & ~n7206;
  assign n7208 = ~n7114 & ~n7128;
  assign n7209 = ~n7123 & n7125;
  assign n7210 = ~n7208 & ~n7209;
  assign n7211 = ~n6699 & n6720;
  assign n7212 = n6699 & ~n6720;
  assign n7213 = ~n7211 & ~n7212;
  assign n7214 = n7210 & ~n7213;
  assign n7215 = ~n7210 & n7213;
  assign n7216 = ~n7214 & ~n7215;
  assign n7217 = ~n7207 & ~n7216;
  assign n7218 = n7207 & n7216;
  assign n7219 = ~n7217 & ~n7218;
  assign n7220 = ~n7131 & ~n7149;
  assign n7221 = ~n7133 & ~n7146;
  assign n7222 = ~n7220 & ~n7221;
  assign n7223 = n7219 & ~n7222;
  assign n7224 = ~n7219 & n7222;
  assign n7225 = ~n7223 & ~n7224;
  assign n7226 = n7204 & n7225;
  assign n7227 = ~n7204 & ~n7225;
  assign n7228 = ~n7226 & ~n7227;
  assign n7229 = n7202 & ~n7228;
  assign n7230 = ~n7202 & n7228;
  assign n7231 = ~n7229 & ~n7230;
  assign n7232 = n7166 & ~n7231;
  assign n7233 = ~n7166 & n7231;
  assign n7234 = ~n7232 & ~n7233;
  assign n7235 = ~n7164 & ~n7234;
  assign n7236 = g74 & g93;
  assign n7237 = g80 & g87;
  assign n7238 = n7236 & n7237;
  assign n7239 = g81 & g86;
  assign n7240 = ~n7236 & ~n7237;
  assign n7241 = ~n7238 & ~n7240;
  assign n7242 = n7239 & n7241;
  assign n7243 = ~n7238 & ~n7242;
  assign n7244 = g70 & g97;
  assign n7245 = g73 & g94;
  assign n7246 = n7244 & n7245;
  assign n7247 = g79 & g88;
  assign n7248 = ~n7244 & ~n7245;
  assign n7249 = ~n7246 & ~n7248;
  assign n7250 = n7247 & n7249;
  assign n7251 = ~n7246 & ~n7250;
  assign n7252 = n7243 & ~n7251;
  assign n7253 = ~n7243 & n7251;
  assign n7254 = ~n7252 & ~n7253;
  assign n7255 = n6951 & ~n6953;
  assign n7256 = ~n6951 & n6953;
  assign n7257 = ~n7255 & ~n7256;
  assign n7258 = n7254 & ~n7257;
  assign n7259 = ~n7254 & n7257;
  assign n7260 = ~n7258 & ~n7259;
  assign n7261 = g76 & g91;
  assign n7262 = g75 & g92;
  assign n7263 = g71 & g96;
  assign n7264 = n7262 & ~n7263;
  assign n7265 = ~n7262 & n7263;
  assign n7266 = ~n7264 & ~n7265;
  assign n7267 = n7261 & ~n7266;
  assign n7268 = n7262 & n7263;
  assign n7269 = ~n7267 & ~n7268;
  assign n7270 = ~g4 & n6942;
  assign n7271 = g4 & ~n6942;
  assign n7272 = ~n7270 & ~n7271;
  assign n7273 = g78 & g89;
  assign n7274 = g72 & g95;
  assign n7275 = g77 & g90;
  assign n7276 = ~n7274 & n7275;
  assign n7277 = n7274 & ~n7275;
  assign n7278 = ~n7276 & ~n7277;
  assign n7279 = n7273 & ~n7278;
  assign n7280 = n7274 & n7275;
  assign n7281 = ~n7279 & ~n7280;
  assign n7282 = n7272 & ~n7281;
  assign n7283 = ~n7272 & n7281;
  assign n7284 = ~n7282 & ~n7283;
  assign n7285 = ~n7269 & n7284;
  assign n7286 = n7269 & ~n7284;
  assign n7287 = ~n7285 & ~n7286;
  assign n7288 = ~n7261 & ~n7266;
  assign n7289 = n7261 & n7266;
  assign n7290 = ~n7288 & ~n7289;
  assign n7291 = g80 & g88;
  assign n7292 = g74 & g94;
  assign n7293 = g71 & g97;
  assign n7294 = ~n7292 & n7293;
  assign n7295 = n7292 & ~n7293;
  assign n7296 = ~n7294 & ~n7295;
  assign n7297 = n7291 & ~n7296;
  assign n7298 = n7292 & n7293;
  assign n7299 = ~n7297 & ~n7298;
  assign n7300 = ~n7239 & n7241;
  assign n7301 = n7239 & ~n7241;
  assign n7302 = ~n7300 & ~n7301;
  assign n7303 = ~n7299 & n7302;
  assign n7304 = n7299 & ~n7302;
  assign n7305 = ~n7303 & ~n7304;
  assign n7306 = ~n7290 & ~n7305;
  assign n7307 = ~n7299 & ~n7302;
  assign n7308 = ~n7306 & ~n7307;
  assign n7309 = ~n7287 & n7308;
  assign n7310 = n7287 & ~n7308;
  assign n7311 = ~n7309 & ~n7310;
  assign n7312 = ~n7260 & ~n7311;
  assign n7313 = ~n7287 & ~n7308;
  assign n7314 = ~n7312 & ~n7313;
  assign n7315 = ~n6760 & n6781;
  assign n7316 = n6760 & ~n6781;
  assign n7317 = ~n7315 & ~n7316;
  assign n7318 = g82 & g86;
  assign n7319 = g75 & g93;
  assign n7320 = g81 & g87;
  assign n7321 = ~n7319 & n7320;
  assign n7322 = n7319 & ~n7320;
  assign n7323 = ~n7321 & ~n7322;
  assign n7324 = n7318 & ~n7323;
  assign n7325 = n7319 & n7320;
  assign n7326 = ~n7324 & ~n7325;
  assign n7327 = g72 & g96;
  assign n7328 = g76 & g92;
  assign n7329 = n7327 & n7328;
  assign n7330 = g77 & g91;
  assign n7331 = ~n7327 & ~n7328;
  assign n7332 = ~n7329 & ~n7331;
  assign n7333 = n7330 & n7332;
  assign n7334 = ~n7329 & ~n7333;
  assign n7335 = g73 & g95;
  assign n7336 = g78 & g90;
  assign n7337 = n7335 & n7336;
  assign n7338 = g79 & g89;
  assign n7339 = ~n7335 & ~n7336;
  assign n7340 = ~n7337 & ~n7339;
  assign n7341 = n7338 & n7340;
  assign n7342 = ~n7337 & ~n7341;
  assign n7343 = n7334 & ~n7342;
  assign n7344 = ~n7334 & n7342;
  assign n7345 = ~n7343 & ~n7344;
  assign n7346 = ~n7326 & ~n7345;
  assign n7347 = ~n7334 & ~n7342;
  assign n7348 = ~n7346 & ~n7347;
  assign n7349 = g82 & g85;
  assign n7350 = g5 & ~n6785;
  assign n7351 = ~g5 & n6785;
  assign n7352 = ~n7350 & ~n7351;
  assign n7353 = n7349 & ~n7352;
  assign n7354 = g70 & g98;
  assign n7355 = g6 & n7354;
  assign n7356 = ~n7349 & n7352;
  assign n7357 = ~n7353 & ~n7356;
  assign n7358 = n7355 & n7357;
  assign n7359 = ~n7353 & ~n7358;
  assign n7360 = ~n6786 & ~n6791;
  assign n7361 = n6786 & n6791;
  assign n7362 = ~n7360 & ~n7361;
  assign n7363 = n7359 & ~n7362;
  assign n7364 = ~n7359 & n7362;
  assign n7365 = ~n7363 & ~n7364;
  assign n7366 = ~n7348 & ~n7365;
  assign n7367 = ~n7359 & ~n7362;
  assign n7368 = ~n7366 & ~n7367;
  assign n7369 = n7317 & ~n7368;
  assign n7370 = ~n7317 & n7368;
  assign n7371 = ~n7369 & ~n7370;
  assign n7372 = ~n7314 & ~n7371;
  assign n7373 = ~n7317 & ~n7368;
  assign n7374 = ~n7372 & ~n7373;
  assign n7375 = n6941 & ~n6976;
  assign n7376 = ~n6941 & n6976;
  assign n7377 = ~n7375 & ~n7376;
  assign n7378 = n6852 & ~n6854;
  assign n7379 = ~n6855 & ~n7378;
  assign n7380 = ~n7377 & ~n7379;
  assign n7381 = n7377 & n7379;
  assign n7382 = ~n7380 & ~n7381;
  assign n7383 = ~n7374 & n7382;
  assign n7384 = n7374 & ~n7382;
  assign n7385 = ~n7383 & ~n7384;
  assign n7386 = ~n7254 & ~n7257;
  assign n7387 = ~n7243 & ~n7251;
  assign n7388 = ~n7386 & ~n7387;
  assign n7389 = ~n7009 & n7030;
  assign n7390 = n7009 & ~n7030;
  assign n7391 = ~n7389 & ~n7390;
  assign n7392 = ~n7388 & ~n7391;
  assign n7393 = ~n6794 & n6815;
  assign n7394 = n6794 & ~n6815;
  assign n7395 = ~n7393 & ~n7394;
  assign n7396 = ~n7388 & n7391;
  assign n7397 = n7388 & ~n7391;
  assign n7398 = ~n7396 & ~n7397;
  assign n7399 = ~n7395 & ~n7398;
  assign n7400 = ~n7392 & ~n7399;
  assign n7401 = ~n7001 & ~n7006;
  assign n7402 = n7001 & n7006;
  assign n7403 = ~n7401 & ~n7402;
  assign n7404 = ~n7010 & n7015;
  assign n7405 = ~n7016 & ~n7404;
  assign n7406 = ~n7403 & n7405;
  assign n7407 = n7019 & n7024;
  assign n7408 = ~n7019 & ~n7024;
  assign n7409 = ~n7407 & ~n7408;
  assign n7410 = ~n7403 & ~n7405;
  assign n7411 = n7403 & n7405;
  assign n7412 = ~n7410 & ~n7411;
  assign n7413 = ~n7409 & ~n7412;
  assign n7414 = ~n7406 & ~n7413;
  assign n7415 = n6955 & ~n6958;
  assign n7416 = ~n6955 & n6958;
  assign n7417 = ~n7415 & ~n7416;
  assign n7418 = ~n7269 & ~n7284;
  assign n7419 = ~n7272 & ~n7281;
  assign n7420 = ~n7418 & ~n7419;
  assign n7421 = ~n7417 & n7420;
  assign n7422 = n7417 & ~n7420;
  assign n7423 = ~n7421 & ~n7422;
  assign n7424 = ~n7414 & ~n7423;
  assign n7425 = ~n7417 & ~n7420;
  assign n7426 = ~n7424 & ~n7425;
  assign n7427 = n7000 & ~n7033;
  assign n7428 = ~n7000 & n7033;
  assign n7429 = ~n7427 & ~n7428;
  assign n7430 = ~n7426 & n7429;
  assign n7431 = n7426 & ~n7429;
  assign n7432 = ~n7430 & ~n7431;
  assign n7433 = ~n7400 & n7432;
  assign n7434 = n7400 & ~n7432;
  assign n7435 = ~n7433 & ~n7434;
  assign n7436 = ~n7348 & n7365;
  assign n7437 = n7348 & ~n7365;
  assign n7438 = ~n7436 & ~n7437;
  assign n7439 = ~n7247 & n7249;
  assign n7440 = n7247 & ~n7249;
  assign n7441 = ~n7439 & ~n7440;
  assign n7442 = ~n7273 & n7278;
  assign n7443 = ~n7279 & ~n7442;
  assign n7444 = ~n7441 & n7443;
  assign n7445 = n7441 & ~n7443;
  assign n7446 = ~n7444 & ~n7445;
  assign n7447 = n7355 & ~n7357;
  assign n7448 = ~n7355 & n7357;
  assign n7449 = ~n7447 & ~n7448;
  assign n7450 = n7446 & ~n7449;
  assign n7451 = ~n7444 & ~n7450;
  assign n7452 = n7409 & n7412;
  assign n7453 = ~n7413 & ~n7452;
  assign n7454 = ~n7451 & ~n7453;
  assign n7455 = n7451 & n7453;
  assign n7456 = ~n7454 & ~n7455;
  assign n7457 = ~n7438 & ~n7456;
  assign n7458 = ~n7451 & n7453;
  assign n7459 = ~n7457 & ~n7458;
  assign n7460 = n7414 & n7423;
  assign n7461 = ~n7424 & ~n7460;
  assign n7462 = ~n7395 & n7398;
  assign n7463 = n7395 & ~n7398;
  assign n7464 = ~n7462 & ~n7463;
  assign n7465 = n7461 & n7464;
  assign n7466 = ~n7461 & ~n7464;
  assign n7467 = ~n7465 & ~n7466;
  assign n7468 = ~n7459 & ~n7467;
  assign n7469 = n7461 & ~n7464;
  assign n7470 = ~n7468 & ~n7469;
  assign n7471 = ~n7435 & n7470;
  assign n7472 = n7435 & ~n7470;
  assign n7473 = ~n7471 & ~n7472;
  assign n7474 = n7385 & ~n7473;
  assign n7475 = ~n7385 & n7473;
  assign n7476 = ~n7474 & ~n7475;
  assign n7477 = n7314 & ~n7371;
  assign n7478 = ~n7314 & n7371;
  assign n7479 = ~n7477 & ~n7478;
  assign n7480 = n7459 & ~n7467;
  assign n7481 = ~n7459 & n7467;
  assign n7482 = ~n7480 & ~n7481;
  assign n7483 = ~n7479 & ~n7482;
  assign n7484 = ~n7260 & n7311;
  assign n7485 = n7260 & ~n7311;
  assign n7486 = ~n7484 & ~n7485;
  assign n7487 = ~n7291 & n7296;
  assign n7488 = ~n7297 & ~n7487;
  assign n7489 = ~n7330 & ~n7332;
  assign n7490 = ~n7333 & ~n7489;
  assign n7491 = ~n7338 & n7340;
  assign n7492 = n7338 & ~n7340;
  assign n7493 = ~n7491 & ~n7492;
  assign n7494 = n7490 & n7493;
  assign n7495 = ~n7490 & ~n7493;
  assign n7496 = ~n7494 & ~n7495;
  assign n7497 = n7488 & ~n7496;
  assign n7498 = n7490 & ~n7493;
  assign n7499 = ~n7497 & ~n7498;
  assign n7500 = g71 & g98;
  assign n7501 = g7 & n7500;
  assign n7502 = ~g6 & ~n7354;
  assign n7503 = ~n7355 & ~n7502;
  assign n7504 = n7501 & n7503;
  assign n7505 = g73 & g96;
  assign n7506 = g77 & g92;
  assign n7507 = n7505 & n7506;
  assign n7508 = g78 & g91;
  assign n7509 = ~n7505 & ~n7506;
  assign n7510 = ~n7507 & ~n7509;
  assign n7511 = n7508 & n7510;
  assign n7512 = ~n7507 & ~n7511;
  assign n7513 = ~n7501 & ~n7503;
  assign n7514 = ~n7504 & ~n7513;
  assign n7515 = ~n7512 & n7514;
  assign n7516 = ~n7504 & ~n7515;
  assign n7517 = n7499 & ~n7516;
  assign n7518 = ~n7499 & n7516;
  assign n7519 = ~n7517 & ~n7518;
  assign n7520 = n7318 & n7323;
  assign n7521 = ~n7318 & ~n7323;
  assign n7522 = ~n7520 & ~n7521;
  assign n7523 = g81 & g88;
  assign n7524 = g75 & g94;
  assign n7525 = g72 & g97;
  assign n7526 = ~n7524 & n7525;
  assign n7527 = n7524 & ~n7525;
  assign n7528 = ~n7526 & ~n7527;
  assign n7529 = n7523 & ~n7528;
  assign n7530 = n7524 & n7525;
  assign n7531 = ~n7529 & ~n7530;
  assign n7532 = g80 & g89;
  assign n7533 = g74 & g95;
  assign n7534 = g79 & g90;
  assign n7535 = ~n7533 & n7534;
  assign n7536 = n7533 & ~n7534;
  assign n7537 = ~n7535 & ~n7536;
  assign n7538 = n7532 & ~n7537;
  assign n7539 = n7533 & n7534;
  assign n7540 = ~n7538 & ~n7539;
  assign n7541 = ~n7531 & n7540;
  assign n7542 = n7531 & ~n7540;
  assign n7543 = ~n7541 & ~n7542;
  assign n7544 = ~n7522 & ~n7543;
  assign n7545 = ~n7531 & ~n7540;
  assign n7546 = ~n7544 & ~n7545;
  assign n7547 = ~n7519 & ~n7546;
  assign n7548 = ~n7499 & ~n7516;
  assign n7549 = ~n7547 & ~n7548;
  assign n7550 = n7486 & ~n7549;
  assign n7551 = ~n7486 & n7549;
  assign n7552 = ~n7550 & ~n7551;
  assign n7553 = ~n7512 & ~n7514;
  assign n7554 = n7512 & n7514;
  assign n7555 = ~n7553 & ~n7554;
  assign n7556 = ~g7 & n7500;
  assign n7557 = g7 & ~n7500;
  assign n7558 = ~n7556 & ~n7557;
  assign n7559 = g76 & g93;
  assign n7560 = g82 & g87;
  assign n7561 = n7559 & ~n7560;
  assign n7562 = ~n7559 & n7560;
  assign n7563 = ~n7561 & ~n7562;
  assign n7564 = ~n7558 & ~n7563;
  assign n7565 = n7559 & n7560;
  assign n7566 = ~n7564 & ~n7565;
  assign n7567 = g72 & g98;
  assign n7568 = g8 & n7567;
  assign n7569 = g81 & g89;
  assign n7570 = g75 & g95;
  assign n7571 = g80 & g90;
  assign n7572 = ~n7570 & n7571;
  assign n7573 = n7570 & ~n7571;
  assign n7574 = ~n7572 & ~n7573;
  assign n7575 = n7569 & ~n7574;
  assign n7576 = n7570 & n7571;
  assign n7577 = ~n7575 & ~n7576;
  assign n7578 = n7568 & ~n7577;
  assign n7579 = g82 & g88;
  assign n7580 = g73 & g97;
  assign n7581 = g76 & g94;
  assign n7582 = ~n7580 & n7581;
  assign n7583 = n7580 & ~n7581;
  assign n7584 = ~n7582 & ~n7583;
  assign n7585 = n7579 & ~n7584;
  assign n7586 = n7580 & n7581;
  assign n7587 = ~n7585 & ~n7586;
  assign n7588 = ~n7568 & n7577;
  assign n7589 = ~n7578 & ~n7588;
  assign n7590 = ~n7587 & n7589;
  assign n7591 = ~n7578 & ~n7590;
  assign n7592 = n7566 & ~n7591;
  assign n7593 = ~n7566 & n7591;
  assign n7594 = ~n7592 & ~n7593;
  assign n7595 = ~n7555 & ~n7594;
  assign n7596 = ~n7566 & ~n7591;
  assign n7597 = ~n7595 & ~n7596;
  assign n7598 = ~n7326 & n7345;
  assign n7599 = n7326 & ~n7345;
  assign n7600 = ~n7598 & ~n7599;
  assign n7601 = ~n7290 & n7305;
  assign n7602 = n7290 & ~n7305;
  assign n7603 = ~n7601 & ~n7602;
  assign n7604 = ~n7600 & n7603;
  assign n7605 = n7600 & ~n7603;
  assign n7606 = ~n7604 & ~n7605;
  assign n7607 = ~n7597 & ~n7606;
  assign n7608 = ~n7600 & ~n7603;
  assign n7609 = ~n7607 & ~n7608;
  assign n7610 = ~n7552 & ~n7609;
  assign n7611 = ~n7486 & ~n7549;
  assign n7612 = ~n7610 & ~n7611;
  assign n7613 = n7479 & n7482;
  assign n7614 = ~n7483 & ~n7613;
  assign n7615 = ~n7612 & n7614;
  assign n7616 = ~n7483 & ~n7615;
  assign n7617 = n7476 & n7616;
  assign n7618 = ~n7377 & n7379;
  assign n7619 = ~n7374 & ~n7382;
  assign n7620 = ~n7618 & ~n7619;
  assign n7621 = ~n7400 & ~n7432;
  assign n7622 = ~n7426 & ~n7429;
  assign n7623 = ~n7621 & ~n7622;
  assign n7624 = ~n7620 & ~n7623;
  assign n7625 = n7620 & n7623;
  assign n7626 = ~n7624 & ~n7625;
  assign n7627 = n6928 & ~n7068;
  assign n7628 = ~n6928 & n7068;
  assign n7629 = ~n7627 & ~n7628;
  assign n7630 = ~n7626 & ~n7629;
  assign n7631 = n7626 & n7629;
  assign n7632 = ~n7630 & ~n7631;
  assign n7633 = ~n7385 & ~n7473;
  assign n7634 = ~n7435 & ~n7470;
  assign n7635 = ~n7633 & ~n7634;
  assign n7636 = n7632 & n7635;
  assign n7637 = ~n7617 & ~n7636;
  assign n7638 = n7597 & ~n7606;
  assign n7639 = ~n7597 & n7606;
  assign n7640 = ~n7638 & ~n7639;
  assign n7641 = ~n7508 & ~n7510;
  assign n7642 = ~n7511 & ~n7641;
  assign n7643 = g77 & g93;
  assign n7644 = g8 & ~n7567;
  assign n7645 = ~g8 & n7567;
  assign n7646 = ~n7644 & ~n7645;
  assign n7647 = n7643 & ~n7646;
  assign n7648 = g73 & g98;
  assign n7649 = g9 & n7648;
  assign n7650 = ~n7643 & n7646;
  assign n7651 = ~n7647 & ~n7650;
  assign n7652 = n7649 & n7651;
  assign n7653 = ~n7647 & ~n7652;
  assign n7654 = n7642 & ~n7653;
  assign n7655 = n7558 & ~n7563;
  assign n7656 = ~n7558 & n7563;
  assign n7657 = ~n7655 & ~n7656;
  assign n7658 = ~n7642 & ~n7653;
  assign n7659 = n7642 & n7653;
  assign n7660 = ~n7658 & ~n7659;
  assign n7661 = ~n7657 & ~n7660;
  assign n7662 = ~n7654 & ~n7661;
  assign n7663 = ~n7587 & ~n7589;
  assign n7664 = n7587 & n7589;
  assign n7665 = ~n7663 & ~n7664;
  assign n7666 = g82 & g89;
  assign n7667 = g81 & g90;
  assign n7668 = g76 & g95;
  assign n7669 = n7667 & ~n7668;
  assign n7670 = ~n7667 & n7668;
  assign n7671 = ~n7669 & ~n7670;
  assign n7672 = n7666 & ~n7671;
  assign n7673 = n7667 & n7668;
  assign n7674 = ~n7672 & ~n7673;
  assign n7675 = g80 & g91;
  assign n7676 = g75 & g96;
  assign n7677 = g79 & g92;
  assign n7678 = ~n7676 & n7677;
  assign n7679 = n7676 & ~n7677;
  assign n7680 = ~n7678 & ~n7679;
  assign n7681 = n7675 & ~n7680;
  assign n7682 = n7676 & n7677;
  assign n7683 = ~n7681 & ~n7682;
  assign n7684 = g77 & g94;
  assign n7685 = g74 & g97;
  assign n7686 = n7684 & n7685;
  assign n7687 = g78 & g93;
  assign n7688 = ~n7684 & ~n7685;
  assign n7689 = ~n7686 & ~n7688;
  assign n7690 = n7687 & n7689;
  assign n7691 = ~n7686 & ~n7690;
  assign n7692 = n7683 & ~n7691;
  assign n7693 = ~n7683 & n7691;
  assign n7694 = ~n7692 & ~n7693;
  assign n7695 = ~n7674 & ~n7694;
  assign n7696 = ~n7683 & ~n7691;
  assign n7697 = ~n7695 & ~n7696;
  assign n7698 = g74 & g96;
  assign n7699 = g78 & g92;
  assign n7700 = ~n7698 & n7699;
  assign n7701 = n7698 & ~n7699;
  assign n7702 = ~n7700 & ~n7701;
  assign n7703 = g79 & g91;
  assign n7704 = ~n7702 & n7703;
  assign n7705 = n7702 & ~n7703;
  assign n7706 = ~n7704 & ~n7705;
  assign n7707 = n7569 & n7574;
  assign n7708 = ~n7569 & ~n7574;
  assign n7709 = ~n7707 & ~n7708;
  assign n7710 = ~n7579 & ~n7584;
  assign n7711 = n7579 & n7584;
  assign n7712 = ~n7710 & ~n7711;
  assign n7713 = ~n7709 & n7712;
  assign n7714 = n7709 & ~n7712;
  assign n7715 = ~n7713 & ~n7714;
  assign n7716 = n7706 & ~n7715;
  assign n7717 = ~n7709 & ~n7712;
  assign n7718 = ~n7716 & ~n7717;
  assign n7719 = n7697 & ~n7718;
  assign n7720 = ~n7697 & n7718;
  assign n7721 = ~n7719 & ~n7720;
  assign n7722 = ~n7665 & ~n7721;
  assign n7723 = ~n7697 & ~n7718;
  assign n7724 = ~n7722 & ~n7723;
  assign n7725 = ~n7662 & ~n7724;
  assign n7726 = n7555 & ~n7594;
  assign n7727 = ~n7555 & n7594;
  assign n7728 = ~n7726 & ~n7727;
  assign n7729 = n7662 & n7724;
  assign n7730 = ~n7725 & ~n7729;
  assign n7731 = ~n7728 & n7730;
  assign n7732 = ~n7725 & ~n7731;
  assign n7733 = ~n7640 & ~n7732;
  assign n7734 = ~n7519 & n7546;
  assign n7735 = n7519 & ~n7546;
  assign n7736 = ~n7734 & ~n7735;
  assign n7737 = n7488 & n7496;
  assign n7738 = ~n7488 & ~n7496;
  assign n7739 = ~n7737 & ~n7738;
  assign n7740 = n7532 & n7537;
  assign n7741 = ~n7532 & ~n7537;
  assign n7742 = ~n7740 & ~n7741;
  assign n7743 = n7698 & n7699;
  assign n7744 = ~n7704 & ~n7743;
  assign n7745 = ~n7523 & ~n7528;
  assign n7746 = n7523 & n7528;
  assign n7747 = ~n7745 & ~n7746;
  assign n7748 = ~n7744 & n7747;
  assign n7749 = n7744 & ~n7747;
  assign n7750 = ~n7748 & ~n7749;
  assign n7751 = ~n7742 & ~n7750;
  assign n7752 = ~n7744 & ~n7747;
  assign n7753 = ~n7751 & ~n7752;
  assign n7754 = n7522 & ~n7543;
  assign n7755 = ~n7522 & n7543;
  assign n7756 = ~n7754 & ~n7755;
  assign n7757 = n7753 & ~n7756;
  assign n7758 = ~n7753 & n7756;
  assign n7759 = ~n7757 & ~n7758;
  assign n7760 = ~n7739 & ~n7759;
  assign n7761 = ~n7753 & ~n7756;
  assign n7762 = ~n7760 & ~n7761;
  assign n7763 = ~n7446 & ~n7449;
  assign n7764 = n7446 & n7449;
  assign n7765 = ~n7763 & ~n7764;
  assign n7766 = ~n7762 & ~n7765;
  assign n7767 = n7762 & n7765;
  assign n7768 = ~n7766 & ~n7767;
  assign n7769 = ~n7736 & ~n7768;
  assign n7770 = n7736 & n7768;
  assign n7771 = ~n7769 & ~n7770;
  assign n7772 = n7640 & n7732;
  assign n7773 = ~n7733 & ~n7772;
  assign n7774 = ~n7771 & n7773;
  assign n7775 = ~n7733 & ~n7774;
  assign n7776 = ~n7736 & n7768;
  assign n7777 = ~n7766 & ~n7776;
  assign n7778 = n7438 & ~n7456;
  assign n7779 = ~n7438 & n7456;
  assign n7780 = ~n7778 & ~n7779;
  assign n7781 = n7777 & ~n7780;
  assign n7782 = ~n7777 & n7780;
  assign n7783 = ~n7781 & ~n7782;
  assign n7784 = ~n7552 & n7609;
  assign n7785 = n7552 & ~n7609;
  assign n7786 = ~n7784 & ~n7785;
  assign n7787 = ~n7783 & n7786;
  assign n7788 = n7783 & ~n7786;
  assign n7789 = ~n7787 & ~n7788;
  assign n7790 = ~n7775 & ~n7789;
  assign n7791 = n7612 & n7614;
  assign n7792 = ~n7612 & ~n7614;
  assign n7793 = ~n7791 & ~n7792;
  assign n7794 = ~n7783 & ~n7786;
  assign n7795 = ~n7777 & ~n7780;
  assign n7796 = ~n7794 & ~n7795;
  assign n7797 = n7793 & n7796;
  assign n7798 = n7790 & ~n7797;
  assign n7799 = ~n7793 & ~n7796;
  assign n7800 = ~n7798 & ~n7799;
  assign n7801 = n7164 & n7234;
  assign n7802 = ~n7071 & n7161;
  assign n7803 = n7071 & ~n7161;
  assign n7804 = ~n7802 & ~n7803;
  assign n7805 = n7626 & ~n7629;
  assign n7806 = ~n7624 & ~n7805;
  assign n7807 = n7804 & n7806;
  assign n7808 = ~n7801 & ~n7807;
  assign n7809 = ~n7800 & n7808;
  assign n7810 = n7637 & n7809;
  assign n7811 = ~n7476 & ~n7616;
  assign n7812 = ~n7636 & n7811;
  assign n7813 = ~n7632 & ~n7635;
  assign n7814 = ~n7812 & ~n7813;
  assign n7815 = ~n7807 & ~n7814;
  assign n7816 = ~n7804 & ~n7806;
  assign n7817 = ~n7815 & ~n7816;
  assign n7818 = ~n7801 & ~n7817;
  assign n7819 = ~n7810 & ~n7818;
  assign n7820 = ~n7235 & n7819;
  assign n7821 = n7637 & ~n7807;
  assign n7822 = n7775 & n7789;
  assign n7823 = ~n7771 & ~n7773;
  assign n7824 = n7771 & n7773;
  assign n7825 = ~n7823 & ~n7824;
  assign n7826 = n7728 & ~n7730;
  assign n7827 = ~n7731 & ~n7826;
  assign n7828 = ~n7674 & n7694;
  assign n7829 = n7674 & ~n7694;
  assign n7830 = ~n7828 & ~n7829;
  assign n7831 = n7649 & ~n7651;
  assign n7832 = ~n7649 & n7651;
  assign n7833 = ~n7831 & ~n7832;
  assign n7834 = g75 & g97;
  assign n7835 = g77 & g95;
  assign n7836 = g82 & g90;
  assign n7837 = ~n7835 & n7836;
  assign n7838 = n7835 & ~n7836;
  assign n7839 = ~n7837 & ~n7838;
  assign n7840 = n7834 & ~n7839;
  assign n7841 = n7835 & n7836;
  assign n7842 = ~n7840 & ~n7841;
  assign n7843 = g74 & g98;
  assign n7844 = g10 & n7843;
  assign n7845 = ~g9 & n7648;
  assign n7846 = g9 & ~n7648;
  assign n7847 = ~n7845 & ~n7846;
  assign n7848 = ~n7844 & ~n7847;
  assign n7849 = n7844 & n7847;
  assign n7850 = ~n7848 & ~n7849;
  assign n7851 = ~n7842 & ~n7850;
  assign n7852 = n7844 & ~n7847;
  assign n7853 = ~n7851 & ~n7852;
  assign n7854 = n7833 & ~n7853;
  assign n7855 = ~n7833 & n7853;
  assign n7856 = ~n7854 & ~n7855;
  assign n7857 = ~n7830 & ~n7856;
  assign n7858 = ~n7833 & ~n7853;
  assign n7859 = ~n7857 & ~n7858;
  assign n7860 = ~n7742 & n7750;
  assign n7861 = n7742 & ~n7750;
  assign n7862 = ~n7860 & ~n7861;
  assign n7863 = ~n7657 & n7660;
  assign n7864 = n7657 & ~n7660;
  assign n7865 = ~n7863 & ~n7864;
  assign n7866 = ~n7862 & n7865;
  assign n7867 = n7862 & ~n7865;
  assign n7868 = ~n7866 & ~n7867;
  assign n7869 = ~n7859 & ~n7868;
  assign n7870 = ~n7862 & ~n7865;
  assign n7871 = ~n7869 & ~n7870;
  assign n7872 = ~n7739 & n7759;
  assign n7873 = n7739 & ~n7759;
  assign n7874 = ~n7872 & ~n7873;
  assign n7875 = n7871 & ~n7874;
  assign n7876 = ~n7871 & n7874;
  assign n7877 = ~n7875 & ~n7876;
  assign n7878 = n7827 & ~n7877;
  assign n7879 = ~n7871 & ~n7874;
  assign n7880 = ~n7878 & ~n7879;
  assign n7881 = ~n7825 & ~n7880;
  assign n7882 = ~n7687 & ~n7689;
  assign n7883 = ~n7690 & ~n7882;
  assign n7884 = ~n7675 & ~n7680;
  assign n7885 = n7675 & n7680;
  assign n7886 = ~n7884 & ~n7885;
  assign n7887 = g81 & g91;
  assign n7888 = g76 & g96;
  assign n7889 = g80 & g92;
  assign n7890 = ~n7888 & n7889;
  assign n7891 = n7888 & ~n7889;
  assign n7892 = ~n7890 & ~n7891;
  assign n7893 = n7887 & ~n7892;
  assign n7894 = n7888 & n7889;
  assign n7895 = ~n7893 & ~n7894;
  assign n7896 = n7886 & ~n7895;
  assign n7897 = ~n7886 & n7895;
  assign n7898 = ~n7896 & ~n7897;
  assign n7899 = n7883 & ~n7898;
  assign n7900 = ~n7886 & ~n7895;
  assign n7901 = ~n7899 & ~n7900;
  assign n7902 = ~n7706 & ~n7715;
  assign n7903 = n7706 & n7715;
  assign n7904 = ~n7902 & ~n7903;
  assign n7905 = ~n7901 & ~n7904;
  assign n7906 = n7842 & ~n7850;
  assign n7907 = ~n7842 & n7850;
  assign n7908 = ~n7906 & ~n7907;
  assign n7909 = ~n7666 & n7671;
  assign n7910 = ~n7672 & ~n7909;
  assign n7911 = g79 & g93;
  assign n7912 = g78 & g94;
  assign n7913 = n7911 & n7912;
  assign n7914 = g10 & ~n7843;
  assign n7915 = ~g10 & n7843;
  assign n7916 = ~n7914 & ~n7915;
  assign n7917 = ~n7911 & ~n7912;
  assign n7918 = ~n7913 & ~n7917;
  assign n7919 = ~n7916 & n7918;
  assign n7920 = ~n7913 & ~n7919;
  assign n7921 = ~n7910 & ~n7920;
  assign n7922 = n7910 & n7920;
  assign n7923 = ~n7921 & ~n7922;
  assign n7924 = ~n7908 & ~n7923;
  assign n7925 = n7910 & ~n7920;
  assign n7926 = ~n7924 & ~n7925;
  assign n7927 = n7901 & n7904;
  assign n7928 = ~n7905 & ~n7927;
  assign n7929 = ~n7926 & n7928;
  assign n7930 = ~n7905 & ~n7929;
  assign n7931 = ~n7665 & n7721;
  assign n7932 = n7665 & ~n7721;
  assign n7933 = ~n7931 & ~n7932;
  assign n7934 = ~n7930 & ~n7933;
  assign n7935 = ~n7859 & n7868;
  assign n7936 = n7859 & ~n7868;
  assign n7937 = ~n7935 & ~n7936;
  assign n7938 = n7930 & n7933;
  assign n7939 = ~n7934 & ~n7938;
  assign n7940 = ~n7937 & n7939;
  assign n7941 = ~n7934 & ~n7940;
  assign n7942 = n7827 & n7877;
  assign n7943 = ~n7827 & ~n7877;
  assign n7944 = ~n7942 & ~n7943;
  assign n7945 = n7941 & n7944;
  assign n7946 = ~n7830 & n7856;
  assign n7947 = n7830 & ~n7856;
  assign n7948 = ~n7946 & ~n7947;
  assign n7949 = g82 & g91;
  assign n7950 = g77 & g96;
  assign n7951 = g81 & g92;
  assign n7952 = ~n7950 & n7951;
  assign n7953 = n7950 & ~n7951;
  assign n7954 = ~n7952 & ~n7953;
  assign n7955 = n7949 & ~n7954;
  assign n7956 = n7950 & n7951;
  assign n7957 = ~n7955 & ~n7956;
  assign n7958 = g75 & g98;
  assign n7959 = g11 & n7958;
  assign n7960 = g79 & g94;
  assign n7961 = g78 & g95;
  assign n7962 = g76 & g97;
  assign n7963 = ~n7961 & n7962;
  assign n7964 = n7961 & ~n7962;
  assign n7965 = ~n7963 & ~n7964;
  assign n7966 = n7960 & ~n7965;
  assign n7967 = n7961 & n7962;
  assign n7968 = ~n7966 & ~n7967;
  assign n7969 = n7959 & n7968;
  assign n7970 = ~n7959 & ~n7968;
  assign n7971 = ~n7969 & ~n7970;
  assign n7972 = ~n7957 & ~n7971;
  assign n7973 = n7959 & ~n7968;
  assign n7974 = ~n7972 & ~n7973;
  assign n7975 = ~n7883 & n7898;
  assign n7976 = ~n7899 & ~n7975;
  assign n7977 = ~n7974 & n7976;
  assign n7978 = g80 & g93;
  assign n7979 = ~g11 & n7958;
  assign n7980 = g11 & ~n7958;
  assign n7981 = ~n7979 & ~n7980;
  assign n7982 = n7978 & ~n7981;
  assign n7983 = g76 & g98;
  assign n7984 = g12 & n7983;
  assign n7985 = ~n7978 & ~n7981;
  assign n7986 = n7978 & n7981;
  assign n7987 = ~n7985 & ~n7986;
  assign n7988 = n7984 & ~n7987;
  assign n7989 = ~n7982 & ~n7988;
  assign n7990 = ~n7834 & ~n7839;
  assign n7991 = n7834 & n7839;
  assign n7992 = ~n7990 & ~n7991;
  assign n7993 = ~n7887 & n7892;
  assign n7994 = ~n7893 & ~n7993;
  assign n7995 = n7992 & n7994;
  assign n7996 = ~n7992 & ~n7994;
  assign n7997 = ~n7995 & ~n7996;
  assign n7998 = ~n7989 & ~n7997;
  assign n7999 = ~n7992 & n7994;
  assign n8000 = ~n7998 & ~n7999;
  assign n8001 = n7974 & ~n7976;
  assign n8002 = ~n7977 & ~n8001;
  assign n8003 = ~n8000 & n8002;
  assign n8004 = ~n7977 & ~n8003;
  assign n8005 = ~n7948 & ~n8004;
  assign n8006 = n7926 & ~n7928;
  assign n8007 = ~n7929 & ~n8006;
  assign n8008 = n7948 & n8004;
  assign n8009 = ~n8005 & ~n8008;
  assign n8010 = n8007 & n8009;
  assign n8011 = ~n8005 & ~n8010;
  assign n8012 = n7937 & n7939;
  assign n8013 = ~n7937 & ~n7939;
  assign n8014 = ~n8012 & ~n8013;
  assign n8015 = n8011 & n8014;
  assign n8016 = n8000 & n8002;
  assign n8017 = ~n8000 & ~n8002;
  assign n8018 = ~n8016 & ~n8017;
  assign n8019 = ~n7908 & n7923;
  assign n8020 = n7908 & ~n7923;
  assign n8021 = ~n8019 & ~n8020;
  assign n8022 = ~n7960 & ~n7965;
  assign n8023 = n7960 & n7965;
  assign n8024 = ~n8022 & ~n8023;
  assign n8025 = g81 & g93;
  assign n8026 = g80 & g94;
  assign n8027 = g77 & g97;
  assign n8028 = ~n8026 & n8027;
  assign n8029 = n8026 & ~n8027;
  assign n8030 = ~n8028 & ~n8029;
  assign n8031 = n8025 & ~n8030;
  assign n8032 = n8026 & n8027;
  assign n8033 = ~n8031 & ~n8032;
  assign n8034 = g79 & g95;
  assign n8035 = g78 & g96;
  assign n8036 = g82 & g92;
  assign n8037 = ~n8035 & n8036;
  assign n8038 = n8035 & ~n8036;
  assign n8039 = ~n8037 & ~n8038;
  assign n8040 = n8034 & ~n8039;
  assign n8041 = n8035 & n8036;
  assign n8042 = ~n8040 & ~n8041;
  assign n8043 = n8033 & ~n8042;
  assign n8044 = ~n8033 & n8042;
  assign n8045 = ~n8043 & ~n8044;
  assign n8046 = ~n8024 & ~n8045;
  assign n8047 = ~n8033 & ~n8042;
  assign n8048 = ~n8046 & ~n8047;
  assign n8049 = n7916 & n7918;
  assign n8050 = ~n7916 & ~n7918;
  assign n8051 = ~n8049 & ~n8050;
  assign n8052 = n7957 & ~n7971;
  assign n8053 = ~n7957 & n7971;
  assign n8054 = ~n8052 & ~n8053;
  assign n8055 = n8051 & ~n8054;
  assign n8056 = ~n8051 & n8054;
  assign n8057 = ~n8055 & ~n8056;
  assign n8058 = ~n8048 & ~n8057;
  assign n8059 = ~n8051 & ~n8054;
  assign n8060 = ~n8058 & ~n8059;
  assign n8061 = ~n8021 & n8060;
  assign n8062 = n8021 & ~n8060;
  assign n8063 = ~n8061 & ~n8062;
  assign n8064 = ~n8018 & ~n8063;
  assign n8065 = ~n8021 & ~n8060;
  assign n8066 = ~n8064 & ~n8065;
  assign n8067 = ~n8007 & n8009;
  assign n8068 = n8007 & ~n8009;
  assign n8069 = ~n8067 & ~n8068;
  assign n8070 = n8066 & n8069;
  assign n8071 = n8048 & ~n8057;
  assign n8072 = ~n8048 & n8057;
  assign n8073 = ~n8071 & ~n8072;
  assign n8074 = g78 & g97;
  assign n8075 = g79 & g96;
  assign n8076 = g80 & g95;
  assign n8077 = ~n8075 & n8076;
  assign n8078 = n8075 & ~n8076;
  assign n8079 = ~n8077 & ~n8078;
  assign n8080 = n8074 & ~n8079;
  assign n8081 = n8075 & n8076;
  assign n8082 = ~n8080 & ~n8081;
  assign n8083 = g77 & g98;
  assign n8084 = g13 & n8083;
  assign n8085 = ~g12 & n7983;
  assign n8086 = g12 & ~n7983;
  assign n8087 = ~n8085 & ~n8086;
  assign n8088 = ~n8084 & ~n8087;
  assign n8089 = n8084 & n8087;
  assign n8090 = ~n8088 & ~n8089;
  assign n8091 = ~n8082 & ~n8090;
  assign n8092 = n8084 & ~n8087;
  assign n8093 = ~n8091 & ~n8092;
  assign n8094 = n7949 & n7954;
  assign n8095 = ~n7949 & ~n7954;
  assign n8096 = ~n8094 & ~n8095;
  assign n8097 = ~n8093 & ~n8096;
  assign n8098 = n7984 & n7987;
  assign n8099 = ~n7984 & ~n7987;
  assign n8100 = ~n8098 & ~n8099;
  assign n8101 = n8093 & n8096;
  assign n8102 = ~n8097 & ~n8101;
  assign n8103 = ~n8100 & n8102;
  assign n8104 = ~n8097 & ~n8103;
  assign n8105 = n7989 & n7997;
  assign n8106 = ~n7998 & ~n8105;
  assign n8107 = n8104 & n8106;
  assign n8108 = ~n8104 & ~n8106;
  assign n8109 = ~n8107 & ~n8108;
  assign n8110 = ~n8073 & ~n8109;
  assign n8111 = ~n8104 & n8106;
  assign n8112 = ~n8110 & ~n8111;
  assign n8113 = ~n8018 & n8063;
  assign n8114 = n8018 & ~n8063;
  assign n8115 = ~n8113 & ~n8114;
  assign n8116 = n8112 & n8115;
  assign n8117 = n8073 & ~n8109;
  assign n8118 = ~n8073 & n8109;
  assign n8119 = ~n8117 & ~n8118;
  assign n8120 = n8100 & n8102;
  assign n8121 = ~n8100 & ~n8102;
  assign n8122 = ~n8120 & ~n8121;
  assign n8123 = g82 & g93;
  assign n8124 = g81 & g94;
  assign n8125 = n8123 & n8124;
  assign n8126 = g78 & g98;
  assign n8127 = g14 & n8126;
  assign n8128 = ~n8123 & ~n8124;
  assign n8129 = ~n8125 & ~n8128;
  assign n8130 = n8127 & n8129;
  assign n8131 = ~n8125 & ~n8130;
  assign n8132 = ~n8034 & n8039;
  assign n8133 = ~n8040 & ~n8132;
  assign n8134 = ~n8025 & n8030;
  assign n8135 = ~n8031 & ~n8134;
  assign n8136 = n8133 & ~n8135;
  assign n8137 = ~n8133 & n8135;
  assign n8138 = ~n8136 & ~n8137;
  assign n8139 = ~n8131 & ~n8138;
  assign n8140 = n8133 & n8135;
  assign n8141 = ~n8139 & ~n8140;
  assign n8142 = ~n8024 & n8045;
  assign n8143 = n8024 & ~n8045;
  assign n8144 = ~n8142 & ~n8143;
  assign n8145 = n8141 & ~n8144;
  assign n8146 = ~n8141 & n8144;
  assign n8147 = ~n8145 & ~n8146;
  assign n8148 = ~n8122 & ~n8147;
  assign n8149 = ~n8141 & ~n8144;
  assign n8150 = ~n8148 & ~n8149;
  assign n8151 = n8119 & n8150;
  assign n8152 = ~n8074 & ~n8079;
  assign n8153 = n8074 & n8079;
  assign n8154 = ~n8152 & ~n8153;
  assign n8155 = ~g13 & ~n8083;
  assign n8156 = ~n8084 & ~n8155;
  assign n8157 = g79 & g97;
  assign n8158 = g80 & g96;
  assign n8159 = g81 & g95;
  assign n8160 = ~n8158 & n8159;
  assign n8161 = n8158 & ~n8159;
  assign n8162 = ~n8160 & ~n8161;
  assign n8163 = n8157 & ~n8162;
  assign n8164 = n8158 & n8159;
  assign n8165 = ~n8163 & ~n8164;
  assign n8166 = ~n8156 & ~n8165;
  assign n8167 = n8156 & n8165;
  assign n8168 = ~n8166 & ~n8167;
  assign n8169 = ~n8154 & ~n8168;
  assign n8170 = n8156 & ~n8165;
  assign n8171 = ~n8169 & ~n8170;
  assign n8172 = n8082 & ~n8090;
  assign n8173 = ~n8082 & n8090;
  assign n8174 = ~n8172 & ~n8173;
  assign n8175 = ~n8171 & ~n8174;
  assign n8176 = ~n8131 & n8138;
  assign n8177 = n8131 & ~n8138;
  assign n8178 = ~n8176 & ~n8177;
  assign n8179 = n8171 & n8174;
  assign n8180 = ~n8175 & ~n8179;
  assign n8181 = ~n8178 & n8180;
  assign n8182 = ~n8175 & ~n8181;
  assign n8183 = n8122 & n8147;
  assign n8184 = ~n8148 & ~n8183;
  assign n8185 = n8182 & ~n8184;
  assign n8186 = n8127 & ~n8129;
  assign n8187 = ~n8127 & n8129;
  assign n8188 = ~n8186 & ~n8187;
  assign n8189 = g82 & g94;
  assign n8190 = ~g14 & n8126;
  assign n8191 = g14 & ~n8126;
  assign n8192 = ~n8190 & ~n8191;
  assign n8193 = n8189 & ~n8192;
  assign n8194 = g80 & g97;
  assign n8195 = g81 & g96;
  assign n8196 = g82 & g95;
  assign n8197 = ~n8195 & n8196;
  assign n8198 = n8195 & ~n8196;
  assign n8199 = ~n8197 & ~n8198;
  assign n8200 = n8194 & ~n8199;
  assign n8201 = n8195 & n8196;
  assign n8202 = ~n8200 & ~n8201;
  assign n8203 = ~n8189 & n8192;
  assign n8204 = ~n8193 & ~n8203;
  assign n8205 = ~n8202 & n8204;
  assign n8206 = ~n8193 & ~n8205;
  assign n8207 = n8188 & ~n8206;
  assign n8208 = ~n8188 & n8206;
  assign n8209 = ~n8207 & ~n8208;
  assign n8210 = ~n8154 & n8168;
  assign n8211 = n8154 & ~n8168;
  assign n8212 = ~n8210 & ~n8211;
  assign n8213 = ~n8209 & ~n8212;
  assign n8214 = ~n8188 & ~n8206;
  assign n8215 = ~n8213 & ~n8214;
  assign n8216 = n8178 & n8180;
  assign n8217 = ~n8178 & ~n8180;
  assign n8218 = ~n8216 & ~n8217;
  assign n8219 = ~n8215 & ~n8218;
  assign n8220 = n8215 & n8218;
  assign n8221 = g79 & g98;
  assign n8222 = ~g15 & ~n8221;
  assign n8223 = n8157 & n8162;
  assign n8224 = ~n8157 & ~n8162;
  assign n8225 = ~n8223 & ~n8224;
  assign n8226 = n8222 & ~n8225;
  assign n8227 = ~n8222 & n8225;
  assign n8228 = ~n8226 & ~n8227;
  assign n8229 = ~n8202 & ~n8204;
  assign n8230 = n8202 & n8204;
  assign n8231 = ~n8229 & ~n8230;
  assign n8232 = ~n8228 & ~n8231;
  assign n8233 = ~n8222 & ~n8225;
  assign n8234 = ~n8232 & ~n8233;
  assign n8235 = n8209 & ~n8212;
  assign n8236 = ~n8209 & n8212;
  assign n8237 = ~n8235 & ~n8236;
  assign n8238 = ~n8234 & ~n8237;
  assign n8239 = n8234 & n8237;
  assign n8240 = g15 & ~n8221;
  assign n8241 = ~g15 & n8221;
  assign n8242 = ~n8240 & ~n8241;
  assign n8243 = g80 & g98;
  assign n8244 = g16 & n8243;
  assign n8245 = ~n8242 & n8244;
  assign n8246 = n8242 & ~n8244;
  assign n8247 = ~n8245 & ~n8246;
  assign n8248 = ~n8194 & n8199;
  assign n8249 = ~n8200 & ~n8248;
  assign n8250 = ~n8247 & n8249;
  assign n8251 = n8242 & n8244;
  assign n8252 = ~n8250 & ~n8251;
  assign n8253 = ~n8228 & n8231;
  assign n8254 = n8228 & ~n8231;
  assign n8255 = ~n8253 & ~n8254;
  assign n8256 = ~n8252 & ~n8255;
  assign n8257 = n8252 & n8255;
  assign n8258 = n8247 & n8249;
  assign n8259 = ~n8247 & ~n8249;
  assign n8260 = ~n8258 & ~n8259;
  assign n8261 = g82 & g96;
  assign n8262 = g81 & g97;
  assign n8263 = n8261 & n8262;
  assign n8264 = ~g16 & ~n8243;
  assign n8265 = ~n8244 & ~n8264;
  assign n8266 = ~n8261 & ~n8262;
  assign n8267 = ~n8263 & ~n8266;
  assign n8268 = n8265 & n8267;
  assign n8269 = ~n8263 & ~n8268;
  assign n8270 = n8260 & n8269;
  assign n8271 = g82 & g98;
  assign n8272 = g18 & n8271;
  assign n8273 = g81 & g98;
  assign n8274 = n8272 & n8273;
  assign n8275 = g82 & g97;
  assign n8276 = ~g17 & n8275;
  assign n8277 = g17 & ~n8275;
  assign n8278 = ~n8276 & ~n8277;
  assign n8279 = ~n8272 & ~n8273;
  assign n8280 = ~n8274 & ~n8279;
  assign n8281 = ~n8278 & n8280;
  assign n8282 = ~n8274 & ~n8281;
  assign n8283 = g17 & n8275;
  assign n8284 = ~n8282 & n8283;
  assign n8285 = n8265 & ~n8267;
  assign n8286 = ~n8265 & n8267;
  assign n8287 = ~n8285 & ~n8286;
  assign n8288 = n8282 & ~n8283;
  assign n8289 = ~n8284 & ~n8288;
  assign n8290 = ~n8287 & n8289;
  assign n8291 = ~n8284 & ~n8290;
  assign n8292 = ~n8270 & ~n8291;
  assign n8293 = ~n8260 & ~n8269;
  assign n8294 = ~n8292 & ~n8293;
  assign n8295 = ~n8257 & ~n8294;
  assign n8296 = ~n8256 & ~n8295;
  assign n8297 = ~n8239 & ~n8296;
  assign n8298 = ~n8238 & ~n8297;
  assign n8299 = ~n8220 & ~n8298;
  assign n8300 = ~n8219 & ~n8299;
  assign n8301 = ~n8185 & ~n8300;
  assign n8302 = ~n8182 & n8184;
  assign n8303 = ~n8301 & ~n8302;
  assign n8304 = ~n8151 & ~n8303;
  assign n8305 = ~n8119 & ~n8150;
  assign n8306 = ~n8304 & ~n8305;
  assign n8307 = ~n8116 & ~n8306;
  assign n8308 = ~n8112 & ~n8115;
  assign n8309 = ~n8307 & ~n8308;
  assign n8310 = ~n8070 & ~n8309;
  assign n8311 = ~n8066 & ~n8069;
  assign n8312 = ~n8310 & ~n8311;
  assign n8313 = ~n8015 & ~n8312;
  assign n8314 = ~n8011 & ~n8014;
  assign n8315 = ~n8313 & ~n8314;
  assign n8316 = ~n7945 & ~n8315;
  assign n8317 = ~n7941 & ~n7944;
  assign n8318 = ~n8316 & ~n8317;
  assign n8319 = n7825 & n7880;
  assign n8320 = ~n7881 & ~n8319;
  assign n8321 = ~n8318 & n8320;
  assign n8322 = ~n7881 & ~n8321;
  assign n8323 = ~n7822 & ~n8322;
  assign n8324 = ~n7797 & n8323;
  assign n8325 = n7821 & n8324;
  assign n8326 = ~n7801 & n8325;
  assign n8327 = n7820 & ~n8326;
  assign n8328 = ~n6738 & n6747;
  assign n8329 = n6738 & ~n6747;
  assign n8330 = ~n8328 & ~n8329;
  assign n8331 = n6584 & ~n6591;
  assign n8332 = ~n6584 & n6591;
  assign n8333 = ~n8331 & ~n8332;
  assign n8334 = ~n7183 & n7191;
  assign n8335 = ~n7189 & ~n8334;
  assign n8336 = ~n8333 & n8335;
  assign n8337 = n8333 & ~n8335;
  assign n8338 = ~n8336 & ~n8337;
  assign n8339 = ~n7168 & ~n7177;
  assign n8340 = ~n7171 & ~n7174;
  assign n8341 = ~n8339 & ~n8340;
  assign n8342 = n8338 & ~n8341;
  assign n8343 = ~n8338 & n8341;
  assign n8344 = ~n8342 & ~n8343;
  assign n8345 = ~n7210 & ~n7213;
  assign n8346 = ~n7217 & ~n8345;
  assign n8347 = n6691 & n6729;
  assign n8348 = ~n6730 & ~n8347;
  assign n8349 = n8346 & n8348;
  assign n8350 = ~n8346 & ~n8348;
  assign n8351 = ~n8349 & ~n8350;
  assign n8352 = ~n8344 & ~n8351;
  assign n8353 = ~n8346 & n8348;
  assign n8354 = ~n8352 & ~n8353;
  assign n8355 = ~n6685 & n6735;
  assign n8356 = n6685 & ~n6735;
  assign n8357 = ~n8355 & ~n8356;
  assign n8358 = ~n8338 & ~n8341;
  assign n8359 = ~n8333 & ~n8335;
  assign n8360 = ~n8358 & ~n8359;
  assign n8361 = n8357 & ~n8360;
  assign n8362 = ~n8357 & n8360;
  assign n8363 = ~n8361 & ~n8362;
  assign n8364 = ~n8354 & ~n8363;
  assign n8365 = ~n8357 & ~n8360;
  assign n8366 = ~n8364 & ~n8365;
  assign n8367 = n8330 & n8366;
  assign n8368 = ~n7166 & ~n7231;
  assign n8369 = ~n7202 & ~n7228;
  assign n8370 = ~n8368 & ~n8369;
  assign n8371 = ~n8344 & n8351;
  assign n8372 = n8344 & ~n8351;
  assign n8373 = ~n8371 & ~n8372;
  assign n8374 = ~n7197 & ~n7199;
  assign n8375 = ~n7180 & ~n7194;
  assign n8376 = ~n8374 & ~n8375;
  assign n8377 = ~n8373 & n8376;
  assign n8378 = n8373 & ~n8376;
  assign n8379 = ~n8377 & ~n8378;
  assign n8380 = ~n7204 & n7225;
  assign n8381 = ~n7223 & ~n8380;
  assign n8382 = ~n8379 & n8381;
  assign n8383 = n8379 & ~n8381;
  assign n8384 = ~n8382 & ~n8383;
  assign n8385 = n8370 & n8384;
  assign n8386 = n8354 & ~n8363;
  assign n8387 = ~n8354 & n8363;
  assign n8388 = ~n8386 & ~n8387;
  assign n8389 = ~n8379 & ~n8381;
  assign n8390 = ~n8373 & ~n8376;
  assign n8391 = ~n8389 & ~n8390;
  assign n8392 = n8388 & n8391;
  assign n8393 = ~n8385 & ~n8392;
  assign n8394 = ~n8367 & n8393;
  assign n8395 = ~n8327 & n8394;
  assign n8396 = ~n6751 & n8395;
  assign n8397 = ~n8370 & ~n8384;
  assign n8398 = ~n8392 & n8397;
  assign n8399 = ~n8388 & ~n8391;
  assign n8400 = ~n8398 & ~n8399;
  assign n8401 = ~n8367 & ~n8400;
  assign n8402 = ~n8330 & ~n8366;
  assign n8403 = ~n8401 & ~n8402;
  assign n8404 = ~n6751 & ~n8403;
  assign n8405 = ~n6682 & ~n6750;
  assign n8406 = ~n8404 & ~n8405;
  assign n8407 = ~n8396 & n8406;
  assign n8408 = ~n6679 & ~n8407;
  assign n8409 = ~n6576 & ~n6678;
  assign n8410 = ~n8408 & ~n8409;
  assign n8411 = n6573 & ~n8410;
  assign n8412 = n6527 & n8411;
  assign n8413 = n6562 & ~n6565;
  assign n8414 = ~n6560 & n8413;
  assign n8415 = ~n6544 & ~n6559;
  assign n8416 = ~n8414 & ~n8415;
  assign n8417 = ~n6436 & ~n6524;
  assign n8418 = ~n6433 & n8417;
  assign n8419 = ~n6313 & ~n6432;
  assign n8420 = ~n8418 & ~n8419;
  assign n8421 = ~n6310 & ~n8420;
  assign n8422 = ~n6236 & ~n6309;
  assign n8423 = ~n8421 & ~n8422;
  assign n8424 = n6567 & ~n8423;
  assign n8425 = n8416 & ~n8424;
  assign n8426 = ~n6572 & ~n8425;
  assign n8427 = n6568 & ~n6571;
  assign n8428 = ~n8426 & ~n8427;
  assign n8429 = ~n8412 & n8428;
  assign n8430 = ~g0 & ~n8429;
  assign n8431 = ~n6042 & ~n8430;
  assign n8432 = n6436 & ~n6524;
  assign n8433 = ~n6436 & n6524;
  assign n8434 = ~n8432 & ~n8433;
  assign n8435 = ~n6236 & n6309;
  assign n8436 = n6236 & ~n6309;
  assign n8437 = ~n8435 & ~n8436;
  assign n8438 = ~n6313 & n6432;
  assign n8439 = n6313 & ~n6432;
  assign n8440 = ~n8438 & ~n8439;
  assign n8441 = ~n8437 & ~n8440;
  assign n8442 = ~n8434 & n8441;
  assign n8443 = ~n8410 & n8442;
  assign n8444 = n8423 & ~n8443;
  assign n8445 = ~n6566 & ~n8444;
  assign n8446 = ~n8413 & ~n8445;
  assign n8447 = n6544 & ~n6559;
  assign n8448 = ~n6544 & n6559;
  assign n8449 = ~n8447 & ~n8448;
  assign n8450 = ~n8446 & ~n8449;
  assign n8451 = ~n8415 & ~n8450;
  assign n8452 = ~n8427 & n8451;
  assign n8453 = ~g0 & ~n6572;
  assign n8454 = ~n8452 & n8453;
  assign n8455 = ~n6164 & ~n8454;
  assign n8456 = n8431 & ~n8455;
  assign n8457 = ~n8431 & n8455;
  assign n8458 = ~n8456 & ~n8457;
  assign n8459 = n6167 & n8458;
  assign n8460 = n6167 & n8459;
  assign n8461 = n6167 & n8460;
  assign n8462 = n6167 & n8461;
  assign n8463 = ~n6572 & ~n8427;
  assign n8464 = ~n8451 & n8463;
  assign n8465 = n8451 & ~n8463;
  assign n8466 = ~n8464 & ~n8465;
  assign n8467 = ~g0 & n8466;
  assign n8468 = ~n6042 & ~n8467;
  assign n8469 = ~n6164 & ~n8467;
  assign n8470 = n8468 & ~n8469;
  assign n8471 = ~n8468 & n8469;
  assign n8472 = ~n8470 & ~n8471;
  assign n8473 = n8446 & n8449;
  assign n8474 = ~g0 & ~n8450;
  assign n8475 = ~n8473 & n8474;
  assign n8476 = n5475 & n5704;
  assign n8477 = ~n5701 & ~n6036;
  assign n8478 = n6035 & n8477;
  assign n8479 = n8476 & n8478;
  assign n8480 = n5702 & ~n6039;
  assign n8481 = n5516 & n8480;
  assign n8482 = n5663 & n8481;
  assign n8483 = ~n8479 & ~n8482;
  assign n8484 = g0 & ~n8483;
  assign n8485 = ~n8475 & ~n8484;
  assign n8486 = g0 & n6152;
  assign n8487 = n6154 & n8486;
  assign n8488 = ~n8475 & ~n8487;
  assign n8489 = ~n6164 & n8488;
  assign n8490 = n8485 & ~n8489;
  assign n8491 = ~n8485 & n8489;
  assign n8492 = ~n8490 & ~n8491;
  assign n8493 = n8472 & n8492;
  assign n8494 = n5663 & ~n6035;
  assign n8495 = n8476 & ~n8494;
  assign n8496 = n5516 & ~n8495;
  assign n8497 = ~n5452 & n5701;
  assign n8498 = ~n6036 & ~n8497;
  assign n8499 = n8496 & ~n8498;
  assign n8500 = g0 & ~n8499;
  assign n8501 = ~n8496 & n8498;
  assign n8502 = n8500 & ~n8501;
  assign n8503 = ~n6566 & ~n8413;
  assign n8504 = n8444 & ~n8503;
  assign n8505 = ~n8444 & n8503;
  assign n8506 = ~n8504 & ~n8505;
  assign n8507 = ~g0 & n8506;
  assign n8508 = ~n8502 & ~n8507;
  assign n8509 = ~n6078 & ~n6099;
  assign n8510 = n6078 & n6099;
  assign n8511 = ~n8509 & ~n8510;
  assign n8512 = n6092 & ~n6099;
  assign n8513 = ~n6092 & n6099;
  assign n8514 = ~n8512 & ~n8513;
  assign n8515 = ~n6124 & n6131;
  assign n8516 = n6124 & ~n6131;
  assign n8517 = ~n8515 & ~n8516;
  assign n8518 = ~n8515 & ~n8517;
  assign n8519 = ~n5732 & ~n5802;
  assign n8520 = ~n5748 & ~n5776;
  assign n8521 = n5736 & ~n8520;
  assign n8522 = n8519 & ~n8521;
  assign n8523 = ~n5870 & n5882;
  assign n8524 = n5870 & ~n5882;
  assign n8525 = ~n8523 & ~n8524;
  assign n8526 = ~n6022 & ~n8525;
  assign n8527 = ~n5883 & ~n8526;
  assign n8528 = ~n5889 & n8527;
  assign n8529 = n5839 & ~n5893;
  assign n8530 = ~n5839 & n5893;
  assign n8531 = ~n8529 & ~n8530;
  assign n8532 = ~n5886 & ~n8531;
  assign n8533 = ~n8528 & n8532;
  assign n8534 = ~n5827 & ~n5894;
  assign n8535 = ~n8533 & n8534;
  assign n8536 = n5782 & ~n5796;
  assign n8537 = ~n5782 & n5796;
  assign n8538 = ~n8536 & ~n8537;
  assign n8539 = ~n5844 & ~n8538;
  assign n8540 = ~n8535 & n8539;
  assign n8541 = ~n5797 & ~n8540;
  assign n8542 = ~n5749 & ~n5778;
  assign n8543 = n8541 & n8542;
  assign n8544 = n8522 & ~n8543;
  assign n8545 = n5625 & n5655;
  assign n8546 = n5636 & ~n8545;
  assign n8547 = ~n5732 & ~n8546;
  assign n8548 = ~n8544 & n8547;
  assign n8549 = ~n5625 & ~n5655;
  assign n8550 = ~n5636 & ~n8549;
  assign n8551 = ~n8548 & ~n8550;
  assign n8552 = n5609 & n5636;
  assign n8553 = ~n6138 & ~n8552;
  assign n8554 = n8551 & ~n8553;
  assign n8555 = n5567 & ~n5609;
  assign n8556 = n5609 & ~n5636;
  assign n8557 = ~n8555 & ~n8556;
  assign n8558 = ~n8554 & n8557;
  assign n8559 = ~n5567 & n6131;
  assign n8560 = ~n6158 & ~n8559;
  assign n8561 = ~n5709 & ~n8560;
  assign n8562 = ~n8558 & n8561;
  assign n8563 = ~n5567 & ~n6131;
  assign n8564 = ~n8515 & ~n8563;
  assign n8565 = ~n8562 & n8564;
  assign n8566 = ~n8518 & ~n8565;
  assign n8567 = ~n6092 & n6106;
  assign n8568 = ~n6106 & n6119;
  assign n8569 = ~n6119 & n6124;
  assign n8570 = ~n8568 & ~n8569;
  assign n8571 = ~n8567 & n8570;
  assign n8572 = ~n8566 & n8571;
  assign n8573 = n6119 & ~n6124;
  assign n8574 = ~n8569 & ~n8573;
  assign n8575 = n8570 & ~n8574;
  assign n8576 = n6106 & ~n6119;
  assign n8577 = ~n8575 & ~n8576;
  assign n8578 = n6092 & ~n8577;
  assign n8579 = n6092 & ~n6106;
  assign n8580 = ~n8578 & ~n8579;
  assign n8581 = ~n8572 & n8580;
  assign n8582 = n8514 & n8581;
  assign n8583 = ~n8512 & ~n8582;
  assign n8584 = ~n8511 & ~n8583;
  assign n8585 = ~n6078 & n6099;
  assign n8586 = ~n8584 & ~n8585;
  assign n8587 = n6078 & ~n6085;
  assign n8588 = n8586 & ~n8587;
  assign n8589 = ~n6086 & ~n8588;
  assign n8590 = n6085 & ~n6152;
  assign n8591 = ~n6153 & ~n8590;
  assign n8592 = ~n8589 & n8591;
  assign n8593 = g0 & n8592;
  assign n8594 = n8589 & ~n8591;
  assign n8595 = g0 & n8594;
  assign n8596 = ~n8507 & ~n8595;
  assign n8597 = ~n8593 & n8596;
  assign n8598 = n8508 & ~n8597;
  assign n8599 = ~n8508 & n8597;
  assign n8600 = ~n8598 & ~n8599;
  assign n8601 = n6526 & n8409;
  assign n8602 = n8420 & ~n8601;
  assign n8603 = n6526 & ~n6679;
  assign n8604 = ~n8407 & n8603;
  assign n8605 = n8602 & ~n8604;
  assign n8606 = ~n8437 & ~n8605;
  assign n8607 = n8437 & n8605;
  assign n8608 = ~g0 & ~n8607;
  assign n8609 = ~n8606 & n8608;
  assign n8610 = ~n5453 & ~n5473;
  assign n8611 = ~n5474 & ~n5513;
  assign n8612 = ~n5471 & ~n8611;
  assign n8613 = ~n5474 & ~n8494;
  assign n8614 = n5704 & n8613;
  assign n8615 = n8612 & ~n8614;
  assign n8616 = g0 & ~n8615;
  assign n8617 = ~n8610 & n8616;
  assign n8618 = g0 & n8610;
  assign n8619 = n8612 & n8618;
  assign n8620 = ~n8614 & n8619;
  assign n8621 = ~n8617 & ~n8620;
  assign n8622 = ~n8609 & n8621;
  assign n8623 = n6078 & n6085;
  assign n8624 = ~n6078 & ~n6085;
  assign n8625 = ~n8623 & ~n8624;
  assign n8626 = ~n8586 & ~n8625;
  assign n8627 = n8586 & n8625;
  assign n8628 = ~n8626 & ~n8627;
  assign n8629 = g0 & n8628;
  assign n8630 = ~n8609 & ~n8629;
  assign n8631 = n8622 & ~n8630;
  assign n8632 = ~n8622 & n8630;
  assign n8633 = ~n8631 & ~n8632;
  assign n8634 = ~n5663 & n5704;
  assign n8635 = n5513 & ~n8634;
  assign n8636 = n5704 & n6035;
  assign n8637 = n8635 & ~n8636;
  assign n8638 = ~n5471 & ~n5474;
  assign n8639 = g0 & ~n8638;
  assign n8640 = ~n8637 & n8639;
  assign n8641 = ~n8410 & ~n8434;
  assign n8642 = ~n8417 & ~n8641;
  assign n8643 = n8440 & n8642;
  assign n8644 = ~n8440 & ~n8642;
  assign n8645 = ~g0 & ~n8644;
  assign n8646 = ~n8643 & n8645;
  assign n8647 = g0 & n8635;
  assign n8648 = n8638 & n8647;
  assign n8649 = ~n8636 & n8648;
  assign n8650 = ~n8646 & ~n8649;
  assign n8651 = ~n8640 & n8650;
  assign n8652 = ~n8511 & n8583;
  assign n8653 = n8511 & ~n8583;
  assign n8654 = ~n8652 & ~n8653;
  assign n8655 = g0 & ~n8654;
  assign n8656 = ~n8646 & ~n8655;
  assign n8657 = n8651 & ~n8656;
  assign n8658 = ~n8651 & n8656;
  assign n8659 = ~n8657 & ~n8658;
  assign n8660 = n8633 & n8659;
  assign n8661 = n8600 & n8660;
  assign n8662 = n8493 & n8661;
  assign n8663 = ~n8410 & n8434;
  assign n8664 = n8410 & ~n8434;
  assign n8665 = ~n8663 & ~n8664;
  assign n8666 = ~g0 & ~n8665;
  assign n8667 = ~n5703 & n6035;
  assign n8668 = ~n5510 & ~n8667;
  assign n8669 = ~n5491 & ~n5512;
  assign n8670 = ~n8668 & n8669;
  assign n8671 = g0 & ~n8670;
  assign n8672 = ~n5663 & ~n5703;
  assign n8673 = ~n8669 & ~n8672;
  assign n8674 = n8668 & n8673;
  assign n8675 = n8671 & ~n8674;
  assign n8676 = ~n8634 & n8675;
  assign n8677 = ~n8666 & ~n8676;
  assign n8678 = n8514 & ~n8581;
  assign n8679 = ~n8514 & n8581;
  assign n8680 = ~n8678 & ~n8679;
  assign n8681 = g0 & ~n8680;
  assign n8682 = ~n8666 & ~n8681;
  assign n8683 = n8677 & ~n8682;
  assign n8684 = ~n8677 & n8682;
  assign n8685 = ~n8683 & ~n8684;
  assign n8686 = ~n5510 & ~n5703;
  assign n8687 = g0 & ~n8686;
  assign n8688 = ~n8494 & n8687;
  assign n8689 = g0 & n8686;
  assign n8690 = n8494 & n8689;
  assign n8691 = ~n6576 & n6678;
  assign n8692 = n6576 & ~n6678;
  assign n8693 = ~n8691 & ~n8692;
  assign n8694 = ~n8407 & ~n8693;
  assign n8695 = n8407 & n8693;
  assign n8696 = ~g0 & ~n8695;
  assign n8697 = ~n8694 & n8696;
  assign n8698 = ~n8690 & ~n8697;
  assign n8699 = ~n8688 & n8698;
  assign n8700 = ~n8566 & n8570;
  assign n8701 = n8577 & ~n8700;
  assign n8702 = ~n6092 & ~n6106;
  assign n8703 = ~n6107 & ~n8702;
  assign n8704 = ~n8701 & n8703;
  assign n8705 = n8701 & ~n8703;
  assign n8706 = ~n8704 & ~n8705;
  assign n8707 = g0 & n8706;
  assign n8708 = ~n8697 & ~n8707;
  assign n8709 = n8699 & ~n8708;
  assign n8710 = ~n8699 & n8708;
  assign n8711 = ~n8709 & ~n8710;
  assign n8712 = n5711 & ~n6032;
  assign n8713 = n5594 & n8712;
  assign n8714 = ~n5547 & n8713;
  assign n8715 = n5594 & n5659;
  assign n8716 = ~n5547 & n8715;
  assign n8717 = ~n5547 & n5585;
  assign n8718 = ~n8716 & ~n8717;
  assign n8719 = ~n8714 & n8718;
  assign n8720 = ~n5589 & n8719;
  assign n8721 = ~n5535 & ~n5548;
  assign n8722 = ~n8720 & n8721;
  assign n8723 = n8718 & ~n8721;
  assign n8724 = ~n8714 & n8723;
  assign n8725 = ~n5589 & n8724;
  assign n8726 = ~n8722 & ~n8725;
  assign n8727 = g0 & n8726;
  assign n8728 = n6682 & ~n6750;
  assign n8729 = ~n6682 & n6750;
  assign n8730 = ~n8728 & ~n8729;
  assign n8731 = n8330 & ~n8366;
  assign n8732 = ~n8330 & n8366;
  assign n8733 = ~n8731 & ~n8732;
  assign n8734 = ~n8388 & n8391;
  assign n8735 = n8388 & ~n8391;
  assign n8736 = ~n8734 & ~n8735;
  assign n8737 = ~n8370 & n8384;
  assign n8738 = n8370 & ~n8384;
  assign n8739 = ~n8737 & ~n8738;
  assign n8740 = ~n8327 & ~n8739;
  assign n8741 = ~n8397 & ~n8740;
  assign n8742 = ~n8736 & ~n8741;
  assign n8743 = ~n8399 & ~n8742;
  assign n8744 = ~n8733 & ~n8743;
  assign n8745 = ~n8402 & ~n8744;
  assign n8746 = n8730 & ~n8745;
  assign n8747 = ~n8730 & n8745;
  assign n8748 = ~n8746 & ~n8747;
  assign n8749 = ~g0 & ~n8748;
  assign n8750 = ~n8727 & ~n8749;
  assign n8751 = n8566 & n8574;
  assign n8752 = ~n8569 & ~n8751;
  assign n8753 = n6106 & n6119;
  assign n8754 = ~n6106 & ~n6119;
  assign n8755 = ~n8753 & ~n8754;
  assign n8756 = ~n8752 & ~n8755;
  assign n8757 = n8752 & n8755;
  assign n8758 = ~n8756 & ~n8757;
  assign n8759 = g0 & n8758;
  assign n8760 = ~n8749 & ~n8759;
  assign n8761 = n8750 & ~n8760;
  assign n8762 = ~n8750 & n8760;
  assign n8763 = ~n8761 & ~n8762;
  assign n8764 = n8711 & n8763;
  assign n8765 = n8685 & n8764;
  assign n8766 = ~n5547 & ~n5589;
  assign n8767 = ~n5585 & ~n8715;
  assign n8768 = ~n8713 & n8767;
  assign n8769 = g0 & n8768;
  assign n8770 = n8766 & n8769;
  assign n8771 = g0 & ~n8766;
  assign n8772 = ~n8768 & n8771;
  assign n8773 = n8733 & n8743;
  assign n8774 = ~g0 & ~n8744;
  assign n8775 = ~n8773 & n8774;
  assign n8776 = ~n8772 & ~n8775;
  assign n8777 = ~n8770 & n8776;
  assign n8778 = ~n8566 & ~n8574;
  assign n8779 = ~n8751 & ~n8778;
  assign n8780 = g0 & n8779;
  assign n8781 = ~n8775 & ~n8780;
  assign n8782 = n8777 & ~n8781;
  assign n8783 = ~n8777 & n8781;
  assign n8784 = ~n8782 & ~n8783;
  assign n8785 = ~n5546 & ~n5583;
  assign n8786 = n5546 & n5583;
  assign n8787 = ~n8785 & ~n8786;
  assign n8788 = ~n5659 & ~n8712;
  assign n8789 = ~n5593 & ~n8788;
  assign n8790 = ~n5567 & n5583;
  assign n8791 = ~n8789 & ~n8790;
  assign n8792 = ~n8787 & ~n8791;
  assign n8793 = n8787 & n8791;
  assign n8794 = g0 & ~n8793;
  assign n8795 = ~n8792 & n8794;
  assign n8796 = n8736 & ~n8741;
  assign n8797 = ~n8736 & n8741;
  assign n8798 = ~n8796 & ~n8797;
  assign n8799 = ~g0 & ~n8798;
  assign n8800 = ~n8795 & ~n8799;
  assign n8801 = ~n8562 & ~n8563;
  assign n8802 = ~n8517 & n8801;
  assign n8803 = n8517 & ~n8801;
  assign n8804 = ~n8802 & ~n8803;
  assign n8805 = g0 & n8804;
  assign n8806 = ~n8799 & ~n8805;
  assign n8807 = n8800 & ~n8806;
  assign n8808 = ~n8800 & n8806;
  assign n8809 = ~n8807 & ~n8808;
  assign n8810 = ~n5593 & ~n8790;
  assign n8811 = ~n8788 & n8810;
  assign n8812 = n8788 & ~n8810;
  assign n8813 = g0 & ~n8812;
  assign n8814 = ~n8811 & n8813;
  assign n8815 = ~n8327 & n8739;
  assign n8816 = n8327 & ~n8739;
  assign n8817 = ~n8815 & ~n8816;
  assign n8818 = ~g0 & ~n8817;
  assign n8819 = ~n8814 & ~n8818;
  assign n8820 = n8560 & ~n8788;
  assign n8821 = ~n8560 & n8788;
  assign n8822 = ~n8820 & ~n8821;
  assign n8823 = g0 & ~n8822;
  assign n8824 = ~n8818 & ~n8823;
  assign n8825 = n8819 & ~n8824;
  assign n8826 = ~n8819 & n8824;
  assign n8827 = ~n8825 & ~n8826;
  assign n8828 = n8809 & n8827;
  assign n8829 = n8784 & n8828;
  assign n8830 = n8765 & n8829;
  assign n8831 = n8662 & n8830;
  assign n8832 = n8462 & n8831;
  assign n8833 = n6167 & n8832;
  assign n8834 = ~n8651 & ~n8677;
  assign n8835 = ~n8508 & n8834;
  assign n8836 = ~n8622 & n8835;
  assign n8837 = ~n8699 & ~n8750;
  assign n8838 = ~n8777 & n8837;
  assign n8839 = ~n8800 & n8838;
  assign n8840 = ~n8551 & n8553;
  assign n8841 = ~n8554 & ~n8840;
  assign n8842 = g0 & n8841;
  assign n8843 = n7804 & ~n7806;
  assign n8844 = ~n7804 & n7806;
  assign n8845 = ~n8843 & ~n8844;
  assign n8846 = ~n7632 & n7635;
  assign n8847 = n7632 & ~n7635;
  assign n8848 = ~n8846 & ~n8847;
  assign n8849 = ~n7476 & n7616;
  assign n8850 = n7476 & ~n7616;
  assign n8851 = ~n8849 & ~n8850;
  assign n8852 = ~n7793 & n7796;
  assign n8853 = n7793 & ~n7796;
  assign n8854 = ~n8852 & ~n8853;
  assign n8855 = ~n7775 & n7789;
  assign n8856 = n7775 & ~n7789;
  assign n8857 = ~n8855 & ~n8856;
  assign n8858 = ~n8322 & ~n8857;
  assign n8859 = ~n7790 & ~n8858;
  assign n8860 = ~n8854 & ~n8859;
  assign n8861 = ~n7799 & ~n8860;
  assign n8862 = ~n8851 & ~n8861;
  assign n8863 = ~n7811 & ~n8862;
  assign n8864 = ~n8848 & ~n8863;
  assign n8865 = ~n7813 & ~n8864;
  assign n8866 = n8845 & ~n8865;
  assign n8867 = ~n8845 & n8865;
  assign n8868 = ~n8866 & ~n8867;
  assign n8869 = ~g0 & ~n8868;
  assign n8870 = ~n8842 & ~n8869;
  assign n8871 = ~n5567 & ~n5609;
  assign n8872 = n5567 & n5609;
  assign n8873 = ~n8871 & ~n8872;
  assign n8874 = ~n5708 & n8551;
  assign n8875 = ~n8556 & ~n8874;
  assign n8876 = ~n8873 & ~n8875;
  assign n8877 = n8873 & n8875;
  assign n8878 = g0 & ~n8877;
  assign n8879 = ~n8876 & n8878;
  assign n8880 = ~n7164 & n7234;
  assign n8881 = n7164 & ~n7234;
  assign n8882 = ~n8880 & ~n8881;
  assign n8883 = n7816 & ~n8882;
  assign n8884 = n7807 & n8882;
  assign n8885 = ~n8883 & ~n8884;
  assign n8886 = ~g0 & n8885;
  assign n8887 = ~n7816 & n8882;
  assign n8888 = n8865 & n8887;
  assign n8889 = ~n8865 & ~n8882;
  assign n8890 = ~n7807 & n8889;
  assign n8891 = ~n8888 & ~n8890;
  assign n8892 = n8886 & n8891;
  assign n8893 = ~n8879 & ~n8892;
  assign n8894 = ~n5705 & ~n6032;
  assign n8895 = ~n5625 & n5655;
  assign n8896 = ~n8894 & ~n8895;
  assign n8897 = ~n5636 & ~n5655;
  assign n8898 = ~n5656 & ~n8897;
  assign n8899 = g0 & n8898;
  assign n8900 = ~n8896 & n8899;
  assign n8901 = g0 & ~n8898;
  assign n8902 = ~n8894 & n8901;
  assign n8903 = ~n8895 & n8902;
  assign n8904 = n8848 & n8863;
  assign n8905 = ~g0 & ~n8904;
  assign n8906 = ~n8864 & n8905;
  assign n8907 = ~n8903 & ~n8906;
  assign n8908 = ~n8900 & n8907;
  assign n8909 = n8854 & ~n8859;
  assign n8910 = ~n8854 & n8859;
  assign n8911 = ~n8909 & ~n8910;
  assign n8912 = ~g0 & ~n8911;
  assign n8913 = n5805 & ~n6028;
  assign n8914 = ~n5777 & n8913;
  assign n8915 = ~n5749 & ~n5800;
  assign n8916 = ~n8519 & n8915;
  assign n8917 = ~n8914 & n8916;
  assign n8918 = g0 & ~n8544;
  assign n8919 = ~n8917 & n8918;
  assign n8920 = ~n8912 & ~n8919;
  assign n8921 = n8851 & ~n8861;
  assign n8922 = ~n8851 & n8861;
  assign n8923 = ~n8921 & ~n8922;
  assign n8924 = ~g0 & ~n8923;
  assign n8925 = ~n5705 & ~n8895;
  assign n8926 = n6032 & ~n8925;
  assign n8927 = ~n6032 & n8925;
  assign n8928 = ~n8926 & ~n8927;
  assign n8929 = g0 & n8928;
  assign n8930 = ~n8924 & ~n8929;
  assign n8931 = ~n5776 & ~n5778;
  assign n8932 = n8541 & ~n8931;
  assign n8933 = g0 & ~n8932;
  assign n8934 = ~n8541 & n8931;
  assign n8935 = n8933 & ~n8934;
  assign n8936 = ~n8318 & ~n8320;
  assign n8937 = n8318 & n8320;
  assign n8938 = ~n8936 & ~n8937;
  assign n8939 = ~g0 & ~n8938;
  assign n8940 = ~n8935 & ~n8939;
  assign n8941 = ~n5749 & ~n5777;
  assign n8942 = n5805 & ~n5897;
  assign n8943 = n5805 & n6027;
  assign n8944 = ~n5776 & ~n5798;
  assign n8945 = ~n8943 & ~n8944;
  assign n8946 = ~n8942 & n8945;
  assign n8947 = n8941 & ~n8946;
  assign n8948 = g0 & ~n8947;
  assign n8949 = ~n8941 & n8946;
  assign n8950 = n8948 & ~n8949;
  assign n8951 = ~n8322 & n8857;
  assign n8952 = n8322 & ~n8857;
  assign n8953 = ~n8951 & ~n8952;
  assign n8954 = ~g0 & ~n8953;
  assign n8955 = ~n8950 & ~n8954;
  assign n8956 = ~n8940 & ~n8955;
  assign n8957 = ~n8930 & n8956;
  assign n8958 = ~n8920 & n8957;
  assign n8959 = ~n7941 & n7944;
  assign n8960 = n7941 & ~n7944;
  assign n8961 = ~n8959 & ~n8960;
  assign n8962 = n8315 & ~n8961;
  assign n8963 = ~n8315 & n8961;
  assign n8964 = ~n8962 & ~n8963;
  assign n8965 = ~g0 & ~n8964;
  assign n8966 = g0 & ~n8538;
  assign n8967 = n6028 & n8966;
  assign n8968 = g0 & n8538;
  assign n8969 = ~n6028 & n8968;
  assign n8970 = ~n8967 & ~n8969;
  assign n8971 = ~n8965 & n8970;
  assign n8972 = n8066 & ~n8069;
  assign n8973 = ~n8066 & n8069;
  assign n8974 = ~n8972 & ~n8973;
  assign n8975 = ~n8309 & n8974;
  assign n8976 = n8309 & ~n8974;
  assign n8977 = ~n8975 & ~n8976;
  assign n8978 = ~g0 & ~n8977;
  assign n8979 = n5890 & ~n6025;
  assign n8980 = n8531 & n8979;
  assign n8981 = g0 & ~n8533;
  assign n8982 = ~n8980 & n8981;
  assign n8983 = ~n8978 & ~n8982;
  assign n8984 = n6022 & n8525;
  assign n8985 = g0 & ~n8526;
  assign n8986 = ~n8984 & n8985;
  assign n8987 = ~n8119 & n8150;
  assign n8988 = n8119 & ~n8150;
  assign n8989 = ~n8987 & ~n8988;
  assign n8990 = ~n8303 & ~n8989;
  assign n8991 = n8303 & n8989;
  assign n8992 = ~n8990 & ~n8991;
  assign n8993 = ~g0 & n8992;
  assign n8994 = ~n8986 & ~n8993;
  assign n8995 = g15 & ~n8994;
  assign n8996 = ~g15 & n8994;
  assign n8997 = ~g92 & n5929;
  assign n8998 = g92 & ~n5929;
  assign n8999 = ~n8997 & ~n8998;
  assign n9000 = n5912 & n8999;
  assign n9001 = ~n5912 & ~n8999;
  assign n9002 = ~n9000 & ~n9001;
  assign n9003 = n5937 & ~n5948;
  assign n9004 = ~n5937 & n5948;
  assign n9005 = ~n9003 & ~n9004;
  assign n9006 = ~g94 & n5948;
  assign n9007 = g94 & ~n5948;
  assign n9008 = ~n9006 & ~n9007;
  assign n9009 = n6013 & ~n9008;
  assign n9010 = ~n6014 & ~n9009;
  assign n9011 = ~n9005 & n9010;
  assign n9012 = ~n5949 & ~n9011;
  assign n9013 = n9002 & ~n9012;
  assign n9014 = ~n5933 & ~n9013;
  assign n9015 = ~g91 & n5913;
  assign n9016 = g91 & ~n5913;
  assign n9017 = ~n9015 & ~n9016;
  assign n9018 = n5881 & n9017;
  assign n9019 = ~n5881 & ~n9017;
  assign n9020 = ~n9018 & ~n9019;
  assign n9021 = ~n9014 & n9020;
  assign n9022 = n9014 & ~n9020;
  assign n9023 = g0 & ~n9022;
  assign n9024 = ~n9021 & n9023;
  assign n9025 = ~n8182 & ~n8184;
  assign n9026 = n8182 & n8184;
  assign n9027 = ~n9025 & ~n9026;
  assign n9028 = n8300 & n9027;
  assign n9029 = ~n8300 & ~n9027;
  assign n9030 = ~g0 & ~n9029;
  assign n9031 = ~n9028 & n9030;
  assign n9032 = ~n9024 & ~n9031;
  assign n9033 = ~g16 & n9032;
  assign n9034 = ~n8238 & ~n8239;
  assign n9035 = n8296 & n9034;
  assign n9036 = ~n8296 & ~n9034;
  assign n9037 = ~n9035 & ~n9036;
  assign n9038 = ~g0 & ~n9037;
  assign n9039 = n9005 & ~n9010;
  assign n9040 = ~n9011 & ~n9039;
  assign n9041 = g0 & n9040;
  assign n9042 = ~n9038 & ~n9041;
  assign n9043 = g18 & ~n9042;
  assign n9044 = g17 & n9043;
  assign n9045 = g0 & ~n9012;
  assign n9046 = ~n9002 & n9045;
  assign n9047 = ~n8219 & ~n8220;
  assign n9048 = ~n8298 & n9047;
  assign n9049 = n8298 & ~n9047;
  assign n9050 = ~g0 & ~n9049;
  assign n9051 = ~n9048 & n9050;
  assign n9052 = g0 & n9012;
  assign n9053 = n9002 & n9052;
  assign n9054 = ~n9051 & ~n9053;
  assign n9055 = ~n9046 & n9054;
  assign n9056 = ~g17 & ~n9043;
  assign n9057 = ~n9055 & ~n9056;
  assign n9058 = ~n9044 & ~n9057;
  assign n9059 = ~n9033 & ~n9058;
  assign n9060 = g16 & ~n9032;
  assign n9061 = ~n9059 & ~n9060;
  assign n9062 = ~n8996 & ~n9061;
  assign n9063 = ~n8995 & ~n9062;
  assign n9064 = ~n5886 & ~n5889;
  assign n9065 = ~n8527 & n9064;
  assign n9066 = n8527 & ~n9064;
  assign n9067 = g0 & ~n9066;
  assign n9068 = ~n9065 & n9067;
  assign n9069 = ~n8112 & n8115;
  assign n9070 = n8112 & ~n8115;
  assign n9071 = ~n9069 & ~n9070;
  assign n9072 = ~n8306 & n9071;
  assign n9073 = n8306 & ~n9071;
  assign n9074 = ~n9072 & ~n9073;
  assign n9075 = ~g0 & ~n9074;
  assign n9076 = ~n9068 & ~n9075;
  assign n9077 = ~g14 & n9076;
  assign n9078 = ~n9063 & ~n9077;
  assign n9079 = ~n8983 & n9078;
  assign n9080 = g14 & ~n9076;
  assign n9081 = ~n8983 & n9080;
  assign n9082 = ~n9079 & ~n9081;
  assign n9083 = ~n5842 & ~n8979;
  assign n9084 = ~n5894 & ~n9083;
  assign n9085 = ~n5827 & ~n5844;
  assign n9086 = g0 & ~n9085;
  assign n9087 = ~n9084 & n9086;
  assign n9088 = n8011 & ~n8014;
  assign n9089 = ~n8011 & n8014;
  assign n9090 = ~n9088 & ~n9089;
  assign n9091 = ~n8312 & n9090;
  assign n9092 = n8312 & ~n9090;
  assign n9093 = ~n9091 & ~n9092;
  assign n9094 = ~g0 & ~n9093;
  assign n9095 = g0 & n9085;
  assign n9096 = n9084 & n9095;
  assign n9097 = ~n9094 & ~n9096;
  assign n9098 = ~n9087 & n9097;
  assign n9099 = ~n9082 & ~n9098;
  assign n9100 = ~n8971 & n9099;
  assign n9101 = n8958 & n9100;
  assign n9102 = ~n8908 & n9101;
  assign n9103 = ~n8819 & n9102;
  assign n9104 = ~n8893 & n9103;
  assign n9105 = ~n8870 & n9104;
  assign n9106 = n8839 & n9105;
  assign n9107 = n8836 & n9106;
  assign n9108 = ~g0 & ~g2;
  assign n9109 = g0 & g2;
  assign n9110 = ~n9108 & ~n9109;
  assign n9111 = ~g1 & n9110;
  assign n9112 = g1 & ~n9110;
  assign n9113 = ~n9111 & ~n9112;
  assign n9114 = n6042 & ~n9113;
  assign n9115 = ~n9107 & n9114;
  assign n9116 = ~n8870 & ~n8908;
  assign n9117 = n9101 & n9116;
  assign n9118 = ~n8824 & n9117;
  assign n9119 = ~n8893 & n9118;
  assign n9120 = ~n8781 & n9119;
  assign n9121 = ~n8806 & n9120;
  assign n9122 = ~n8708 & ~n8760;
  assign n9123 = n9121 & n9122;
  assign n9124 = ~n8682 & n9123;
  assign n9125 = ~n8656 & n9124;
  assign n9126 = ~n8630 & n9125;
  assign n9127 = ~n8597 & n9126;
  assign n9128 = n6164 & ~n9127;
  assign n9129 = ~n9113 & n9128;
  assign n9130 = ~n9115 & n9129;
  assign n9131 = n9115 & ~n9129;
  assign n9132 = ~n9130 & ~n9131;
  assign n9133 = ~n8870 & ~n9113;
  assign n9134 = ~n8819 & ~n8893;
  assign n9135 = ~n8908 & n8958;
  assign n9136 = n9100 & n9135;
  assign n9137 = n9134 & n9136;
  assign n9138 = n9133 & n9137;
  assign n9139 = n8839 & n9138;
  assign n9140 = n6042 & n9139;
  assign n9141 = n8836 & n9140;
  assign n9142 = n6164 & ~n9113;
  assign n9143 = n9127 & n9142;
  assign n9144 = ~n9141 & n9143;
  assign n9145 = n9141 & ~n9143;
  assign n9146 = ~n9144 & ~n9145;
  assign n9147 = n9132 & n9146;
  assign n9148 = n9132 & n9147;
  assign n9149 = n9132 & n9148;
  assign n9150 = n9132 & n9149;
  assign n9151 = g36 & ~n110;
  assign n9152 = n758 & ~n762;
  assign n9153 = ~n110 & ~n9152;
  assign n9154 = ~n154 & ~n9153;
  assign n9155 = n154 & n9153;
  assign n9156 = ~n9154 & ~n9155;
  assign n9157 = ~n9151 & ~n9156;
  assign n9158 = n9151 & n9156;
  assign n9159 = ~n9157 & ~n9158;
  assign n9160 = n155 & n762;
  assign n9161 = ~n110 & ~n758;
  assign n9162 = ~n9160 & ~n9161;
  assign n9163 = ~n9151 & ~n9162;
  assign n9164 = n9151 & n9162;
  assign n9165 = ~n9163 & ~n9164;
  assign n9166 = ~g36 & n110;
  assign n9167 = ~n9151 & ~n9166;
  assign n9168 = n762 & n9167;
  assign n9169 = n155 & ~n758;
  assign n9170 = ~n9168 & ~n9169;
  assign n9171 = ~n730 & ~n733;
  assign n9172 = ~n126 & ~n9171;
  assign n9173 = ~n9170 & n9172;
  assign n9174 = n9170 & ~n9172;
  assign n9175 = ~n9173 & ~n9174;
  assign n9176 = n112 & ~n9175;
  assign n9177 = ~n9170 & ~n9172;
  assign n9178 = ~n9176 & ~n9177;
  assign n9179 = n9165 & ~n9178;
  assign n9180 = ~n9163 & ~n9179;
  assign n9181 = n9159 & ~n9180;
  assign n9182 = ~n9159 & n9180;
  assign n9183 = ~n9181 & ~n9182;
  assign n9184 = g39 & ~n110;
  assign n9185 = ~n698 & ~n700;
  assign n9186 = ~n198 & ~n9185;
  assign n9187 = g36 & n126;
  assign n9188 = ~g36 & ~n126;
  assign n9189 = ~n9187 & ~n9188;
  assign n9190 = n733 & ~n9189;
  assign n9191 = ~n129 & n730;
  assign n9192 = ~n9190 & ~n9191;
  assign n9193 = ~n9186 & n9192;
  assign n9194 = n9186 & ~n9192;
  assign n9195 = ~n9193 & ~n9194;
  assign n9196 = n9184 & ~n9195;
  assign n9197 = ~n9186 & ~n9192;
  assign n9198 = ~n9196 & ~n9197;
  assign n9199 = ~n129 & n733;
  assign n9200 = ~n126 & n730;
  assign n9201 = ~n9199 & ~n9200;
  assign n9202 = g38 & ~n110;
  assign n9203 = n113 & n762;
  assign n9204 = ~n758 & n9167;
  assign n9205 = ~n9203 & ~n9204;
  assign n9206 = n9202 & n9205;
  assign n9207 = ~n9202 & ~n9205;
  assign n9208 = ~n9206 & ~n9207;
  assign n9209 = n9201 & ~n9208;
  assign n9210 = ~n9201 & n9208;
  assign n9211 = ~n9209 & ~n9210;
  assign n9212 = n9198 & n9211;
  assign n9213 = ~n9198 & ~n9211;
  assign n9214 = ~n9212 & ~n9213;
  assign n9215 = n201 & n700;
  assign n9216 = ~n198 & n698;
  assign n9217 = ~n9215 & ~n9216;
  assign n9218 = ~g38 & n110;
  assign n9219 = ~n9202 & ~n9218;
  assign n9220 = n762 & n9219;
  assign n9221 = n113 & ~n758;
  assign n9222 = ~n9220 & ~n9221;
  assign n9223 = ~n9217 & n9222;
  assign n9224 = n9217 & ~n9222;
  assign n9225 = ~n9223 & ~n9224;
  assign n9226 = ~n758 & n9219;
  assign n9227 = ~n179 & n762;
  assign n9228 = ~n9226 & ~n9227;
  assign n9229 = ~n208 & n733;
  assign n9230 = n730 & ~n9189;
  assign n9231 = ~n9229 & ~n9230;
  assign n9232 = g40 & ~n110;
  assign n9233 = n9231 & n9232;
  assign n9234 = ~n9231 & ~n9232;
  assign n9235 = ~n9233 & ~n9234;
  assign n9236 = ~n9228 & ~n9235;
  assign n9237 = ~n9231 & n9232;
  assign n9238 = ~n9236 & ~n9237;
  assign n9239 = ~n9225 & ~n9238;
  assign n9240 = ~n9217 & ~n9222;
  assign n9241 = ~n9239 & ~n9240;
  assign n9242 = n9214 & ~n9241;
  assign n9243 = ~n9214 & n9241;
  assign n9244 = ~n9242 & ~n9243;
  assign n9245 = ~n9228 & n9235;
  assign n9246 = n9228 & ~n9235;
  assign n9247 = ~n9245 & ~n9246;
  assign n9248 = ~g40 & n110;
  assign n9249 = ~n9232 & ~n9248;
  assign n9250 = n762 & n9249;
  assign n9251 = ~n179 & ~n758;
  assign n9252 = ~n9250 & ~n9251;
  assign n9253 = g36 & n198;
  assign n9254 = ~g36 & ~n198;
  assign n9255 = ~n9253 & ~n9254;
  assign n9256 = n700 & ~n9255;
  assign n9257 = n201 & n698;
  assign n9258 = ~n9256 & ~n9257;
  assign n9259 = ~n710 & ~n715;
  assign n9260 = n314 & ~n9259;
  assign n9261 = ~n9258 & n9260;
  assign n9262 = n9258 & ~n9260;
  assign n9263 = ~n9261 & ~n9262;
  assign n9264 = ~n9252 & ~n9263;
  assign n9265 = ~n9258 & ~n9260;
  assign n9266 = ~n9264 & ~n9265;
  assign n9267 = n9217 & n9266;
  assign n9268 = ~n9217 & ~n9266;
  assign n9269 = ~n9267 & ~n9268;
  assign n9270 = ~n9247 & ~n9269;
  assign n9271 = n9217 & ~n9266;
  assign n9272 = ~n9270 & ~n9271;
  assign n9273 = n9184 & n9195;
  assign n9274 = ~n9184 & ~n9195;
  assign n9275 = ~n9273 & ~n9274;
  assign n9276 = ~n9225 & n9238;
  assign n9277 = n9225 & ~n9238;
  assign n9278 = ~n9276 & ~n9277;
  assign n9279 = ~n9275 & n9278;
  assign n9280 = n9275 & ~n9278;
  assign n9281 = ~n9279 & ~n9280;
  assign n9282 = ~n9272 & ~n9281;
  assign n9283 = ~n9275 & ~n9278;
  assign n9284 = ~n9282 & ~n9283;
  assign n9285 = n9244 & n9284;
  assign n9286 = n9202 & ~n9205;
  assign n9287 = ~n9209 & ~n9286;
  assign n9288 = ~n112 & ~n9175;
  assign n9289 = n112 & n9175;
  assign n9290 = ~n9288 & ~n9289;
  assign n9291 = ~n9201 & n9290;
  assign n9292 = n9201 & ~n9290;
  assign n9293 = ~n9291 & ~n9292;
  assign n9294 = ~n9287 & n9293;
  assign n9295 = n9287 & ~n9293;
  assign n9296 = ~n9294 & ~n9295;
  assign n9297 = ~n9214 & ~n9241;
  assign n9298 = ~n9198 & n9211;
  assign n9299 = ~n9297 & ~n9298;
  assign n9300 = n9296 & n9299;
  assign n9301 = ~n9285 & ~n9300;
  assign n9302 = n9165 & n9178;
  assign n9303 = ~n9165 & ~n9178;
  assign n9304 = ~n9302 & ~n9303;
  assign n9305 = ~n9287 & ~n9293;
  assign n9306 = ~n9201 & ~n9290;
  assign n9307 = ~n9305 & ~n9306;
  assign n9308 = n9304 & n9307;
  assign n9309 = ~n3398 & ~n3401;
  assign n9310 = ~n3392 & ~n3395;
  assign n9311 = ~n9309 & ~n9310;
  assign n9312 = ~n3376 & n3377;
  assign n9313 = ~n3370 & ~n3373;
  assign n9314 = ~n9312 & ~n9313;
  assign n9315 = ~n379 & n700;
  assign n9316 = n698 & ~n9255;
  assign n9317 = ~n9315 & ~n9316;
  assign n9318 = ~n339 & n733;
  assign n9319 = g38 & ~n126;
  assign n9320 = ~g38 & n126;
  assign n9321 = ~n9319 & ~n9320;
  assign n9322 = n730 & n9321;
  assign n9323 = ~n9318 & ~n9322;
  assign n9324 = n9317 & ~n9323;
  assign n9325 = ~n9317 & n9323;
  assign n9326 = ~n9324 & ~n9325;
  assign n9327 = n9314 & n9326;
  assign n9328 = ~n9314 & ~n9326;
  assign n9329 = ~n9327 & ~n9328;
  assign n9330 = ~n3358 & ~n3361;
  assign n9331 = ~n3353 & ~n3355;
  assign n9332 = ~n9330 & ~n9331;
  assign n9333 = n314 & n710;
  assign n9334 = n317 & n715;
  assign n9335 = ~n9333 & ~n9334;
  assign n9336 = ~n302 & n762;
  assign n9337 = ~n758 & n9249;
  assign n9338 = ~n9336 & ~n9337;
  assign n9339 = n1029 & n9338;
  assign n9340 = ~n1029 & ~n9338;
  assign n9341 = ~n9339 & ~n9340;
  assign n9342 = n9335 & ~n9341;
  assign n9343 = ~n9335 & n9341;
  assign n9344 = ~n9342 & ~n9343;
  assign n9345 = n9332 & ~n9344;
  assign n9346 = ~n9332 & n9344;
  assign n9347 = ~n9345 & ~n9346;
  assign n9348 = ~n9329 & n9347;
  assign n9349 = n9329 & ~n9347;
  assign n9350 = ~n9348 & ~n9349;
  assign n9351 = ~n3380 & n3386;
  assign n9352 = ~n3384 & ~n9351;
  assign n9353 = ~n9350 & n9352;
  assign n9354 = n9350 & ~n9352;
  assign n9355 = ~n9353 & ~n9354;
  assign n9356 = ~n3367 & ~n3389;
  assign n9357 = ~n3350 & ~n3364;
  assign n9358 = ~n9356 & ~n9357;
  assign n9359 = ~n9355 & n9358;
  assign n9360 = n9355 & ~n9358;
  assign n9361 = ~n9359 & ~n9360;
  assign n9362 = n9311 & n9361;
  assign n9363 = n3408 & ~n9362;
  assign n9364 = ~n9311 & ~n9361;
  assign n9365 = ~n9363 & ~n9364;
  assign n9366 = ~n9329 & ~n9347;
  assign n9367 = ~n9332 & ~n9344;
  assign n9368 = ~n9366 & ~n9367;
  assign n9369 = ~n9314 & n9326;
  assign n9370 = ~n9324 & ~n9369;
  assign n9371 = n733 & n9321;
  assign n9372 = ~n208 & n730;
  assign n9373 = ~n9371 & ~n9372;
  assign n9374 = g41 & ~n110;
  assign n9375 = n9373 & n9374;
  assign n9376 = ~n9373 & ~n9374;
  assign n9377 = ~n9375 & ~n9376;
  assign n9378 = ~n9317 & ~n9377;
  assign n9379 = n9317 & n9377;
  assign n9380 = ~n9378 & ~n9379;
  assign n9381 = n9252 & ~n9263;
  assign n9382 = ~n9252 & n9263;
  assign n9383 = ~n9381 & ~n9382;
  assign n9384 = ~n9335 & ~n9341;
  assign n9385 = n1029 & ~n9338;
  assign n9386 = ~n9384 & ~n9385;
  assign n9387 = n9383 & ~n9386;
  assign n9388 = ~n9383 & n9386;
  assign n9389 = ~n9387 & ~n9388;
  assign n9390 = ~n9380 & ~n9389;
  assign n9391 = n9380 & n9389;
  assign n9392 = ~n9390 & ~n9391;
  assign n9393 = ~n9370 & n9392;
  assign n9394 = n9370 & ~n9392;
  assign n9395 = ~n9393 & ~n9394;
  assign n9396 = n9368 & ~n9395;
  assign n9397 = ~n9368 & n9395;
  assign n9398 = ~n9396 & ~n9397;
  assign n9399 = ~n9355 & ~n9358;
  assign n9400 = ~n9350 & ~n9352;
  assign n9401 = ~n9399 & ~n9400;
  assign n9402 = n9398 & n9401;
  assign n9403 = ~n9365 & ~n9402;
  assign n9404 = ~n9398 & ~n9401;
  assign n9405 = ~n9403 & ~n9404;
  assign n9406 = ~n9362 & ~n9402;
  assign n9407 = ~n2034 & ~n3409;
  assign n9408 = n9406 & n9407;
  assign n9409 = n9405 & ~n9408;
  assign n9410 = n9272 & ~n9281;
  assign n9411 = ~n9272 & n9281;
  assign n9412 = ~n9410 & ~n9411;
  assign n9413 = n9380 & ~n9389;
  assign n9414 = ~n9383 & ~n9386;
  assign n9415 = ~n9413 & ~n9414;
  assign n9416 = ~n9373 & n9374;
  assign n9417 = ~n9378 & ~n9416;
  assign n9418 = n9247 & ~n9269;
  assign n9419 = ~n9247 & n9269;
  assign n9420 = ~n9418 & ~n9419;
  assign n9421 = ~n9417 & n9420;
  assign n9422 = n9417 & ~n9420;
  assign n9423 = ~n9421 & ~n9422;
  assign n9424 = ~n9415 & ~n9423;
  assign n9425 = ~n9417 & ~n9420;
  assign n9426 = ~n9424 & ~n9425;
  assign n9427 = n9412 & n9426;
  assign n9428 = n9415 & ~n9423;
  assign n9429 = ~n9415 & n9423;
  assign n9430 = ~n9428 & ~n9429;
  assign n9431 = ~n9368 & ~n9395;
  assign n9432 = ~n9370 & ~n9392;
  assign n9433 = ~n9431 & ~n9432;
  assign n9434 = n9430 & n9433;
  assign n9435 = ~n9427 & ~n9434;
  assign n9436 = ~n9409 & n9435;
  assign n9437 = ~n9308 & n9436;
  assign n9438 = n9301 & n9437;
  assign n9439 = ~n9430 & ~n9433;
  assign n9440 = ~n9427 & n9439;
  assign n9441 = ~n9412 & ~n9426;
  assign n9442 = ~n9440 & ~n9441;
  assign n9443 = n9301 & ~n9442;
  assign n9444 = ~n9244 & ~n9284;
  assign n9445 = ~n9300 & n9444;
  assign n9446 = ~n9296 & ~n9299;
  assign n9447 = ~n9445 & ~n9446;
  assign n9448 = ~n9443 & n9447;
  assign n9449 = ~n9308 & ~n9448;
  assign n9450 = ~n9304 & ~n9307;
  assign n9451 = ~n9449 & ~n9450;
  assign n9452 = ~n9438 & n9451;
  assign n9453 = ~n9183 & ~n9452;
  assign n9454 = n9183 & n9452;
  assign n9455 = n9113 & ~n9454;
  assign n9456 = ~n9453 & n9455;
  assign n9457 = ~n9115 & ~n9456;
  assign n9458 = ~n9129 & ~n9456;
  assign n9459 = n9457 & ~n9458;
  assign n9460 = ~n9457 & n9458;
  assign n9461 = ~n9459 & ~n9460;
  assign n9462 = ~n9304 & n9307;
  assign n9463 = n9304 & ~n9307;
  assign n9464 = ~n9462 & ~n9463;
  assign n9465 = n9301 & n9464;
  assign n9466 = n9435 & n9465;
  assign n9467 = ~n9405 & n9466;
  assign n9468 = n9412 & ~n9426;
  assign n9469 = ~n9412 & n9426;
  assign n9470 = ~n9468 & ~n9469;
  assign n9471 = ~n9430 & n9433;
  assign n9472 = n9430 & ~n9433;
  assign n9473 = ~n9471 & ~n9472;
  assign n9474 = ~n9409 & ~n9473;
  assign n9475 = ~n9439 & ~n9474;
  assign n9476 = ~n9470 & ~n9475;
  assign n9477 = ~n9441 & ~n9476;
  assign n9478 = n9301 & ~n9477;
  assign n9479 = n9447 & ~n9464;
  assign n9480 = ~n9478 & n9479;
  assign n9481 = ~n9442 & n9465;
  assign n9482 = ~n9447 & n9464;
  assign n9483 = ~n9481 & ~n9482;
  assign n9484 = n9408 & n9466;
  assign n9485 = n9483 & ~n9484;
  assign n9486 = ~n9480 & n9485;
  assign n9487 = ~n9467 & n9486;
  assign n9488 = n9113 & ~n9487;
  assign n9489 = ~n9115 & ~n9488;
  assign n9490 = ~n9129 & ~n9488;
  assign n9491 = n9489 & ~n9490;
  assign n9492 = ~n9489 & n9490;
  assign n9493 = ~n9491 & ~n9492;
  assign n9494 = n9461 & n9493;
  assign n9495 = n9132 & n9494;
  assign n9496 = ~n8431 & ~n8485;
  assign n9497 = ~n8468 & n8839;
  assign n9498 = n8836 & n9105;
  assign n9499 = n9497 & n9498;
  assign n9500 = n9496 & n9499;
  assign n9501 = n9114 & ~n9500;
  assign n9502 = ~n9296 & n9299;
  assign n9503 = n9296 & ~n9299;
  assign n9504 = ~n9502 & ~n9503;
  assign n9505 = ~n9244 & n9284;
  assign n9506 = n9244 & ~n9284;
  assign n9507 = ~n9505 & ~n9506;
  assign n9508 = n9477 & ~n9507;
  assign n9509 = ~n9285 & ~n9508;
  assign n9510 = ~n9504 & ~n9509;
  assign n9511 = n9504 & n9509;
  assign n9512 = ~n9510 & ~n9511;
  assign n9513 = n9113 & ~n9512;
  assign n9514 = ~n9501 & ~n9513;
  assign n9515 = ~n9129 & ~n9513;
  assign n9516 = n9514 & ~n9515;
  assign n9517 = ~n9514 & n9515;
  assign n9518 = ~n9516 & ~n9517;
  assign n9519 = ~n8468 & ~n8699;
  assign n9520 = ~n8777 & ~n8800;
  assign n9521 = ~n8750 & n9520;
  assign n9522 = n9105 & n9521;
  assign n9523 = ~n8485 & n9522;
  assign n9524 = n8431 & ~n9113;
  assign n9525 = n8836 & n9524;
  assign n9526 = n9523 & n9525;
  assign n9527 = n9519 & n9526;
  assign n9528 = n9519 & n9523;
  assign n9529 = n8836 & n9528;
  assign n9530 = ~n9113 & ~n9529;
  assign n9531 = ~n8431 & n9530;
  assign n9532 = ~n9477 & ~n9507;
  assign n9533 = n9477 & n9507;
  assign n9534 = n9113 & ~n9533;
  assign n9535 = ~n9532 & n9534;
  assign n9536 = ~n9531 & ~n9535;
  assign n9537 = ~n9527 & n9536;
  assign n9538 = ~n8455 & ~n9113;
  assign n9539 = ~n8507 & ~n8593;
  assign n9540 = ~n8489 & ~n9539;
  assign n9541 = n9538 & ~n9540;
  assign n9542 = ~n8469 & n9126;
  assign n9543 = n9538 & ~n9542;
  assign n9544 = n8455 & ~n9113;
  assign n9545 = n9126 & n9540;
  assign n9546 = n9544 & n9545;
  assign n9547 = ~n8469 & n9546;
  assign n9548 = ~n9543 & ~n9547;
  assign n9549 = ~n9541 & n9548;
  assign n9550 = ~n9535 & n9549;
  assign n9551 = n9537 & ~n9550;
  assign n9552 = ~n9537 & n9550;
  assign n9553 = ~n9551 & ~n9552;
  assign n9554 = n9470 & n9475;
  assign n9555 = n9113 & ~n9554;
  assign n9556 = ~n9476 & n9555;
  assign n9557 = ~n8508 & n8839;
  assign n9558 = ~n8485 & n9557;
  assign n9559 = ~n8622 & n9558;
  assign n9560 = ~n8468 & ~n9113;
  assign n9561 = ~n9559 & n9560;
  assign n9562 = n8468 & ~n9113;
  assign n9563 = ~n8651 & n9105;
  assign n9564 = ~n8677 & n9563;
  assign n9565 = ~n9562 & n9564;
  assign n9566 = n9559 & ~n9565;
  assign n9567 = ~n9561 & ~n9566;
  assign n9568 = ~n9560 & ~n9564;
  assign n9569 = ~n9567 & ~n9568;
  assign n9570 = ~n9556 & ~n9569;
  assign n9571 = ~n8469 & ~n9113;
  assign n9572 = ~n9545 & n9571;
  assign n9573 = n8469 & ~n9113;
  assign n9574 = n9540 & n9573;
  assign n9575 = n9126 & n9574;
  assign n9576 = ~n9572 & ~n9575;
  assign n9577 = ~n9556 & n9576;
  assign n9578 = n9570 & ~n9577;
  assign n9579 = ~n9570 & n9577;
  assign n9580 = ~n9578 & ~n9579;
  assign n9581 = n9553 & n9580;
  assign n9582 = n9518 & n9581;
  assign n9583 = n9495 & n9582;
  assign n9584 = n9132 & n9583;
  assign n9585 = n8485 & ~n9113;
  assign n9586 = n9106 & n9585;
  assign n9587 = n8836 & n9586;
  assign n9588 = n9409 & n9473;
  assign n9589 = n9113 & ~n9474;
  assign n9590 = ~n9588 & n9589;
  assign n9591 = ~n8485 & ~n9113;
  assign n9592 = ~n9107 & n9591;
  assign n9593 = ~n9590 & ~n9592;
  assign n9594 = ~n9587 & n9593;
  assign n9595 = n8489 & ~n9127;
  assign n9596 = ~n9113 & ~n9595;
  assign n9597 = ~n9545 & n9596;
  assign n9598 = ~n9590 & ~n9597;
  assign n9599 = n9594 & ~n9598;
  assign n9600 = ~n9594 & n9598;
  assign n9601 = ~n9599 & ~n9600;
  assign n9602 = n8839 & n9564;
  assign n9603 = n8508 & n9602;
  assign n9604 = ~n8622 & n9603;
  assign n9605 = ~n9113 & n9604;
  assign n9606 = ~n2034 & n3410;
  assign n9607 = ~n3408 & ~n9606;
  assign n9608 = n9398 & ~n9401;
  assign n9609 = ~n9398 & n9401;
  assign n9610 = ~n9608 & ~n9609;
  assign n9611 = ~n9364 & ~n9610;
  assign n9612 = n9607 & n9611;
  assign n9613 = ~n9362 & ~n9607;
  assign n9614 = n9610 & n9613;
  assign n9615 = ~n9612 & ~n9614;
  assign n9616 = ~n9364 & n9610;
  assign n9617 = ~n9362 & ~n9610;
  assign n9618 = ~n9616 & ~n9617;
  assign n9619 = n9615 & ~n9618;
  assign n9620 = n9113 & ~n9619;
  assign n9621 = ~n8622 & n9602;
  assign n9622 = ~n9113 & ~n9621;
  assign n9623 = ~n8508 & n9622;
  assign n9624 = ~n9620 & ~n9623;
  assign n9625 = ~n9605 & n9624;
  assign n9626 = n8597 & ~n9126;
  assign n9627 = ~n9113 & ~n9127;
  assign n9628 = ~n9626 & n9627;
  assign n9629 = ~n9620 & ~n9628;
  assign n9630 = n9625 & ~n9629;
  assign n9631 = ~n9625 & n9629;
  assign n9632 = ~n9630 & ~n9631;
  assign n9633 = n9601 & n9632;
  assign n9634 = ~n9311 & n9361;
  assign n9635 = n9311 & ~n9361;
  assign n9636 = ~n9634 & ~n9635;
  assign n9637 = ~n9607 & ~n9636;
  assign n9638 = n9607 & n9636;
  assign n9639 = ~n9637 & ~n9638;
  assign n9640 = n9113 & n9639;
  assign n9641 = n8622 & ~n9113;
  assign n9642 = n9602 & n9641;
  assign n9643 = ~n8622 & ~n9113;
  assign n9644 = ~n9602 & n9643;
  assign n9645 = ~n9642 & ~n9644;
  assign n9646 = ~n9640 & n9645;
  assign n9647 = n8630 & ~n9125;
  assign n9648 = ~n9113 & ~n9647;
  assign n9649 = ~n9126 & n9648;
  assign n9650 = ~n9640 & ~n9649;
  assign n9651 = n9646 & ~n9650;
  assign n9652 = ~n9646 & n9650;
  assign n9653 = ~n9651 & ~n9652;
  assign n9654 = ~n8677 & n9106;
  assign n9655 = ~n8651 & n9654;
  assign n9656 = n8651 & ~n9654;
  assign n9657 = ~n9113 & ~n9656;
  assign n9658 = ~n9655 & n9657;
  assign n9659 = n2034 & n3410;
  assign n9660 = ~n2034 & ~n3410;
  assign n9661 = ~n9659 & ~n9660;
  assign n9662 = n9113 & ~n9661;
  assign n9663 = ~n9658 & ~n9662;
  assign n9664 = n8656 & ~n9124;
  assign n9665 = ~n9113 & ~n9664;
  assign n9666 = ~n9125 & n9665;
  assign n9667 = ~n9662 & ~n9666;
  assign n9668 = n9663 & ~n9667;
  assign n9669 = ~n9663 & n9667;
  assign n9670 = ~n9668 & ~n9669;
  assign n9671 = n991 & ~n1062;
  assign n9672 = ~n991 & n1062;
  assign n9673 = ~n9671 & ~n9672;
  assign n9674 = ~n1442 & ~n2021;
  assign n9675 = ~n2013 & n9674;
  assign n9676 = n2011 & n9675;
  assign n9677 = n2017 & ~n2020;
  assign n9678 = ~n2017 & n2020;
  assign n9679 = ~n9677 & ~n9678;
  assign n9680 = ~n1556 & ~n9679;
  assign n9681 = n9674 & ~n9680;
  assign n9682 = ~n1441 & ~n9681;
  assign n9683 = ~n9676 & n9682;
  assign n9684 = n1239 & ~n1346;
  assign n9685 = ~n1239 & n1346;
  assign n9686 = ~n9684 & ~n9685;
  assign n9687 = n9683 & ~n9686;
  assign n9688 = ~n1347 & ~n9687;
  assign n9689 = n1143 & ~n1235;
  assign n9690 = ~n1143 & n1235;
  assign n9691 = ~n9689 & ~n9690;
  assign n9692 = ~n9688 & ~n9691;
  assign n9693 = ~n1349 & ~n9692;
  assign n9694 = ~n1359 & n9693;
  assign n9695 = n9673 & n9694;
  assign n9696 = ~n1357 & ~n9693;
  assign n9697 = ~n9673 & n9696;
  assign n9698 = n1357 & n9673;
  assign n9699 = n1359 & ~n9673;
  assign n9700 = n9113 & ~n9699;
  assign n9701 = ~n9698 & n9700;
  assign n9702 = ~n9697 & n9701;
  assign n9703 = ~n9695 & n9702;
  assign n9704 = n8677 & ~n9106;
  assign n9705 = ~n9113 & ~n9704;
  assign n9706 = ~n9654 & n9705;
  assign n9707 = ~n9703 & ~n9706;
  assign n9708 = n8682 & ~n9123;
  assign n9709 = ~n9113 & ~n9708;
  assign n9710 = ~n9124 & n9709;
  assign n9711 = ~n9703 & ~n9710;
  assign n9712 = n9707 & ~n9711;
  assign n9713 = ~n9707 & n9711;
  assign n9714 = ~n9712 & ~n9713;
  assign n9715 = n9670 & n9714;
  assign n9716 = n9653 & n9715;
  assign n9717 = n9633 & n9716;
  assign n9718 = n878 & ~n1353;
  assign n9719 = ~n878 & n1353;
  assign n9720 = ~n9718 & ~n9719;
  assign n9721 = n988 & ~n9720;
  assign n9722 = ~n988 & n9720;
  assign n9723 = ~n9721 & ~n9722;
  assign n9724 = n9693 & n9723;
  assign n9725 = ~n9693 & ~n9723;
  assign n9726 = ~n9724 & ~n9725;
  assign n9727 = n9113 & n9726;
  assign n9728 = n8699 & ~n9113;
  assign n9729 = n9105 & n9728;
  assign n9730 = n9521 & n9729;
  assign n9731 = ~n8699 & ~n9113;
  assign n9732 = ~n9522 & n9731;
  assign n9733 = ~n9730 & ~n9732;
  assign n9734 = ~n9727 & n9733;
  assign n9735 = ~n8760 & n9121;
  assign n9736 = n8708 & ~n9735;
  assign n9737 = ~n9123 & ~n9736;
  assign n9738 = ~n9113 & n9737;
  assign n9739 = ~n9727 & ~n9738;
  assign n9740 = n9734 & ~n9739;
  assign n9741 = ~n9734 & n9739;
  assign n9742 = ~n9740 & ~n9741;
  assign n9743 = n9688 & ~n9691;
  assign n9744 = ~n9688 & n9691;
  assign n9745 = ~n9743 & ~n9744;
  assign n9746 = n9113 & ~n9745;
  assign n9747 = ~n8777 & ~n8870;
  assign n9748 = ~n8800 & n9747;
  assign n9749 = ~n8750 & n9102;
  assign n9750 = n9748 & n9749;
  assign n9751 = n9134 & n9750;
  assign n9752 = n8750 & ~n9102;
  assign n9753 = n9134 & n9748;
  assign n9754 = n8750 & ~n9753;
  assign n9755 = ~n9113 & ~n9754;
  assign n9756 = ~n9752 & n9755;
  assign n9757 = ~n9751 & n9756;
  assign n9758 = ~n9746 & ~n9757;
  assign n9759 = n8760 & ~n9121;
  assign n9760 = ~n9735 & ~n9759;
  assign n9761 = ~n9113 & n9760;
  assign n9762 = ~n9746 & ~n9761;
  assign n9763 = n9758 & ~n9762;
  assign n9764 = ~n9758 & n9762;
  assign n9765 = ~n9763 & ~n9764;
  assign n9766 = n8777 & ~n9113;
  assign n9767 = n9105 & n9766;
  assign n9768 = ~n8800 & n9767;
  assign n9769 = ~n8800 & n9105;
  assign n9770 = ~n9113 & ~n9769;
  assign n9771 = ~n8777 & n9770;
  assign n9772 = ~n9683 & ~n9686;
  assign n9773 = n9683 & n9686;
  assign n9774 = ~n9772 & ~n9773;
  assign n9775 = n9113 & ~n9774;
  assign n9776 = ~n9771 & ~n9775;
  assign n9777 = ~n9768 & n9776;
  assign n9778 = ~n8806 & n9119;
  assign n9779 = n8781 & ~n9778;
  assign n9780 = ~n9113 & ~n9779;
  assign n9781 = ~n9121 & n9780;
  assign n9782 = ~n9775 & ~n9781;
  assign n9783 = n9777 & ~n9782;
  assign n9784 = ~n9777 & n9782;
  assign n9785 = ~n9783 & ~n9784;
  assign n9786 = n9765 & n9785;
  assign n9787 = n9742 & n9786;
  assign n9788 = ~n8800 & ~n9105;
  assign n9789 = n8800 & n9105;
  assign n9790 = ~n9788 & ~n9789;
  assign n9791 = ~n9113 & n9790;
  assign n9792 = ~n1364 & ~n2024;
  assign n9793 = n1440 & n9792;
  assign n9794 = n1364 & ~n2024;
  assign n9795 = ~n1440 & n9794;
  assign n9796 = ~n1364 & n1440;
  assign n9797 = n1364 & ~n1440;
  assign n9798 = ~n9796 & ~n9797;
  assign n9799 = n2024 & n9798;
  assign n9800 = ~n9795 & ~n9799;
  assign n9801 = ~n9793 & n9800;
  assign n9802 = n9113 & n9801;
  assign n9803 = ~n9791 & ~n9802;
  assign n9804 = ~n8893 & n9117;
  assign n9805 = ~n8824 & n9804;
  assign n9806 = n8806 & ~n9805;
  assign n9807 = ~n9113 & ~n9806;
  assign n9808 = ~n9778 & n9807;
  assign n9809 = n9113 & ~n9801;
  assign n9810 = ~n9808 & ~n9809;
  assign n9811 = ~n9803 & ~n9810;
  assign n9812 = n9803 & n9810;
  assign n9813 = ~n9811 & ~n9812;
  assign n9814 = ~n2014 & n9679;
  assign n9815 = n2014 & ~n9679;
  assign n9816 = ~n9814 & ~n9815;
  assign n9817 = n9113 & ~n9816;
  assign n9818 = ~n8870 & n8958;
  assign n9819 = n9100 & n9818;
  assign n9820 = ~n8908 & n9819;
  assign n9821 = n8819 & ~n9113;
  assign n9822 = n9820 & n9821;
  assign n9823 = ~n8893 & n9822;
  assign n9824 = ~n8893 & n9820;
  assign n9825 = ~n8819 & ~n9113;
  assign n9826 = ~n9824 & n9825;
  assign n9827 = ~n9823 & ~n9826;
  assign n9828 = ~n9817 & n9827;
  assign n9829 = n8824 & ~n9804;
  assign n9830 = ~n9113 & ~n9829;
  assign n9831 = ~n9805 & n9830;
  assign n9832 = ~n9817 & ~n9831;
  assign n9833 = n9828 & ~n9832;
  assign n9834 = ~n9828 & n9832;
  assign n9835 = ~n9833 & ~n9834;
  assign n9836 = n6167 & n9835;
  assign n9837 = n9813 & n9836;
  assign n9838 = n9787 & n9837;
  assign n9839 = n9717 & n9838;
  assign n9840 = n9584 & n9839;
  assign n9841 = n9150 & n9840;
  assign miter = ~n8833 | ~n9841;
endmodule


