module top (out_0, out_1, out_2, out_3, out_4, out_5, out_6, out_7, out_8, out_9, out_10, out_11, out_12, out_13, out_14, out_15, out_16, out_17, out_18, out_19, out_20, out_21, in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, in_17, in_18, in_19, in_20, in_21);
	input in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, in_17, in_18, in_19, in_20, in_21;
	output out_0, out_1, out_2, out_3, out_4, out_5, out_6, out_7, out_8, out_9, out_10, out_11, out_12, out_13, out_14, out_15, out_16, out_17, out_18, out_19, out_20, out_21;
	wire gm_n100, gm_n1000, gm_n1001, gm_n1002, gm_n1003, gm_n1004, gm_n1005, gm_n1006, gm_n1007, gm_n1008, gm_n1009, gm_n101, gm_n1010, gm_n1011, gm_n1012, gm_n1013, gm_n1014, gm_n1015, gm_n1016, gm_n1017, gm_n1018, gm_n1019, gm_n102, gm_n1020, gm_n1021, gm_n1022, gm_n1023, gm_n1024, gm_n1025, gm_n1026, gm_n1027, gm_n1028, gm_n1029, gm_n103, gm_n1030, gm_n1031, gm_n1032, gm_n1033, gm_n1034, gm_n1035, gm_n1036, gm_n1037, gm_n1038, gm_n1039, gm_n104, gm_n1040, gm_n1041, gm_n1042, gm_n1043, gm_n1044, gm_n1045, gm_n1046, gm_n1047, gm_n1048, gm_n1049, gm_n105, gm_n1050, gm_n1051, gm_n1052, gm_n1053, gm_n1054, gm_n1055, gm_n1056, gm_n1057, gm_n1058, gm_n1059, gm_n106, gm_n1060, gm_n1061, gm_n1062, gm_n1063, gm_n1064, gm_n1065, gm_n1066, gm_n1067, gm_n1068, gm_n1069, gm_n107, gm_n1070, gm_n1071, gm_n1072, gm_n1073, gm_n1074, gm_n1075, gm_n1076, gm_n1077, gm_n1078, gm_n1079, gm_n108, gm_n1080, gm_n1081, gm_n1082, gm_n1083, gm_n1084, gm_n1085, gm_n1086, gm_n1087, gm_n1088, gm_n1089, gm_n109, gm_n1090, gm_n1091, gm_n1092, gm_n1093, gm_n1094, gm_n1095, gm_n1096, gm_n1097, gm_n1098, gm_n1099, gm_n110, gm_n1100, gm_n1101, gm_n1102, gm_n1103, gm_n1104, gm_n1105, gm_n1106, gm_n1107, gm_n1108, gm_n1109, gm_n111, gm_n1110, gm_n1112, gm_n1113, gm_n1114, gm_n1115, gm_n1116, gm_n1117, gm_n1118, gm_n1119, gm_n112, gm_n1120, gm_n1121, gm_n1122, gm_n1123, gm_n1124, gm_n1125, gm_n1126, gm_n1127, gm_n1128, gm_n1129, gm_n113, gm_n1130, gm_n1131, gm_n1132, gm_n1133, gm_n1134, gm_n1135, gm_n1136, gm_n1137, gm_n1138, gm_n1139, gm_n114, gm_n1140, gm_n1141, gm_n1142, gm_n1143, gm_n1144, gm_n1145, gm_n1146, gm_n1147, gm_n1148, gm_n1149, gm_n115, gm_n1150, gm_n1151, gm_n1152, gm_n1153, gm_n1154, gm_n1155, gm_n1156, gm_n1157, gm_n1158, gm_n1159, gm_n116, gm_n1160, gm_n1161, gm_n1162, gm_n1163, gm_n1164, gm_n1165, gm_n1166, gm_n1167, gm_n1168, gm_n1169, gm_n117, gm_n1170, gm_n1171, gm_n1172, gm_n1173, gm_n1174, gm_n1175, gm_n1176, gm_n1177, gm_n1178, gm_n1179, gm_n118, gm_n1180, gm_n1181, gm_n1182, gm_n1183, gm_n1184, gm_n1185, gm_n1186, gm_n1187, gm_n1188, gm_n1189, gm_n119, gm_n1190, gm_n1191, gm_n1192, gm_n1193, gm_n1194, gm_n1195, gm_n1196, gm_n1197, gm_n1198, gm_n1199, gm_n120, gm_n1200, gm_n1201, gm_n1202, gm_n1203, gm_n1204, gm_n1205, gm_n1206, gm_n1207, gm_n1208, gm_n1209, gm_n121, gm_n1210, gm_n1211, gm_n1212, gm_n1213, gm_n1214, gm_n1215, gm_n1216, gm_n1217, gm_n1218, gm_n1219, gm_n122, gm_n1220, gm_n1221, gm_n1222, gm_n1223, gm_n1224, gm_n1225, gm_n1226, gm_n1227, gm_n1228, gm_n1229, gm_n123, gm_n1230, gm_n1231, gm_n1232, gm_n1233, gm_n1234, gm_n1235, gm_n1236, gm_n1237, gm_n1238, gm_n1239, gm_n124, gm_n1240, gm_n1241, gm_n1242, gm_n1243, gm_n1244, gm_n1245, gm_n1246, gm_n1247, gm_n1248, gm_n1249, gm_n125, gm_n1250, gm_n1251, gm_n1252, gm_n1253, gm_n1254, gm_n1255, gm_n1256, gm_n1257, gm_n1258, gm_n1259, gm_n126, gm_n1260, gm_n1261, gm_n1262, gm_n1263, gm_n1264, gm_n1265, gm_n1266, gm_n1267, gm_n1268, gm_n1269, gm_n127, gm_n1270, gm_n1271, gm_n1272, gm_n1273, gm_n1274, gm_n1275, gm_n1276, gm_n1277, gm_n1278, gm_n1279, gm_n128, gm_n1280, gm_n1281, gm_n1282, gm_n1283, gm_n1284, gm_n1285, gm_n1286, gm_n1287, gm_n1288, gm_n1289, gm_n129, gm_n1290, gm_n1291, gm_n1292, gm_n1293, gm_n1294, gm_n1295, gm_n1296, gm_n1297, gm_n1298, gm_n1299, gm_n130, gm_n1300, gm_n1301, gm_n1302, gm_n1303, gm_n1304, gm_n1305, gm_n1306, gm_n1307, gm_n1308, gm_n1309, gm_n131, gm_n1310, gm_n1311, gm_n1312, gm_n1313, gm_n1314, gm_n1315, gm_n1316, gm_n1317, gm_n1318, gm_n1319, gm_n132, gm_n1320, gm_n1321, gm_n1322, gm_n1323, gm_n1324, gm_n1325, gm_n1326, gm_n1327, gm_n1328, gm_n1329, gm_n133, gm_n1330, gm_n1331, gm_n1332, gm_n1333, gm_n1334, gm_n1335, gm_n1336, gm_n1337, gm_n1338, gm_n1339, gm_n134, gm_n1340, gm_n1341, gm_n1342, gm_n1343, gm_n1344, gm_n1345, gm_n1346, gm_n1347, gm_n1348, gm_n1349, gm_n135, gm_n1350, gm_n1351, gm_n1352, gm_n1353, gm_n1354, gm_n1355, gm_n1356, gm_n1357, gm_n1358, gm_n1359, gm_n136, gm_n1360, gm_n1361, gm_n1362, gm_n1363, gm_n1364, gm_n1365, gm_n1366, gm_n1367, gm_n1368, gm_n1369, gm_n137, gm_n1370, gm_n1371, gm_n1372, gm_n1373, gm_n1374, gm_n1375, gm_n1376, gm_n1377, gm_n1378, gm_n1379, gm_n138, gm_n1380, gm_n1381, gm_n1382, gm_n1383, gm_n1384, gm_n1385, gm_n1386, gm_n1387, gm_n1388, gm_n1389, gm_n139, gm_n1390, gm_n1391, gm_n1392, gm_n1393, gm_n1394, gm_n1395, gm_n1396, gm_n1397, gm_n1398, gm_n1399, gm_n140, gm_n1400, gm_n1401, gm_n1402, gm_n1403, gm_n1404, gm_n1405, gm_n1406, gm_n1407, gm_n1408, gm_n1409, gm_n141, gm_n1410, gm_n1411, gm_n1412, gm_n1413, gm_n1414, gm_n1415, gm_n1416, gm_n1417, gm_n1418, gm_n1419, gm_n142, gm_n1420, gm_n1421, gm_n1422, gm_n1423, gm_n1424, gm_n1425, gm_n1426, gm_n1427, gm_n1428, gm_n1429, gm_n143, gm_n1430, gm_n1431, gm_n1432, gm_n1433, gm_n1434, gm_n1435, gm_n1436, gm_n1437, gm_n1438, gm_n1439, gm_n144, gm_n1440, gm_n1441, gm_n1442, gm_n1443, gm_n1444, gm_n1445, gm_n1446, gm_n1447, gm_n1448, gm_n1449, gm_n145, gm_n1450, gm_n1451, gm_n1452, gm_n1453, gm_n1454, gm_n1455, gm_n1456, gm_n1457, gm_n1458, gm_n1459, gm_n146, gm_n1460, gm_n1461, gm_n1462, gm_n1463, gm_n1464, gm_n1465, gm_n1466, gm_n1467, gm_n1468, gm_n1469, gm_n147, gm_n1470, gm_n1471, gm_n1472, gm_n1473, gm_n1474, gm_n1475, gm_n1476, gm_n1477, gm_n1478, gm_n1479, gm_n148, gm_n1480, gm_n1481, gm_n1482, gm_n1483, gm_n1484, gm_n1485, gm_n1486, gm_n1487, gm_n1488, gm_n1489, gm_n149, gm_n1490, gm_n1491, gm_n1492, gm_n1493, gm_n1494, gm_n1495, gm_n1496, gm_n1497, gm_n1498, gm_n1499, gm_n150, gm_n1500, gm_n1501, gm_n1502, gm_n1503, gm_n1504, gm_n1505, gm_n1506, gm_n1508, gm_n1509, gm_n151, gm_n1510, gm_n1511, gm_n1512, gm_n1513, gm_n1514, gm_n1515, gm_n1516, gm_n1517, gm_n1518, gm_n1519, gm_n152, gm_n1520, gm_n1521, gm_n1522, gm_n1523, gm_n1524, gm_n1525, gm_n1526, gm_n1527, gm_n1528, gm_n1529, gm_n153, gm_n1530, gm_n1531, gm_n1532, gm_n1533, gm_n1534, gm_n1535, gm_n1536, gm_n1537, gm_n1538, gm_n1539, gm_n154, gm_n1540, gm_n1541, gm_n1542, gm_n1543, gm_n1544, gm_n1545, gm_n1546, gm_n1547, gm_n1548, gm_n1549, gm_n155, gm_n1550, gm_n1551, gm_n1552, gm_n1553, gm_n1554, gm_n1555, gm_n1556, gm_n1557, gm_n1558, gm_n1559, gm_n156, gm_n1560, gm_n1561, gm_n1562, gm_n1563, gm_n1564, gm_n1565, gm_n1566, gm_n1567, gm_n1568, gm_n1569, gm_n157, gm_n1570, gm_n1571, gm_n1572, gm_n1573, gm_n1574, gm_n1575, gm_n1576, gm_n1577, gm_n1578, gm_n1579, gm_n158, gm_n1580, gm_n1581, gm_n1582, gm_n1583, gm_n1584, gm_n1585, gm_n1586, gm_n1587, gm_n1588, gm_n1589, gm_n159, gm_n1590, gm_n1591, gm_n1592, gm_n1593, gm_n1594, gm_n1595, gm_n1596, gm_n1597, gm_n1598, gm_n1599, gm_n160, gm_n1600, gm_n1601, gm_n1602, gm_n1603, gm_n1604, gm_n1605, gm_n1606, gm_n1607, gm_n1608, gm_n1609, gm_n161, gm_n1610, gm_n1611, gm_n1612, gm_n1613, gm_n1614, gm_n1615, gm_n1616, gm_n1617, gm_n1618, gm_n1619, gm_n162, gm_n1620, gm_n1621, gm_n1622, gm_n1623, gm_n1624, gm_n1625, gm_n1626, gm_n1627, gm_n1628, gm_n1629, gm_n163, gm_n1630, gm_n1631, gm_n1632, gm_n1633, gm_n1634, gm_n1635, gm_n1636, gm_n1637, gm_n1638, gm_n1639, gm_n164, gm_n1640, gm_n1641, gm_n1642, gm_n1643, gm_n1644, gm_n1645, gm_n1646, gm_n1647, gm_n1648, gm_n1649, gm_n165, gm_n1650, gm_n1651, gm_n1652, gm_n1653, gm_n1654, gm_n1655, gm_n1656, gm_n1657, gm_n1658, gm_n1659, gm_n166, gm_n1660, gm_n1661, gm_n1662, gm_n1663, gm_n1664, gm_n1665, gm_n1666, gm_n1667, gm_n1668, gm_n1669, gm_n167, gm_n1670, gm_n1671, gm_n1672, gm_n1673, gm_n1674, gm_n1675, gm_n1676, gm_n1677, gm_n1678, gm_n1679, gm_n168, gm_n1680, gm_n1681, gm_n1682, gm_n1683, gm_n1684, gm_n1685, gm_n1686, gm_n1687, gm_n1688, gm_n1689, gm_n169, gm_n1690, gm_n1691, gm_n1692, gm_n1693, gm_n1694, gm_n1695, gm_n1696, gm_n1697, gm_n1698, gm_n1699, gm_n170, gm_n1700, gm_n1701, gm_n1702, gm_n1703, gm_n1704, gm_n1705, gm_n1706, gm_n1707, gm_n1708, gm_n1709, gm_n171, gm_n1710, gm_n1711, gm_n1712, gm_n1713, gm_n1714, gm_n1715, gm_n1716, gm_n1717, gm_n1718, gm_n1719, gm_n172, gm_n1720, gm_n1721, gm_n1722, gm_n1723, gm_n1724, gm_n1725, gm_n1726, gm_n1727, gm_n1728, gm_n1729, gm_n173, gm_n1730, gm_n1731, gm_n1732, gm_n1733, gm_n1734, gm_n1735, gm_n1736, gm_n1737, gm_n1738, gm_n1739, gm_n174, gm_n1740, gm_n1741, gm_n1742, gm_n1743, gm_n1744, gm_n1745, gm_n1746, gm_n1747, gm_n1748, gm_n1749, gm_n175, gm_n1750, gm_n1751, gm_n1752, gm_n1753, gm_n1754, gm_n1755, gm_n1756, gm_n1757, gm_n1758, gm_n1759, gm_n176, gm_n1760, gm_n1761, gm_n1762, gm_n1763, gm_n1764, gm_n1765, gm_n1766, gm_n1767, gm_n1768, gm_n1769, gm_n177, gm_n1770, gm_n1771, gm_n1772, gm_n1773, gm_n1774, gm_n1775, gm_n1776, gm_n1777, gm_n1778, gm_n1779, gm_n178, gm_n1780, gm_n1781, gm_n1782, gm_n1783, gm_n1784, gm_n1785, gm_n1786, gm_n1787, gm_n1788, gm_n1789, gm_n179, gm_n1790, gm_n1791, gm_n1792, gm_n1793, gm_n1794, gm_n1795, gm_n1796, gm_n1797, gm_n1798, gm_n1799, gm_n180, gm_n1800, gm_n1801, gm_n1802, gm_n1803, gm_n1804, gm_n1805, gm_n1806, gm_n1807, gm_n1808, gm_n1809, gm_n181, gm_n1810, gm_n1811, gm_n1812, gm_n1813, gm_n1814, gm_n1815, gm_n1816, gm_n1817, gm_n1818, gm_n1819, gm_n182, gm_n1820, gm_n1821, gm_n1822, gm_n1823, gm_n1824, gm_n1825, gm_n1826, gm_n1827, gm_n1828, gm_n1829, gm_n183, gm_n1830, gm_n1831, gm_n1832, gm_n1833, gm_n1834, gm_n1835, gm_n1836, gm_n1837, gm_n1838, gm_n1839, gm_n184, gm_n1840, gm_n1841, gm_n1842, gm_n1843, gm_n1844, gm_n1845, gm_n1846, gm_n1847, gm_n1848, gm_n1849, gm_n185, gm_n1850, gm_n1851, gm_n1852, gm_n1853, gm_n1854, gm_n1855, gm_n1856, gm_n1857, gm_n1858, gm_n1859, gm_n186, gm_n1860, gm_n1861, gm_n1862, gm_n1863, gm_n1864, gm_n1865, gm_n1866, gm_n1867, gm_n1868, gm_n1869, gm_n187, gm_n1870, gm_n1871, gm_n1872, gm_n1873, gm_n1874, gm_n1875, gm_n1876, gm_n1877, gm_n1878, gm_n1879, gm_n188, gm_n1880, gm_n1881, gm_n1882, gm_n1883, gm_n1884, gm_n1885, gm_n1886, gm_n1887, gm_n1888, gm_n1889, gm_n189, gm_n1890, gm_n1891, gm_n1893, gm_n1894, gm_n1895, gm_n1896, gm_n1897, gm_n1898, gm_n1899, gm_n190, gm_n1900, gm_n1901, gm_n1902, gm_n1903, gm_n1904, gm_n1905, gm_n1906, gm_n1907, gm_n1908, gm_n1909, gm_n191, gm_n1910, gm_n1911, gm_n1912, gm_n1913, gm_n1914, gm_n1915, gm_n1916, gm_n1917, gm_n1918, gm_n1919, gm_n192, gm_n1920, gm_n1921, gm_n1922, gm_n1923, gm_n1924, gm_n1925, gm_n1926, gm_n1927, gm_n1928, gm_n1929, gm_n193, gm_n1930, gm_n1931, gm_n1932, gm_n1933, gm_n1934, gm_n1935, gm_n1936, gm_n1937, gm_n1938, gm_n1939, gm_n194, gm_n1940, gm_n1941, gm_n1942, gm_n1943, gm_n1944, gm_n1945, gm_n1946, gm_n1947, gm_n1948, gm_n1949, gm_n195, gm_n1950, gm_n1951, gm_n1952, gm_n1953, gm_n1954, gm_n1955, gm_n1956, gm_n1957, gm_n1958, gm_n1959, gm_n196, gm_n1960, gm_n1961, gm_n1962, gm_n1963, gm_n1964, gm_n1965, gm_n1966, gm_n1967, gm_n1968, gm_n1969, gm_n197, gm_n1970, gm_n1971, gm_n1972, gm_n1973, gm_n1974, gm_n1975, gm_n1976, gm_n1977, gm_n1978, gm_n1979, gm_n198, gm_n1980, gm_n1981, gm_n1982, gm_n1983, gm_n1984, gm_n1985, gm_n1986, gm_n1987, gm_n1988, gm_n1989, gm_n199, gm_n1990, gm_n1991, gm_n1992, gm_n1993, gm_n1994, gm_n1995, gm_n1996, gm_n1997, gm_n1998, gm_n1999, gm_n200, gm_n2000, gm_n2001, gm_n2002, gm_n2003, gm_n2004, gm_n2005, gm_n2006, gm_n2007, gm_n2008, gm_n2009, gm_n201, gm_n2010, gm_n2011, gm_n2012, gm_n2013, gm_n2014, gm_n2015, gm_n2016, gm_n2017, gm_n2018, gm_n2019, gm_n202, gm_n2020, gm_n2021, gm_n2022, gm_n2023, gm_n2024, gm_n2025, gm_n2026, gm_n2027, gm_n2028, gm_n2029, gm_n203, gm_n2030, gm_n2031, gm_n2032, gm_n2033, gm_n2034, gm_n2035, gm_n2036, gm_n2037, gm_n2038, gm_n2039, gm_n204, gm_n2040, gm_n2041, gm_n2042, gm_n2043, gm_n2044, gm_n2045, gm_n2046, gm_n2047, gm_n2048, gm_n2049, gm_n205, gm_n2050, gm_n2051, gm_n2052, gm_n2053, gm_n2054, gm_n2055, gm_n2056, gm_n2057, gm_n2058, gm_n2059, gm_n206, gm_n2060, gm_n2061, gm_n2062, gm_n2063, gm_n2064, gm_n2065, gm_n2066, gm_n2067, gm_n2068, gm_n2069, gm_n207, gm_n2070, gm_n2071, gm_n2072, gm_n2073, gm_n2074, gm_n2075, gm_n2076, gm_n2077, gm_n2078, gm_n2079, gm_n208, gm_n2080, gm_n2081, gm_n2082, gm_n2083, gm_n2084, gm_n2085, gm_n2086, gm_n2087, gm_n2088, gm_n2089, gm_n209, gm_n2090, gm_n2091, gm_n2092, gm_n2093, gm_n2094, gm_n2095, gm_n2096, gm_n2097, gm_n2098, gm_n2099, gm_n210, gm_n2100, gm_n2101, gm_n2102, gm_n2103, gm_n2104, gm_n2105, gm_n2106, gm_n2107, gm_n2108, gm_n2109, gm_n211, gm_n2110, gm_n2111, gm_n2112, gm_n2113, gm_n2114, gm_n2115, gm_n2116, gm_n2117, gm_n2118, gm_n2119, gm_n212, gm_n2120, gm_n2121, gm_n2122, gm_n2123, gm_n2124, gm_n2125, gm_n2126, gm_n2127, gm_n2128, gm_n2129, gm_n213, gm_n2130, gm_n2131, gm_n2132, gm_n2133, gm_n2134, gm_n2135, gm_n2136, gm_n2137, gm_n2138, gm_n2139, gm_n214, gm_n2140, gm_n2141, gm_n2142, gm_n2143, gm_n2144, gm_n2145, gm_n2146, gm_n2147, gm_n2148, gm_n2149, gm_n215, gm_n2150, gm_n2151, gm_n2152, gm_n2153, gm_n2154, gm_n2155, gm_n2156, gm_n2157, gm_n2158, gm_n2159, gm_n216, gm_n2160, gm_n2161, gm_n2162, gm_n2163, gm_n2164, gm_n2165, gm_n2166, gm_n2167, gm_n2168, gm_n2169, gm_n217, gm_n2170, gm_n2171, gm_n2172, gm_n2173, gm_n2174, gm_n2175, gm_n2176, gm_n2177, gm_n2178, gm_n2179, gm_n218, gm_n2180, gm_n2181, gm_n2182, gm_n2183, gm_n2184, gm_n2185, gm_n2186, gm_n2187, gm_n2188, gm_n2189, gm_n219, gm_n2190, gm_n2191, gm_n2192, gm_n2193, gm_n2194, gm_n2195, gm_n2196, gm_n2197, gm_n2198, gm_n2199, gm_n220, gm_n2200, gm_n2201, gm_n2202, gm_n2203, gm_n2204, gm_n2205, gm_n2206, gm_n2207, gm_n2208, gm_n2209, gm_n221, gm_n2210, gm_n2211, gm_n2212, gm_n2213, gm_n2214, gm_n2215, gm_n2216, gm_n2217, gm_n2218, gm_n2219, gm_n222, gm_n2220, gm_n2221, gm_n2222, gm_n2223, gm_n2224, gm_n2225, gm_n2226, gm_n2227, gm_n2228, gm_n2229, gm_n223, gm_n2230, gm_n2231, gm_n2232, gm_n2233, gm_n2234, gm_n2235, gm_n2236, gm_n2237, gm_n2238, gm_n2239, gm_n224, gm_n2240, gm_n2241, gm_n2242, gm_n2243, gm_n2244, gm_n2245, gm_n2246, gm_n2247, gm_n2248, gm_n2249, gm_n225, gm_n2250, gm_n2251, gm_n2252, gm_n2253, gm_n2254, gm_n2255, gm_n2256, gm_n2257, gm_n2258, gm_n2259, gm_n226, gm_n2260, gm_n2261, gm_n2262, gm_n2263, gm_n2264, gm_n2265, gm_n2266, gm_n2267, gm_n2268, gm_n2269, gm_n227, gm_n2270, gm_n2271, gm_n2272, gm_n2273, gm_n2274, gm_n2276, gm_n2277, gm_n2278, gm_n2279, gm_n228, gm_n2280, gm_n2281, gm_n2282, gm_n2283, gm_n2284, gm_n2285, gm_n2286, gm_n2287, gm_n2288, gm_n2289, gm_n229, gm_n2290, gm_n2291, gm_n2292, gm_n2293, gm_n2294, gm_n2295, gm_n2296, gm_n2297, gm_n2298, gm_n2299, gm_n230, gm_n2300, gm_n2301, gm_n2302, gm_n2303, gm_n2304, gm_n2305, gm_n2306, gm_n2307, gm_n2308, gm_n2309, gm_n231, gm_n2310, gm_n2311, gm_n2312, gm_n2313, gm_n2314, gm_n2315, gm_n2316, gm_n2317, gm_n2318, gm_n2319, gm_n232, gm_n2320, gm_n2321, gm_n2322, gm_n2323, gm_n2324, gm_n2325, gm_n2326, gm_n2327, gm_n2328, gm_n2329, gm_n233, gm_n2330, gm_n2331, gm_n2332, gm_n2333, gm_n2334, gm_n2335, gm_n2336, gm_n2337, gm_n2338, gm_n2339, gm_n234, gm_n2340, gm_n2341, gm_n2342, gm_n2343, gm_n2344, gm_n2345, gm_n2346, gm_n2347, gm_n2348, gm_n2349, gm_n235, gm_n2350, gm_n2351, gm_n2352, gm_n2353, gm_n2354, gm_n2355, gm_n2356, gm_n2357, gm_n2358, gm_n2359, gm_n236, gm_n2360, gm_n2361, gm_n2362, gm_n2363, gm_n2364, gm_n2365, gm_n2366, gm_n2367, gm_n2368, gm_n2369, gm_n237, gm_n2370, gm_n2371, gm_n2372, gm_n2373, gm_n2374, gm_n2375, gm_n2376, gm_n2377, gm_n2378, gm_n2379, gm_n238, gm_n2380, gm_n2381, gm_n2382, gm_n2383, gm_n2384, gm_n2385, gm_n2386, gm_n2387, gm_n2388, gm_n2389, gm_n239, gm_n2390, gm_n2391, gm_n2392, gm_n2393, gm_n2394, gm_n2395, gm_n2396, gm_n2397, gm_n2398, gm_n2399, gm_n240, gm_n2400, gm_n2401, gm_n2402, gm_n2403, gm_n2404, gm_n2405, gm_n2406, gm_n2407, gm_n2408, gm_n2409, gm_n241, gm_n2410, gm_n2411, gm_n2412, gm_n2413, gm_n2414, gm_n2415, gm_n2416, gm_n2417, gm_n2418, gm_n2419, gm_n242, gm_n2420, gm_n2421, gm_n2422, gm_n2423, gm_n2424, gm_n2425, gm_n2426, gm_n2427, gm_n2428, gm_n2429, gm_n243, gm_n2430, gm_n2431, gm_n2432, gm_n2433, gm_n2434, gm_n2435, gm_n2436, gm_n2437, gm_n2438, gm_n2439, gm_n244, gm_n2440, gm_n2441, gm_n2442, gm_n2443, gm_n2444, gm_n2445, gm_n2446, gm_n2447, gm_n2448, gm_n2449, gm_n245, gm_n2450, gm_n2451, gm_n2452, gm_n2453, gm_n2454, gm_n2455, gm_n2456, gm_n2457, gm_n2458, gm_n2459, gm_n246, gm_n2460, gm_n2461, gm_n2462, gm_n2463, gm_n2464, gm_n2465, gm_n2466, gm_n2467, gm_n2468, gm_n2469, gm_n247, gm_n2470, gm_n2471, gm_n2472, gm_n2473, gm_n2474, gm_n2475, gm_n2476, gm_n2477, gm_n2478, gm_n2479, gm_n248, gm_n2480, gm_n2481, gm_n2482, gm_n2483, gm_n2484, gm_n2485, gm_n2486, gm_n2487, gm_n2488, gm_n2489, gm_n249, gm_n2490, gm_n2491, gm_n2492, gm_n2493, gm_n2494, gm_n2495, gm_n2496, gm_n2497, gm_n2498, gm_n2499, gm_n250, gm_n2500, gm_n2501, gm_n2502, gm_n2503, gm_n2504, gm_n2505, gm_n2506, gm_n2507, gm_n2508, gm_n2509, gm_n251, gm_n2510, gm_n2511, gm_n2512, gm_n2513, gm_n2514, gm_n2515, gm_n2516, gm_n2517, gm_n2518, gm_n2519, gm_n252, gm_n2520, gm_n2521, gm_n2522, gm_n2523, gm_n2524, gm_n2525, gm_n2526, gm_n2527, gm_n2528, gm_n2529, gm_n253, gm_n2530, gm_n2531, gm_n2532, gm_n2533, gm_n2534, gm_n2535, gm_n2536, gm_n2537, gm_n2538, gm_n2539, gm_n254, gm_n2540, gm_n2541, gm_n2542, gm_n2543, gm_n2544, gm_n2545, gm_n2546, gm_n2547, gm_n2548, gm_n2549, gm_n255, gm_n2550, gm_n2551, gm_n2552, gm_n2553, gm_n2554, gm_n2555, gm_n2556, gm_n2557, gm_n2558, gm_n2559, gm_n256, gm_n2560, gm_n2561, gm_n2562, gm_n2563, gm_n2564, gm_n2565, gm_n2566, gm_n2567, gm_n2568, gm_n2569, gm_n257, gm_n2570, gm_n2571, gm_n2572, gm_n2573, gm_n2574, gm_n2575, gm_n2576, gm_n2577, gm_n2578, gm_n2579, gm_n258, gm_n2580, gm_n2581, gm_n2582, gm_n2583, gm_n2584, gm_n2585, gm_n2586, gm_n2587, gm_n2588, gm_n2589, gm_n259, gm_n2590, gm_n2591, gm_n2592, gm_n2593, gm_n2594, gm_n2595, gm_n2596, gm_n2597, gm_n2598, gm_n2599, gm_n260, gm_n2600, gm_n2601, gm_n2602, gm_n2603, gm_n2604, gm_n2605, gm_n2606, gm_n2607, gm_n2608, gm_n2609, gm_n261, gm_n2610, gm_n2611, gm_n2612, gm_n2613, gm_n2614, gm_n2615, gm_n2616, gm_n2617, gm_n2618, gm_n2619, gm_n262, gm_n2620, gm_n2621, gm_n2622, gm_n2623, gm_n2624, gm_n2625, gm_n2626, gm_n2627, gm_n2628, gm_n2629, gm_n263, gm_n2630, gm_n2631, gm_n2632, gm_n2633, gm_n2634, gm_n2635, gm_n2636, gm_n2637, gm_n2638, gm_n2639, gm_n264, gm_n2640, gm_n2641, gm_n2642, gm_n2643, gm_n2644, gm_n2646, gm_n2647, gm_n2648, gm_n2649, gm_n265, gm_n2650, gm_n2651, gm_n2652, gm_n2653, gm_n2654, gm_n2655, gm_n2656, gm_n2657, gm_n2658, gm_n2659, gm_n266, gm_n2660, gm_n2661, gm_n2662, gm_n2663, gm_n2664, gm_n2665, gm_n2666, gm_n2667, gm_n2668, gm_n2669, gm_n267, gm_n2670, gm_n2671, gm_n2672, gm_n2673, gm_n2674, gm_n2675, gm_n2676, gm_n2677, gm_n2678, gm_n2679, gm_n268, gm_n2680, gm_n2681, gm_n2682, gm_n2683, gm_n2684, gm_n2685, gm_n2686, gm_n2687, gm_n2688, gm_n2689, gm_n269, gm_n2690, gm_n2691, gm_n2692, gm_n2693, gm_n2694, gm_n2695, gm_n2696, gm_n2697, gm_n2698, gm_n2699, gm_n270, gm_n2700, gm_n2701, gm_n2702, gm_n2703, gm_n2704, gm_n2705, gm_n2706, gm_n2707, gm_n2708, gm_n2709, gm_n271, gm_n2710, gm_n2711, gm_n2712, gm_n2713, gm_n2714, gm_n2715, gm_n2716, gm_n2717, gm_n2718, gm_n2719, gm_n272, gm_n2720, gm_n2721, gm_n2722, gm_n2723, gm_n2724, gm_n2725, gm_n2726, gm_n2727, gm_n2728, gm_n2729, gm_n273, gm_n2730, gm_n2731, gm_n2732, gm_n2733, gm_n2734, gm_n2735, gm_n2736, gm_n2737, gm_n2738, gm_n2739, gm_n274, gm_n2740, gm_n2741, gm_n2742, gm_n2743, gm_n2744, gm_n2745, gm_n2746, gm_n2747, gm_n2748, gm_n2749, gm_n275, gm_n2750, gm_n2751, gm_n2752, gm_n2753, gm_n2754, gm_n2755, gm_n2756, gm_n2757, gm_n2758, gm_n2759, gm_n276, gm_n2760, gm_n2761, gm_n2762, gm_n2763, gm_n2764, gm_n2765, gm_n2766, gm_n2767, gm_n2768, gm_n2769, gm_n277, gm_n2770, gm_n2771, gm_n2772, gm_n2773, gm_n2774, gm_n2775, gm_n2776, gm_n2777, gm_n2778, gm_n2779, gm_n278, gm_n2780, gm_n2781, gm_n2782, gm_n2783, gm_n2784, gm_n2785, gm_n2786, gm_n2787, gm_n2788, gm_n2789, gm_n279, gm_n2790, gm_n2791, gm_n2792, gm_n2793, gm_n2794, gm_n2795, gm_n2796, gm_n2797, gm_n2798, gm_n2799, gm_n280, gm_n2800, gm_n2801, gm_n2802, gm_n2803, gm_n2804, gm_n2805, gm_n2806, gm_n2807, gm_n2808, gm_n2809, gm_n281, gm_n2810, gm_n2811, gm_n2812, gm_n2813, gm_n2814, gm_n2815, gm_n2816, gm_n2817, gm_n2818, gm_n2819, gm_n282, gm_n2820, gm_n2821, gm_n2822, gm_n2823, gm_n2824, gm_n2825, gm_n2826, gm_n2827, gm_n2828, gm_n2829, gm_n283, gm_n2830, gm_n2831, gm_n2832, gm_n2833, gm_n2834, gm_n2835, gm_n2836, gm_n2837, gm_n2838, gm_n2839, gm_n284, gm_n2840, gm_n2841, gm_n2842, gm_n2843, gm_n2844, gm_n2845, gm_n2846, gm_n2847, gm_n2848, gm_n2849, gm_n285, gm_n2850, gm_n2851, gm_n2852, gm_n2853, gm_n2854, gm_n2855, gm_n2856, gm_n2857, gm_n2858, gm_n2859, gm_n286, gm_n2860, gm_n2861, gm_n2862, gm_n2863, gm_n2864, gm_n2865, gm_n2866, gm_n2867, gm_n2868, gm_n2869, gm_n287, gm_n2870, gm_n2871, gm_n2872, gm_n2873, gm_n2874, gm_n2875, gm_n2876, gm_n2877, gm_n2878, gm_n2879, gm_n288, gm_n2880, gm_n2881, gm_n2882, gm_n2883, gm_n2884, gm_n2885, gm_n2886, gm_n2887, gm_n2888, gm_n2889, gm_n289, gm_n2890, gm_n2891, gm_n2892, gm_n2893, gm_n2894, gm_n2895, gm_n2896, gm_n2897, gm_n2898, gm_n2899, gm_n290, gm_n2900, gm_n2901, gm_n2902, gm_n2903, gm_n2904, gm_n2905, gm_n2906, gm_n2907, gm_n2908, gm_n2909, gm_n291, gm_n2910, gm_n2911, gm_n2912, gm_n2913, gm_n2914, gm_n2915, gm_n2916, gm_n2917, gm_n2918, gm_n2919, gm_n292, gm_n2920, gm_n2921, gm_n2922, gm_n2923, gm_n2924, gm_n2925, gm_n2926, gm_n2927, gm_n2928, gm_n2929, gm_n293, gm_n2930, gm_n2931, gm_n2932, gm_n2933, gm_n2934, gm_n2935, gm_n2936, gm_n2937, gm_n2938, gm_n2939, gm_n294, gm_n2940, gm_n2941, gm_n2942, gm_n2943, gm_n2944, gm_n2945, gm_n2946, gm_n2947, gm_n2948, gm_n2949, gm_n295, gm_n2950, gm_n2951, gm_n2952, gm_n2953, gm_n2954, gm_n2955, gm_n2956, gm_n2957, gm_n2958, gm_n2959, gm_n296, gm_n2960, gm_n2961, gm_n2962, gm_n2963, gm_n2964, gm_n2965, gm_n2966, gm_n2967, gm_n2968, gm_n2969, gm_n297, gm_n2970, gm_n2971, gm_n2972, gm_n2973, gm_n2974, gm_n2975, gm_n2976, gm_n2977, gm_n2978, gm_n2979, gm_n298, gm_n2980, gm_n2981, gm_n2982, gm_n2983, gm_n2984, gm_n2985, gm_n2986, gm_n2987, gm_n2988, gm_n2989, gm_n299, gm_n2990, gm_n2991, gm_n2992, gm_n2993, gm_n2994, gm_n2995, gm_n2996, gm_n2997, gm_n2998, gm_n2999, gm_n300, gm_n3000, gm_n3001, gm_n3002, gm_n3003, gm_n3004, gm_n3005, gm_n3006, gm_n3007, gm_n3008, gm_n3009, gm_n301, gm_n3010, gm_n3011, gm_n3012, gm_n3013, gm_n3014, gm_n3015, gm_n3016, gm_n3017, gm_n3018, gm_n302, gm_n3020, gm_n3021, gm_n3022, gm_n3023, gm_n3024, gm_n3025, gm_n3026, gm_n3027, gm_n3028, gm_n3029, gm_n303, gm_n3030, gm_n3031, gm_n3032, gm_n3033, gm_n3034, gm_n3035, gm_n3036, gm_n3037, gm_n3038, gm_n3039, gm_n304, gm_n3040, gm_n3041, gm_n3042, gm_n3043, gm_n3044, gm_n3045, gm_n3046, gm_n3047, gm_n3048, gm_n3049, gm_n305, gm_n3050, gm_n3051, gm_n3052, gm_n3053, gm_n3054, gm_n3055, gm_n3056, gm_n3057, gm_n3058, gm_n3059, gm_n306, gm_n3060, gm_n3061, gm_n3062, gm_n3063, gm_n3064, gm_n3065, gm_n3066, gm_n3067, gm_n3068, gm_n3069, gm_n307, gm_n3070, gm_n3071, gm_n3072, gm_n3073, gm_n3074, gm_n3075, gm_n3076, gm_n3077, gm_n3078, gm_n3079, gm_n308, gm_n3080, gm_n3081, gm_n3082, gm_n3083, gm_n3084, gm_n3085, gm_n3086, gm_n3087, gm_n3088, gm_n3089, gm_n309, gm_n3090, gm_n3091, gm_n3092, gm_n3093, gm_n3094, gm_n3095, gm_n3096, gm_n3097, gm_n3098, gm_n3099, gm_n310, gm_n3100, gm_n3101, gm_n3102, gm_n3103, gm_n3104, gm_n3105, gm_n3106, gm_n3107, gm_n3108, gm_n3109, gm_n311, gm_n3110, gm_n3111, gm_n3112, gm_n3113, gm_n3114, gm_n3115, gm_n3116, gm_n3117, gm_n3118, gm_n3119, gm_n312, gm_n3120, gm_n3121, gm_n3122, gm_n3123, gm_n3124, gm_n3125, gm_n3126, gm_n3127, gm_n3128, gm_n3129, gm_n313, gm_n3130, gm_n3131, gm_n3132, gm_n3133, gm_n3134, gm_n3135, gm_n3136, gm_n3137, gm_n3138, gm_n3139, gm_n314, gm_n3140, gm_n3141, gm_n3142, gm_n3143, gm_n3144, gm_n3145, gm_n3146, gm_n3147, gm_n3148, gm_n3149, gm_n315, gm_n3150, gm_n3151, gm_n3152, gm_n3153, gm_n3154, gm_n3155, gm_n3156, gm_n3157, gm_n3158, gm_n3159, gm_n316, gm_n3160, gm_n3161, gm_n3162, gm_n3163, gm_n3164, gm_n3165, gm_n3166, gm_n3167, gm_n3168, gm_n3169, gm_n317, gm_n3170, gm_n3171, gm_n3172, gm_n3173, gm_n3174, gm_n3175, gm_n3176, gm_n3177, gm_n3178, gm_n3179, gm_n318, gm_n3180, gm_n3181, gm_n3182, gm_n3183, gm_n3184, gm_n3185, gm_n3186, gm_n3187, gm_n3188, gm_n3189, gm_n319, gm_n3190, gm_n3191, gm_n3192, gm_n3193, gm_n3194, gm_n3195, gm_n3196, gm_n3197, gm_n3198, gm_n3199, gm_n320, gm_n3200, gm_n3201, gm_n3202, gm_n3203, gm_n3204, gm_n3205, gm_n3206, gm_n3207, gm_n3208, gm_n3209, gm_n321, gm_n3210, gm_n3211, gm_n3212, gm_n3213, gm_n3214, gm_n3215, gm_n3216, gm_n3217, gm_n3218, gm_n3219, gm_n322, gm_n3220, gm_n3221, gm_n3222, gm_n3223, gm_n3224, gm_n3225, gm_n3226, gm_n3227, gm_n3228, gm_n3229, gm_n323, gm_n3230, gm_n3231, gm_n3232, gm_n3233, gm_n3234, gm_n3235, gm_n3236, gm_n3237, gm_n3238, gm_n3239, gm_n324, gm_n3240, gm_n3241, gm_n3242, gm_n3243, gm_n3244, gm_n3245, gm_n3246, gm_n3247, gm_n3248, gm_n3249, gm_n325, gm_n3250, gm_n3251, gm_n3252, gm_n3253, gm_n3254, gm_n3255, gm_n3256, gm_n3257, gm_n3258, gm_n3259, gm_n326, gm_n3260, gm_n3261, gm_n3262, gm_n3263, gm_n3264, gm_n3265, gm_n3266, gm_n3267, gm_n3268, gm_n3269, gm_n327, gm_n3270, gm_n3271, gm_n3272, gm_n3273, gm_n3274, gm_n3275, gm_n3276, gm_n3277, gm_n3278, gm_n3279, gm_n328, gm_n3280, gm_n3281, gm_n3282, gm_n3283, gm_n3284, gm_n3285, gm_n3286, gm_n3287, gm_n3288, gm_n3289, gm_n329, gm_n3290, gm_n3291, gm_n3292, gm_n3293, gm_n3294, gm_n3295, gm_n3296, gm_n3297, gm_n3298, gm_n3299, gm_n330, gm_n3300, gm_n3301, gm_n3302, gm_n3303, gm_n3304, gm_n3305, gm_n3306, gm_n3307, gm_n3308, gm_n3309, gm_n331, gm_n3310, gm_n3311, gm_n3312, gm_n3313, gm_n3314, gm_n3315, gm_n3316, gm_n3317, gm_n3318, gm_n3319, gm_n332, gm_n3320, gm_n3321, gm_n3322, gm_n3323, gm_n3324, gm_n3325, gm_n3326, gm_n3327, gm_n3328, gm_n3329, gm_n333, gm_n3330, gm_n3331, gm_n3332, gm_n3333, gm_n3334, gm_n3335, gm_n3336, gm_n3337, gm_n3338, gm_n3339, gm_n334, gm_n3340, gm_n3341, gm_n3342, gm_n3343, gm_n3344, gm_n3345, gm_n3346, gm_n3347, gm_n3348, gm_n3349, gm_n335, gm_n3350, gm_n3351, gm_n3352, gm_n3353, gm_n3354, gm_n3355, gm_n3356, gm_n3357, gm_n3358, gm_n3359, gm_n336, gm_n3360, gm_n3361, gm_n3362, gm_n3363, gm_n3364, gm_n3365, gm_n3366, gm_n3367, gm_n3368, gm_n3369, gm_n337, gm_n3370, gm_n3372, gm_n3373, gm_n3374, gm_n3375, gm_n3376, gm_n3377, gm_n3378, gm_n3379, gm_n338, gm_n3380, gm_n3381, gm_n3382, gm_n3383, gm_n3384, gm_n3385, gm_n3386, gm_n3387, gm_n3388, gm_n3389, gm_n339, gm_n3390, gm_n3391, gm_n3392, gm_n3393, gm_n3394, gm_n3395, gm_n3396, gm_n3397, gm_n3398, gm_n3399, gm_n340, gm_n3400, gm_n3401, gm_n3402, gm_n3403, gm_n3404, gm_n3405, gm_n3406, gm_n3407, gm_n3408, gm_n3409, gm_n341, gm_n3410, gm_n3411, gm_n3412, gm_n3413, gm_n3414, gm_n3415, gm_n3416, gm_n3417, gm_n3418, gm_n3419, gm_n342, gm_n3420, gm_n3421, gm_n3422, gm_n3423, gm_n3424, gm_n3425, gm_n3426, gm_n3427, gm_n3428, gm_n3429, gm_n343, gm_n3430, gm_n3431, gm_n3432, gm_n3433, gm_n3434, gm_n3435, gm_n3436, gm_n3437, gm_n3438, gm_n3439, gm_n344, gm_n3440, gm_n3441, gm_n3442, gm_n3443, gm_n3444, gm_n3445, gm_n3446, gm_n3447, gm_n3448, gm_n3449, gm_n345, gm_n3450, gm_n3451, gm_n3452, gm_n3453, gm_n3454, gm_n3455, gm_n3456, gm_n3457, gm_n3458, gm_n3459, gm_n346, gm_n3460, gm_n3461, gm_n3462, gm_n3463, gm_n3464, gm_n3465, gm_n3466, gm_n3467, gm_n3468, gm_n3469, gm_n347, gm_n3470, gm_n3471, gm_n3472, gm_n3473, gm_n3474, gm_n3475, gm_n3476, gm_n3477, gm_n3478, gm_n3479, gm_n348, gm_n3480, gm_n3481, gm_n3482, gm_n3483, gm_n3484, gm_n3485, gm_n3486, gm_n3487, gm_n3488, gm_n3489, gm_n349, gm_n3490, gm_n3491, gm_n3492, gm_n3493, gm_n3494, gm_n3495, gm_n3496, gm_n3497, gm_n3498, gm_n3499, gm_n350, gm_n3500, gm_n3501, gm_n3502, gm_n3503, gm_n3504, gm_n3505, gm_n3506, gm_n3507, gm_n3508, gm_n3509, gm_n351, gm_n3510, gm_n3511, gm_n3512, gm_n3513, gm_n3514, gm_n3515, gm_n3516, gm_n3517, gm_n3518, gm_n3519, gm_n352, gm_n3520, gm_n3521, gm_n3522, gm_n3523, gm_n3524, gm_n3525, gm_n3526, gm_n3527, gm_n3528, gm_n3529, gm_n353, gm_n3530, gm_n3531, gm_n3532, gm_n3533, gm_n3534, gm_n3535, gm_n3536, gm_n3537, gm_n3538, gm_n3539, gm_n354, gm_n3540, gm_n3541, gm_n3542, gm_n3543, gm_n3544, gm_n3545, gm_n3546, gm_n3547, gm_n3548, gm_n3549, gm_n355, gm_n3550, gm_n3551, gm_n3552, gm_n3553, gm_n3554, gm_n3555, gm_n3556, gm_n3557, gm_n3558, gm_n3559, gm_n356, gm_n3560, gm_n3561, gm_n3562, gm_n3563, gm_n3564, gm_n3565, gm_n3566, gm_n3567, gm_n3568, gm_n3569, gm_n357, gm_n3570, gm_n3571, gm_n3572, gm_n3573, gm_n3574, gm_n3575, gm_n3576, gm_n3577, gm_n3578, gm_n3579, gm_n358, gm_n3580, gm_n3581, gm_n3582, gm_n3583, gm_n3584, gm_n3585, gm_n3586, gm_n3587, gm_n3588, gm_n3589, gm_n359, gm_n3590, gm_n3591, gm_n3592, gm_n3593, gm_n3594, gm_n3595, gm_n3596, gm_n3597, gm_n3598, gm_n3599, gm_n360, gm_n3600, gm_n3601, gm_n3602, gm_n3603, gm_n3604, gm_n3605, gm_n3606, gm_n3607, gm_n3608, gm_n3609, gm_n361, gm_n3610, gm_n3611, gm_n3612, gm_n3613, gm_n3614, gm_n3615, gm_n3616, gm_n3617, gm_n3618, gm_n3619, gm_n362, gm_n3620, gm_n3621, gm_n3622, gm_n3623, gm_n3624, gm_n3625, gm_n3626, gm_n3627, gm_n3628, gm_n3629, gm_n363, gm_n3630, gm_n3631, gm_n3632, gm_n3633, gm_n3634, gm_n3635, gm_n3636, gm_n3637, gm_n3638, gm_n3639, gm_n364, gm_n3640, gm_n3641, gm_n3642, gm_n3643, gm_n3644, gm_n3645, gm_n3646, gm_n3647, gm_n3648, gm_n3649, gm_n365, gm_n3650, gm_n3651, gm_n3652, gm_n3653, gm_n3654, gm_n3655, gm_n3656, gm_n3657, gm_n3658, gm_n3659, gm_n366, gm_n3660, gm_n3661, gm_n3662, gm_n3663, gm_n3664, gm_n3665, gm_n3666, gm_n3667, gm_n3668, gm_n3669, gm_n367, gm_n3670, gm_n3671, gm_n3672, gm_n3673, gm_n3674, gm_n3675, gm_n3676, gm_n3677, gm_n3678, gm_n3679, gm_n368, gm_n3680, gm_n3681, gm_n3682, gm_n3683, gm_n3684, gm_n3685, gm_n3686, gm_n3687, gm_n3688, gm_n3689, gm_n369, gm_n3690, gm_n3691, gm_n3692, gm_n3693, gm_n3694, gm_n3695, gm_n3696, gm_n3697, gm_n3698, gm_n3699, gm_n370, gm_n3700, gm_n3701, gm_n3702, gm_n3703, gm_n3704, gm_n3705, gm_n3706, gm_n3707, gm_n3708, gm_n3709, gm_n371, gm_n3710, gm_n3711, gm_n3712, gm_n3713, gm_n3714, gm_n3715, gm_n3716, gm_n3717, gm_n3718, gm_n3719, gm_n372, gm_n3720, gm_n3721, gm_n3722, gm_n3723, gm_n3724, gm_n3726, gm_n3727, gm_n3728, gm_n3729, gm_n373, gm_n3730, gm_n3731, gm_n3732, gm_n3733, gm_n3734, gm_n3735, gm_n3736, gm_n3737, gm_n3738, gm_n3739, gm_n374, gm_n3740, gm_n3741, gm_n3742, gm_n3743, gm_n3744, gm_n3745, gm_n3746, gm_n3747, gm_n3748, gm_n3749, gm_n375, gm_n3750, gm_n3751, gm_n3752, gm_n3753, gm_n3754, gm_n3755, gm_n3756, gm_n3757, gm_n3758, gm_n3759, gm_n376, gm_n3760, gm_n3761, gm_n3762, gm_n3763, gm_n3764, gm_n3765, gm_n3766, gm_n3767, gm_n3768, gm_n3769, gm_n377, gm_n3770, gm_n3771, gm_n3772, gm_n3773, gm_n3774, gm_n3775, gm_n3776, gm_n3777, gm_n3778, gm_n3779, gm_n378, gm_n3780, gm_n3781, gm_n3782, gm_n3783, gm_n3784, gm_n3785, gm_n3786, gm_n3787, gm_n3788, gm_n3789, gm_n379, gm_n3790, gm_n3791, gm_n3792, gm_n3793, gm_n3794, gm_n3795, gm_n3796, gm_n3797, gm_n3798, gm_n3799, gm_n380, gm_n3800, gm_n3801, gm_n3802, gm_n3803, gm_n3804, gm_n3805, gm_n3806, gm_n3807, gm_n3808, gm_n3809, gm_n381, gm_n3810, gm_n3811, gm_n3812, gm_n3813, gm_n3814, gm_n3815, gm_n3816, gm_n3817, gm_n3818, gm_n3819, gm_n382, gm_n3820, gm_n3821, gm_n3822, gm_n3823, gm_n3824, gm_n3825, gm_n3826, gm_n3827, gm_n3828, gm_n3829, gm_n383, gm_n3830, gm_n3831, gm_n3832, gm_n3833, gm_n3834, gm_n3835, gm_n3836, gm_n3837, gm_n3838, gm_n3839, gm_n384, gm_n3840, gm_n3841, gm_n3842, gm_n3843, gm_n3844, gm_n3845, gm_n3846, gm_n3847, gm_n3848, gm_n385, gm_n3850, gm_n3851, gm_n3852, gm_n3853, gm_n3854, gm_n3855, gm_n3856, gm_n3857, gm_n3858, gm_n3859, gm_n386, gm_n3860, gm_n3861, gm_n3862, gm_n3863, gm_n3864, gm_n3865, gm_n3866, gm_n3867, gm_n3868, gm_n3869, gm_n387, gm_n3870, gm_n3871, gm_n3872, gm_n3873, gm_n3874, gm_n3875, gm_n3876, gm_n3877, gm_n3878, gm_n3879, gm_n388, gm_n3880, gm_n3881, gm_n3882, gm_n3883, gm_n3884, gm_n3885, gm_n3886, gm_n3887, gm_n3888, gm_n3889, gm_n389, gm_n3890, gm_n3891, gm_n3892, gm_n3893, gm_n3894, gm_n3895, gm_n3896, gm_n3897, gm_n3898, gm_n3899, gm_n390, gm_n3900, gm_n3901, gm_n3902, gm_n3903, gm_n3904, gm_n3905, gm_n3906, gm_n3907, gm_n3908, gm_n3909, gm_n391, gm_n3910, gm_n3911, gm_n3912, gm_n3913, gm_n3914, gm_n3915, gm_n3916, gm_n3917, gm_n3918, gm_n3919, gm_n392, gm_n3920, gm_n3921, gm_n3922, gm_n3923, gm_n3924, gm_n3925, gm_n3926, gm_n3927, gm_n3928, gm_n3929, gm_n393, gm_n3930, gm_n3931, gm_n3932, gm_n3933, gm_n3934, gm_n3935, gm_n3936, gm_n3937, gm_n3938, gm_n3939, gm_n394, gm_n3940, gm_n3941, gm_n3942, gm_n3943, gm_n3944, gm_n3945, gm_n3946, gm_n3947, gm_n3948, gm_n3949, gm_n395, gm_n3950, gm_n3951, gm_n3952, gm_n3953, gm_n3954, gm_n3955, gm_n3956, gm_n3957, gm_n3958, gm_n3959, gm_n396, gm_n3960, gm_n3961, gm_n3962, gm_n3963, gm_n3964, gm_n3965, gm_n3966, gm_n3967, gm_n3968, gm_n3969, gm_n397, gm_n3970, gm_n3971, gm_n3972, gm_n3973, gm_n3974, gm_n3975, gm_n3976, gm_n3977, gm_n3978, gm_n3979, gm_n398, gm_n3980, gm_n3981, gm_n3982, gm_n3983, gm_n3984, gm_n3985, gm_n3986, gm_n3987, gm_n3988, gm_n3989, gm_n399, gm_n3990, gm_n3991, gm_n3992, gm_n3993, gm_n3994, gm_n3995, gm_n3996, gm_n3997, gm_n3998, gm_n3999, gm_n400, gm_n4000, gm_n4001, gm_n4002, gm_n4003, gm_n4004, gm_n4005, gm_n4006, gm_n4007, gm_n4008, gm_n4009, gm_n401, gm_n4010, gm_n4011, gm_n4012, gm_n4013, gm_n4014, gm_n4015, gm_n4016, gm_n4017, gm_n4018, gm_n4019, gm_n402, gm_n4020, gm_n4021, gm_n4022, gm_n4023, gm_n4024, gm_n4025, gm_n4026, gm_n4027, gm_n4028, gm_n4029, gm_n403, gm_n4030, gm_n4031, gm_n4032, gm_n4033, gm_n4034, gm_n4035, gm_n4036, gm_n4037, gm_n4038, gm_n4039, gm_n404, gm_n4040, gm_n4041, gm_n4042, gm_n4043, gm_n4044, gm_n4045, gm_n4046, gm_n4047, gm_n4048, gm_n4049, gm_n405, gm_n4050, gm_n4051, gm_n4052, gm_n4053, gm_n4054, gm_n4055, gm_n4056, gm_n4057, gm_n4058, gm_n4059, gm_n406, gm_n4060, gm_n4061, gm_n4062, gm_n4063, gm_n4064, gm_n4065, gm_n4066, gm_n4067, gm_n4068, gm_n4069, gm_n407, gm_n4070, gm_n4071, gm_n4072, gm_n4073, gm_n4074, gm_n4075, gm_n4076, gm_n4077, gm_n4078, gm_n4079, gm_n408, gm_n4080, gm_n4081, gm_n4082, gm_n4083, gm_n4084, gm_n4085, gm_n4086, gm_n4087, gm_n4088, gm_n4089, gm_n409, gm_n4090, gm_n4091, gm_n4092, gm_n4093, gm_n4094, gm_n4095, gm_n4096, gm_n4097, gm_n4098, gm_n4099, gm_n410, gm_n4100, gm_n4101, gm_n4102, gm_n4103, gm_n4104, gm_n4105, gm_n4106, gm_n4107, gm_n4108, gm_n4109, gm_n411, gm_n4110, gm_n4111, gm_n4112, gm_n4113, gm_n4114, gm_n4115, gm_n4116, gm_n4117, gm_n4118, gm_n4119, gm_n412, gm_n4120, gm_n4121, gm_n4122, gm_n4123, gm_n4124, gm_n4125, gm_n4126, gm_n4127, gm_n4128, gm_n4129, gm_n413, gm_n4130, gm_n4131, gm_n4132, gm_n4133, gm_n4134, gm_n4135, gm_n4136, gm_n4137, gm_n4138, gm_n4139, gm_n414, gm_n4140, gm_n4141, gm_n4142, gm_n4143, gm_n4144, gm_n4145, gm_n4146, gm_n4147, gm_n4148, gm_n4149, gm_n415, gm_n4150, gm_n4151, gm_n4152, gm_n4153, gm_n4154, gm_n4155, gm_n4156, gm_n4157, gm_n4158, gm_n4159, gm_n416, gm_n4160, gm_n4161, gm_n4162, gm_n4163, gm_n4164, gm_n4165, gm_n4166, gm_n4167, gm_n4168, gm_n4169, gm_n417, gm_n4170, gm_n4171, gm_n4172, gm_n4173, gm_n4174, gm_n4175, gm_n4176, gm_n4177, gm_n4178, gm_n4179, gm_n418, gm_n4180, gm_n4181, gm_n4182, gm_n4183, gm_n4184, gm_n4185, gm_n4186, gm_n4187, gm_n4188, gm_n4189, gm_n419, gm_n4190, gm_n4191, gm_n4192, gm_n4193, gm_n4194, gm_n4195, gm_n4196, gm_n4197, gm_n4198, gm_n4199, gm_n420, gm_n4200, gm_n4201, gm_n4203, gm_n4204, gm_n4205, gm_n4206, gm_n4207, gm_n4208, gm_n4209, gm_n421, gm_n4210, gm_n4211, gm_n4212, gm_n4213, gm_n4214, gm_n4215, gm_n4216, gm_n4217, gm_n4218, gm_n4219, gm_n422, gm_n4220, gm_n4221, gm_n4222, gm_n4223, gm_n4224, gm_n4225, gm_n4226, gm_n4227, gm_n4228, gm_n4229, gm_n423, gm_n4230, gm_n4231, gm_n4232, gm_n4233, gm_n4234, gm_n4235, gm_n4236, gm_n4237, gm_n4238, gm_n4239, gm_n424, gm_n4240, gm_n4241, gm_n4242, gm_n4243, gm_n4244, gm_n4245, gm_n4246, gm_n4247, gm_n4248, gm_n4249, gm_n425, gm_n4250, gm_n4251, gm_n4252, gm_n4253, gm_n4254, gm_n4255, gm_n4256, gm_n4257, gm_n4258, gm_n4259, gm_n426, gm_n4260, gm_n4261, gm_n4262, gm_n4263, gm_n4264, gm_n4265, gm_n4266, gm_n4267, gm_n4268, gm_n4269, gm_n427, gm_n4270, gm_n4271, gm_n4272, gm_n4273, gm_n4274, gm_n4275, gm_n4276, gm_n4277, gm_n4278, gm_n4279, gm_n428, gm_n4280, gm_n4281, gm_n4282, gm_n4283, gm_n4284, gm_n4285, gm_n4286, gm_n4287, gm_n4288, gm_n4289, gm_n429, gm_n4290, gm_n4291, gm_n4292, gm_n4293, gm_n4294, gm_n4295, gm_n4296, gm_n4297, gm_n4298, gm_n4299, gm_n430, gm_n4300, gm_n4301, gm_n4302, gm_n4303, gm_n4304, gm_n4305, gm_n4306, gm_n4307, gm_n4308, gm_n4309, gm_n431, gm_n4310, gm_n4311, gm_n4312, gm_n4313, gm_n4314, gm_n4315, gm_n4316, gm_n4317, gm_n4318, gm_n4319, gm_n432, gm_n4320, gm_n4321, gm_n4322, gm_n4323, gm_n4324, gm_n4325, gm_n4326, gm_n4327, gm_n4328, gm_n4329, gm_n433, gm_n4330, gm_n4331, gm_n4332, gm_n4333, gm_n4334, gm_n4335, gm_n4336, gm_n4337, gm_n4338, gm_n4339, gm_n434, gm_n4340, gm_n4341, gm_n4342, gm_n4343, gm_n4344, gm_n4345, gm_n4346, gm_n4347, gm_n4348, gm_n4349, gm_n435, gm_n4350, gm_n4351, gm_n4352, gm_n4353, gm_n4354, gm_n4355, gm_n4356, gm_n4357, gm_n4358, gm_n4359, gm_n436, gm_n4360, gm_n4361, gm_n4362, gm_n4363, gm_n4364, gm_n4365, gm_n4366, gm_n4367, gm_n4368, gm_n4369, gm_n437, gm_n4370, gm_n4371, gm_n4372, gm_n4373, gm_n4374, gm_n4375, gm_n4376, gm_n4377, gm_n4378, gm_n4379, gm_n438, gm_n4380, gm_n4381, gm_n4382, gm_n4383, gm_n4384, gm_n4385, gm_n4386, gm_n4387, gm_n4388, gm_n4389, gm_n439, gm_n4390, gm_n4391, gm_n4392, gm_n4393, gm_n4394, gm_n4395, gm_n4396, gm_n4397, gm_n4398, gm_n4399, gm_n440, gm_n4400, gm_n4401, gm_n4402, gm_n4403, gm_n4404, gm_n4405, gm_n4406, gm_n4407, gm_n4408, gm_n4409, gm_n441, gm_n4410, gm_n4411, gm_n4412, gm_n4413, gm_n4414, gm_n4415, gm_n4416, gm_n4417, gm_n4418, gm_n4419, gm_n442, gm_n4420, gm_n4421, gm_n4422, gm_n4423, gm_n4424, gm_n4425, gm_n4426, gm_n4427, gm_n4428, gm_n4429, gm_n443, gm_n4430, gm_n4431, gm_n4432, gm_n4433, gm_n4434, gm_n4435, gm_n4436, gm_n4437, gm_n4438, gm_n4439, gm_n444, gm_n4440, gm_n4441, gm_n4442, gm_n4443, gm_n4444, gm_n4445, gm_n4446, gm_n4447, gm_n4448, gm_n4449, gm_n445, gm_n4450, gm_n4451, gm_n4452, gm_n4453, gm_n4454, gm_n4455, gm_n4456, gm_n4457, gm_n4458, gm_n4459, gm_n446, gm_n4460, gm_n4461, gm_n4462, gm_n4463, gm_n4464, gm_n4465, gm_n4466, gm_n4467, gm_n4468, gm_n4469, gm_n447, gm_n4470, gm_n4471, gm_n4472, gm_n4473, gm_n4474, gm_n4475, gm_n4476, gm_n4477, gm_n4478, gm_n4479, gm_n448, gm_n4480, gm_n4481, gm_n4482, gm_n4483, gm_n4484, gm_n4485, gm_n4486, gm_n4487, gm_n4488, gm_n4489, gm_n449, gm_n4490, gm_n4491, gm_n4492, gm_n4493, gm_n4494, gm_n4495, gm_n4496, gm_n4497, gm_n4498, gm_n4499, gm_n450, gm_n4500, gm_n4501, gm_n4502, gm_n4503, gm_n4504, gm_n4505, gm_n4506, gm_n4507, gm_n4508, gm_n4509, gm_n451, gm_n4510, gm_n4511, gm_n4512, gm_n4513, gm_n4514, gm_n4515, gm_n4516, gm_n4517, gm_n4518, gm_n4519, gm_n452, gm_n4520, gm_n4521, gm_n4522, gm_n4523, gm_n4524, gm_n4525, gm_n4526, gm_n4527, gm_n4528, gm_n4529, gm_n453, gm_n4530, gm_n4531, gm_n4532, gm_n4533, gm_n4534, gm_n4535, gm_n4536, gm_n4537, gm_n4538, gm_n4539, gm_n454, gm_n4540, gm_n4541, gm_n4542, gm_n4543, gm_n4544, gm_n4545, gm_n4546, gm_n4547, gm_n4548, gm_n455, gm_n4550, gm_n4551, gm_n4552, gm_n4553, gm_n4554, gm_n4555, gm_n4556, gm_n4557, gm_n4558, gm_n4559, gm_n456, gm_n4560, gm_n4561, gm_n4562, gm_n4563, gm_n4564, gm_n4565, gm_n4566, gm_n4567, gm_n4568, gm_n4569, gm_n457, gm_n4570, gm_n4571, gm_n4572, gm_n4573, gm_n4574, gm_n4575, gm_n4576, gm_n4577, gm_n4578, gm_n4579, gm_n458, gm_n4580, gm_n4581, gm_n4582, gm_n4583, gm_n4584, gm_n4585, gm_n4586, gm_n4587, gm_n4588, gm_n4589, gm_n459, gm_n4590, gm_n4591, gm_n4592, gm_n4593, gm_n4594, gm_n4595, gm_n4596, gm_n4597, gm_n4598, gm_n4599, gm_n460, gm_n4600, gm_n4601, gm_n4602, gm_n4603, gm_n4604, gm_n4605, gm_n4606, gm_n4607, gm_n4608, gm_n4609, gm_n461, gm_n4610, gm_n4611, gm_n4612, gm_n4613, gm_n4614, gm_n4615, gm_n4616, gm_n4617, gm_n4618, gm_n4619, gm_n462, gm_n4620, gm_n4621, gm_n4622, gm_n4623, gm_n4624, gm_n4625, gm_n4626, gm_n4627, gm_n4628, gm_n4629, gm_n463, gm_n4630, gm_n4631, gm_n4632, gm_n4633, gm_n4634, gm_n4635, gm_n4636, gm_n4637, gm_n4638, gm_n4639, gm_n464, gm_n4640, gm_n4641, gm_n4642, gm_n4643, gm_n4644, gm_n4645, gm_n4646, gm_n4647, gm_n4648, gm_n4649, gm_n465, gm_n4650, gm_n4651, gm_n4652, gm_n4653, gm_n4654, gm_n4655, gm_n4656, gm_n4657, gm_n4658, gm_n4659, gm_n466, gm_n4660, gm_n4661, gm_n4662, gm_n4663, gm_n4664, gm_n4665, gm_n4666, gm_n4667, gm_n4668, gm_n4669, gm_n467, gm_n4670, gm_n4671, gm_n4672, gm_n4673, gm_n4674, gm_n4675, gm_n4676, gm_n4677, gm_n4678, gm_n4679, gm_n468, gm_n4680, gm_n4681, gm_n4682, gm_n4683, gm_n4684, gm_n4685, gm_n4686, gm_n4687, gm_n4688, gm_n4689, gm_n469, gm_n4690, gm_n4691, gm_n4692, gm_n4693, gm_n4694, gm_n4695, gm_n4696, gm_n4697, gm_n4698, gm_n4699, gm_n470, gm_n4700, gm_n4701, gm_n4702, gm_n4703, gm_n4704, gm_n4705, gm_n4706, gm_n4707, gm_n4708, gm_n4709, gm_n471, gm_n4710, gm_n4711, gm_n4712, gm_n4713, gm_n4714, gm_n4715, gm_n4716, gm_n4717, gm_n4718, gm_n4719, gm_n472, gm_n4720, gm_n4721, gm_n4722, gm_n4723, gm_n4724, gm_n4725, gm_n4726, gm_n4727, gm_n4728, gm_n4729, gm_n473, gm_n4730, gm_n4731, gm_n4732, gm_n4733, gm_n4734, gm_n4735, gm_n4736, gm_n4737, gm_n4738, gm_n4739, gm_n474, gm_n4740, gm_n4741, gm_n4742, gm_n4743, gm_n4744, gm_n4745, gm_n4746, gm_n4747, gm_n4748, gm_n4749, gm_n475, gm_n4750, gm_n4751, gm_n4752, gm_n4753, gm_n4754, gm_n4755, gm_n4756, gm_n4757, gm_n4758, gm_n4759, gm_n476, gm_n4760, gm_n4761, gm_n4762, gm_n4763, gm_n4764, gm_n4765, gm_n4766, gm_n4767, gm_n4768, gm_n4769, gm_n477, gm_n4770, gm_n4771, gm_n4772, gm_n4773, gm_n4774, gm_n4775, gm_n4776, gm_n4777, gm_n4778, gm_n4779, gm_n478, gm_n4780, gm_n4781, gm_n4782, gm_n4783, gm_n4784, gm_n4785, gm_n4786, gm_n4787, gm_n4788, gm_n4789, gm_n479, gm_n4790, gm_n4791, gm_n4792, gm_n4793, gm_n4794, gm_n4795, gm_n4796, gm_n4797, gm_n4798, gm_n4799, gm_n480, gm_n4800, gm_n4801, gm_n4802, gm_n4803, gm_n4804, gm_n4805, gm_n4806, gm_n4807, gm_n4808, gm_n4809, gm_n481, gm_n4810, gm_n4811, gm_n4812, gm_n4813, gm_n4814, gm_n4815, gm_n4816, gm_n4817, gm_n4818, gm_n4819, gm_n482, gm_n4820, gm_n4821, gm_n4822, gm_n4823, gm_n4824, gm_n4825, gm_n4826, gm_n4827, gm_n4828, gm_n4829, gm_n483, gm_n4830, gm_n4831, gm_n4832, gm_n4833, gm_n4834, gm_n4835, gm_n4836, gm_n4837, gm_n4838, gm_n4839, gm_n484, gm_n4840, gm_n4841, gm_n4842, gm_n4843, gm_n4844, gm_n4845, gm_n4846, gm_n4847, gm_n4848, gm_n4849, gm_n485, gm_n4850, gm_n4851, gm_n4852, gm_n4853, gm_n4854, gm_n4855, gm_n4856, gm_n4857, gm_n4858, gm_n4859, gm_n486, gm_n4860, gm_n4861, gm_n4862, gm_n4863, gm_n4864, gm_n4865, gm_n4866, gm_n4867, gm_n4868, gm_n4869, gm_n487, gm_n4870, gm_n4871, gm_n4872, gm_n4873, gm_n4874, gm_n4875, gm_n4876, gm_n4877, gm_n4878, gm_n4879, gm_n488, gm_n4880, gm_n4881, gm_n4882, gm_n4883, gm_n4884, gm_n4885, gm_n4886, gm_n4887, gm_n4888, gm_n4889, gm_n489, gm_n4891, gm_n4892, gm_n4893, gm_n4894, gm_n4895, gm_n4896, gm_n4897, gm_n4898, gm_n4899, gm_n490, gm_n4900, gm_n4901, gm_n4902, gm_n4903, gm_n4904, gm_n4905, gm_n4906, gm_n4907, gm_n4908, gm_n4909, gm_n491, gm_n4910, gm_n4911, gm_n4912, gm_n4913, gm_n4914, gm_n4915, gm_n4916, gm_n4917, gm_n4918, gm_n4919, gm_n492, gm_n4920, gm_n4921, gm_n4922, gm_n4923, gm_n4924, gm_n4925, gm_n4926, gm_n4927, gm_n4928, gm_n4929, gm_n493, gm_n4930, gm_n4931, gm_n4932, gm_n4933, gm_n4934, gm_n4935, gm_n4936, gm_n4937, gm_n4938, gm_n4939, gm_n494, gm_n4940, gm_n4941, gm_n4942, gm_n4943, gm_n4944, gm_n4945, gm_n4946, gm_n4947, gm_n4948, gm_n4949, gm_n495, gm_n4950, gm_n4951, gm_n4952, gm_n4953, gm_n4954, gm_n4955, gm_n4956, gm_n4957, gm_n4958, gm_n4959, gm_n496, gm_n4960, gm_n4961, gm_n4962, gm_n4963, gm_n4964, gm_n4965, gm_n4966, gm_n4967, gm_n4968, gm_n4969, gm_n497, gm_n4970, gm_n4971, gm_n4972, gm_n4973, gm_n4974, gm_n4975, gm_n4976, gm_n4977, gm_n4978, gm_n4979, gm_n498, gm_n4980, gm_n4981, gm_n4982, gm_n4983, gm_n4984, gm_n4985, gm_n4986, gm_n4987, gm_n4988, gm_n4989, gm_n499, gm_n4990, gm_n4991, gm_n4992, gm_n4993, gm_n4994, gm_n4995, gm_n4996, gm_n4997, gm_n4998, gm_n4999, gm_n500, gm_n5000, gm_n5001, gm_n5002, gm_n5003, gm_n5004, gm_n5005, gm_n5006, gm_n5007, gm_n5008, gm_n5009, gm_n501, gm_n5010, gm_n5011, gm_n5012, gm_n5013, gm_n5014, gm_n5015, gm_n5016, gm_n5017, gm_n5018, gm_n5019, gm_n502, gm_n5020, gm_n5021, gm_n5022, gm_n5023, gm_n5024, gm_n5025, gm_n5026, gm_n5027, gm_n5028, gm_n5029, gm_n503, gm_n5030, gm_n5031, gm_n5032, gm_n5033, gm_n5034, gm_n5035, gm_n5036, gm_n5037, gm_n5038, gm_n5039, gm_n504, gm_n5040, gm_n5041, gm_n5042, gm_n5043, gm_n5044, gm_n5045, gm_n5046, gm_n5047, gm_n5048, gm_n5049, gm_n505, gm_n5050, gm_n5051, gm_n5052, gm_n5053, gm_n5054, gm_n5055, gm_n5056, gm_n5057, gm_n5058, gm_n5059, gm_n506, gm_n5060, gm_n5061, gm_n5062, gm_n5063, gm_n5064, gm_n5065, gm_n5066, gm_n5067, gm_n5068, gm_n5069, gm_n507, gm_n5070, gm_n5071, gm_n5072, gm_n5073, gm_n5074, gm_n5075, gm_n5076, gm_n5077, gm_n5078, gm_n5079, gm_n508, gm_n5080, gm_n5081, gm_n5082, gm_n5083, gm_n5084, gm_n5085, gm_n5086, gm_n5087, gm_n5088, gm_n5089, gm_n509, gm_n5090, gm_n5091, gm_n5092, gm_n5093, gm_n5094, gm_n5095, gm_n5096, gm_n5097, gm_n5098, gm_n5099, gm_n510, gm_n5100, gm_n5101, gm_n5102, gm_n5103, gm_n5104, gm_n5105, gm_n5106, gm_n5107, gm_n5108, gm_n5109, gm_n511, gm_n5110, gm_n5111, gm_n5112, gm_n5113, gm_n5114, gm_n5115, gm_n5116, gm_n5117, gm_n5118, gm_n5119, gm_n512, gm_n5120, gm_n5121, gm_n5122, gm_n5123, gm_n5124, gm_n5125, gm_n5126, gm_n5127, gm_n5128, gm_n5129, gm_n513, gm_n5130, gm_n5131, gm_n5132, gm_n5133, gm_n5134, gm_n5135, gm_n5136, gm_n5137, gm_n5138, gm_n5139, gm_n514, gm_n5140, gm_n5141, gm_n5142, gm_n5143, gm_n5144, gm_n5145, gm_n5146, gm_n5147, gm_n5148, gm_n5149, gm_n515, gm_n5150, gm_n5151, gm_n5152, gm_n5153, gm_n5154, gm_n5155, gm_n5156, gm_n5157, gm_n5158, gm_n5159, gm_n516, gm_n5160, gm_n5161, gm_n5162, gm_n5163, gm_n5164, gm_n5165, gm_n5166, gm_n5167, gm_n5168, gm_n5169, gm_n517, gm_n5170, gm_n5171, gm_n5172, gm_n5173, gm_n5174, gm_n5175, gm_n5176, gm_n5177, gm_n5178, gm_n5179, gm_n518, gm_n5180, gm_n5181, gm_n5182, gm_n5183, gm_n5184, gm_n5185, gm_n5186, gm_n5187, gm_n5188, gm_n5189, gm_n519, gm_n5190, gm_n5191, gm_n5192, gm_n5193, gm_n5194, gm_n5195, gm_n5196, gm_n5197, gm_n5198, gm_n5199, gm_n520, gm_n5200, gm_n5201, gm_n5202, gm_n5203, gm_n5204, gm_n5205, gm_n5206, gm_n5207, gm_n5208, gm_n5209, gm_n521, gm_n5210, gm_n5211, gm_n5212, gm_n5213, gm_n5214, gm_n5215, gm_n5216, gm_n5217, gm_n5218, gm_n5219, gm_n522, gm_n5220, gm_n5221, gm_n5222, gm_n5223, gm_n5224, gm_n5225, gm_n5226, gm_n5227, gm_n5228, gm_n5229, gm_n523, gm_n5230, gm_n5231, gm_n5232, gm_n5233, gm_n5234, gm_n5235, gm_n5237, gm_n5238, gm_n5239, gm_n524, gm_n5240, gm_n5241, gm_n5242, gm_n5243, gm_n5244, gm_n5245, gm_n5246, gm_n5247, gm_n5248, gm_n5249, gm_n525, gm_n5250, gm_n5251, gm_n5252, gm_n5253, gm_n5254, gm_n5255, gm_n5256, gm_n5257, gm_n5258, gm_n5259, gm_n526, gm_n5260, gm_n5261, gm_n5262, gm_n5263, gm_n5264, gm_n5265, gm_n5266, gm_n5267, gm_n5268, gm_n5269, gm_n527, gm_n5270, gm_n5271, gm_n5272, gm_n5273, gm_n5274, gm_n5275, gm_n5276, gm_n5277, gm_n5278, gm_n5279, gm_n528, gm_n5280, gm_n5281, gm_n5282, gm_n5283, gm_n5284, gm_n5285, gm_n5286, gm_n5287, gm_n5288, gm_n5289, gm_n529, gm_n5290, gm_n5291, gm_n5292, gm_n5293, gm_n5294, gm_n5295, gm_n5296, gm_n5297, gm_n5298, gm_n5299, gm_n530, gm_n5300, gm_n5301, gm_n5302, gm_n5303, gm_n5304, gm_n5305, gm_n5306, gm_n5307, gm_n5308, gm_n5309, gm_n531, gm_n5310, gm_n5311, gm_n5312, gm_n5313, gm_n5314, gm_n5315, gm_n5316, gm_n5317, gm_n5318, gm_n5319, gm_n532, gm_n5320, gm_n5321, gm_n5322, gm_n5323, gm_n5324, gm_n5325, gm_n5326, gm_n5327, gm_n5328, gm_n5329, gm_n533, gm_n5330, gm_n5331, gm_n5332, gm_n5333, gm_n5334, gm_n5335, gm_n5336, gm_n5337, gm_n5338, gm_n5339, gm_n534, gm_n5340, gm_n5341, gm_n5342, gm_n5343, gm_n5344, gm_n5345, gm_n5346, gm_n5347, gm_n5348, gm_n5349, gm_n535, gm_n5350, gm_n5351, gm_n5352, gm_n5353, gm_n5354, gm_n5355, gm_n5356, gm_n5357, gm_n5358, gm_n5359, gm_n536, gm_n5360, gm_n5361, gm_n5362, gm_n5363, gm_n5364, gm_n5365, gm_n5366, gm_n5367, gm_n5368, gm_n5369, gm_n537, gm_n5370, gm_n5371, gm_n5372, gm_n5373, gm_n5374, gm_n5375, gm_n5376, gm_n5377, gm_n5378, gm_n5379, gm_n538, gm_n5380, gm_n5381, gm_n5382, gm_n5383, gm_n5384, gm_n5385, gm_n5386, gm_n5387, gm_n5388, gm_n5389, gm_n539, gm_n5390, gm_n5391, gm_n5392, gm_n5393, gm_n5394, gm_n5395, gm_n5396, gm_n5397, gm_n5398, gm_n5399, gm_n540, gm_n5400, gm_n5401, gm_n5402, gm_n5403, gm_n5404, gm_n5405, gm_n5406, gm_n5407, gm_n5408, gm_n5409, gm_n541, gm_n5410, gm_n5411, gm_n5412, gm_n5413, gm_n5414, gm_n5415, gm_n5416, gm_n5417, gm_n5418, gm_n5419, gm_n542, gm_n5420, gm_n5421, gm_n5422, gm_n5423, gm_n5424, gm_n5425, gm_n5426, gm_n5427, gm_n5428, gm_n5429, gm_n543, gm_n5430, gm_n5431, gm_n5432, gm_n5433, gm_n5434, gm_n5435, gm_n5436, gm_n5437, gm_n5438, gm_n544, gm_n5440, gm_n5441, gm_n5442, gm_n5443, gm_n5444, gm_n5445, gm_n5446, gm_n5447, gm_n5448, gm_n5449, gm_n545, gm_n5450, gm_n5451, gm_n5452, gm_n5453, gm_n5454, gm_n5455, gm_n5456, gm_n5457, gm_n5458, gm_n5459, gm_n546, gm_n5460, gm_n5461, gm_n5462, gm_n5463, gm_n5464, gm_n5465, gm_n5466, gm_n5467, gm_n5468, gm_n5469, gm_n547, gm_n5470, gm_n5471, gm_n5472, gm_n5473, gm_n5474, gm_n5475, gm_n5476, gm_n5478, gm_n5479, gm_n548, gm_n5480, gm_n5481, gm_n5482, gm_n5483, gm_n5484, gm_n5485, gm_n5486, gm_n5487, gm_n5488, gm_n5489, gm_n549, gm_n5490, gm_n5491, gm_n5492, gm_n5493, gm_n5494, gm_n5495, gm_n5496, gm_n5497, gm_n5498, gm_n5499, gm_n55, gm_n550, gm_n5500, gm_n5501, gm_n5502, gm_n5503, gm_n5504, gm_n5505, gm_n5506, gm_n5507, gm_n5508, gm_n5509, gm_n551, gm_n5510, gm_n5511, gm_n5512, gm_n5513, gm_n5514, gm_n5515, gm_n5516, gm_n5517, gm_n5518, gm_n5519, gm_n552, gm_n5520, gm_n5521, gm_n5522, gm_n5523, gm_n5524, gm_n5525, gm_n5526, gm_n5527, gm_n5528, gm_n5529, gm_n553, gm_n5530, gm_n5531, gm_n5532, gm_n5533, gm_n5534, gm_n5535, gm_n5536, gm_n5537, gm_n5538, gm_n5539, gm_n554, gm_n5540, gm_n5541, gm_n5542, gm_n5543, gm_n5544, gm_n5545, gm_n5546, gm_n5547, gm_n5548, gm_n5549, gm_n555, gm_n5550, gm_n5551, gm_n5552, gm_n5553, gm_n5554, gm_n5555, gm_n5556, gm_n5557, gm_n5558, gm_n5559, gm_n556, gm_n5560, gm_n5561, gm_n5562, gm_n5563, gm_n5564, gm_n5565, gm_n5566, gm_n5567, gm_n5568, gm_n5569, gm_n557, gm_n5570, gm_n5571, gm_n5572, gm_n5573, gm_n5574, gm_n5575, gm_n5576, gm_n5577, gm_n5578, gm_n5579, gm_n558, gm_n5580, gm_n5581, gm_n5582, gm_n5583, gm_n5584, gm_n5585, gm_n5586, gm_n5587, gm_n5588, gm_n5589, gm_n559, gm_n5590, gm_n5591, gm_n5592, gm_n5593, gm_n5594, gm_n5595, gm_n5596, gm_n5597, gm_n5598, gm_n5599, gm_n56, gm_n560, gm_n5600, gm_n5601, gm_n5602, gm_n5603, gm_n5604, gm_n5605, gm_n5606, gm_n5607, gm_n5608, gm_n5609, gm_n561, gm_n5610, gm_n5611, gm_n5612, gm_n5613, gm_n5614, gm_n5615, gm_n5616, gm_n5617, gm_n5618, gm_n5619, gm_n562, gm_n5620, gm_n5621, gm_n5622, gm_n5623, gm_n5624, gm_n5625, gm_n5626, gm_n5627, gm_n5628, gm_n5629, gm_n563, gm_n5630, gm_n5631, gm_n5632, gm_n5633, gm_n5634, gm_n5635, gm_n5636, gm_n5637, gm_n5638, gm_n5639, gm_n564, gm_n5640, gm_n5641, gm_n5642, gm_n5643, gm_n5644, gm_n5645, gm_n5646, gm_n5647, gm_n5648, gm_n5649, gm_n565, gm_n5650, gm_n5651, gm_n5652, gm_n5653, gm_n5654, gm_n5655, gm_n5656, gm_n5657, gm_n5658, gm_n5659, gm_n566, gm_n5660, gm_n5661, gm_n5662, gm_n5663, gm_n5664, gm_n5665, gm_n5666, gm_n5667, gm_n5668, gm_n5669, gm_n567, gm_n5670, gm_n5671, gm_n5672, gm_n5673, gm_n5674, gm_n5675, gm_n5676, gm_n5677, gm_n5678, gm_n5679, gm_n568, gm_n5680, gm_n5681, gm_n5682, gm_n5683, gm_n5684, gm_n5685, gm_n5686, gm_n5687, gm_n5688, gm_n5689, gm_n569, gm_n5690, gm_n5691, gm_n5692, gm_n5693, gm_n5694, gm_n5695, gm_n5696, gm_n5697, gm_n5698, gm_n5699, gm_n57, gm_n570, gm_n5700, gm_n5701, gm_n5702, gm_n5703, gm_n5704, gm_n5705, gm_n5706, gm_n5707, gm_n5708, gm_n5709, gm_n571, gm_n5710, gm_n5711, gm_n5712, gm_n5713, gm_n5714, gm_n5715, gm_n5716, gm_n5717, gm_n5718, gm_n5719, gm_n572, gm_n5720, gm_n5721, gm_n5722, gm_n5723, gm_n5724, gm_n5725, gm_n5726, gm_n5727, gm_n5728, gm_n5729, gm_n573, gm_n5730, gm_n5731, gm_n5732, gm_n5733, gm_n5734, gm_n5735, gm_n5736, gm_n5737, gm_n5738, gm_n5739, gm_n574, gm_n5740, gm_n5741, gm_n5742, gm_n5743, gm_n5744, gm_n5745, gm_n5746, gm_n5747, gm_n5748, gm_n5749, gm_n575, gm_n5750, gm_n5751, gm_n5752, gm_n5753, gm_n5754, gm_n5755, gm_n5756, gm_n5757, gm_n5758, gm_n5759, gm_n576, gm_n5760, gm_n5761, gm_n5762, gm_n5763, gm_n5764, gm_n5765, gm_n5766, gm_n5767, gm_n5768, gm_n5769, gm_n577, gm_n5770, gm_n5771, gm_n5772, gm_n5773, gm_n5774, gm_n5775, gm_n5776, gm_n5777, gm_n5778, gm_n5779, gm_n578, gm_n5780, gm_n5781, gm_n5782, gm_n5783, gm_n5784, gm_n5785, gm_n5786, gm_n5787, gm_n5788, gm_n5789, gm_n579, gm_n5790, gm_n5791, gm_n5792, gm_n5793, gm_n5794, gm_n5795, gm_n5796, gm_n5797, gm_n5798, gm_n5799, gm_n58, gm_n580, gm_n5800, gm_n5801, gm_n5802, gm_n5803, gm_n5804, gm_n5805, gm_n5806, gm_n5807, gm_n5808, gm_n581, gm_n5810, gm_n5811, gm_n5812, gm_n5813, gm_n5814, gm_n5815, gm_n5816, gm_n5817, gm_n5818, gm_n5819, gm_n582, gm_n5820, gm_n5821, gm_n5822, gm_n5823, gm_n5824, gm_n5825, gm_n5826, gm_n5827, gm_n5828, gm_n5829, gm_n583, gm_n5830, gm_n5831, gm_n5832, gm_n5833, gm_n5834, gm_n5835, gm_n5836, gm_n5837, gm_n5838, gm_n5839, gm_n584, gm_n5840, gm_n5841, gm_n5842, gm_n5843, gm_n5844, gm_n5845, gm_n5846, gm_n5847, gm_n5848, gm_n5849, gm_n585, gm_n5850, gm_n5851, gm_n5852, gm_n5853, gm_n5854, gm_n5855, gm_n5856, gm_n5857, gm_n5858, gm_n5859, gm_n586, gm_n5860, gm_n5861, gm_n5862, gm_n5863, gm_n5864, gm_n5865, gm_n5866, gm_n5867, gm_n5868, gm_n5869, gm_n587, gm_n5870, gm_n5871, gm_n5872, gm_n5873, gm_n5874, gm_n5875, gm_n5876, gm_n5877, gm_n5878, gm_n5879, gm_n588, gm_n5880, gm_n5881, gm_n5882, gm_n5883, gm_n5884, gm_n5885, gm_n5886, gm_n5887, gm_n5888, gm_n5889, gm_n589, gm_n5890, gm_n5891, gm_n5892, gm_n5893, gm_n5894, gm_n5895, gm_n5896, gm_n5897, gm_n5898, gm_n5899, gm_n59, gm_n590, gm_n5900, gm_n5901, gm_n5902, gm_n5903, gm_n5904, gm_n5905, gm_n5906, gm_n5907, gm_n5908, gm_n5909, gm_n591, gm_n5910, gm_n5911, gm_n5912, gm_n5913, gm_n5914, gm_n5915, gm_n5916, gm_n5917, gm_n5918, gm_n5919, gm_n592, gm_n5920, gm_n5921, gm_n5922, gm_n5923, gm_n5924, gm_n5925, gm_n5926, gm_n5927, gm_n5928, gm_n5929, gm_n593, gm_n5930, gm_n5931, gm_n5932, gm_n5933, gm_n5934, gm_n5935, gm_n5936, gm_n5937, gm_n5938, gm_n5939, gm_n594, gm_n5940, gm_n5941, gm_n5942, gm_n5943, gm_n5944, gm_n5945, gm_n5946, gm_n5947, gm_n5948, gm_n5949, gm_n595, gm_n5950, gm_n5951, gm_n5952, gm_n5953, gm_n5954, gm_n5955, gm_n5956, gm_n5957, gm_n5958, gm_n5959, gm_n596, gm_n5960, gm_n5961, gm_n5962, gm_n5963, gm_n5964, gm_n5965, gm_n5966, gm_n5967, gm_n5968, gm_n5969, gm_n597, gm_n5970, gm_n5971, gm_n5972, gm_n5973, gm_n5974, gm_n5975, gm_n5976, gm_n5977, gm_n5978, gm_n5979, gm_n598, gm_n5980, gm_n5981, gm_n5982, gm_n5983, gm_n5984, gm_n5985, gm_n5986, gm_n5987, gm_n5988, gm_n5989, gm_n599, gm_n5990, gm_n5991, gm_n5992, gm_n5993, gm_n5994, gm_n5995, gm_n5996, gm_n5997, gm_n5998, gm_n5999, gm_n60, gm_n600, gm_n6000, gm_n6001, gm_n6002, gm_n6003, gm_n6004, gm_n6005, gm_n6006, gm_n6007, gm_n6008, gm_n6009, gm_n601, gm_n6010, gm_n6011, gm_n6012, gm_n6013, gm_n6014, gm_n6015, gm_n6016, gm_n6017, gm_n6018, gm_n6019, gm_n602, gm_n6020, gm_n6021, gm_n6022, gm_n6023, gm_n6024, gm_n6025, gm_n6026, gm_n6027, gm_n6028, gm_n6029, gm_n603, gm_n6030, gm_n6031, gm_n6032, gm_n6033, gm_n6034, gm_n6035, gm_n6036, gm_n6037, gm_n6038, gm_n6039, gm_n604, gm_n6040, gm_n6041, gm_n6042, gm_n6043, gm_n6044, gm_n6045, gm_n6046, gm_n6047, gm_n6048, gm_n6049, gm_n605, gm_n6050, gm_n6051, gm_n6052, gm_n6053, gm_n6054, gm_n6055, gm_n6056, gm_n6057, gm_n6058, gm_n6059, gm_n606, gm_n6060, gm_n6061, gm_n6062, gm_n6063, gm_n6064, gm_n6065, gm_n6066, gm_n6067, gm_n6068, gm_n6069, gm_n607, gm_n6070, gm_n6071, gm_n6072, gm_n6073, gm_n6074, gm_n6075, gm_n6076, gm_n6077, gm_n6078, gm_n6079, gm_n608, gm_n6080, gm_n6081, gm_n6082, gm_n6083, gm_n6084, gm_n6085, gm_n6086, gm_n6087, gm_n6088, gm_n6089, gm_n609, gm_n6090, gm_n6091, gm_n6092, gm_n6093, gm_n6094, gm_n6095, gm_n6096, gm_n6097, gm_n6098, gm_n6099, gm_n61, gm_n610, gm_n6100, gm_n6101, gm_n6102, gm_n6103, gm_n6104, gm_n6105, gm_n6106, gm_n6107, gm_n6108, gm_n6109, gm_n611, gm_n6110, gm_n6111, gm_n6112, gm_n6113, gm_n6114, gm_n6115, gm_n6116, gm_n6117, gm_n6118, gm_n6119, gm_n612, gm_n6120, gm_n6121, gm_n6122, gm_n6123, gm_n6124, gm_n6125, gm_n6126, gm_n6127, gm_n6128, gm_n6129, gm_n613, gm_n6130, gm_n6131, gm_n6132, gm_n6133, gm_n6134, gm_n6135, gm_n6136, gm_n6137, gm_n6138, gm_n6139, gm_n614, gm_n6140, gm_n6141, gm_n6142, gm_n6143, gm_n6144, gm_n6145, gm_n6147, gm_n6148, gm_n6149, gm_n615, gm_n6150, gm_n6151, gm_n6152, gm_n6153, gm_n6154, gm_n6155, gm_n6156, gm_n6157, gm_n6158, gm_n6159, gm_n616, gm_n6160, gm_n6161, gm_n6162, gm_n6163, gm_n6164, gm_n6165, gm_n6166, gm_n6167, gm_n6168, gm_n6169, gm_n617, gm_n6170, gm_n6171, gm_n6172, gm_n6173, gm_n6174, gm_n6175, gm_n6176, gm_n6177, gm_n6178, gm_n6179, gm_n618, gm_n6180, gm_n6181, gm_n6182, gm_n6183, gm_n6184, gm_n6185, gm_n6186, gm_n6187, gm_n6188, gm_n6189, gm_n619, gm_n6190, gm_n6191, gm_n6192, gm_n6193, gm_n6194, gm_n6195, gm_n6196, gm_n6197, gm_n6198, gm_n6199, gm_n62, gm_n620, gm_n6200, gm_n6201, gm_n6202, gm_n6203, gm_n6204, gm_n6205, gm_n6206, gm_n6207, gm_n6208, gm_n6209, gm_n621, gm_n6210, gm_n6211, gm_n6212, gm_n6213, gm_n6214, gm_n6215, gm_n6216, gm_n6217, gm_n6218, gm_n6219, gm_n622, gm_n6220, gm_n6221, gm_n6222, gm_n6223, gm_n6224, gm_n6225, gm_n6226, gm_n6227, gm_n6228, gm_n6229, gm_n623, gm_n6230, gm_n6231, gm_n6232, gm_n6233, gm_n6234, gm_n6235, gm_n6236, gm_n6237, gm_n6238, gm_n6239, gm_n624, gm_n6240, gm_n6241, gm_n6242, gm_n6243, gm_n6244, gm_n6245, gm_n6246, gm_n6247, gm_n6248, gm_n6249, gm_n625, gm_n6250, gm_n6251, gm_n6252, gm_n6253, gm_n6254, gm_n6255, gm_n6256, gm_n6257, gm_n6258, gm_n6259, gm_n626, gm_n6260, gm_n6261, gm_n6262, gm_n6263, gm_n6264, gm_n6265, gm_n6266, gm_n6267, gm_n6268, gm_n6269, gm_n627, gm_n6270, gm_n6271, gm_n6272, gm_n6273, gm_n6274, gm_n6275, gm_n6276, gm_n6277, gm_n6278, gm_n6279, gm_n628, gm_n6280, gm_n6281, gm_n6282, gm_n6283, gm_n6284, gm_n6285, gm_n6286, gm_n6287, gm_n6288, gm_n6289, gm_n629, gm_n6290, gm_n6291, gm_n6292, gm_n6293, gm_n6294, gm_n6295, gm_n6296, gm_n6297, gm_n6298, gm_n6299, gm_n63, gm_n630, gm_n6300, gm_n6301, gm_n6302, gm_n6303, gm_n6304, gm_n6305, gm_n6306, gm_n6307, gm_n6308, gm_n6309, gm_n631, gm_n6310, gm_n6311, gm_n6312, gm_n6313, gm_n6314, gm_n6315, gm_n6316, gm_n6317, gm_n6318, gm_n6319, gm_n632, gm_n6320, gm_n6321, gm_n6322, gm_n6323, gm_n6324, gm_n6325, gm_n6326, gm_n6327, gm_n6328, gm_n6329, gm_n633, gm_n6330, gm_n6331, gm_n6332, gm_n6333, gm_n6334, gm_n6335, gm_n6336, gm_n6337, gm_n6338, gm_n6339, gm_n634, gm_n6340, gm_n6341, gm_n6342, gm_n6343, gm_n6344, gm_n6345, gm_n6346, gm_n6347, gm_n6348, gm_n6349, gm_n635, gm_n6350, gm_n6351, gm_n6352, gm_n6353, gm_n6354, gm_n6355, gm_n6356, gm_n6357, gm_n6358, gm_n6359, gm_n636, gm_n6360, gm_n6361, gm_n6362, gm_n6363, gm_n6364, gm_n6365, gm_n6366, gm_n6367, gm_n6368, gm_n6369, gm_n637, gm_n6370, gm_n6371, gm_n6372, gm_n6373, gm_n6374, gm_n6375, gm_n6376, gm_n6377, gm_n6378, gm_n6379, gm_n638, gm_n6380, gm_n6381, gm_n6382, gm_n6383, gm_n6384, gm_n6385, gm_n6386, gm_n6387, gm_n6388, gm_n6389, gm_n639, gm_n6390, gm_n6391, gm_n6392, gm_n6393, gm_n6394, gm_n6395, gm_n6396, gm_n6397, gm_n6398, gm_n6399, gm_n64, gm_n640, gm_n6400, gm_n6401, gm_n6402, gm_n6403, gm_n6404, gm_n6405, gm_n6406, gm_n6407, gm_n6408, gm_n6409, gm_n641, gm_n6410, gm_n6411, gm_n6412, gm_n6413, gm_n6414, gm_n6415, gm_n6416, gm_n6417, gm_n6418, gm_n6419, gm_n642, gm_n6420, gm_n6421, gm_n6422, gm_n6423, gm_n6424, gm_n6425, gm_n6426, gm_n6427, gm_n6428, gm_n6429, gm_n643, gm_n6430, gm_n6431, gm_n6432, gm_n6433, gm_n6434, gm_n6435, gm_n6436, gm_n6437, gm_n6438, gm_n6439, gm_n644, gm_n6440, gm_n6441, gm_n6442, gm_n6443, gm_n6444, gm_n6445, gm_n6446, gm_n6447, gm_n6448, gm_n6449, gm_n645, gm_n6450, gm_n6451, gm_n6452, gm_n6453, gm_n6454, gm_n6455, gm_n6456, gm_n6457, gm_n6458, gm_n6459, gm_n646, gm_n6460, gm_n6461, gm_n6462, gm_n6463, gm_n6464, gm_n6465, gm_n6466, gm_n6467, gm_n6468, gm_n6469, gm_n647, gm_n6470, gm_n6471, gm_n6472, gm_n6473, gm_n6474, gm_n6475, gm_n6476, gm_n6477, gm_n6478, gm_n6479, gm_n648, gm_n6480, gm_n6481, gm_n6482, gm_n6483, gm_n6484, gm_n6485, gm_n6486, gm_n6487, gm_n6488, gm_n649, gm_n6490, gm_n6491, gm_n6492, gm_n6493, gm_n6494, gm_n6495, gm_n6496, gm_n6497, gm_n6498, gm_n6499, gm_n65, gm_n650, gm_n6500, gm_n6501, gm_n6502, gm_n6503, gm_n6504, gm_n6505, gm_n6506, gm_n6507, gm_n6508, gm_n6509, gm_n651, gm_n6510, gm_n6511, gm_n6512, gm_n6513, gm_n6514, gm_n6515, gm_n6516, gm_n6517, gm_n6518, gm_n6519, gm_n652, gm_n6520, gm_n6521, gm_n6522, gm_n6523, gm_n6524, gm_n6525, gm_n6526, gm_n6527, gm_n6528, gm_n6529, gm_n653, gm_n6530, gm_n6531, gm_n6532, gm_n6533, gm_n6534, gm_n6535, gm_n6536, gm_n6537, gm_n6538, gm_n6539, gm_n654, gm_n6540, gm_n6541, gm_n6542, gm_n6543, gm_n6544, gm_n6545, gm_n6546, gm_n6547, gm_n6548, gm_n6549, gm_n655, gm_n6550, gm_n6551, gm_n6552, gm_n6553, gm_n6554, gm_n6555, gm_n6556, gm_n6557, gm_n6558, gm_n6559, gm_n656, gm_n6560, gm_n6561, gm_n6562, gm_n6563, gm_n6564, gm_n6565, gm_n6566, gm_n6567, gm_n6568, gm_n6569, gm_n657, gm_n6570, gm_n6571, gm_n6572, gm_n6573, gm_n6574, gm_n6575, gm_n6576, gm_n6577, gm_n6578, gm_n6579, gm_n658, gm_n6580, gm_n6581, gm_n6582, gm_n6583, gm_n6584, gm_n6585, gm_n6586, gm_n6587, gm_n6588, gm_n6589, gm_n659, gm_n6590, gm_n6591, gm_n6592, gm_n6593, gm_n6594, gm_n6595, gm_n6596, gm_n6597, gm_n6598, gm_n6599, gm_n66, gm_n660, gm_n6600, gm_n6601, gm_n6602, gm_n6603, gm_n6604, gm_n6605, gm_n6606, gm_n6607, gm_n6608, gm_n6609, gm_n661, gm_n6610, gm_n6611, gm_n6612, gm_n6613, gm_n6614, gm_n6615, gm_n6616, gm_n6617, gm_n6618, gm_n6619, gm_n662, gm_n6620, gm_n6621, gm_n6622, gm_n6623, gm_n6624, gm_n6625, gm_n6626, gm_n6627, gm_n6628, gm_n6629, gm_n663, gm_n6630, gm_n6631, gm_n6632, gm_n6633, gm_n6634, gm_n6635, gm_n6636, gm_n6637, gm_n6638, gm_n6639, gm_n664, gm_n6640, gm_n6641, gm_n6642, gm_n6643, gm_n6644, gm_n6645, gm_n6646, gm_n6647, gm_n6648, gm_n6649, gm_n665, gm_n6650, gm_n6651, gm_n6652, gm_n6653, gm_n6654, gm_n6655, gm_n6656, gm_n6657, gm_n6658, gm_n6659, gm_n666, gm_n6660, gm_n6661, gm_n6662, gm_n6663, gm_n6664, gm_n6665, gm_n6666, gm_n6667, gm_n6668, gm_n6669, gm_n667, gm_n6670, gm_n6671, gm_n6672, gm_n6673, gm_n6674, gm_n6675, gm_n6676, gm_n6677, gm_n6678, gm_n6679, gm_n668, gm_n6680, gm_n6681, gm_n6682, gm_n6683, gm_n6684, gm_n6685, gm_n6686, gm_n6687, gm_n6688, gm_n6689, gm_n669, gm_n6690, gm_n6691, gm_n6692, gm_n6693, gm_n6694, gm_n6695, gm_n6696, gm_n6697, gm_n6698, gm_n6699, gm_n67, gm_n670, gm_n6700, gm_n6701, gm_n6702, gm_n6703, gm_n6704, gm_n6705, gm_n6706, gm_n6707, gm_n6708, gm_n6709, gm_n671, gm_n6710, gm_n6711, gm_n6712, gm_n6713, gm_n6714, gm_n6715, gm_n6716, gm_n6717, gm_n6718, gm_n6719, gm_n672, gm_n6720, gm_n6721, gm_n6722, gm_n6723, gm_n6724, gm_n6725, gm_n6726, gm_n6727, gm_n6728, gm_n6729, gm_n673, gm_n6730, gm_n6731, gm_n6732, gm_n6733, gm_n6734, gm_n6735, gm_n6736, gm_n6737, gm_n6738, gm_n6739, gm_n674, gm_n6740, gm_n6741, gm_n6742, gm_n6743, gm_n6744, gm_n6745, gm_n6746, gm_n6747, gm_n6748, gm_n6749, gm_n675, gm_n6750, gm_n6751, gm_n6752, gm_n6753, gm_n6754, gm_n6755, gm_n6756, gm_n6757, gm_n6758, gm_n6759, gm_n676, gm_n6760, gm_n6761, gm_n6762, gm_n6763, gm_n6764, gm_n6765, gm_n6766, gm_n6767, gm_n6768, gm_n6769, gm_n677, gm_n6770, gm_n6771, gm_n6772, gm_n6773, gm_n6774, gm_n6775, gm_n6776, gm_n6777, gm_n6778, gm_n6779, gm_n678, gm_n6780, gm_n6781, gm_n6782, gm_n6783, gm_n6784, gm_n6785, gm_n6786, gm_n6787, gm_n6788, gm_n6789, gm_n679, gm_n6790, gm_n6791, gm_n6792, gm_n6793, gm_n6794, gm_n6795, gm_n6796, gm_n6797, gm_n6798, gm_n6799, gm_n68, gm_n680, gm_n6800, gm_n6801, gm_n6802, gm_n6803, gm_n6804, gm_n6805, gm_n6806, gm_n6807, gm_n6808, gm_n6809, gm_n681, gm_n6810, gm_n6811, gm_n6812, gm_n6813, gm_n6814, gm_n6815, gm_n6816, gm_n6817, gm_n6818, gm_n6819, gm_n682, gm_n6820, gm_n6821, gm_n6822, gm_n6823, gm_n6824, gm_n6826, gm_n6827, gm_n6828, gm_n6829, gm_n683, gm_n6830, gm_n6831, gm_n6832, gm_n6833, gm_n6834, gm_n6835, gm_n6836, gm_n6837, gm_n6838, gm_n6839, gm_n684, gm_n6840, gm_n6841, gm_n6842, gm_n6843, gm_n6844, gm_n6845, gm_n6846, gm_n6847, gm_n6848, gm_n6849, gm_n685, gm_n6850, gm_n6851, gm_n6852, gm_n6853, gm_n6854, gm_n6855, gm_n6856, gm_n6857, gm_n6858, gm_n6859, gm_n686, gm_n6860, gm_n6861, gm_n6862, gm_n6863, gm_n6864, gm_n6865, gm_n6866, gm_n6867, gm_n6868, gm_n6869, gm_n687, gm_n6870, gm_n6871, gm_n6872, gm_n6873, gm_n6874, gm_n6875, gm_n6876, gm_n6877, gm_n6878, gm_n6879, gm_n688, gm_n6880, gm_n6881, gm_n6882, gm_n6883, gm_n6884, gm_n6885, gm_n6886, gm_n6887, gm_n6888, gm_n6889, gm_n689, gm_n6890, gm_n6891, gm_n6892, gm_n6893, gm_n6894, gm_n6895, gm_n6896, gm_n6897, gm_n6898, gm_n6899, gm_n69, gm_n690, gm_n6900, gm_n6901, gm_n6902, gm_n6903, gm_n6904, gm_n6905, gm_n6906, gm_n6907, gm_n6908, gm_n6909, gm_n691, gm_n6910, gm_n6911, gm_n6912, gm_n6913, gm_n6914, gm_n6915, gm_n6916, gm_n6917, gm_n6918, gm_n6919, gm_n692, gm_n6920, gm_n6921, gm_n6922, gm_n6923, gm_n6924, gm_n6925, gm_n6926, gm_n6927, gm_n6928, gm_n6929, gm_n693, gm_n6930, gm_n6931, gm_n6932, gm_n6933, gm_n6934, gm_n6935, gm_n6936, gm_n6937, gm_n6938, gm_n6939, gm_n694, gm_n6940, gm_n6941, gm_n6942, gm_n6943, gm_n6944, gm_n6945, gm_n6946, gm_n6947, gm_n6948, gm_n6949, gm_n695, gm_n6950, gm_n6951, gm_n6952, gm_n6953, gm_n6954, gm_n6955, gm_n6956, gm_n6957, gm_n6958, gm_n6959, gm_n696, gm_n6960, gm_n6961, gm_n6962, gm_n6963, gm_n6964, gm_n6965, gm_n6966, gm_n6967, gm_n6968, gm_n6969, gm_n697, gm_n6970, gm_n6971, gm_n6972, gm_n6973, gm_n6974, gm_n6975, gm_n6976, gm_n6977, gm_n6978, gm_n6979, gm_n698, gm_n6980, gm_n6981, gm_n6982, gm_n6983, gm_n6984, gm_n6985, gm_n6986, gm_n6987, gm_n6988, gm_n6989, gm_n699, gm_n6990, gm_n6991, gm_n6992, gm_n6993, gm_n6994, gm_n6995, gm_n6996, gm_n6997, gm_n6998, gm_n6999, gm_n70, gm_n700, gm_n7000, gm_n7001, gm_n7002, gm_n7003, gm_n7004, gm_n7005, gm_n7006, gm_n7007, gm_n7008, gm_n7009, gm_n701, gm_n7010, gm_n7011, gm_n7012, gm_n7013, gm_n7014, gm_n7015, gm_n7016, gm_n7017, gm_n7018, gm_n7019, gm_n702, gm_n7020, gm_n7021, gm_n7022, gm_n7023, gm_n7024, gm_n7025, gm_n7026, gm_n7027, gm_n7028, gm_n7029, gm_n703, gm_n7030, gm_n7031, gm_n7032, gm_n7033, gm_n7034, gm_n7035, gm_n7036, gm_n7037, gm_n7038, gm_n7039, gm_n704, gm_n7040, gm_n7041, gm_n7042, gm_n7043, gm_n7044, gm_n7045, gm_n7046, gm_n7047, gm_n7048, gm_n7049, gm_n705, gm_n7050, gm_n7051, gm_n7052, gm_n7053, gm_n7054, gm_n7055, gm_n7056, gm_n7057, gm_n7058, gm_n7059, gm_n706, gm_n7060, gm_n7061, gm_n7062, gm_n7063, gm_n7064, gm_n7065, gm_n7066, gm_n7067, gm_n7068, gm_n7069, gm_n707, gm_n7070, gm_n7071, gm_n7072, gm_n7073, gm_n7074, gm_n7075, gm_n7076, gm_n7077, gm_n7078, gm_n7079, gm_n708, gm_n7080, gm_n7081, gm_n7082, gm_n7083, gm_n7084, gm_n7085, gm_n7086, gm_n7087, gm_n7088, gm_n7089, gm_n709, gm_n7090, gm_n7091, gm_n7092, gm_n7093, gm_n7094, gm_n7095, gm_n7096, gm_n7097, gm_n7098, gm_n7099, gm_n71, gm_n710, gm_n7100, gm_n7101, gm_n7102, gm_n7103, gm_n7104, gm_n7105, gm_n7106, gm_n7107, gm_n7108, gm_n7109, gm_n711, gm_n7110, gm_n7111, gm_n7112, gm_n7113, gm_n7114, gm_n7115, gm_n7116, gm_n7117, gm_n7118, gm_n7119, gm_n712, gm_n7120, gm_n7121, gm_n7122, gm_n7123, gm_n7124, gm_n7125, gm_n7126, gm_n7127, gm_n7128, gm_n7129, gm_n713, gm_n7130, gm_n7131, gm_n7132, gm_n7133, gm_n7134, gm_n7135, gm_n7136, gm_n7137, gm_n7138, gm_n7139, gm_n714, gm_n7140, gm_n7141, gm_n7142, gm_n7143, gm_n7144, gm_n7145, gm_n7146, gm_n7147, gm_n7148, gm_n7149, gm_n715, gm_n7150, gm_n7151, gm_n7152, gm_n7153, gm_n7154, gm_n7155, gm_n7156, gm_n7157, gm_n7158, gm_n7159, gm_n716, gm_n7160, gm_n7161, gm_n7163, gm_n7164, gm_n7165, gm_n7166, gm_n7167, gm_n7168, gm_n7169, gm_n717, gm_n7170, gm_n7171, gm_n7172, gm_n7173, gm_n7174, gm_n7175, gm_n7176, gm_n7177, gm_n7178, gm_n7179, gm_n718, gm_n7180, gm_n7181, gm_n7182, gm_n7183, gm_n7184, gm_n7185, gm_n7186, gm_n7187, gm_n7188, gm_n7189, gm_n719, gm_n7190, gm_n7191, gm_n7192, gm_n7193, gm_n7194, gm_n7195, gm_n7196, gm_n7197, gm_n7198, gm_n7199, gm_n72, gm_n720, gm_n7200, gm_n7201, gm_n7202, gm_n7203, gm_n7204, gm_n7205, gm_n7206, gm_n7207, gm_n7208, gm_n7209, gm_n721, gm_n7210, gm_n7211, gm_n7212, gm_n7213, gm_n7214, gm_n7215, gm_n7216, gm_n7217, gm_n7218, gm_n7219, gm_n722, gm_n7220, gm_n7221, gm_n7222, gm_n7223, gm_n7224, gm_n7225, gm_n7226, gm_n7227, gm_n7228, gm_n7229, gm_n723, gm_n7230, gm_n7231, gm_n7232, gm_n7233, gm_n7234, gm_n7235, gm_n7236, gm_n7237, gm_n7238, gm_n7239, gm_n724, gm_n7240, gm_n7241, gm_n7242, gm_n7243, gm_n7244, gm_n7245, gm_n7246, gm_n7247, gm_n7248, gm_n7249, gm_n725, gm_n7250, gm_n7251, gm_n7252, gm_n7253, gm_n7254, gm_n7255, gm_n7256, gm_n7257, gm_n7258, gm_n7259, gm_n726, gm_n7260, gm_n7261, gm_n7262, gm_n7263, gm_n7264, gm_n7265, gm_n7266, gm_n7267, gm_n7268, gm_n7269, gm_n727, gm_n7270, gm_n7271, gm_n7272, gm_n7273, gm_n7274, gm_n7275, gm_n7276, gm_n7277, gm_n7278, gm_n7279, gm_n728, gm_n7280, gm_n7281, gm_n7282, gm_n7283, gm_n7284, gm_n7285, gm_n7286, gm_n7287, gm_n7288, gm_n7289, gm_n729, gm_n7290, gm_n7291, gm_n7292, gm_n7293, gm_n7294, gm_n7295, gm_n7296, gm_n7297, gm_n7298, gm_n7299, gm_n73, gm_n730, gm_n7300, gm_n7301, gm_n7302, gm_n7303, gm_n7304, gm_n7305, gm_n7306, gm_n7307, gm_n7308, gm_n7309, gm_n731, gm_n7310, gm_n7311, gm_n7312, gm_n7313, gm_n7314, gm_n7315, gm_n7316, gm_n7317, gm_n7318, gm_n7319, gm_n732, gm_n7320, gm_n7321, gm_n7322, gm_n7323, gm_n7324, gm_n7325, gm_n7326, gm_n7327, gm_n7328, gm_n7329, gm_n733, gm_n7330, gm_n7331, gm_n7332, gm_n7333, gm_n7334, gm_n7335, gm_n7336, gm_n7337, gm_n7338, gm_n7339, gm_n734, gm_n7340, gm_n7341, gm_n7342, gm_n7343, gm_n7344, gm_n7345, gm_n7346, gm_n7347, gm_n7348, gm_n7349, gm_n735, gm_n7350, gm_n7351, gm_n7352, gm_n7353, gm_n7354, gm_n7355, gm_n7356, gm_n7357, gm_n7358, gm_n7359, gm_n736, gm_n7360, gm_n7361, gm_n7362, gm_n7363, gm_n7364, gm_n7365, gm_n7366, gm_n7367, gm_n7368, gm_n7369, gm_n737, gm_n7370, gm_n7371, gm_n7372, gm_n7373, gm_n7374, gm_n7375, gm_n7376, gm_n7377, gm_n7378, gm_n7379, gm_n738, gm_n7380, gm_n7381, gm_n7382, gm_n7383, gm_n7384, gm_n7385, gm_n7386, gm_n7387, gm_n7388, gm_n7389, gm_n739, gm_n7390, gm_n7391, gm_n7392, gm_n7393, gm_n7394, gm_n7395, gm_n7396, gm_n7397, gm_n7398, gm_n7399, gm_n74, gm_n740, gm_n7400, gm_n7401, gm_n7402, gm_n7403, gm_n7404, gm_n7405, gm_n7406, gm_n7407, gm_n7408, gm_n7409, gm_n741, gm_n7410, gm_n7411, gm_n7412, gm_n7413, gm_n7414, gm_n7415, gm_n7416, gm_n7417, gm_n7418, gm_n7419, gm_n742, gm_n7420, gm_n7421, gm_n7422, gm_n7423, gm_n7424, gm_n7425, gm_n7426, gm_n7427, gm_n7428, gm_n7429, gm_n743, gm_n7430, gm_n7431, gm_n7432, gm_n7433, gm_n7434, gm_n7435, gm_n7436, gm_n7437, gm_n7438, gm_n7439, gm_n744, gm_n7440, gm_n7441, gm_n7442, gm_n7443, gm_n7444, gm_n7445, gm_n7446, gm_n7447, gm_n7448, gm_n7449, gm_n745, gm_n7450, gm_n7451, gm_n7452, gm_n7453, gm_n7454, gm_n7455, gm_n7456, gm_n7457, gm_n7458, gm_n7459, gm_n746, gm_n7460, gm_n7461, gm_n7462, gm_n7463, gm_n7464, gm_n7465, gm_n7466, gm_n7467, gm_n7468, gm_n7469, gm_n747, gm_n7470, gm_n7471, gm_n7472, gm_n7473, gm_n7474, gm_n7475, gm_n7476, gm_n7477, gm_n7478, gm_n7479, gm_n748, gm_n7480, gm_n7481, gm_n7482, gm_n7483, gm_n7484, gm_n7485, gm_n7486, gm_n7487, gm_n7488, gm_n7489, gm_n749, gm_n7490, gm_n7491, gm_n7492, gm_n7493, gm_n7494, gm_n7495, gm_n7496, gm_n75, gm_n750, gm_n751, gm_n752, gm_n753, gm_n754, gm_n755, gm_n756, gm_n757, gm_n758, gm_n76, gm_n760, gm_n761, gm_n762, gm_n763, gm_n764, gm_n765, gm_n766, gm_n767, gm_n768, gm_n769, gm_n77, gm_n770, gm_n771, gm_n772, gm_n773, gm_n774, gm_n775, gm_n776, gm_n777, gm_n778, gm_n779, gm_n78, gm_n780, gm_n781, gm_n782, gm_n783, gm_n784, gm_n785, gm_n786, gm_n787, gm_n788, gm_n789, gm_n79, gm_n790, gm_n791, gm_n792, gm_n793, gm_n794, gm_n795, gm_n796, gm_n797, gm_n798, gm_n799, gm_n80, gm_n800, gm_n801, gm_n802, gm_n803, gm_n804, gm_n805, gm_n806, gm_n807, gm_n808, gm_n809, gm_n81, gm_n810, gm_n811, gm_n812, gm_n813, gm_n814, gm_n815, gm_n816, gm_n817, gm_n818, gm_n819, gm_n82, gm_n820, gm_n821, gm_n822, gm_n823, gm_n824, gm_n825, gm_n826, gm_n827, gm_n828, gm_n829, gm_n83, gm_n830, gm_n831, gm_n832, gm_n833, gm_n834, gm_n835, gm_n836, gm_n837, gm_n838, gm_n839, gm_n84, gm_n840, gm_n841, gm_n842, gm_n843, gm_n844, gm_n845, gm_n846, gm_n847, gm_n848, gm_n849, gm_n85, gm_n850, gm_n851, gm_n852, gm_n853, gm_n854, gm_n855, gm_n856, gm_n857, gm_n858, gm_n859, gm_n86, gm_n860, gm_n861, gm_n862, gm_n863, gm_n864, gm_n865, gm_n866, gm_n867, gm_n868, gm_n869, gm_n87, gm_n870, gm_n871, gm_n872, gm_n873, gm_n874, gm_n875, gm_n876, gm_n877, gm_n878, gm_n879, gm_n88, gm_n880, gm_n881, gm_n882, gm_n883, gm_n884, gm_n885, gm_n886, gm_n887, gm_n888, gm_n889, gm_n89, gm_n890, gm_n891, gm_n892, gm_n893, gm_n894, gm_n895, gm_n896, gm_n897, gm_n898, gm_n899, gm_n90, gm_n900, gm_n901, gm_n902, gm_n903, gm_n904, gm_n905, gm_n906, gm_n907, gm_n908, gm_n909, gm_n91, gm_n910, gm_n911, gm_n912, gm_n913, gm_n914, gm_n915, gm_n916, gm_n917, gm_n918, gm_n919, gm_n92, gm_n920, gm_n921, gm_n922, gm_n923, gm_n924, gm_n925, gm_n926, gm_n927, gm_n928, gm_n929, gm_n93, gm_n930, gm_n931, gm_n932, gm_n933, gm_n934, gm_n935, gm_n936, gm_n937, gm_n938, gm_n939, gm_n94, gm_n940, gm_n941, gm_n942, gm_n943, gm_n944, gm_n945, gm_n946, gm_n947, gm_n948, gm_n949, gm_n95, gm_n950, gm_n951, gm_n952, gm_n953, gm_n954, gm_n955, gm_n956, gm_n957, gm_n958, gm_n959, gm_n96, gm_n960, gm_n961, gm_n962, gm_n963, gm_n964, gm_n965, gm_n966, gm_n967, gm_n968, gm_n969, gm_n97, gm_n970, gm_n971, gm_n972, gm_n973, gm_n974, gm_n975, gm_n976, gm_n977, gm_n978, gm_n979, gm_n98, gm_n980, gm_n981, gm_n982, gm_n983, gm_n984, gm_n985, gm_n986, gm_n987, gm_n988, gm_n989, gm_n99, gm_n990, gm_n991, gm_n992, gm_n993, gm_n994, gm_n995, gm_n996, gm_n997, gm_n998, gm_n999;
	wire t_5, t_6, t_8, t_2, t_0, t_7, t_3, t_9, t_1, t_4;
	not (gm_n55, in_17);
	not (gm_n56, in_19);
	nor (gm_n57, gm_n56, in_18, gm_n55);
	not (gm_n58, gm_n57);
	not (gm_n59, in_12);
	not (gm_n60, in_15);
	nor (gm_n61, gm_n60, in_14, in_13);
	not (gm_n62, in_9);
	not (gm_n63, in_11);
	nor (gm_n64, gm_n63, in_10, gm_n62);
	not (gm_n65, in_1);
	not (gm_n66, in_2);
	nand (gm_n67, gm_n66, gm_n65, in_0, in_4, in_3);
	nand (gm_n68, in_7, in_6, in_5);
	nor (gm_n69, gm_n68, gm_n67);
	nand (gm_n70, gm_n61, gm_n59, in_8, gm_n69, gm_n64);
	nor (gm_n71, in_21, in_20, in_16, gm_n70, gm_n58);
	not (gm_n72, in_21);
	not (gm_n73, in_16);
	nand (gm_n74, in_18, in_17, gm_n73);
	not (gm_n75, gm_n74);
	not (gm_n76, in_13);
	nor (gm_n77, gm_n60, in_14, gm_n76);
	not (gm_n78, in_10);
	nor (gm_n79, gm_n63, gm_n78, in_9);
	and (gm_n80, in_2, in_1, in_0, in_4, in_3);
	nor (gm_n81, in_7, in_6, in_5);
	and (gm_n82, gm_n81, gm_n80, in_8);
	and (gm_n83, gm_n79, gm_n77, gm_n59, gm_n82);
	nand (gm_n84, gm_n72, in_20, in_19, gm_n83, gm_n75);
	not (gm_n85, in_20);
	nor (gm_n86, gm_n72, gm_n85, in_19);
	not (gm_n87, gm_n86);
	nor (gm_n88, in_17, in_16, gm_n60);
	not (gm_n89, gm_n88);
	not (gm_n90, in_14);
	and (gm_n91, in_13, in_12, in_11);
	not (gm_n92, gm_n91);
	not (gm_n93, in_7);
	not (gm_n94, in_8);
	nand (gm_n95, in_9, gm_n94, gm_n93);
	not (gm_n96, in_3);
	not (gm_n97, in_5);
	and (gm_n98, in_2, in_1, in_0);
	nand (gm_n99, gm_n97, in_4, gm_n96, gm_n98, in_6);
	or (gm_n100, gm_n92, gm_n90, gm_n78, gm_n99, gm_n95);
	nor (gm_n101, gm_n89, gm_n87, in_18, gm_n100);
	nor (gm_n102, gm_n85, in_19, in_18);
	not (gm_n103, gm_n102);
	nor (gm_n104, in_16, gm_n60, in_14);
	not (gm_n105, gm_n104);
	nor (gm_n106, gm_n59, in_11, in_10);
	nor (gm_n107, gm_n94, in_7, in_6);
	not (gm_n108, in_4);
	and (gm_n109, in_1, in_0);
	and (gm_n110, gm_n108, in_3, gm_n66, gm_n109, gm_n97);
	nand (gm_n111, gm_n106, in_13, in_9, gm_n110, gm_n107);
	nor (gm_n112, gm_n103, in_21, gm_n55, gm_n111, gm_n105);
	and (gm_n113, in_19, in_18, in_17);
	nand (gm_n114, in_15, gm_n90, gm_n76);
	nand (gm_n115, gm_n63, gm_n78, in_9);
	or (gm_n116, gm_n93, in_6, gm_n97, gm_n67, gm_n94);
	nor (gm_n117, gm_n114, gm_n73, gm_n59, gm_n116, gm_n115);
	nand (gm_n118, gm_n113, in_21, in_20, gm_n117);
	not (gm_n119, in_18);
	nor (gm_n120, gm_n85, in_19, gm_n119);
	nand (gm_n121, gm_n73, gm_n60, in_14);
	not (gm_n122, gm_n121);
	nor (gm_n123, in_12, in_11, in_10);
	not (gm_n124, in_6);
	nor (gm_n125, in_8, gm_n93, gm_n124);
	and (gm_n126, in_4, gm_n96, gm_n66, gm_n109, gm_n97);
	and (gm_n127, gm_n123, in_13, gm_n62, gm_n126, gm_n125);
	nand (gm_n128, gm_n120, gm_n72, gm_n55, gm_n127, gm_n122);
	and (gm_n129, in_21, in_20, in_19);
	not (gm_n130, gm_n129);
	nor (gm_n131, gm_n55, gm_n73, in_15);
	not (gm_n132, gm_n131);
	nand (gm_n133, in_13, in_12, gm_n63);
	nor (gm_n134, in_2, in_1, in_0, in_4, in_3);
	nand (gm_n135, gm_n93, gm_n124, in_5, gm_n134, gm_n94);
	or (gm_n136, in_14, gm_n78, gm_n62, gm_n135, gm_n133);
	nor (gm_n137, gm_n132, gm_n130, gm_n119, gm_n136);
	nor (gm_n138, gm_n56, in_18, in_17);
	not (gm_n139, gm_n138);
	not (gm_n140, in_0);
	nand (gm_n141, gm_n66, in_1, gm_n140, in_4, in_3);
	nor (gm_n142, gm_n93, in_6, in_5, gm_n141, gm_n94);
	nor (gm_n143, gm_n63, in_10, in_9);
	nand (gm_n144, gm_n61, in_16, in_12, gm_n143, gm_n142);
	nor (gm_n145, gm_n139, gm_n72, in_20, gm_n144);
	nor (gm_n146, in_21, in_20, gm_n56);
	nand (gm_n147, gm_n76, in_12, in_11);
	or (gm_n148, in_9, in_8, in_7);
	nand (gm_n149, gm_n97, in_4, gm_n96, gm_n98, gm_n124);
	nor (gm_n150, gm_n147, gm_n90, gm_n78, gm_n149, gm_n148);
	nand (gm_n151, gm_n146, gm_n131, in_18, gm_n150);
	nand (gm_n152, gm_n60, gm_n90, in_13);
	nand (gm_n153, in_7, gm_n124, in_5, gm_n80, gm_n94);
	nor (gm_n154, in_11, in_10, in_9);
	not (gm_n155, gm_n154);
	nor (gm_n156, gm_n152, gm_n73, gm_n59, gm_n155, gm_n153);
	nand (gm_n157, gm_n113, gm_n72, in_20, gm_n156);
	nand (gm_n158, in_11, in_10, gm_n62);
	nand (gm_n159, in_14, gm_n76, in_12);
	nor (gm_n160, in_2, in_1, gm_n140, gm_n108, in_3);
	nand (gm_n161, gm_n160, gm_n81);
	or (gm_n162, gm_n158, in_15, gm_n94, gm_n161, gm_n159);
	nor (gm_n163, in_21, gm_n85, gm_n56, gm_n162, gm_n74);
	nor (gm_n164, in_21, gm_n85, gm_n56);
	not (gm_n165, gm_n164);
	nor (gm_n166, in_17, in_16, in_15);
	not (gm_n167, gm_n166);
	nand (gm_n168, gm_n90, gm_n76, in_12);
	and (gm_n169, in_2, in_1, in_0, in_3);
	and (gm_n170, gm_n124, in_5, gm_n108, gm_n169, gm_n93);
	nor (gm_n171, in_10, in_9, in_8);
	nand (gm_n172, gm_n171, gm_n170, in_11);
	nor (gm_n173, gm_n167, gm_n165, in_18, gm_n172, gm_n168);
	nor (gm_n174, in_20, gm_n56, in_18);
	nor (gm_n175, in_2, in_1, in_0, in_3);
	and (gm_n176, in_6, in_5, in_4, gm_n175, in_7);
	and (gm_n177, in_13, gm_n62, in_8, gm_n176, gm_n106);
	nand (gm_n178, gm_n122, in_21, gm_n55, gm_n177, gm_n174);
	nor (gm_n179, gm_n56, gm_n119, in_17);
	nand (gm_n180, in_7, gm_n124, gm_n97, gm_n80, gm_n94);
	nor (gm_n181, gm_n114, in_16, in_12, gm_n180, gm_n158);
	nand (gm_n182, gm_n179, in_21, gm_n85, gm_n181);
	not (gm_n183, gm_n120);
	nand (gm_n184, gm_n73, in_15, in_14);
	nor (gm_n185, in_12, in_11, gm_n78);
	nor (gm_n186, in_8, in_7, in_6);
	and (gm_n187, gm_n108, gm_n96, gm_n66, gm_n109, gm_n97);
	nand (gm_n188, gm_n185, gm_n76, gm_n62, gm_n187, gm_n186);
	nor (gm_n189, gm_n183, gm_n72, in_17, gm_n188, gm_n184);
	nand (gm_n190, in_11, gm_n78, in_9);
	nand (gm_n191, gm_n119, in_17, gm_n73);
	and (gm_n192, in_14, in_13, in_12);
	not (gm_n193, gm_n192);
	nand (gm_n194, gm_n93, gm_n124, in_5);
	nand (gm_n195, gm_n66, gm_n65, in_0, in_4, gm_n96);
	or (gm_n196, gm_n195, gm_n194, gm_n94);
	or (gm_n197, gm_n191, gm_n190, in_15, gm_n196, gm_n193);
	nor (gm_n198, gm_n72, gm_n85, in_19, gm_n197);
	nor (gm_n199, in_21, in_20, in_19);
	and (gm_n200, in_17, in_16, in_15);
	nand (gm_n201, in_2, in_1, gm_n140, gm_n108, gm_n96);
	nand (gm_n202, in_7, in_6, gm_n97);
	or (gm_n203, gm_n202, gm_n201, gm_n94);
	nor (gm_n204, gm_n90, in_10, gm_n62, gm_n203, gm_n147);
	nand (gm_n205, gm_n200, gm_n199, in_18, gm_n204);
	nor (gm_n206, in_20, in_19, gm_n119);
	nand (gm_n207, gm_n76, in_12, gm_n63);
	nand (gm_n208, in_5, in_4, gm_n96, gm_n98, gm_n124);
	nor (gm_n209, gm_n207, gm_n148, in_10, gm_n208);
	nand (gm_n210, gm_n122, gm_n72, gm_n55, gm_n209, gm_n206);
	not (gm_n211, gm_n146);
	nand (gm_n212, gm_n55, in_16, gm_n60);
	nand (gm_n213, gm_n63, in_10, in_9);
	not (gm_n214, gm_n213);
	nand (gm_n215, in_2, gm_n65, in_0, in_4, gm_n96);
	nor (gm_n216, in_7, in_6, in_5, gm_n215, gm_n94);
	nand (gm_n217, in_14, in_13, in_12, gm_n216, gm_n214);
	nor (gm_n218, gm_n212, gm_n211, gm_n119, gm_n217);
	not (gm_n219, gm_n113);
	nand (gm_n220, gm_n60, in_14, in_13);
	not (gm_n221, gm_n220);
	and (gm_n222, in_11, in_10, in_9);
	nand (gm_n223, gm_n66, in_1, gm_n140, gm_n108, in_3);
	nor (gm_n224, gm_n223, gm_n194, gm_n94);
	nand (gm_n225, gm_n221, in_16, in_12, gm_n224, gm_n222);
	nor (gm_n226, gm_n219, in_21, gm_n85, gm_n225);
	nand (gm_n227, in_15, gm_n90, in_13);
	nand (gm_n228, gm_n93, in_6, in_5);
	nand (gm_n229, in_2, in_1, gm_n140, gm_n108, in_3);
	or (gm_n230, gm_n229, gm_n228, in_8);
	nor (gm_n231, gm_n190, in_16, in_12, gm_n230, gm_n227);
	nand (gm_n232, gm_n179, gm_n72, gm_n85, gm_n231);
	nor (gm_n233, in_11, in_10, gm_n62);
	nand (gm_n234, in_2, in_1, gm_n140, in_4, in_3);
	nor (gm_n235, gm_n234, gm_n68, gm_n94);
	and (gm_n236, in_14, gm_n76, gm_n59, gm_n235, gm_n233);
	nand (gm_n237, gm_n166, gm_n164, gm_n119, gm_n236);
	nand (gm_n238, in_2, in_1, gm_n140, in_4, gm_n96);
	or (gm_n239, gm_n238, gm_n228);
	nand (gm_n240, gm_n78, gm_n62, in_8);
	or (gm_n241, gm_n193, gm_n60, gm_n63, gm_n240, gm_n239);
	nor (gm_n242, gm_n72, gm_n85, gm_n56, gm_n241, gm_n74);
	nor (gm_n243, gm_n72, in_20, in_19);
	not (gm_n244, gm_n243);
	nor (gm_n245, gm_n55, in_16, gm_n60);
	not (gm_n246, gm_n245);
	nand (gm_n247, in_9, in_8, gm_n93);
	nand (gm_n248, in_5, gm_n108, gm_n96, gm_n98, in_6);
	or (gm_n249, gm_n207, gm_n90, gm_n78, gm_n248, gm_n247);
	nor (gm_n250, gm_n246, gm_n244, in_18, gm_n249);
	or (gm_n251, gm_n229, gm_n68, gm_n94);
	nor (gm_n252, gm_n191, gm_n159, in_15, gm_n251, gm_n213);
	nand (gm_n253, gm_n72, gm_n85, gm_n56, gm_n252);
	nor (gm_n254, in_20, gm_n56, gm_n119);
	and (gm_n255, in_16, in_15, in_14);
	not (gm_n256, gm_n255);
	nand (gm_n257, in_12, in_11, gm_n78);
	nor (gm_n258, in_2, in_1, in_0);
	nand (gm_n259, in_5, gm_n108, in_3, gm_n258, gm_n124);
	nor (gm_n260, gm_n256, gm_n247, in_13, gm_n259, gm_n257);
	nand (gm_n261, gm_n254, in_21, in_17, gm_n260);
	not (gm_n262, gm_n179);
	nand (gm_n263, gm_n63, in_10, gm_n62);
	not (gm_n264, gm_n263);
	nor (gm_n265, gm_n228, gm_n223, gm_n94);
	nand (gm_n266, gm_n77, in_16, in_12, gm_n265, gm_n264);
	nor (gm_n267, gm_n262, in_21, gm_n85, gm_n266);
	nor (gm_n268, in_18, in_17, in_16);
	not (gm_n269, gm_n268);
	nand (gm_n270, in_6, in_5, gm_n108, gm_n169, in_7);
	nand (gm_n271, in_10, in_9, gm_n94);
	or (gm_n272, gm_n168, in_15, gm_n63, gm_n271, gm_n270);
	nor (gm_n273, in_21, in_20, in_19, gm_n272, gm_n269);
	not (gm_n274, gm_n222);
	and (gm_n275, in_15, in_14, in_13);
	not (gm_n276, gm_n275);
	nand (gm_n277, gm_n66, in_1, gm_n140, in_4, gm_n96);
	or (gm_n278, gm_n277, gm_n194, gm_n94);
	nor (gm_n279, gm_n274, in_16, in_12, gm_n278, gm_n276);
	nand (gm_n280, gm_n138, gm_n72, in_20, gm_n279);
	and (gm_n281, in_18, in_17, in_16);
	nand (gm_n282, gm_n93, in_6, gm_n97, gm_n134);
	nand (gm_n283, gm_n78, in_9, gm_n94);
	nor (gm_n284, gm_n193, in_15, gm_n63, gm_n283, gm_n282);
	nand (gm_n285, gm_n72, in_20, gm_n56, gm_n284, gm_n281);
	nand (gm_n286, in_5, in_4, in_3, gm_n258, gm_n124);
	nand (gm_n287, in_9, gm_n94, in_7);
	or (gm_n288, gm_n133, gm_n90, gm_n78, gm_n287, gm_n286);
	nor (gm_n289, gm_n246, gm_n130, in_18, gm_n288);
	nand (gm_n290, gm_n90, in_13, in_12);
	nor (gm_n291, gm_n93, in_6, gm_n97);
	nand (gm_n292, gm_n160, gm_n291, in_8);
	nand (gm_n293, gm_n119, gm_n55, in_16);
	or (gm_n294, gm_n290, gm_n213, in_15, gm_n293, gm_n292);
	nor (gm_n295, in_21, in_20, in_19, gm_n294);
	nor (gm_n296, in_19, gm_n119, in_17);
	nand (gm_n297, in_11, gm_n78, gm_n62);
	or (gm_n298, in_7, in_6, in_5, gm_n223, gm_n94);
	nor (gm_n299, gm_n114, in_16, in_12, gm_n298, gm_n297);
	nand (gm_n300, gm_n296, gm_n72, in_20, gm_n299);
	and (gm_n301, gm_n61, gm_n73, gm_n59, gm_n224, gm_n143);
	nand (gm_n302, gm_n296, gm_n72, gm_n85, gm_n301);
	nor (gm_n303, in_15, in_14, in_13);
	nor (gm_n304, gm_n93, in_6, in_5);
	nor (gm_n305, in_2, gm_n65, in_0, gm_n108, in_3);
	and (gm_n306, gm_n305, gm_n304, gm_n94);
	nand (gm_n307, gm_n214, gm_n73, in_12, gm_n306, gm_n303);
	nor (gm_n308, gm_n139, in_21, in_20, gm_n307);
	nand (gm_n309, gm_n81, gm_n80, in_8, gm_n222);
	nor (gm_n310, gm_n159, gm_n132, gm_n119, gm_n309, gm_n165);
	nor (gm_n311, in_20, in_19, in_18);
	not (gm_n312, gm_n311);
	nand (gm_n313, in_16, gm_n60, gm_n90);
	and (gm_n314, in_12, in_11, in_10);
	nor (gm_n315, in_1, in_0);
	and (gm_n316, gm_n108, in_3, in_2, gm_n315, gm_n97);
	nand (gm_n317, gm_n125, gm_n76, gm_n62, gm_n316, gm_n314);
	or (gm_n318, gm_n312, gm_n72, in_17, gm_n317, gm_n313);
	nand (gm_n319, in_15, in_14, gm_n76);
	or (gm_n320, gm_n234, gm_n228, gm_n94);
	nor (gm_n321, gm_n155, gm_n73, gm_n59, gm_n320, gm_n319);
	nand (gm_n322, gm_n113, gm_n72, in_20, gm_n321);
	nor (gm_n323, in_17, gm_n73, gm_n60);
	or (gm_n324, gm_n234, gm_n202, in_8);
	nor (gm_n325, in_14, gm_n76, gm_n59, gm_n324, gm_n274);
	nand (gm_n326, gm_n323, gm_n243, in_18, gm_n325);
	nor (gm_n327, gm_n85, gm_n56, in_18);
	nand (gm_n328, in_16, gm_n60, in_14);
	or (gm_n329, gm_n93, in_6, in_5, gm_n215, gm_n94);
	nor (gm_n330, gm_n257, in_13, in_9, gm_n329, gm_n328);
	nand (gm_n331, gm_n327, in_21, gm_n55, gm_n330);
	or (gm_n332, in_2, in_1, in_0);
	nor (gm_n333, gm_n97, gm_n108, gm_n96, gm_n332, in_6);
	nor (gm_n334, in_13, in_12, in_11);
	nor (gm_n335, in_9, gm_n94, in_7);
	and (gm_n336, gm_n334, gm_n333, gm_n78, gm_n335);
	nand (gm_n337, gm_n255, in_21, gm_n55, gm_n336, gm_n327);
	nand (gm_n338, gm_n326, gm_n322, gm_n318, gm_n337, gm_n331);
	nor (gm_n339, in_16, in_15, in_14);
	nor (gm_n340, in_12, gm_n63, in_10);
	and (gm_n341, in_8, in_7, in_6);
	and (gm_n342, gm_n316, gm_n76, gm_n62, gm_n341, gm_n340);
	nand (gm_n343, gm_n102, gm_n72, in_17, gm_n342, gm_n339);
	nand (gm_n344, in_8, gm_n93, in_6);
	nand (gm_n345, in_4, gm_n96, in_2, gm_n315, gm_n97);
	nor (gm_n346, gm_n257, in_13, in_9, gm_n345, gm_n344);
	nand (gm_n347, gm_n122, gm_n72, in_17, gm_n346, gm_n327);
	nor (gm_n348, in_21, gm_n85, in_19);
	nand (gm_n349, gm_n62, in_8, gm_n93);
	nand (gm_n350, in_5, gm_n108, in_3, gm_n258, in_6);
	nor (gm_n351, gm_n92, gm_n90, gm_n78, gm_n350, gm_n349);
	nand (gm_n352, gm_n348, gm_n200, in_18, gm_n351);
	nand (gm_n353, gm_n352, gm_n347, gm_n343);
	nand (gm_n354, gm_n60, in_14, gm_n76);
	or (gm_n355, gm_n141, gm_n68, gm_n94);
	nor (gm_n356, gm_n155, gm_n73, gm_n59, gm_n355, gm_n354);
	nand (gm_n357, gm_n138, in_21, in_20, gm_n356);
	not (gm_n358, gm_n123);
	nand (gm_n359, gm_n108, in_3, gm_n66, gm_n109, in_5);
	nor (gm_n360, gm_n358, in_13, gm_n62, gm_n359, gm_n344);
	nand (gm_n361, gm_n102, in_21, in_17, gm_n360, gm_n339);
	nand (gm_n362, gm_n76, gm_n59, in_11);
	nor (gm_n363, in_14, gm_n78, in_9, gm_n362, gm_n355);
	nand (gm_n364, gm_n129, gm_n88, gm_n119, gm_n363);
	nand (gm_n365, gm_n364, gm_n361, gm_n357);
	nor (gm_n366, gm_n338, gm_n310, gm_n308, gm_n365, gm_n353);
	nor (gm_n367, gm_n72, in_20, gm_n56);
	not (gm_n368, gm_n367);
	nand (gm_n369, in_13, gm_n59, in_11);
	nand (gm_n370, gm_n62, in_8, in_7);
	or (gm_n371, gm_n99, gm_n90, in_10, gm_n370, gm_n369);
	nor (gm_n372, gm_n368, gm_n132, in_18, gm_n371);
	and (gm_n373, in_20, in_19, in_18);
	not (gm_n374, gm_n373);
	nand (gm_n375, in_16, in_15, gm_n90);
	nand (gm_n376, gm_n97, gm_n108, gm_n96, gm_n98, gm_n124);
	or (gm_n377, gm_n358, gm_n95, in_13, gm_n376, gm_n375);
	nor (gm_n378, gm_n374, gm_n72, gm_n55, gm_n377);
	not (gm_n379, gm_n191);
	nand (gm_n380, gm_n379, gm_n154, gm_n60, gm_n265, gm_n192);
	nor (gm_n381, in_21, gm_n85, in_19, gm_n380);
	nor (gm_n382, gm_n381, gm_n378, gm_n372);
	nor (gm_n383, in_19, gm_n119, gm_n55);
	not (gm_n384, gm_n383);
	not (gm_n385, gm_n303);
	or (gm_n386, gm_n158, in_16, gm_n59, gm_n385, gm_n203);
	nor (gm_n387, gm_n384, gm_n72, gm_n85, gm_n386);
	not (gm_n388, gm_n254);
	nand (gm_n389, gm_n97, in_4, in_3, gm_n258, in_6);
	or (gm_n390, gm_n370, gm_n92, in_10, gm_n389);
	nor (gm_n391, gm_n184, gm_n72, in_17, gm_n390, gm_n388);
	not (gm_n392, gm_n159);
	nand (gm_n393, gm_n119, in_17, in_16);
	not (gm_n394, gm_n393);
	nand (gm_n395, gm_n222, gm_n392, gm_n60, gm_n394, gm_n265);
	nor (gm_n396, in_21, in_20, gm_n56, gm_n395);
	nor (gm_n397, gm_n396, gm_n391, gm_n387);
	nand (gm_n398, gm_n366, gm_n302, gm_n300, gm_n397, gm_n382);
	or (gm_n399, gm_n228, gm_n141, in_8);
	nor (gm_n400, in_14, in_10, in_9, gm_n399, gm_n362);
	nand (gm_n401, gm_n245, gm_n243, in_18, gm_n400);
	nor (gm_n402, in_12, gm_n63, gm_n78);
	and (gm_n403, gm_n126, in_13, in_9, gm_n402, gm_n186);
	nand (gm_n404, gm_n255, gm_n72, in_17, gm_n403, gm_n373);
	not (gm_n405, gm_n313);
	nand (gm_n406, gm_n59, in_11, gm_n78);
	nand (gm_n407, in_6, gm_n97, in_4, gm_n175, gm_n93);
	nor (gm_n408, gm_n76, in_9, in_8, gm_n407, gm_n406);
	nand (gm_n409, gm_n102, gm_n72, gm_n55, gm_n408, gm_n405);
	nand (gm_n410, gm_n409, gm_n404, gm_n401);
	nor (gm_n411, gm_n223, gm_n202, gm_n94);
	and (gm_n412, gm_n214, gm_n76, in_12, gm_n411);
	nand (gm_n413, gm_n174, gm_n72, gm_n55, gm_n412, gm_n255);
	nand (gm_n414, gm_n97, gm_n108, gm_n96, gm_n98, in_6);
	nor (gm_n415, gm_n287, gm_n358, in_13, gm_n414);
	nand (gm_n416, gm_n104, in_21, gm_n55, gm_n415, gm_n311);
	or (gm_n417, gm_n195, gm_n68);
	nor (gm_n418, gm_n297, in_12, in_8, gm_n417, gm_n220);
	nand (gm_n419, gm_n72, in_20, gm_n73, gm_n418, gm_n138);
	nand (gm_n420, gm_n419, gm_n416, gm_n413);
	nor (gm_n421, gm_n398, gm_n295, gm_n289, gm_n420, gm_n410);
	not (gm_n422, gm_n290);
	and (gm_n423, gm_n134, gm_n81, gm_n94);
	nand (gm_n424, gm_n268, gm_n233, in_15, gm_n423, gm_n422);
	nor (gm_n425, in_21, in_20, in_19, gm_n424);
	nor (gm_n426, gm_n66, in_1, gm_n140, gm_n108, gm_n96);
	and (gm_n427, in_7, in_6, gm_n97, gm_n426, gm_n94);
	nand (gm_n428, gm_n222, in_16, gm_n59, gm_n427, gm_n275);
	nor (gm_n429, gm_n262, in_21, in_20, gm_n428);
	not (gm_n430, gm_n186);
	not (gm_n431, gm_n314);
	nand (gm_n432, gm_n108, gm_n96, in_2, gm_n315, in_5);
	or (gm_n433, gm_n430, in_13, gm_n62, gm_n432, gm_n431);
	nor (gm_n434, gm_n388, gm_n72, in_17, gm_n433, gm_n313);
	nor (gm_n435, gm_n434, gm_n429, gm_n425);
	nor (gm_n436, gm_n55, in_16, in_15);
	not (gm_n437, gm_n436);
	nand (gm_n438, gm_n62, gm_n94, in_7);
	or (gm_n439, gm_n92, in_14, gm_n78, gm_n438, gm_n208);
	nor (gm_n440, gm_n437, gm_n165, gm_n119, gm_n439);
	not (gm_n441, gm_n174);
	nand (gm_n442, in_12, gm_n63, in_10);
	nand (gm_n443, gm_n94, gm_n93, in_6);
	or (gm_n444, gm_n359, in_13, in_9, gm_n443, gm_n442);
	nor (gm_n445, gm_n441, in_21, gm_n55, gm_n444, gm_n184);
	nor (gm_n446, gm_n229, gm_n68, gm_n94);
	nand (gm_n447, in_18, gm_n55, in_16);
	not (gm_n448, gm_n447);
	nor (gm_n449, in_14, in_13, in_12);
	nand (gm_n450, gm_n264, gm_n446, gm_n60, gm_n449, gm_n448);
	nor (gm_n451, in_21, in_20, in_19, gm_n450);
	nor (gm_n452, gm_n451, gm_n445, gm_n440);
	nand (gm_n453, gm_n421, gm_n285, gm_n280, gm_n452, gm_n435);
	nor (gm_n454, in_2, in_1, gm_n140, in_4, in_3);
	and (gm_n455, in_7, in_6, in_5, gm_n454);
	and (gm_n456, gm_n392, gm_n60, in_8, gm_n455, gm_n222);
	nand (gm_n457, in_21, in_20, gm_n56, gm_n456, gm_n75);
	or (gm_n458, gm_n229, gm_n194, in_8);
	nor (gm_n459, gm_n90, gm_n78, gm_n62, gm_n458, gm_n362);
	nand (gm_n460, gm_n323, gm_n129, in_18, gm_n459);
	nand (gm_n461, gm_n59, gm_n63, in_10);
	nand (gm_n462, gm_n108, gm_n96, in_2, gm_n315, gm_n97);
	nand (gm_n463, in_8, in_7, gm_n124);
	nor (gm_n464, gm_n461, in_13, in_9, gm_n463, gm_n462);
	nand (gm_n465, gm_n104, gm_n72, in_17, gm_n464, gm_n373);
	nand (gm_n466, gm_n465, gm_n460, gm_n457);
	nand (gm_n467, in_13, gm_n59, gm_n63);
	nand (gm_n468, gm_n454, gm_n304, gm_n94);
	nor (gm_n469, in_14, gm_n78, gm_n62, gm_n468, gm_n467);
	nand (gm_n470, gm_n166, gm_n86, in_18, gm_n469);
	nor (gm_n471, gm_n228, gm_n67, in_8);
	and (gm_n472, gm_n339, in_13, in_9, gm_n471, gm_n402);
	nand (gm_n473, gm_n102, gm_n72, gm_n55, gm_n472);
	nand (gm_n474, gm_n93, gm_n124, in_5, gm_n80, gm_n94);
	nor (gm_n475, gm_n115, in_16, in_12, gm_n474, gm_n319);
	nand (gm_n476, gm_n296, gm_n72, gm_n85, gm_n475);
	nand (gm_n477, gm_n476, gm_n473, gm_n470);
	nor (gm_n478, gm_n453, gm_n273, gm_n267, gm_n477, gm_n466);
	not (gm_n479, gm_n206);
	nand (gm_n480, gm_n59, in_11, in_10);
	nand (gm_n481, in_4, in_3, gm_n66, gm_n109, gm_n97);
	or (gm_n482, gm_n480, in_13, gm_n62, gm_n481, gm_n443);
	nor (gm_n483, gm_n184, gm_n72, in_17, gm_n482, gm_n479);
	not (gm_n484, gm_n168);
	nand (gm_n485, in_18, gm_n55, gm_n73);
	not (gm_n486, gm_n485);
	nor (gm_n487, gm_n215, gm_n202, in_8);
	nand (gm_n488, gm_n484, gm_n154, gm_n60, gm_n487, gm_n486);
	nor (gm_n489, in_21, gm_n85, gm_n56, gm_n488);
	and (gm_n490, in_9, in_8, in_7);
	not (gm_n491, gm_n490);
	or (gm_n492, gm_n92, gm_n90, gm_n78, gm_n491, gm_n248);
	nor (gm_n493, gm_n167, gm_n87, gm_n119, gm_n492);
	nor (gm_n494, gm_n493, gm_n489, gm_n483);
	nor (gm_n495, in_19, in_18, in_17);
	not (gm_n496, gm_n495);
	or (gm_n497, gm_n116, in_16, gm_n59, gm_n385, gm_n263);
	nor (gm_n498, gm_n496, gm_n72, gm_n85, gm_n497);
	or (gm_n499, gm_n93, in_6, in_5, gm_n229, gm_n94);
	or (gm_n500, gm_n159, gm_n190, in_15, gm_n499, gm_n447);
	nor (gm_n501, in_21, in_20, gm_n56, gm_n500);
	nand (gm_n502, gm_n94, in_7, gm_n124);
	nand (gm_n503, in_4, gm_n96, in_2, gm_n315, in_5);
	or (gm_n504, gm_n442, in_13, gm_n62, gm_n503, gm_n502);
	nor (gm_n505, gm_n256, gm_n72, gm_n55, gm_n504, gm_n312);
	nor (gm_n506, gm_n505, gm_n501, gm_n498);
	nand (gm_n507, gm_n478, gm_n261, gm_n253, gm_n506, gm_n494);
	or (gm_n508, gm_n201, gm_n68);
	nor (gm_n509, gm_n78, gm_n62, in_8, gm_n508, gm_n92);
	nand (gm_n510, gm_n131, gm_n119, gm_n90, gm_n509, gm_n367);
	or (gm_n511, gm_n223, gm_n202, in_8);
	nor (gm_n512, gm_n115, gm_n74, in_15, gm_n511, gm_n193);
	nand (gm_n513, gm_n72, in_20, in_19, gm_n512);
	nand (gm_n514, in_12, gm_n63, gm_n78);
	or (gm_n515, gm_n195, gm_n194, in_8);
	nor (gm_n516, gm_n514, in_13, gm_n62, gm_n515, gm_n375);
	nand (gm_n517, gm_n373, gm_n72, gm_n55, gm_n516);
	nand (gm_n518, gm_n517, gm_n513, gm_n510);
	nor (gm_n519, in_2, gm_n65, in_0, in_4, in_3);
	nand (gm_n520, in_7, in_6, in_5, gm_n519, gm_n94);
	nor (gm_n521, gm_n155, gm_n73, in_12, gm_n520, gm_n220);
	nand (gm_n522, gm_n495, in_21, in_20, gm_n521);
	nor (gm_n523, in_16, gm_n60, gm_n90);
	nor (gm_n524, gm_n257, in_13, gm_n62, gm_n345, gm_n344);
	nand (gm_n525, gm_n523, gm_n72, gm_n55, gm_n524, gm_n206);
	nand (gm_n526, in_5, in_4, in_3, gm_n258, in_6);
	nor (gm_n527, gm_n207, in_14, gm_n78, gm_n526, gm_n247);
	nand (gm_n528, gm_n131, gm_n86, in_18, gm_n527);
	nand (gm_n529, gm_n528, gm_n525, gm_n522);
	nor (gm_n530, gm_n507, gm_n250, gm_n242, gm_n529, gm_n518);
	not (gm_n531, gm_n348);
	nor (gm_n532, in_13, gm_n59, gm_n63);
	nand (gm_n533, gm_n107, gm_n78, in_9, gm_n532, gm_n126);
	nor (gm_n534, gm_n89, gm_n119, in_14, gm_n533, gm_n531);
	and (gm_n535, in_7, in_6, gm_n97, gm_n454, in_8);
	nand (gm_n536, gm_n339, in_13, gm_n62, gm_n535, gm_n340);
	nor (gm_n537, gm_n312, gm_n72, in_17, gm_n536);
	or (gm_n538, gm_n92, in_14, in_10, gm_n438, gm_n414);
	nor (gm_n539, gm_n437, gm_n165, in_18, gm_n538);
	nor (gm_n540, gm_n539, gm_n537, gm_n534);
	nand (gm_n541, in_10, in_9, in_8);
	or (gm_n542, gm_n159, gm_n60, in_11, gm_n541, gm_n270);
	nor (gm_n543, in_21, in_20, gm_n56, gm_n542, gm_n393);
	and (gm_n544, t_8, gm_n72);
	nor (gm_n545, in_14, gm_n76, in_12);
	nor (gm_n546, gm_n66, in_1, gm_n140, in_4, in_3);
	and (gm_n547, gm_n546, gm_n81, gm_n94);
	nand (gm_n548, gm_n233, gm_n75, in_15, gm_n547, gm_n545);
	nor (gm_n549, gm_n72, gm_n85, in_19, gm_n548);
	nor (gm_n550, gm_n549, gm_n544, gm_n543);
	nand (gm_n551, gm_n530, gm_n237, gm_n232, gm_n550, gm_n540);
	nand (gm_n552, gm_n160, gm_n304, gm_n94);
	nor (gm_n553, gm_n158, gm_n73, in_12, gm_n552, gm_n354);
	nand (gm_n554, gm_n138, in_21, gm_n85, gm_n553);
	not (gm_n555, gm_n541);
	and (gm_n556, in_6, gm_n97, in_4, gm_n175, in_7);
	and (gm_n557, gm_n422, gm_n60, gm_n63, gm_n556, gm_n555);
	nand (gm_n558, gm_n72, in_20, gm_n56, gm_n557, gm_n268);
	nor (gm_n559, gm_n92, in_14, gm_n78, gm_n350, gm_n148);
	nand (gm_n560, gm_n245, gm_n146, in_18, gm_n559);
	nand (gm_n561, gm_n560, gm_n558, gm_n554);
	or (gm_n562, in_7, in_6, in_5, gm_n215, in_8);
	nor (gm_n563, gm_n158, gm_n73, in_12, gm_n562, gm_n152);
	nand (gm_n564, gm_n138, gm_n72, gm_n85, gm_n563);
	nor (gm_n565, gm_n149, gm_n95, gm_n76, gm_n313, gm_n461);
	nand (gm_n566, gm_n373, gm_n72, gm_n55, gm_n565);
	nor (gm_n567, gm_n247, gm_n149, gm_n78, gm_n369);
	nand (gm_n568, gm_n255, in_21, in_17, gm_n567, gm_n327);
	nand (gm_n569, gm_n568, gm_n566, gm_n564);
	nor (gm_n570, gm_n551, gm_n226, gm_n218, gm_n569, gm_n561);
	not (gm_n571, gm_n354);
	nand (gm_n572, gm_n93, in_6, gm_n97);
	nor (gm_n573, gm_n274, in_12, in_8, gm_n572, gm_n234);
	and (gm_n574, gm_n119, gm_n55, in_16, gm_n573, gm_n571);
	and (gm_n575, gm_n574, gm_n243);
	and (gm_n576, gm_n124, gm_n97, gm_n108, gm_n169, gm_n93);
	nand (gm_n577, in_13, gm_n62, in_8, gm_n576, gm_n314);
	nor (gm_n578, gm_n103, gm_n72, in_17, gm_n577, gm_n375);
	nor (gm_n579, gm_n59, gm_n63, in_10);
	and (gm_n580, gm_n426, gm_n291);
	nand (gm_n581, in_13, gm_n62, in_8, gm_n580, gm_n579);
	nor (gm_n582, gm_n183, gm_n72, in_17, gm_n581, gm_n184);
	nor (gm_n583, gm_n582, gm_n578, gm_n575);
	nand (gm_n584, gm_n125, gm_n76, in_9, gm_n402, gm_n126);
	nor (gm_n585, gm_n388, in_21, gm_n55, gm_n584, gm_n328);
	nor (gm_n586, gm_n93, in_6, in_5, gm_n223, in_8);
	nand (gm_n587, gm_n106, gm_n76, in_9, gm_n586);
	nor (gm_n588, gm_n183, in_21, in_17, gm_n587, gm_n121);
	nand (gm_n589, in_5, in_4, gm_n96, gm_n98, in_6);
	or (gm_n590, gm_n247, in_11, in_10, gm_n589);
	or (gm_n591, gm_n193, in_19, gm_n60, gm_n590, gm_n269);
	nor (gm_n592, gm_n591, in_21, gm_n85);
	nor (gm_n593, gm_n592, gm_n588, gm_n585);
	nand (gm_n594, gm_n570, gm_n210, gm_n205, gm_n593, gm_n583);
	not (gm_n595, gm_n328);
	not (gm_n596, gm_n341);
	nand (gm_n597, in_4, in_3, gm_n66, gm_n109, in_5);
	nor (gm_n598, gm_n461, gm_n76, in_9, gm_n597, gm_n596);
	nand (gm_n599, gm_n327, gm_n72, gm_n55, gm_n598, gm_n595);
	nor (gm_n600, in_13, gm_n59, in_11);
	and (gm_n601, gm_n124, in_5, gm_n108, gm_n169, in_7);
	nor (gm_n602, in_10, gm_n62, gm_n94);
	and (gm_n603, gm_n600, gm_n131, gm_n90, gm_n602, gm_n601);
	nand (gm_n604, gm_n603, gm_n199, in_18);
	nand (gm_n605, in_10, gm_n62, in_8);
	nor (gm_n606, gm_n147, gm_n141, gm_n194, gm_n605);
	nand (gm_n607, gm_n104, gm_n72, gm_n55, gm_n606, gm_n120);
	nand (gm_n608, gm_n607, gm_n604, gm_n599);
	nand (gm_n609, in_8, gm_n93, gm_n124);
	nor (gm_n610, gm_n609, in_13, gm_n62, gm_n432, gm_n406);
	nand (gm_n611, gm_n122, gm_n72, gm_n55, gm_n610, gm_n206);
	and (gm_n612, gm_n93, gm_n124, in_5, gm_n134, in_8);
	and (gm_n613, gm_n545, gm_n143, gm_n60, gm_n612);
	nand (gm_n614, gm_n72, in_20, in_19, gm_n613, gm_n486);
	nor (gm_n615, gm_n93, in_6, in_5, gm_n201, in_8);
	and (gm_n616, gm_n77, gm_n73, gm_n59, gm_n615, gm_n154);
	nand (gm_n617, gm_n57, in_21, gm_n85, gm_n616);
	nand (gm_n618, gm_n617, gm_n614, gm_n611);
	nor (gm_n619, gm_n594, gm_n198, gm_n189, gm_n618, gm_n608);
	not (gm_n620, gm_n327);
	nand (gm_n621, in_4, in_3, in_2, gm_n315, in_5);
	or (gm_n622, gm_n461, gm_n76, gm_n62, gm_n621, gm_n443);
	nor (gm_n623, gm_n620, in_21, gm_n55, gm_n622, gm_n328);
	nor (gm_n624, gm_n76, gm_n59, in_11);
	nand (gm_n625, in_2, gm_n65, in_0, gm_n108, in_3);
	nor (gm_n626, gm_n625, gm_n194, gm_n94);
	nand (gm_n627, gm_n90, in_10, in_9, gm_n626, gm_n624);
	nor (gm_n628, gm_n368, gm_n212, gm_n119, gm_n627);
	or (gm_n629, gm_n256, gm_n148, gm_n76, gm_n286, gm_n257);
	nor (gm_n630, gm_n388, gm_n72, gm_n55, gm_n629);
	nor (gm_n631, gm_n630, gm_n628, gm_n623);
	or (gm_n632, gm_n93, in_6, gm_n97, gm_n223, in_8);
	nand (gm_n633, in_14, gm_n76, gm_n59);
	or (gm_n634, gm_n447, gm_n274, in_15, gm_n633, gm_n632);
	nor (gm_n635, in_21, in_20, in_19, gm_n634);
	nor (gm_n636, gm_n625, gm_n68, in_8);
	nand (gm_n637, gm_n264, in_16, in_12, gm_n636, gm_n303);
	nor (gm_n638, gm_n58, in_21, gm_n85, gm_n637);
	nand (gm_n639, gm_n90, gm_n78, gm_n62, gm_n626, gm_n334);
	nor (gm_n640, gm_n531, gm_n132, gm_n119, gm_n639);
	nor (gm_n641, gm_n640, gm_n638, gm_n635);
	nand (gm_n642, gm_n619, gm_n182, gm_n178, gm_n641, gm_n631);
	not (gm_n643, gm_n449);
	nor (gm_n644, gm_n239, gm_n60, gm_n63, gm_n643, gm_n240);
	nand (gm_n645, in_21, gm_n85, in_19, gm_n644, gm_n281);
	or (gm_n646, gm_n431, gm_n76, gm_n62, gm_n432, gm_n344);
	or (gm_n647, gm_n388, gm_n72, in_17, gm_n646, gm_n328);
	or (gm_n648, gm_n572, gm_n215, gm_n94);
	nor (gm_n649, gm_n297, gm_n73, in_12, gm_n648, gm_n152);
	nand (gm_n650, gm_n383, gm_n72, in_20, gm_n649);
	nand (gm_n651, gm_n650, gm_n647, gm_n645);
	nor (gm_n652, gm_n328, gm_n208, in_13, gm_n491, gm_n406);
	nand (gm_n653, gm_n102, in_21, gm_n55, gm_n652);
	nand (gm_n654, gm_n454, gm_n81, in_8);
	nor (gm_n655, in_14, in_13, gm_n59, gm_n654, gm_n158);
	nand (gm_n656, gm_n243, gm_n200, gm_n119, gm_n655);
	nand (gm_n657, gm_n93, in_6, gm_n97, gm_n426, in_8);
	nor (gm_n658, gm_n191, gm_n158, in_15, gm_n657, gm_n193);
	nand (gm_n659, in_21, in_20, gm_n56, gm_n658);
	nand (gm_n660, gm_n659, gm_n656, gm_n653);
	nor (gm_n661, gm_n642, gm_n173, gm_n163, gm_n660, gm_n651);
	not (gm_n662, gm_n339);
	nand (gm_n663, gm_n110, in_13, in_9, gm_n314, gm_n186);
	nor (gm_n664, gm_n662, in_21, gm_n55, gm_n663, gm_n374);
	or (gm_n665, gm_n461, in_13, in_9, gm_n503, gm_n443);
	nor (gm_n666, gm_n183, gm_n72, gm_n55, gm_n665, gm_n313);
	nand (gm_n667, gm_n94, in_7, in_6);
	or (gm_n668, gm_n667, in_13, gm_n62, gm_n481, gm_n431);
	nor (gm_n669, gm_n313, gm_n72, gm_n55, gm_n668, gm_n374);
	nor (gm_n670, gm_n669, gm_n666, gm_n664);
	nand (gm_n671, gm_n66, gm_n65, in_0, gm_n108, in_3);
	nor (gm_n672, gm_n93, in_6, gm_n97, gm_n671, in_8);
	nand (gm_n673, gm_n233, gm_n73, gm_n59, gm_n672, gm_n571);
	nor (gm_n674, gm_n262, gm_n72, gm_n85, gm_n673);
	nand (gm_n675, gm_n546, gm_n291, gm_n94);
	or (gm_n676, gm_n115, gm_n76, gm_n59, gm_n675, gm_n184);
	nor (gm_n677, gm_n103, gm_n72, gm_n55, gm_n676);
	nor (gm_n678, gm_n671, gm_n228, gm_n94);
	nand (gm_n679, gm_n233, in_16, in_12, gm_n678, gm_n275);
	nor (gm_n680, gm_n262, in_21, gm_n85, gm_n679);
	nor (gm_n681, gm_n680, gm_n677, gm_n674);
	nand (gm_n682, gm_n661, gm_n157, gm_n151, gm_n681, gm_n670);
	nor (gm_n683, gm_n95, in_14, in_10, gm_n389, gm_n207);
	nand (gm_n684, gm_n323, gm_n86, in_18, gm_n683);
	and (gm_n685, in_7, gm_n124, in_5, gm_n80, in_8);
	and (gm_n686, gm_n402, gm_n76, in_9, gm_n685);
	nand (gm_n687, gm_n122, in_21, gm_n55, gm_n686, gm_n373);
	nor (gm_n688, gm_n430, in_13, in_9, gm_n621, gm_n431);
	nand (gm_n689, gm_n174, in_21, gm_n55, gm_n688, gm_n255);
	nand (gm_n690, gm_n689, gm_n687, gm_n684);
	nor (gm_n691, gm_n609, in_13, in_9, gm_n462, gm_n257);
	nand (gm_n692, gm_n523, in_21, gm_n55, gm_n691, gm_n327);
	nor (gm_n693, gm_n358, gm_n76, gm_n62, gm_n481, gm_n443);
	nand (gm_n694, gm_n102, gm_n72, in_17, gm_n693, gm_n104);
	or (gm_n695, gm_n572, gm_n238, gm_n94);
	nor (gm_n696, gm_n190, in_16, gm_n59, gm_n695, gm_n276);
	nor (gm_n697, in_19, in_18, gm_n55);
	nand (gm_n698, gm_n696, gm_n72, gm_n85, gm_n697);
	nand (gm_n699, gm_n698, gm_n694, gm_n692);
	nor (gm_n700, gm_n682, gm_n145, gm_n137, gm_n699, gm_n690);
	or (gm_n701, gm_n115, in_16, in_12, gm_n648, gm_n354);
	nor (gm_n702, gm_n262, in_21, in_20, gm_n701);
	nand (gm_n703, gm_n64, in_16, gm_n59, gm_n571, gm_n142);
	nor (gm_n704, gm_n262, in_21, in_20, gm_n703);
	nand (gm_n705, in_7, in_6, gm_n97, gm_n519, in_8);
	or (gm_n706, gm_n227, gm_n73, in_12, gm_n705, gm_n213);
	nor (gm_n707, gm_n219, gm_n72, in_20, gm_n706);
	nor (gm_n708, gm_n707, gm_n704, gm_n702);
	or (gm_n709, gm_n480, gm_n76, in_9, gm_n503, gm_n443);
	nor (gm_n710, gm_n121, gm_n72, in_17, gm_n709, gm_n441);
	nand (gm_n711, gm_n123, in_13, in_9, gm_n471, gm_n405);
	nor (gm_n712, gm_n183, gm_n72, in_17, gm_n711);
	not (gm_n713, gm_n362);
	nor (gm_n714, gm_n228, gm_n215);
	nand (gm_n715, in_10, in_9, in_8, gm_n714, gm_n713);
	nor (gm_n716, gm_n211, gm_n119, in_14, gm_n715, gm_n246);
	nor (gm_n717, gm_n716, gm_n712, gm_n710);
	nand (gm_n718, gm_n700, gm_n128, gm_n118, gm_n717, gm_n708);
	nor (gm_n719, gm_n480, gm_n76, in_9, gm_n502, gm_n432);
	nand (gm_n720, gm_n255, in_21, in_17, gm_n719, gm_n327);
	not (gm_n721, gm_n438);
	nor (gm_n722, in_5, in_4, gm_n96, gm_n332, gm_n124);
	and (gm_n723, gm_n600, in_14, gm_n78, gm_n722, gm_n721);
	nand (gm_n724, gm_n243, gm_n88, gm_n119, gm_n723);
	nor (gm_n725, gm_n609, in_13, gm_n62, gm_n432, gm_n358);
	nand (gm_n726, gm_n102, in_21, in_17, gm_n725, gm_n104);
	nand (gm_n727, gm_n726, gm_n724, gm_n720);
	nor (gm_n728, gm_n514, gm_n76, gm_n62, gm_n481, gm_n443);
	nand (gm_n729, gm_n405, gm_n72, in_17, gm_n728, gm_n327);
	nand (gm_n730, in_7, gm_n124, gm_n97, gm_n134, gm_n94);
	nor (gm_n731, gm_n263, in_16, in_12, gm_n730, gm_n385);
	nand (gm_n732, gm_n179, gm_n72, gm_n85, gm_n731);
	nor (gm_n733, in_15, in_14, gm_n76);
	nor (gm_n734, gm_n202, gm_n141, gm_n94);
	and (gm_n735, gm_n214, gm_n733, gm_n59, gm_n734);
	nand (gm_n736, gm_n72, gm_n85, gm_n56, gm_n735, gm_n486);
	nand (gm_n737, gm_n736, gm_n732, gm_n729);
	nor (gm_n738, gm_n718, gm_n112, gm_n101, gm_n737, gm_n727);
	nor (gm_n739, gm_n609, gm_n76, gm_n62, gm_n621, gm_n442);
	nand (gm_n740, gm_n405, in_21, in_17, gm_n739, gm_n327);
	nor (gm_n741, gm_n227, in_16, gm_n59, gm_n153, gm_n115);
	nand (gm_n742, gm_n57, in_21, gm_n85, gm_n741);
	nand (gm_n743, in_4, gm_n96, gm_n66, gm_n109, in_5);
	nor (gm_n744, gm_n609, in_13, in_9, gm_n743, gm_n442);
	nand (gm_n745, gm_n102, gm_n72, in_17, gm_n744, gm_n339);
	nand (gm_n746, gm_n740, gm_n738, gm_n84, gm_n745, gm_n742);
	nor (gm_n747, gm_n376, in_14, in_10, gm_n467, gm_n438);
	nand (gm_n748, gm_n323, gm_n243, gm_n119, gm_n747);
	nor (gm_n749, gm_n286, in_14, gm_n78, gm_n491, gm_n467);
	nand (gm_n750, gm_n131, gm_n129, gm_n119, gm_n749);
	nor (gm_n751, gm_n93, in_6, gm_n97, gm_n201, gm_n94);
	and (gm_n752, gm_n233, in_16, in_12, gm_n751, gm_n571);
	nand (gm_n753, gm_n138, gm_n72, gm_n85, gm_n752);
	nand (gm_n754, gm_n753, gm_n750, gm_n748);
	not (gm_n755, gm_n240);
	and (gm_n756, gm_n124, gm_n97, in_4, gm_n175, in_7);
	nand (gm_n757, gm_n755, in_15, gm_n63, gm_n756, gm_n449);
	nor (gm_n758, in_21, gm_n85, gm_n56, gm_n757, gm_n191);
	nor (out_0, gm_n754, gm_n746, gm_n71, gm_n758);
	nand (gm_n760, in_14, in_13, gm_n59);
	nand (gm_n761, gm_n124, gm_n97, in_4, gm_n175, gm_n93);
	or (gm_n762, gm_n283, gm_n60, in_11, gm_n761, gm_n760);
	nor (gm_n763, in_21, gm_n85, in_19, gm_n762, gm_n293);
	nand (gm_n764, gm_n90, in_13, gm_n59);
	or (gm_n765, gm_n215, gm_n202, gm_n94);
	nor (gm_n766, gm_n269, gm_n158, in_15, gm_n765, gm_n764);
	nand (gm_n767, in_21, gm_n85, gm_n56, gm_n766);
	or (gm_n768, gm_n514, gm_n76, in_9, gm_n481, gm_n443);
	nor (gm_n769, gm_n441, in_21, gm_n55, gm_n768, gm_n313);
	nand (gm_n770, gm_n124, in_5, in_4, gm_n175, gm_n93);
	or (gm_n771, gm_n643, gm_n60, gm_n63, gm_n770, gm_n605);
	nor (gm_n772, gm_n72, gm_n85, in_19, gm_n771, gm_n269);
	and (gm_n773, gm_n107, gm_n76, in_9, gm_n402, gm_n110);
	nand (gm_n774, gm_n255, gm_n72, gm_n55, gm_n773, gm_n373);
	nand (gm_n775, in_5, gm_n108, gm_n96, gm_n98, gm_n124);
	nor (gm_n776, gm_n207, in_14, in_10, gm_n775, gm_n287);
	nand (gm_n777, gm_n200, gm_n86, in_18, gm_n776);
	nor (gm_n778, gm_n572, gm_n195, in_8);
	nand (gm_n779, gm_n268, gm_n143, in_15, gm_n778, gm_n422);
	nor (gm_n780, gm_n72, gm_n85, in_19, gm_n779);
	not (gm_n781, gm_n296);
	nand (gm_n782, gm_n61, in_16, gm_n59, gm_n778, gm_n264);
	nor (gm_n783, gm_n781, gm_n72, in_20, gm_n782);
	nand (gm_n784, in_14, gm_n76, in_12, gm_n626, gm_n64);
	or (gm_n785, gm_n132, gm_n130, in_18, gm_n784);
	nor (gm_n786, gm_n114, gm_n73, gm_n59, gm_n274, gm_n180);
	nand (gm_n787, gm_n113, in_21, gm_n85, gm_n786);
	not (gm_n788, gm_n442);
	nand (gm_n789, gm_n76, gm_n62, in_8, gm_n788, gm_n176);
	nor (gm_n790, gm_n105, in_21, gm_n55, gm_n789, gm_n388);
	nand (gm_n791, gm_n79, in_16, in_12, gm_n446, gm_n221);
	nor (gm_n792, gm_n384, in_21, in_20, gm_n791);
	nor (gm_n793, in_5, gm_n108, gm_n96, gm_n332, in_6);
	and (gm_n794, gm_n713, in_14, gm_n78, gm_n793, gm_n721);
	nand (gm_n795, gm_n367, gm_n200, gm_n119, gm_n794);
	nand (gm_n796, gm_n108, gm_n96, gm_n66, gm_n109, gm_n97);
	nor (gm_n797, gm_n796, gm_n76, in_9, gm_n480, gm_n344);
	nand (gm_n798, gm_n174, in_21, gm_n55, gm_n797, gm_n405);
	or (gm_n799, gm_n671, gm_n202, gm_n94);
	or (gm_n800, in_14, in_10, in_9, gm_n799, gm_n92);
	nor (gm_n801, gm_n437, gm_n165, in_18, gm_n800);
	nor (gm_n802, gm_n66, gm_n65, in_0, gm_n108, gm_n96);
	and (gm_n803, gm_n802, gm_n304, gm_n94);
	and (gm_n804, gm_n106, gm_n76, in_9, gm_n803);
	and (gm_n805, gm_n311, gm_n72, gm_n55, gm_n804, gm_n339);
	not (gm_n806, gm_n212);
	not (gm_n807, gm_n334);
	or (gm_n808, gm_n234, gm_n194, in_8);
	nor (gm_n809, in_14, gm_n78, in_9, gm_n808, gm_n807);
	nand (gm_n810, gm_n806, gm_n164, in_18, gm_n809);
	and (gm_n811, in_13, gm_n62, gm_n94, gm_n576, gm_n314);
	nand (gm_n812, gm_n255, gm_n72, in_17, gm_n811, gm_n373);
	or (gm_n813, gm_n431, gm_n184, gm_n76, gm_n370, gm_n350);
	nor (gm_n814, gm_n388, gm_n72, gm_n55, gm_n813);
	or (gm_n815, gm_n93, in_6, in_5, gm_n223, gm_n94);
	or (gm_n816, gm_n274, gm_n168, gm_n60, gm_n815, gm_n293);
	nor (gm_n817, in_21, in_20, in_19, gm_n816);
	nand (gm_n818, gm_n108, in_3, gm_n66, gm_n109, gm_n97);
	nor (gm_n819, gm_n818, gm_n76, gm_n62, gm_n430, gm_n461);
	nand (gm_n820, gm_n104, gm_n72, in_17, gm_n819, gm_n206);
	or (gm_n821, gm_n671, gm_n68, in_8);
	nor (gm_n822, gm_n168, gm_n158, in_15, gm_n821, gm_n485);
	nand (gm_n823, gm_n72, gm_n85, in_19, gm_n822);
	not (gm_n824, gm_n199);
	nor (gm_n825, gm_n93, in_6, in_5, gm_n67, in_8);
	nand (gm_n826, in_14, gm_n78, in_9, gm_n825, gm_n624);
	nor (gm_n827, gm_n824, gm_n167, gm_n119, gm_n826);
	not (gm_n828, gm_n95);
	nor (gm_n829, in_5, in_4, gm_n96, gm_n332, in_6);
	nand (gm_n830, gm_n828, gm_n90, gm_n78, gm_n829, gm_n532);
	nor (gm_n831, gm_n132, gm_n130, gm_n119, gm_n830);
	nand (gm_n832, gm_n546, gm_n291, in_8);
	nor (gm_n833, gm_n263, in_16, gm_n59, gm_n832, gm_n319);
	nand (gm_n834, gm_n57, in_21, in_20, gm_n833);
	nand (gm_n835, gm_n93, in_6, in_5, gm_n134, in_8);
	nor (gm_n836, gm_n213, gm_n73, in_12, gm_n835, gm_n354);
	nand (gm_n837, gm_n495, in_21, in_20, gm_n836);
	nor (gm_n838, gm_n215, gm_n68, gm_n94);
	nand (gm_n839, gm_n713, gm_n78, gm_n62, gm_n838);
	nor (gm_n840, gm_n441, in_21, gm_n55, gm_n839, gm_n313);
	not (gm_n841, gm_n200);
	nand (gm_n842, in_6, in_5, in_4, gm_n175, gm_n93);
	or (gm_n843, gm_n207, gm_n841, gm_n90, gm_n842, gm_n240);
	nor (gm_n844, gm_n843, gm_n87, in_18);
	nor (gm_n845, gm_n95, in_14, gm_n78, gm_n526, gm_n362);
	nand (gm_n846, gm_n199, gm_n88, gm_n119, gm_n845);
	nor (gm_n847, gm_n430, gm_n76, in_9, gm_n743, gm_n431);
	nand (gm_n848, gm_n327, in_21, gm_n55, gm_n847, gm_n595);
	or (gm_n849, gm_n234, gm_n202, gm_n94);
	nor (gm_n850, gm_n274, gm_n74, in_15, gm_n849, gm_n760);
	nand (gm_n851, in_21, in_20, gm_n56, gm_n850);
	nor (gm_n852, gm_n329, gm_n76, in_9, gm_n480);
	nand (gm_n853, gm_n104, gm_n72, in_17, gm_n852, gm_n174);
	nand (gm_n854, gm_n848, gm_n846, t_0, gm_n853, gm_n851);
	nand (gm_n855, gm_n81, gm_n80, gm_n94);
	nor (gm_n856, gm_n227, in_16, gm_n59, gm_n855, gm_n263);
	nand (gm_n857, gm_n57, gm_n72, in_20, gm_n856);
	nor (gm_n858, gm_n148, gm_n90, in_10, gm_n369, gm_n248);
	nand (gm_n859, gm_n245, gm_n243, in_18, gm_n858);
	or (gm_n860, in_7, in_6, in_5, gm_n671, in_8);
	nor (gm_n861, gm_n293, gm_n155, gm_n60, gm_n860, gm_n760);
	nand (gm_n862, in_21, in_20, in_19, gm_n861);
	nand (gm_n863, gm_n862, gm_n859, gm_n857);
	nor (gm_n864, gm_n376, in_14, gm_n78, gm_n467, gm_n438);
	nand (gm_n865, gm_n243, gm_n806, in_18, gm_n864);
	not (gm_n866, gm_n316);
	nor (gm_n867, gm_n667, in_13, gm_n62, gm_n442, gm_n866);
	nand (gm_n868, gm_n254, in_21, in_17, gm_n867, gm_n405);
	not (gm_n869, gm_n760);
	nor (gm_n870, gm_n572, gm_n277, in_8);
	and (gm_n871, gm_n394, gm_n64, in_15, gm_n870, gm_n869);
	nand (gm_n872, in_21, in_20, in_19, gm_n871);
	nand (gm_n873, gm_n872, gm_n868, gm_n865);
	nor (gm_n874, gm_n854, gm_n844, gm_n840, gm_n873, gm_n863);
	and (gm_n875, gm_n519, gm_n291, in_8);
	nand (gm_n876, gm_n123, in_13, gm_n62, gm_n875);
	nor (gm_n877, gm_n183, gm_n72, gm_n55, gm_n876, gm_n328);
	nand (gm_n878, in_14, gm_n78, in_9, gm_n334, gm_n216);
	nor (gm_n879, gm_n841, gm_n824, gm_n119, gm_n878);
	nor (gm_n880, gm_n201, gm_n194, gm_n94);
	nand (gm_n881, gm_n64, in_16, in_12, gm_n880, gm_n303);
	nor (gm_n882, gm_n262, gm_n72, gm_n85, gm_n881);
	nor (gm_n883, gm_n882, gm_n879, gm_n877);
	and (gm_n884, gm_n93, gm_n124, in_5, gm_n80, in_8);
	nand (gm_n885, gm_n579, gm_n76, in_9, gm_n884);
	nor (gm_n886, gm_n103, in_21, in_17, gm_n885, gm_n375);
	nand (gm_n887, gm_n93, in_6, in_5, gm_n80, in_8);
	or (gm_n888, gm_n213, gm_n73, in_12, gm_n887, gm_n354);
	nor (gm_n889, gm_n384, in_21, in_20, gm_n888);
	or (gm_n890, gm_n227, gm_n73, gm_n59, gm_n196, gm_n115);
	nor (gm_n891, gm_n58, in_21, in_20, gm_n890);
	nor (gm_n892, gm_n891, gm_n889, gm_n886);
	nand (gm_n893, gm_n874, gm_n837, gm_n834, gm_n892, gm_n883);
	nor (gm_n894, gm_n148, gm_n90, gm_n78, gm_n467, gm_n350);
	nand (gm_n895, gm_n436, gm_n86, in_18, gm_n894);
	nor (gm_n896, gm_n105, in_13, in_9, gm_n468, gm_n461);
	nand (gm_n897, gm_n174, in_21, in_17, gm_n896);
	and (gm_n898, in_13, in_12, gm_n94, gm_n264, gm_n69);
	nand (gm_n899, gm_n122, in_21, in_17, gm_n898, gm_n206);
	nand (gm_n900, gm_n899, gm_n897, gm_n895);
	nor (gm_n901, gm_n818, in_13, gm_n62, gm_n442, gm_n667);
	nand (gm_n902, gm_n339, gm_n72, in_17, gm_n901, gm_n373);
	nor (gm_n903, gm_n147, gm_n90, gm_n78, gm_n414, gm_n370);
	nand (gm_n904, gm_n806, gm_n164, in_18, gm_n903);
	nor (gm_n905, gm_n461, gm_n76, gm_n62, gm_n743, gm_n463);
	nand (gm_n906, gm_n254, gm_n72, gm_n55, gm_n905, gm_n405);
	nand (gm_n907, gm_n906, gm_n904, gm_n902);
	nor (gm_n908, gm_n893, gm_n831, gm_n827, gm_n907, gm_n900);
	nand (gm_n909, gm_n124, in_5, gm_n108, gm_n169, gm_n93);
	or (gm_n910, gm_n909, gm_n92, gm_n90, gm_n605);
	nor (gm_n911, gm_n246, gm_n87, in_18, gm_n910);
	not (gm_n912, gm_n697);
	or (gm_n913, gm_n141, gm_n194);
	or (gm_n914, gm_n155, in_12, in_8, gm_n913, gm_n385);
	nor (gm_n915, in_21, in_20, in_16, gm_n914, gm_n912);
	nor (gm_n916, gm_n447, gm_n297, in_15, gm_n887, gm_n760);
	and (gm_n917, gm_n72, in_20, in_19, gm_n916);
	nor (gm_n918, gm_n917, gm_n915, gm_n911);
	and (gm_n919, gm_n93, in_6, in_5, gm_n134, gm_n94);
	nand (gm_n920, gm_n222, gm_n379, gm_n60, gm_n919, gm_n422);
	nor (gm_n921, gm_n72, gm_n85, gm_n56, gm_n920);
	or (gm_n922, gm_n514, gm_n76, in_9, gm_n503, gm_n502);
	nor (gm_n923, gm_n388, gm_n72, gm_n55, gm_n922, gm_n256);
	or (gm_n924, gm_n297, in_16, gm_n59, gm_n520, gm_n152);
	nor (gm_n925, gm_n384, in_21, in_20, gm_n924);
	nor (gm_n926, gm_n925, gm_n923, gm_n921);
	nand (gm_n927, gm_n908, gm_n823, gm_n820, gm_n926, gm_n918);
	nor (gm_n928, gm_n461, in_13, in_9, gm_n503, gm_n344);
	nand (gm_n929, gm_n102, gm_n72, in_17, gm_n928, gm_n405);
	nor (gm_n930, gm_n227, in_16, gm_n59, gm_n860, gm_n297);
	nand (gm_n931, gm_n697, gm_n72, gm_n85, gm_n930);
	or (gm_n932, gm_n572, gm_n223, gm_n94);
	nor (gm_n933, in_14, gm_n78, gm_n62, gm_n932, gm_n207);
	nand (gm_n934, gm_n200, gm_n164, gm_n119, gm_n933);
	nand (gm_n935, gm_n934, gm_n931, gm_n929);
	nor (gm_n936, gm_n229, gm_n202, in_8);
	and (gm_n937, gm_n61, in_16, gm_n59, gm_n936, gm_n222);
	nand (gm_n938, gm_n697, in_21, in_20, gm_n937);
	or (gm_n939, gm_n238, gm_n68);
	nor (gm_n940, gm_n227, gm_n59, in_8, gm_n939, gm_n263);
	nand (gm_n941, gm_n72, gm_n85, in_16, gm_n940, gm_n57);
	nor (gm_n942, gm_n149, gm_n90, in_10, gm_n491, gm_n807);
	nand (gm_n943, gm_n243, gm_n88, in_18, gm_n942);
	nand (gm_n944, gm_n943, gm_n941, gm_n938);
	nor (gm_n945, gm_n927, gm_n817, gm_n814, gm_n944, gm_n935);
	nor (gm_n946, gm_n93, in_6, in_5, gm_n67, gm_n94);
	nand (gm_n947, gm_n185, gm_n76, in_9, gm_n946, gm_n339);
	nor (gm_n948, gm_n312, gm_n72, in_17, gm_n947);
	not (gm_n949, gm_n319);
	and (gm_n950, gm_n93, gm_n124, in_5, gm_n546, gm_n94);
	nand (gm_n951, gm_n949, gm_n79, in_12, gm_n950);
	nor (gm_n952, in_21, in_20, gm_n56, gm_n951, gm_n393);
	nor (gm_n953, gm_n572, gm_n201, gm_n94);
	nand (gm_n954, gm_n264, in_16, gm_n59, gm_n953, gm_n571);
	nor (gm_n955, gm_n496, gm_n72, gm_n85, gm_n954);
	nor (gm_n956, gm_n955, gm_n952, gm_n948);
	and (gm_n957, gm_n304, gm_n79, in_8, gm_n422, gm_n160);
	nand (gm_n958, gm_n72, in_19, gm_n60, gm_n957, gm_n448);
	nor (gm_n959, gm_n958, in_20);
	or (gm_n960, gm_n514, gm_n76, in_9, gm_n462, gm_n344);
	nor (gm_n961, gm_n103, gm_n72, in_17, gm_n960, gm_n256);
	and (gm_n962, in_7, in_6, gm_n97, gm_n454, gm_n94);
	nand (gm_n963, gm_n255, gm_n76, gm_n62, gm_n962, gm_n314);
	nor (gm_n964, gm_n388, gm_n72, gm_n55, gm_n963);
	nor (gm_n965, gm_n964, gm_n961, gm_n959);
	nand (gm_n966, gm_n945, gm_n812, gm_n810, gm_n965, gm_n956);
	nor (gm_n967, gm_n605, in_15, gm_n63, gm_n761, gm_n633);
	nand (gm_n968, in_21, in_20, in_19, gm_n967, gm_n448);
	and (gm_n969, gm_n93, in_6, gm_n97, gm_n454, in_8);
	and (gm_n970, gm_n64, gm_n76, in_12, gm_n969, gm_n339);
	nand (gm_n971, gm_n254, in_21, gm_n55, gm_n970);
	nor (gm_n972, gm_n90, gm_n78, gm_n62, gm_n807, gm_n320);
	nand (gm_n973, gm_n146, gm_n131, in_18, gm_n972);
	nand (gm_n974, gm_n973, gm_n971, gm_n968);
	nor (gm_n975, gm_n213, gm_n73, gm_n59, gm_n648, gm_n276);
	nand (gm_n976, gm_n179, gm_n72, gm_n85, gm_n975);
	not (gm_n977, gm_n171);
	nor (gm_n978, gm_n977, gm_n133, gm_n90, gm_n572, gm_n215);
	nand (gm_n979, gm_n367, gm_n323, gm_n119, gm_n978);
	not (gm_n980, gm_n602);
	nand (gm_n981, in_6, in_5, gm_n108, gm_n169, gm_n93);
	nor (gm_n982, gm_n980, gm_n60, in_11, gm_n981, gm_n633);
	nand (gm_n983, in_21, gm_n85, in_19, gm_n982, gm_n379);
	nand (gm_n984, gm_n983, gm_n979, gm_n976);
	nor (gm_n985, gm_n966, gm_n805, gm_n801, gm_n984, gm_n974);
	nor (gm_n986, gm_n155, gm_n76, in_12, gm_n695);
	and (gm_n987, gm_n120, gm_n72, in_17, gm_n986, gm_n523);
	nand (gm_n988, gm_n108, in_3, in_2, gm_n315, in_5);
	or (gm_n989, gm_n406, in_13, gm_n62, gm_n988, gm_n344);
	nor (gm_n990, gm_n183, in_21, in_17, gm_n989, gm_n121);
	and (gm_n991, in_7, in_6, gm_n97, gm_n134, in_8);
	nand (gm_n992, gm_n392, gm_n79, in_15, gm_n991, gm_n448);
	nor (gm_n993, in_21, gm_n85, gm_n56, gm_n992);
	nor (gm_n994, gm_n993, gm_n990, gm_n987);
	nor (gm_n995, gm_n62, gm_n94, in_7);
	nand (gm_n996, gm_n91, gm_n90, in_10, gm_n793, gm_n995);
	nor (gm_n997, gm_n531, gm_n167, gm_n119, gm_n996);
	and (gm_n998, gm_n802, gm_n291, in_8);
	nand (gm_n999, in_14, in_10, in_9, gm_n998, gm_n91);
	nor (gm_n1000, gm_n531, gm_n246, gm_n119, gm_n999);
	nor (gm_n1001, gm_n234, gm_n68, in_8);
	nand (gm_n1002, gm_n90, in_10, in_9, gm_n1001, gm_n624);
	nor (gm_n1003, gm_n246, gm_n824, gm_n119, gm_n1002);
	nor (gm_n1004, gm_n1003, gm_n1000, gm_n997);
	nand (gm_n1005, gm_n985, gm_n798, gm_n795, gm_n1004, gm_n994);
	or (gm_n1006, gm_n93, in_6, gm_n97, gm_n671, in_8);
	nor (gm_n1007, gm_n90, gm_n78, gm_n62, gm_n1006, gm_n369);
	nand (gm_n1008, gm_n243, gm_n200, in_18, gm_n1007);
	and (gm_n1009, gm_n61, in_16, gm_n59, gm_n685, gm_n79);
	nand (gm_n1010, gm_n57, in_21, gm_n85, gm_n1009);
	nor (gm_n1011, gm_n76, in_12, gm_n63);
	nor (gm_n1012, gm_n572, gm_n238, in_8);
	and (gm_n1013, gm_n90, gm_n78, gm_n62, gm_n1012, gm_n1011);
	nand (gm_n1014, gm_n323, gm_n164, gm_n119, gm_n1013);
	nand (gm_n1015, gm_n1014, gm_n1010, gm_n1008);
	nand (gm_n1016, in_7, in_6, in_5, gm_n80, gm_n94);
	nor (gm_n1017, gm_n263, gm_n168, gm_n60, gm_n1016, gm_n447);
	nand (gm_n1018, gm_n72, in_20, gm_n56, gm_n1017);
	nand (gm_n1019, in_10, in_9, gm_n94, gm_n160, gm_n81);
	nor (gm_n1020, gm_n1019, gm_n369, gm_n90);
	nand (gm_n1021, gm_n367, gm_n88, gm_n119, gm_n1020);
	nor (gm_n1022, gm_n344, in_13, in_9, gm_n462, gm_n480);
	nand (gm_n1023, gm_n311, gm_n72, gm_n55, gm_n1022, gm_n595);
	nand (gm_n1024, gm_n1023, gm_n1021, gm_n1018);
	nor (gm_n1025, gm_n1005, gm_n792, gm_n790, gm_n1024, gm_n1015);
	or (gm_n1026, in_14, in_10, in_9, gm_n815, gm_n369);
	nor (gm_n1027, gm_n824, gm_n132, gm_n119, gm_n1026);
	or (gm_n1028, gm_n133, in_14, gm_n78, gm_n389, gm_n349);
	nor (gm_n1029, gm_n437, gm_n130, gm_n119, gm_n1028);
	nor (gm_n1030, gm_n277, gm_n202, in_8);
	nand (gm_n1031, in_14, gm_n78, in_9, gm_n1030, gm_n532);
	nor (gm_n1032, gm_n244, gm_n212, gm_n119, gm_n1031);
	nor (gm_n1033, gm_n1032, gm_n1029, gm_n1027);
	nor (gm_n1034, gm_n430, in_13, in_9, gm_n503, gm_n257);
	and (gm_n1035, gm_n174, in_21, in_17, gm_n1034, gm_n405);
	or (gm_n1036, gm_n92, in_10, in_9, gm_n503, gm_n463);
	nor (gm_n1037, gm_n89, gm_n119, in_14, gm_n1036, gm_n244);
	or (gm_n1038, gm_n274, in_16, gm_n59, gm_n399, gm_n385);
	nor (gm_n1039, gm_n139, gm_n72, in_20, gm_n1038);
	nor (gm_n1040, gm_n1039, gm_n1037, gm_n1035);
	nand (gm_n1041, gm_n1025, gm_n787, gm_n785, gm_n1040, gm_n1033);
	and (gm_n1042, gm_n595, in_13, gm_n62, gm_n535, gm_n402);
	nand (gm_n1043, gm_n120, in_21, in_17, gm_n1042);
	nor (gm_n1044, gm_n480, in_13, in_9, gm_n443, gm_n432);
	nand (gm_n1045, gm_n255, gm_n72, in_17, gm_n1044, gm_n373);
	nor (gm_n1046, gm_n514, in_13, in_9, gm_n432, gm_n609);
	nand (gm_n1047, gm_n523, gm_n72, in_17, gm_n1046, gm_n373);
	nand (gm_n1048, gm_n1047, gm_n1045, gm_n1043);
	nor (gm_n1049, in_8, in_7, gm_n124);
	and (gm_n1050, gm_n185, in_13, gm_n62, gm_n1049, gm_n316);
	nand (gm_n1051, gm_n102, in_21, in_17, gm_n1050, gm_n405);
	or (gm_n1052, gm_n277, gm_n68, gm_n94);
	nor (gm_n1053, gm_n290, gm_n213, gm_n60, gm_n1052, gm_n293);
	nand (gm_n1054, gm_n72, in_20, in_19, gm_n1053);
	and (gm_n1055, gm_n90, in_13, gm_n59, gm_n838, gm_n79);
	nand (gm_n1056, gm_n164, gm_n131, gm_n119, gm_n1055);
	nand (gm_n1057, gm_n1056, gm_n1054, gm_n1051);
	nor (gm_n1058, gm_n1041, gm_n783, gm_n780, gm_n1057, gm_n1048);
	nand (gm_n1059, gm_n104, in_13, in_9, gm_n946, gm_n106);
	nor (gm_n1060, gm_n103, gm_n72, in_17, gm_n1059);
	or (gm_n1061, gm_n207, in_14, in_10, gm_n775, gm_n491);
	nor (gm_n1062, gm_n437, gm_n244, gm_n119, gm_n1061);
	nand (gm_n1063, gm_n110, in_13, in_9, gm_n1049, gm_n579);
	nor (gm_n1064, gm_n256, in_21, in_17, gm_n1063, gm_n374);
	nor (gm_n1065, gm_n1064, gm_n1062, gm_n1060);
	nor (gm_n1066, gm_n256, in_21, gm_n55, gm_n960, gm_n312);
	nor (gm_n1067, gm_n66, in_1, gm_n140, in_4, gm_n96);
	and (gm_n1068, gm_n171, gm_n304, gm_n63, gm_n1067);
	and (gm_n1069, gm_n1068, in_13, in_12);
	and (gm_n1070, gm_n174, in_21, in_17, gm_n1069, gm_n523);
	and (gm_n1071, in_7, in_6, in_5, gm_n546, in_8);
	nand (gm_n1072, gm_n154, in_16, in_12, gm_n1071, gm_n221);
	nor (gm_n1073, gm_n262, gm_n72, in_20, gm_n1072);
	nor (gm_n1074, gm_n1073, gm_n1070, gm_n1066);
	nand (gm_n1075, gm_n1058, gm_n777, gm_n774, gm_n1074, gm_n1065);
	not (gm_n1076, gm_n375);
	and (gm_n1077, gm_n106, gm_n76, gm_n62, gm_n316, gm_n186);
	nand (gm_n1078, gm_n254, gm_n72, in_17, gm_n1077, gm_n1076);
	nor (gm_n1079, gm_n201, gm_n194, in_8);
	and (gm_n1080, gm_n624, in_10, gm_n62, gm_n1079, gm_n523);
	nand (gm_n1081, gm_n327, in_21, in_17, gm_n1080);
	nor (gm_n1082, gm_n406, gm_n328, in_13, gm_n775, gm_n370);
	nand (gm_n1083, gm_n120, in_21, in_17, gm_n1082);
	nand (gm_n1084, gm_n1083, gm_n1081, gm_n1078);
	nor (gm_n1085, gm_n461, in_13, gm_n62, gm_n481, gm_n443);
	nand (gm_n1086, gm_n120, gm_n72, in_17, gm_n1085, gm_n339);
	and (gm_n1087, gm_n104, in_13, gm_n62, gm_n306, gm_n106);
	nand (gm_n1088, gm_n254, gm_n72, gm_n55, gm_n1087);
	nor (gm_n1089, gm_n78, in_9, in_8, gm_n467, gm_n270);
	nand (gm_n1090, gm_n199, gm_n119, in_14, gm_n1089, gm_n436);
	nand (gm_n1091, gm_n1090, gm_n1088, gm_n1086);
	nor (gm_n1092, gm_n1075, gm_n772, gm_n769, gm_n1091, gm_n1084);
	nor (gm_n1093, gm_n90, in_10, gm_n62, gm_n1016, gm_n369);
	nand (gm_n1094, gm_n348, gm_n200, gm_n119, gm_n1093);
	nor (gm_n1095, gm_n625, gm_n228, gm_n94);
	and (gm_n1096, gm_n281, gm_n64, in_15, gm_n1095, gm_n449);
	nand (gm_n1097, gm_n72, in_20, in_19, gm_n1096);
	nor (gm_n1098, gm_n406, gm_n76, gm_n62, gm_n597, gm_n502);
	nand (gm_n1099, gm_n327, in_21, gm_n55, gm_n1098, gm_n595);
	nand (gm_n1100, gm_n1094, gm_n1092, gm_n767, gm_n1099, gm_n1097);
	not (gm_n1101, gm_n293);
	nor (gm_n1102, gm_n643, in_15, in_11, gm_n842, gm_n980);
	nand (gm_n1103, gm_n72, in_20, in_19, gm_n1102, gm_n1101);
	nor (gm_n1104, gm_n115, in_12, gm_n94, gm_n939, gm_n354);
	nand (gm_n1105, gm_n72, in_20, gm_n73, gm_n1104, gm_n179);
	and (gm_n1106, gm_n600, gm_n90, in_10, gm_n793, gm_n995);
	nand (gm_n1107, gm_n88, gm_n86, gm_n119, gm_n1106);
	nand (gm_n1108, gm_n1107, gm_n1105, gm_n1103);
	or (gm_n1109, gm_n406, in_13, gm_n62, gm_n503, gm_n502);
	nor (gm_n1110, gm_n256, in_21, gm_n55, gm_n1109, gm_n312);
	nor (out_1, gm_n1108, gm_n1100, gm_n763, gm_n1110);
	or (gm_n1112, gm_n841, gm_n147, in_14, gm_n981, gm_n271);
	nor (gm_n1113, gm_n1112, gm_n87, in_18);
	nor (gm_n1114, gm_n149, in_14, gm_n78, gm_n807, gm_n247);
	nand (gm_n1115, gm_n348, gm_n245, gm_n119, gm_n1114);
	or (gm_n1116, gm_n190, gm_n73, in_12, gm_n835, gm_n276);
	nor (gm_n1117, gm_n781, in_21, in_20, gm_n1116);
	nand (gm_n1118, gm_n90, gm_n78, in_9, gm_n825, gm_n532);
	nor (gm_n1119, gm_n89, gm_n87, gm_n119, gm_n1118);
	and (gm_n1120, in_6, gm_n97, gm_n108, gm_n169, in_7);
	and (gm_n1121, gm_n78, gm_n62, in_8, gm_n1120, gm_n334);
	nand (gm_n1122, gm_n164, gm_n119, gm_n90, gm_n1121, gm_n245);
	nor (gm_n1123, gm_n153, gm_n190, gm_n60, gm_n485, gm_n193);
	nand (gm_n1124, gm_n72, in_20, in_19, gm_n1123);
	or (gm_n1125, gm_n229, gm_n194, gm_n94);
	or (gm_n1126, gm_n90, gm_n78, in_9, gm_n1125, gm_n467);
	nor (gm_n1127, gm_n437, gm_n211, in_18, gm_n1126);
	or (gm_n1128, gm_n155, in_16, gm_n59, gm_n855, gm_n276);
	nor (gm_n1129, gm_n496, in_21, in_20, gm_n1128);
	nor (gm_n1130, gm_n431, in_13, in_9, gm_n432, gm_n344);
	nand (gm_n1131, gm_n174, gm_n72, in_17, gm_n1130, gm_n1076);
	nand (gm_n1132, in_4, in_3, in_2, gm_n315, gm_n97);
	nor (gm_n1133, gm_n514, in_13, in_9, gm_n1132, gm_n609);
	nand (gm_n1134, gm_n405, gm_n72, in_17, gm_n1133, gm_n327);
	and (gm_n1135, gm_n802, gm_n81, gm_n94);
	nand (gm_n1136, gm_n64, gm_n73, gm_n59, gm_n1135, gm_n303);
	nor (gm_n1137, gm_n58, gm_n72, in_20, gm_n1136);
	or (gm_n1138, gm_n263, in_16, in_12, gm_n855, gm_n385);
	nor (gm_n1139, gm_n781, gm_n72, in_20, gm_n1138);
	nor (gm_n1140, gm_n609, gm_n76, gm_n62, gm_n345, gm_n431);
	nand (gm_n1141, gm_n523, gm_n72, in_17, gm_n1140, gm_n373);
	nor (gm_n1142, gm_n344, gm_n76, gm_n62, gm_n743, gm_n480);
	nand (gm_n1143, gm_n174, gm_n72, in_17, gm_n1142, gm_n339);
	not (gm_n1144, gm_n283);
	nand (gm_n1145, gm_n484, in_15, in_11, gm_n601, gm_n1144);
	nor (gm_n1146, in_21, gm_n85, gm_n56, gm_n1145, gm_n485);
	nor (gm_n1147, gm_n625, gm_n194, in_8);
	nand (gm_n1148, gm_n222, gm_n192, in_15, gm_n1147, gm_n394);
	nor (gm_n1149, in_21, gm_n85, in_19, gm_n1148);
	or (gm_n1150, gm_n625, gm_n68, gm_n94);
	nor (gm_n1151, gm_n184, in_13, in_9, gm_n1150, gm_n406);
	nand (gm_n1152, gm_n174, in_21, in_17, gm_n1151);
	nor (gm_n1153, gm_n485, gm_n274, in_15, gm_n552, gm_n764);
	nand (gm_n1154, gm_n72, gm_n85, in_19, gm_n1153);
	nor (gm_n1155, gm_n461, in_13, gm_n62, gm_n743, gm_n443);
	and (gm_n1156, gm_n255, in_21, in_17, gm_n1155, gm_n311);
	not (gm_n1157, gm_n148);
	not (gm_n1158, gm_n467);
	nand (gm_n1159, gm_n1157, in_14, gm_n78, gm_n829, gm_n1158);
	nor (gm_n1160, gm_n841, gm_n824, in_18, gm_n1159);
	nor (gm_n1161, gm_n215, gm_n194, in_8);
	and (gm_n1162, gm_n192, gm_n143, gm_n60, gm_n1161, gm_n486);
	nand (gm_n1163, in_21, gm_n85, in_19, gm_n1162);
	nor (gm_n1164, gm_n609, in_10, in_9, gm_n503, gm_n362);
	nand (gm_n1165, gm_n146, gm_n119, in_14, gm_n1164, gm_n806);
	or (gm_n1166, gm_n190, gm_n73, in_12, gm_n799, gm_n152);
	nor (gm_n1167, gm_n219, gm_n72, gm_n85, gm_n1166);
	or (gm_n1168, gm_n349, gm_n90, in_10, gm_n467, gm_n389);
	nor (gm_n1169, gm_n212, gm_n824, in_18, gm_n1168);
	nand (gm_n1170, in_7, in_6, in_5, gm_n519, in_8);
	nor (gm_n1171, gm_n213, gm_n76, in_12, gm_n1170);
	nand (gm_n1172, gm_n120, in_21, gm_n55, gm_n1171, gm_n1076);
	nand (gm_n1173, gm_n93, in_6, gm_n97, gm_n546, gm_n94);
	nor (gm_n1174, in_14, gm_n78, in_9, gm_n1173, gm_n369);
	nand (gm_n1175, gm_n323, gm_n199, in_18, gm_n1174);
	or (gm_n1176, gm_n572, gm_n277, gm_n94);
	or (gm_n1177, gm_n227, in_16, in_12, gm_n1176, gm_n213);
	nor (gm_n1178, gm_n219, gm_n72, gm_n85, gm_n1177);
	and (gm_n1179, gm_n305, gm_n291, in_8);
	nand (gm_n1180, gm_n281, gm_n79, gm_n60, gm_n1179, gm_n449);
	nor (gm_n1181, gm_n72, gm_n85, in_19, gm_n1180);
	nor (gm_n1182, gm_n286, gm_n461, in_13, gm_n375, gm_n370);
	nand (gm_n1183, gm_n120, in_21, in_17, gm_n1182);
	and (gm_n1184, gm_n449, gm_n79, in_15, gm_n1095, gm_n486);
	nand (gm_n1185, gm_n72, in_20, gm_n56, gm_n1184);
	and (gm_n1186, gm_n93, in_6, gm_n97, gm_n519, in_8);
	nand (gm_n1187, gm_n379, gm_n143, in_15, gm_n1186, gm_n192);
	nor (gm_n1188, gm_n72, in_20, gm_n56, gm_n1187);
	nor (gm_n1189, gm_n208, gm_n461, in_13, gm_n313, gm_n287);
	nand (gm_n1190, gm_n102, gm_n72, gm_n55, gm_n1189);
	nand (gm_n1191, gm_n93, in_6, in_5, gm_n519, in_8);
	nor (gm_n1192, gm_n152, gm_n115, gm_n59, gm_n1191);
	nand (gm_n1193, gm_n72, gm_n85, in_19, gm_n1192, gm_n268);
	or (gm_n1194, gm_n344, in_13, gm_n62, gm_n1132, gm_n442);
	nor (gm_n1195, gm_n121, in_21, in_17, gm_n1194, gm_n374);
	nand (gm_n1196, gm_n222, in_16, gm_n59, gm_n1079, gm_n303);
	nor (gm_n1197, gm_n384, in_21, gm_n85, gm_n1196);
	nor (gm_n1198, gm_n234, gm_n228, in_8);
	nand (gm_n1199, gm_n532, gm_n78, gm_n62, gm_n1198);
	or (gm_n1200, gm_n312, in_21, gm_n55, gm_n1199, gm_n662);
	nor (gm_n1201, gm_n159, gm_n74, gm_n60, gm_n263, gm_n251);
	nand (gm_n1202, in_21, in_20, gm_n56, gm_n1201);
	or (gm_n1203, gm_n234, gm_n228, in_8);
	nor (gm_n1204, gm_n158, gm_n73, gm_n59, gm_n1203, gm_n354);
	nand (gm_n1205, gm_n113, in_21, gm_n85, gm_n1204);
	nor (gm_n1206, gm_n92, in_14, gm_n78, gm_n287, gm_n286);
	nand (gm_n1207, gm_n436, gm_n199, gm_n119, gm_n1206);
	or (gm_n1208, gm_n572, gm_n195, gm_n94);
	nor (gm_n1209, gm_n92, in_10, gm_n62, gm_n1208);
	nand (gm_n1210, gm_n122, in_21, in_17, gm_n1209, gm_n174);
	nand (gm_n1211, gm_n1205, gm_n1202, gm_n1200, gm_n1210, gm_n1207);
	nor (gm_n1212, gm_n263, gm_n73, in_12, gm_n832, gm_n354);
	nand (gm_n1213, gm_n57, in_21, gm_n85, gm_n1212);
	nor (gm_n1214, gm_n193, in_15, in_11, gm_n761, gm_n283);
	nand (gm_n1215, gm_n72, gm_n85, gm_n56, gm_n1214, gm_n75);
	nor (gm_n1216, gm_n135, in_16, in_12, gm_n276, gm_n263);
	nand (gm_n1217, gm_n296, in_21, in_20, gm_n1216);
	nand (gm_n1218, gm_n1217, gm_n1215, gm_n1213);
	and (gm_n1219, gm_n79, gm_n73, gm_n59, gm_n265, gm_n733);
	nand (gm_n1220, gm_n138, in_21, in_20, gm_n1219);
	nor (gm_n1221, gm_n609, in_13, in_9, gm_n621, gm_n431);
	nand (gm_n1222, gm_n174, in_21, gm_n55, gm_n1221, gm_n1076);
	nand (gm_n1223, gm_n93, in_6, gm_n97, gm_n134, in_8);
	nor (gm_n1224, gm_n155, gm_n76, in_12, gm_n1223);
	nand (gm_n1225, gm_n523, gm_n72, in_17, gm_n1224, gm_n206);
	nand (gm_n1226, gm_n1225, gm_n1222, gm_n1220);
	nor (gm_n1227, gm_n1211, gm_n1197, gm_n1195, gm_n1226, gm_n1218);
	or (gm_n1228, gm_n596, in_13, in_9, gm_n621, gm_n442);
	nor (gm_n1229, gm_n256, gm_n72, in_17, gm_n1228, gm_n374);
	nor (gm_n1230, gm_n228, gm_n201, gm_n94);
	nand (gm_n1231, gm_n1158, gm_n78, in_9, gm_n1230);
	nor (gm_n1232, gm_n662, in_21, in_17, gm_n1231, gm_n374);
	or (gm_n1233, gm_n461, gm_n76, gm_n62, gm_n597, gm_n502);
	nor (gm_n1234, gm_n620, in_21, gm_n55, gm_n1233, gm_n662);
	nor (gm_n1235, gm_n1234, gm_n1232, gm_n1229);
	or (gm_n1236, gm_n358, gm_n76, gm_n62, gm_n988, gm_n443);
	nor (gm_n1237, gm_n183, gm_n72, gm_n55, gm_n1236, gm_n256);
	nor (gm_n1238, gm_n105, gm_n72, gm_n55, gm_n390, gm_n374);
	nor (gm_n1239, in_7, in_6, in_5, gm_n67, gm_n94);
	nand (gm_n1240, gm_n64, in_16, gm_n59, gm_n1239, gm_n571);
	nor (gm_n1241, gm_n139, gm_n72, in_20, gm_n1240);
	nor (gm_n1242, gm_n1241, gm_n1238, gm_n1237);
	nand (gm_n1243, gm_n1227, gm_n1193, gm_n1190, gm_n1242, gm_n1235);
	nor (gm_n1244, gm_n290, gm_n158, in_15, gm_n1016, gm_n293);
	nand (gm_n1245, gm_n72, in_20, in_19, gm_n1244);
	or (gm_n1246, gm_n229, gm_n202, gm_n94);
	nor (gm_n1247, gm_n193, gm_n191, gm_n60, gm_n1246, gm_n213);
	nand (gm_n1248, in_21, gm_n85, in_19, gm_n1247);
	nor (gm_n1249, gm_n430, gm_n76, in_9, gm_n359, gm_n431);
	nand (gm_n1250, gm_n122, in_21, in_17, gm_n1249, gm_n206);
	nand (gm_n1251, gm_n1250, gm_n1248, gm_n1245);
	nor (gm_n1252, gm_n293, gm_n297, in_15, gm_n855, gm_n760);
	nand (gm_n1253, in_21, gm_n85, in_19, gm_n1252);
	nor (gm_n1254, gm_n358, gm_n76, in_9, gm_n621, gm_n430);
	nand (gm_n1255, gm_n102, in_21, gm_n55, gm_n1254, gm_n523);
	nor (gm_n1256, gm_n190, in_16, in_12, gm_n1006, gm_n319);
	nand (gm_n1257, gm_n57, in_21, gm_n85, gm_n1256);
	nand (gm_n1258, gm_n1257, gm_n1255, gm_n1253);
	nor (gm_n1259, gm_n1243, gm_n1188, t_6, gm_n1258, gm_n1251);
	or (gm_n1260, gm_n572, gm_n234, gm_n94);
	or (gm_n1261, gm_n147, in_10, gm_n62, gm_n1260);
	nor (gm_n1262, gm_n121, in_21, in_17, gm_n1261, gm_n312);
	nor (gm_n1263, in_7, in_6, in_5, gm_n229);
	nand (gm_n1264, gm_n78, in_9, in_8, gm_n1263, gm_n1158);
	nor (gm_n1265, gm_n824, gm_n119, in_14, gm_n1264, gm_n246);
	or (gm_n1266, gm_n115, gm_n73, gm_n59, gm_n468, gm_n319);
	nor (gm_n1267, gm_n384, in_21, gm_n85, gm_n1266);
	nor (gm_n1268, gm_n1267, gm_n1265, gm_n1262);
	or (gm_n1269, gm_n191, gm_n159, in_15, gm_n552, gm_n274);
	nor (gm_n1270, in_21, gm_n85, in_19, gm_n1269);
	or (gm_n1271, gm_n90, in_13, in_12, gm_n855, gm_n158);
	nor (gm_n1272, gm_n531, gm_n212, gm_n119, gm_n1271);
	or (gm_n1273, gm_n480, in_13, in_9, gm_n621, gm_n443);
	nor (gm_n1274, gm_n103, gm_n72, in_17, gm_n1273, gm_n313);
	nor (gm_n1275, gm_n1274, gm_n1272, gm_n1270);
	nand (gm_n1276, gm_n1259, gm_n1185, gm_n1183, gm_n1275, gm_n1268);
	and (gm_n1277, gm_n579, gm_n76, in_9, gm_n1049, gm_n316);
	nand (gm_n1278, gm_n104, gm_n72, gm_n55, gm_n1277, gm_n373);
	and (gm_n1279, gm_n106, in_13, in_9, gm_n187, gm_n107);
	nand (gm_n1280, gm_n523, gm_n72, gm_n55, gm_n1279, gm_n254);
	nor (gm_n1281, gm_n92, in_14, gm_n78, gm_n389, gm_n349);
	nand (gm_n1282, gm_n367, gm_n166, gm_n119, gm_n1281);
	nand (gm_n1283, gm_n1282, gm_n1280, gm_n1278);
	nand (gm_n1284, gm_n426, gm_n304, gm_n94);
	nor (gm_n1285, in_14, gm_n78, in_9, gm_n1284, gm_n467);
	nand (gm_n1286, gm_n243, gm_n200, gm_n119, gm_n1285);
	nor (gm_n1287, gm_n480, gm_n76, in_9, gm_n481, gm_n463);
	nand (gm_n1288, gm_n255, in_21, in_17, gm_n1287, gm_n373);
	nor (gm_n1289, gm_n358, gm_n76, in_9, gm_n503, gm_n667);
	nand (gm_n1290, gm_n104, in_21, in_17, gm_n1289, gm_n174);
	nand (gm_n1291, gm_n1290, gm_n1288, gm_n1286);
	nor (gm_n1292, gm_n1276, gm_n1181, gm_n1178, gm_n1291, gm_n1283);
	or (gm_n1293, gm_n358, gm_n76, in_9, gm_n481, gm_n596);
	nor (gm_n1294, gm_n183, gm_n72, gm_n55, gm_n1293, gm_n375);
	not (gm_n1295, gm_n126);
	or (gm_n1296, gm_n1295, gm_n76, gm_n62, gm_n344, gm_n406);
	nor (gm_n1297, gm_n441, gm_n72, gm_n55, gm_n1296, gm_n375);
	or (gm_n1298, gm_n431, in_13, gm_n62, gm_n344, gm_n866);
	nor (gm_n1299, gm_n256, in_21, in_17, gm_n1298, gm_n620);
	nor (gm_n1300, gm_n1299, gm_n1297, gm_n1294);
	or (gm_n1301, gm_n191, gm_n190, gm_n60, gm_n855, gm_n290);
	nor (gm_n1302, in_21, gm_n85, in_19, gm_n1301);
	or (gm_n1303, gm_n257, gm_n76, in_9, gm_n621, gm_n443);
	nor (gm_n1304, gm_n313, in_21, in_17, gm_n1303, gm_n620);
	or (gm_n1305, gm_n190, gm_n73, in_12, gm_n319, gm_n116);
	nor (gm_n1306, gm_n781, gm_n72, in_20, gm_n1305);
	nor (gm_n1307, gm_n1306, gm_n1304, gm_n1302);
	nand (gm_n1308, gm_n1292, gm_n1175, gm_n1172, gm_n1307, gm_n1300);
	nor (gm_n1309, gm_n208, gm_n90, in_10, gm_n370, gm_n362);
	nand (gm_n1310, gm_n348, gm_n166, in_18, gm_n1309);
	and (gm_n1311, in_14, gm_n78, gm_n62, gm_n803, gm_n532);
	nand (gm_n1312, gm_n367, gm_n200, in_18, gm_n1311);
	nor (gm_n1313, gm_n158, gm_n76, in_12, gm_n520);
	nand (gm_n1314, gm_n523, gm_n72, in_17, gm_n1313, gm_n206);
	nand (gm_n1315, gm_n1314, gm_n1312, gm_n1310);
	or (gm_n1316, gm_n103, gm_n72, in_17, gm_n1109, gm_n256);
	nor (gm_n1317, gm_n442, in_13, gm_n62, gm_n988, gm_n502);
	nand (gm_n1318, gm_n102, gm_n72, gm_n55, gm_n1317, gm_n104);
	or (gm_n1319, gm_n228, gm_n67, gm_n94);
	nor (gm_n1320, gm_n152, in_16, gm_n59, gm_n1319, gm_n274);
	nand (gm_n1321, gm_n113, in_21, gm_n85, gm_n1320);
	nand (gm_n1322, gm_n1321, gm_n1318, gm_n1316);
	nor (gm_n1323, gm_n1308, gm_n1169, gm_n1167, gm_n1322, gm_n1315);
	or (gm_n1324, in_7, in_6, in_5, gm_n67, in_8);
	or (gm_n1325, gm_n274, gm_n74, in_15, gm_n1324, gm_n633);
	nor (gm_n1326, in_21, gm_n85, gm_n56, gm_n1325);
	nand (gm_n1327, in_14, in_10, gm_n62, gm_n626, gm_n1011);
	nor (gm_n1328, gm_n531, gm_n89, in_18, gm_n1327);
	and (gm_n1329, in_21, in_20, gm_n56, gm_n1192, gm_n281);
	nor (gm_n1330, gm_n1329, gm_n1328, gm_n1326);
	not (gm_n1331, gm_n281);
	nand (gm_n1332, gm_n134, gm_n81, in_8);
	or (gm_n1333, gm_n213, gm_n193, gm_n60, gm_n1332, gm_n1331);
	nor (gm_n1334, gm_n72, in_20, gm_n56, gm_n1333);
	or (gm_n1335, gm_n133, gm_n90, in_10, gm_n775, gm_n247);
	nor (gm_n1336, gm_n437, gm_n824, gm_n119, gm_n1335);
	nand (gm_n1337, gm_n126, gm_n76, in_9, gm_n1049, gm_n314);
	nor (gm_n1338, gm_n183, in_21, gm_n55, gm_n1337, gm_n662);
	nor (gm_n1339, gm_n1338, gm_n1336, gm_n1334);
	nand (gm_n1340, gm_n1323, gm_n1165, gm_n1163, gm_n1339, gm_n1330);
	nor (gm_n1341, gm_n358, in_13, in_9, gm_n597, gm_n430);
	nand (gm_n1342, gm_n174, gm_n72, in_17, gm_n1341, gm_n339);
	nor (gm_n1343, gm_n207, in_14, in_10, gm_n589, gm_n491);
	nand (gm_n1344, gm_n348, gm_n88, gm_n119, gm_n1343);
	not (gm_n1345, gm_n370);
	and (gm_n1346, gm_n532, in_14, in_10, gm_n793, gm_n1345);
	nand (gm_n1347, gm_n323, gm_n164, in_18, gm_n1346);
	nand (gm_n1348, gm_n1347, gm_n1344, gm_n1342);
	nor (gm_n1349, gm_n667, in_13, in_9, gm_n743, gm_n442);
	nand (gm_n1350, gm_n206, gm_n72, in_17, gm_n1349, gm_n405);
	nor (gm_n1351, gm_n115, in_12, gm_n94, gm_n508, gm_n152);
	nand (gm_n1352, in_21, gm_n85, in_16, gm_n1351, gm_n138);
	nor (gm_n1353, gm_n609, in_13, in_9, gm_n481, gm_n358);
	nand (gm_n1354, gm_n327, in_21, in_17, gm_n1353, gm_n339);
	nand (gm_n1355, gm_n1354, gm_n1352, gm_n1350);
	nor (gm_n1356, gm_n1340, gm_n1160, gm_n1156, gm_n1355, gm_n1348);
	nand (gm_n1357, in_13, in_9, gm_n94, gm_n576, gm_n579);
	nor (gm_n1358, gm_n105, gm_n72, in_17, gm_n1357, gm_n183);
	and (gm_n1359, in_7, in_6, gm_n97, gm_n134, gm_n94);
	and (gm_n1360, gm_n90, gm_n76, in_12, gm_n1359, gm_n264);
	and (gm_n1361, gm_n131, gm_n129, gm_n119, gm_n1360);
	nor (gm_n1362, gm_n90, gm_n78, in_9, gm_n499, gm_n362);
	and (gm_n1363, gm_n243, gm_n88, in_18, gm_n1362);
	nor (gm_n1364, gm_n1363, gm_n1361, gm_n1358);
	nor (gm_n1365, gm_n103, in_21, in_17, gm_n587, gm_n313);
	or (gm_n1366, gm_n866, gm_n78, gm_n62, gm_n502, gm_n467);
	nor (gm_n1367, gm_n244, gm_n119, in_14, gm_n1366, gm_n246);
	or (gm_n1368, gm_n406, gm_n76, in_9, gm_n621, gm_n596);
	nor (gm_n1369, gm_n121, in_21, in_17, gm_n1368, gm_n441);
	nor (gm_n1370, gm_n1369, gm_n1367, gm_n1365);
	nand (gm_n1371, gm_n1356, gm_n1154, gm_n1152, gm_n1370, gm_n1364);
	nor (gm_n1372, in_14, gm_n78, gm_n62, gm_n657, gm_n147);
	nand (gm_n1373, gm_n166, gm_n164, gm_n119, gm_n1372);
	nor (gm_n1374, gm_n514, in_13, in_9, gm_n597, gm_n344);
	nand (gm_n1375, gm_n174, gm_n72, in_17, gm_n1374, gm_n595);
	nor (gm_n1376, gm_n431, gm_n76, gm_n62, gm_n481, gm_n596);
	nand (gm_n1377, gm_n327, in_21, in_17, gm_n1376, gm_n1076);
	nand (gm_n1378, gm_n1377, gm_n1375, gm_n1373);
	nor (gm_n1379, gm_n229, gm_n68);
	and (gm_n1380, gm_n64, in_12, gm_n94, gm_n949, gm_n1379);
	nand (gm_n1381, in_21, gm_n85, in_16, gm_n1380, gm_n57);
	or (gm_n1382, gm_n572, gm_n229);
	nor (gm_n1383, gm_n158, gm_n59, in_8, gm_n1382, gm_n152);
	nand (gm_n1384, gm_n119, gm_n55, gm_n73, gm_n1383, gm_n146);
	nor (gm_n1385, gm_n807, gm_n90, in_10, gm_n438, gm_n414);
	nand (gm_n1386, gm_n348, gm_n166, in_18, gm_n1385);
	nand (gm_n1387, gm_n1386, gm_n1384, gm_n1381);
	nor (gm_n1388, gm_n1371, gm_n1149, gm_n1146, gm_n1387, gm_n1378);
	nor (gm_n1389, gm_n496, gm_n72, gm_n85, gm_n706);
	or (gm_n1390, gm_n667, in_13, gm_n62, gm_n345, gm_n431);
	nor (gm_n1391, gm_n103, gm_n72, in_17, gm_n1390, gm_n328);
	and (gm_n1392, gm_n546, gm_n304, in_8);
	nand (gm_n1393, gm_n268, gm_n64, in_15, gm_n1392, gm_n422);
	nor (gm_n1394, gm_n72, in_20, gm_n56, gm_n1393);
	nor (gm_n1395, gm_n1394, gm_n1391, gm_n1389);
	or (gm_n1396, gm_n461, gm_n76, in_9, gm_n1132, gm_n596);
	nor (gm_n1397, gm_n105, gm_n72, gm_n55, gm_n1396, gm_n620);
	not (gm_n1398, gm_n633);
	nand (gm_n1399, gm_n264, gm_n75, gm_n60, gm_n1398, gm_n615);
	nor (gm_n1400, in_21, in_20, in_19, gm_n1399);
	and (gm_n1401, in_7, gm_n124, in_5, gm_n134, in_8);
	nand (gm_n1402, gm_n571, gm_n264, gm_n59, gm_n1401);
	nor (gm_n1403, in_21, gm_n85, in_19, gm_n1402, gm_n393);
	nor (gm_n1404, gm_n1403, gm_n1400, gm_n1397);
	nand (gm_n1405, gm_n1388, gm_n1143, gm_n1141, gm_n1404, gm_n1395);
	nand (gm_n1406, gm_n93, gm_n124, in_5, gm_n426, in_8);
	nor (gm_n1407, gm_n114, gm_n73, gm_n59, gm_n1406, gm_n213);
	nand (gm_n1408, gm_n138, in_21, gm_n85, gm_n1407);
	nor (gm_n1409, gm_n514, gm_n76, gm_n62, gm_n988, gm_n596);
	nand (gm_n1410, gm_n327, gm_n72, gm_n55, gm_n1409, gm_n595);
	nor (gm_n1411, gm_n514, in_13, gm_n62, gm_n359, gm_n430);
	nand (gm_n1412, gm_n122, in_21, gm_n55, gm_n1411, gm_n174);
	nand (gm_n1413, gm_n1412, gm_n1410, gm_n1408);
	nor (gm_n1414, gm_n212, gm_n977, gm_n90, gm_n761, gm_n369);
	nand (gm_n1415, gm_n1414, gm_n348, in_18);
	and (gm_n1416, gm_n426, gm_n81, in_8);
	and (gm_n1417, gm_n733, gm_n73, in_12, gm_n1416, gm_n222);
	nand (gm_n1418, gm_n113, in_21, in_20, gm_n1417);
	nor (gm_n1419, gm_n514, gm_n76, in_9, gm_n596, gm_n818);
	nand (gm_n1420, gm_n311, gm_n72, gm_n55, gm_n1419, gm_n1076);
	nand (gm_n1421, gm_n1420, gm_n1418, gm_n1415);
	nor (gm_n1422, gm_n1405, gm_n1139, gm_n1137, gm_n1421, gm_n1413);
	or (gm_n1423, gm_n431, in_13, gm_n62, gm_n1132, gm_n502);
	nor (gm_n1424, gm_n183, in_21, in_17, gm_n1423, gm_n375);
	or (gm_n1425, gm_n257, gm_n76, in_9, gm_n503, gm_n596);
	nor (gm_n1426, gm_n388, in_21, in_17, gm_n1425, gm_n313);
	and (gm_n1427, in_7, gm_n124, in_5, gm_n134, gm_n94);
	nand (gm_n1428, gm_n523, in_13, in_9, gm_n1427, gm_n185);
	nor (gm_n1429, gm_n441, gm_n72, in_17, gm_n1428);
	nor (gm_n1430, gm_n1429, gm_n1426, gm_n1424);
	or (gm_n1431, gm_n78, in_9, in_8, gm_n807, gm_n270);
	nor (gm_n1432, gm_n165, gm_n119, gm_n90, gm_n1431, gm_n212);
	or (gm_n1433, gm_n430, gm_n76, in_9, gm_n481, gm_n257);
	nor (gm_n1434, gm_n103, gm_n72, gm_n55, gm_n1433, gm_n105);
	nand (gm_n1435, gm_n143, gm_n73, in_12, gm_n1359, gm_n221);
	nor (gm_n1436, gm_n912, in_21, gm_n85, gm_n1435);
	nor (gm_n1437, gm_n1436, gm_n1434, gm_n1432);
	nand (gm_n1438, gm_n1422, gm_n1134, gm_n1131, gm_n1437, gm_n1430);
	and (gm_n1439, gm_n828, in_14, in_10, gm_n829, gm_n600);
	nand (gm_n1440, gm_n323, gm_n199, gm_n119, gm_n1439);
	and (gm_n1441, gm_n79, in_16, gm_n59, gm_n411, gm_n571);
	nand (gm_n1442, gm_n113, in_21, in_20, gm_n1441);
	and (gm_n1443, gm_n532, gm_n104, gm_n78, gm_n490, gm_n333);
	nand (gm_n1444, gm_n311, in_21, gm_n55, gm_n1443);
	nand (gm_n1445, gm_n1444, gm_n1442, gm_n1440);
	nor (gm_n1446, gm_n238, gm_n202, gm_n94);
	and (gm_n1447, gm_n154, in_16, in_12, gm_n1446, gm_n221);
	nand (gm_n1448, gm_n113, gm_n72, in_20, gm_n1447);
	or (gm_n1449, gm_n115, in_16, in_12, gm_n657, gm_n385);
	or (gm_n1450, gm_n244, in_18, gm_n55, gm_n1449);
	nor (gm_n1451, gm_n625, gm_n572, in_8);
	and (gm_n1452, gm_n233, gm_n73, in_12, gm_n1451, gm_n949);
	nand (gm_n1453, gm_n296, gm_n72, gm_n85, gm_n1452);
	nand (gm_n1454, gm_n1453, gm_n1450, gm_n1448);
	nor (gm_n1455, gm_n1438, gm_n1129, gm_n1127, gm_n1454, gm_n1445);
	and (gm_n1456, gm_n93, in_6, in_5, gm_n546, gm_n94);
	nand (gm_n1457, gm_n233, gm_n73, in_12, gm_n1456, gm_n303);
	nor (gm_n1458, gm_n384, gm_n72, gm_n85, gm_n1457);
	or (gm_n1459, gm_n375, gm_n461, in_13, gm_n491, gm_n414);
	nor (gm_n1460, gm_n620, in_21, gm_n55, gm_n1459);
	nand (gm_n1461, gm_n76, in_9, gm_n94, gm_n756, gm_n402);
	nor (gm_n1462, gm_n313, in_21, in_17, gm_n1461, gm_n620);
	nor (gm_n1463, gm_n1462, gm_n1460, gm_n1458);
	nand (gm_n1464, gm_n77, gm_n73, gm_n59, gm_n1079, gm_n222);
	nor (gm_n1465, gm_n384, in_21, gm_n85, gm_n1464);
	nand (gm_n1466, gm_n154, gm_n75, in_15, gm_n1359, gm_n1398);
	nor (gm_n1467, gm_n72, gm_n85, in_19, gm_n1466);
	or (gm_n1468, gm_n1295, gm_n76, gm_n62, gm_n442, gm_n344);
	nor (gm_n1469, gm_n183, gm_n72, in_17, gm_n1468, gm_n121);
	nor (gm_n1470, gm_n1469, gm_n1467, gm_n1465);
	nand (gm_n1471, gm_n1455, gm_n1124, gm_n1122, gm_n1470, gm_n1463);
	nand (gm_n1472, gm_n311, in_21, gm_n55, gm_n1069, gm_n339);
	nor (gm_n1473, gm_n807, in_14, in_10, gm_n589, gm_n438);
	nand (gm_n1474, gm_n243, gm_n88, gm_n119, gm_n1473);
	or (gm_n1475, gm_n277, gm_n228, in_8);
	nor (gm_n1476, gm_n90, gm_n78, in_9, gm_n1475, gm_n807);
	nand (gm_n1477, gm_n245, gm_n86, in_18, gm_n1476);
	nand (gm_n1478, gm_n1477, gm_n1474, gm_n1472);
	and (gm_n1479, gm_n79, gm_n59, gm_n94, gm_n455, gm_n275);
	nand (gm_n1480, in_21, gm_n85, in_16, gm_n1479, gm_n383);
	nand (gm_n1481, in_7, in_6, in_5, gm_n426, gm_n94);
	nor (gm_n1482, gm_n190, in_13, in_12, gm_n1481);
	nand (gm_n1483, gm_n122, gm_n72, gm_n55, gm_n1482, gm_n206);
	or (gm_n1484, gm_n215, gm_n202, in_8);
	nor (gm_n1485, gm_n213, gm_n76, gm_n59, gm_n1484);
	nand (gm_n1486, gm_n254, gm_n72, in_17, gm_n1485, gm_n405);
	nand (gm_n1487, gm_n1486, gm_n1483, gm_n1480);
	nor (gm_n1488, gm_n1471, gm_n1119, gm_n1117, gm_n1487, gm_n1478);
	nor (gm_n1489, gm_n278, gm_n190, in_15, gm_n447, gm_n290);
	nand (gm_n1490, in_21, gm_n85, in_19, gm_n1489);
	and (gm_n1491, gm_n222, gm_n73, in_12, gm_n1456, gm_n949);
	nand (gm_n1492, gm_n113, in_21, gm_n85, gm_n1491);
	nor (gm_n1493, gm_n78, in_9, gm_n94, gm_n417, gm_n362);
	nand (gm_n1494, gm_n199, gm_n119, gm_n90, gm_n1493, gm_n323);
	nand (gm_n1495, gm_n1490, gm_n1488, gm_n1115, gm_n1494, gm_n1492);
	nor (gm_n1496, in_7, in_6, in_5, gm_n201);
	and (gm_n1497, gm_n76, gm_n59, gm_n94, gm_n1496, gm_n264);
	nand (gm_n1498, gm_n122, gm_n72, in_17, gm_n1497, gm_n206);
	nor (gm_n1499, gm_n240, gm_n207, gm_n90, gm_n270);
	nand (gm_n1500, gm_n166, gm_n164, gm_n119, gm_n1499);
	nor (gm_n1501, gm_n228, gm_n195, in_8);
	and (gm_n1502, gm_n64, in_16, gm_n59, gm_n1501, gm_n77);
	nand (gm_n1503, gm_n296, gm_n72, gm_n85, gm_n1502);
	nand (gm_n1504, gm_n1503, gm_n1500, gm_n1498);
	or (gm_n1505, gm_n796, gm_n76, in_9, gm_n463, gm_n257);
	nor (gm_n1506, gm_n620, gm_n72, gm_n55, gm_n1505, gm_n662);
	nor (out_2, gm_n1504, gm_n1495, gm_n1113, gm_n1506);
	or (gm_n1508, in_14, in_10, in_9, gm_n832, gm_n147);
	nor (gm_n1509, gm_n368, gm_n841, in_18, gm_n1508);
	nor (gm_n1510, gm_n147, in_14, in_10, gm_n775, gm_n438);
	nand (gm_n1511, gm_n323, gm_n129, in_18, gm_n1510);
	and (gm_n1512, gm_n624, in_14, in_10, gm_n722, gm_n490);
	nand (gm_n1513, gm_n367, gm_n245, gm_n119, gm_n1512);
	or (gm_n1514, gm_n625, gm_n202, in_8);
	or (gm_n1515, gm_n257, in_13, gm_n62, gm_n1514, gm_n328);
	nor (gm_n1516, gm_n183, gm_n72, in_17, gm_n1515);
	or (gm_n1517, gm_n193, gm_n158, in_15, gm_n765, gm_n1331);
	nor (gm_n1518, in_21, in_20, gm_n56, gm_n1517);
	or (gm_n1519, gm_n202, gm_n201, in_8);
	nor (gm_n1520, gm_n159, gm_n74, in_15, gm_n1519, gm_n274);
	nand (gm_n1521, gm_n72, gm_n85, in_19, gm_n1520);
	nor (gm_n1522, gm_n514, gm_n76, in_9, gm_n443, gm_n818);
	nand (gm_n1523, gm_n327, gm_n72, gm_n55, gm_n1522, gm_n339);
	and (gm_n1524, in_7, in_6, in_5, gm_n80, in_8);
	and (gm_n1525, gm_n733, gm_n64, in_12, gm_n1524);
	and (gm_n1526, gm_n72, in_20, in_19, gm_n1525, gm_n1101);
	or (gm_n1527, gm_n159, in_15, gm_n63, gm_n605, gm_n270);
	nor (gm_n1528, in_21, in_20, gm_n56, gm_n1527, gm_n485);
	and (gm_n1529, gm_n90, gm_n78, in_9, gm_n216, gm_n532);
	nand (gm_n1530, gm_n323, gm_n199, in_18, gm_n1529);
	nor (gm_n1531, gm_n93, in_6, in_5, gm_n238, in_8);
	nand (gm_n1532, gm_n79, gm_n73, in_12, gm_n1531, gm_n571);
	or (gm_n1533, gm_n374, in_21, gm_n55, gm_n1532);
	nand (gm_n1534, in_10, gm_n62, in_8, gm_n1158, gm_n455);
	nor (gm_n1535, gm_n132, gm_n119, gm_n90, gm_n1534, gm_n165);
	nand (gm_n1536, gm_n222, in_12, in_8, gm_n580, gm_n303);
	nor (gm_n1537, gm_n72, gm_n85, in_16, gm_n1536, gm_n219);
	nor (gm_n1538, in_14, in_10, gm_n62, gm_n458, gm_n362);
	nand (gm_n1539, gm_n164, gm_n131, in_18, gm_n1538);
	nand (gm_n1540, gm_n154, in_13, in_12, gm_n953);
	or (gm_n1541, gm_n620, in_21, in_17, gm_n1540, gm_n375);
	nand (gm_n1542, gm_n93, gm_n124, in_5, gm_n546, in_8);
	or (gm_n1543, gm_n290, gm_n274, in_15, gm_n1542, gm_n393);
	nor (gm_n1544, gm_n72, in_20, gm_n56, gm_n1543);
	or (gm_n1545, gm_n643, gm_n60, in_11, gm_n761, gm_n605);
	nor (gm_n1546, in_21, gm_n85, gm_n56, gm_n1545, gm_n447);
	nor (gm_n1547, gm_n442, in_13, gm_n62, gm_n743, gm_n443);
	nand (gm_n1548, gm_n120, in_21, gm_n55, gm_n1547, gm_n595);
	and (gm_n1549, gm_n154, in_16, gm_n59, gm_n423, gm_n275);
	nand (gm_n1550, gm_n296, in_21, in_20, gm_n1549);
	or (gm_n1551, gm_n313, gm_n257, gm_n76, gm_n414, gm_n349);
	nor (gm_n1552, gm_n441, in_21, in_17, gm_n1551);
	nand (gm_n1553, in_14, in_10, in_9, gm_n991, gm_n532);
	nor (gm_n1554, gm_n437, gm_n211, in_18, gm_n1553);
	nor (gm_n1555, gm_n95, in_14, gm_n78, gm_n350, gm_n207);
	nand (gm_n1556, gm_n245, gm_n199, in_18, gm_n1555);
	nor (gm_n1557, gm_n92, gm_n90, in_10, gm_n370, gm_n248);
	nand (gm_n1558, gm_n806, gm_n129, in_18, gm_n1557);
	or (gm_n1559, gm_n358, in_13, gm_n62, gm_n503, gm_n430);
	nor (gm_n1560, gm_n441, gm_n72, in_17, gm_n1559, gm_n256);
	or (gm_n1561, gm_n609, gm_n76, gm_n62, gm_n432, gm_n257);
	nor (gm_n1562, gm_n388, gm_n72, gm_n55, gm_n1561, gm_n328);
	nor (gm_n1563, gm_n287, gm_n90, in_10, gm_n589, gm_n807);
	nand (gm_n1564, gm_n243, gm_n166, gm_n119, gm_n1563);
	nor (gm_n1565, gm_n349, gm_n257, gm_n76, gm_n589);
	nand (gm_n1566, gm_n311, in_21, gm_n55, gm_n1565, gm_n595);
	or (gm_n1567, gm_n158, gm_n73, gm_n59, gm_n799, gm_n354);
	nor (gm_n1568, gm_n384, in_21, in_20, gm_n1567);
	nor (gm_n1569, gm_n202, gm_n195, in_8);
	nand (gm_n1570, gm_n154, gm_n73, in_12, gm_n1569, gm_n571);
	nor (gm_n1571, gm_n58, in_21, in_20, gm_n1570);
	nor (gm_n1572, gm_n263, gm_n73, gm_n59, gm_n1332, gm_n319);
	nand (gm_n1573, gm_n57, in_21, in_20, gm_n1572);
	nor (gm_n1574, gm_n115, gm_n73, gm_n59, gm_n385, gm_n230);
	nand (gm_n1575, gm_n697, gm_n72, gm_n85, gm_n1574);
	or (gm_n1576, gm_n431, gm_n76, in_9, gm_n463, gm_n359);
	nor (gm_n1577, gm_n183, in_21, gm_n55, gm_n1576, gm_n184);
	nor (gm_n1578, gm_n89, gm_n87, in_18, gm_n172, gm_n168);
	and (gm_n1579, gm_n61, in_16, in_12, gm_n919, gm_n154);
	nand (gm_n1580, gm_n495, in_21, gm_n85, gm_n1579);
	nor (gm_n1581, gm_n406, in_13, gm_n62, gm_n597, gm_n443);
	nand (gm_n1582, gm_n102, gm_n72, gm_n55, gm_n1581, gm_n1076);
	nand (gm_n1583, gm_n108, gm_n96, gm_n66, gm_n109, in_5);
	or (gm_n1584, gm_n667, in_13, gm_n62, gm_n1583, gm_n480);
	nor (gm_n1585, gm_n479, gm_n72, gm_n55, gm_n1584, gm_n328);
	nor (gm_n1586, gm_n184, gm_n514, gm_n76, gm_n414, gm_n287);
	nand (gm_n1587, gm_n373, gm_n72, gm_n55, gm_n1586);
	nor (gm_n1588, gm_n461, gm_n76, gm_n62, gm_n502, gm_n345);
	nand (gm_n1589, gm_n104, in_21, gm_n55, gm_n1588, gm_n311);
	or (gm_n1590, gm_n183, in_21, in_17, gm_n960, gm_n375);
	nor (gm_n1591, gm_n514, gm_n76, gm_n62, gm_n432, gm_n596);
	nand (gm_n1592, gm_n174, in_21, in_17, gm_n1591, gm_n255);
	nor (gm_n1593, gm_n406, in_13, in_9, gm_n481, gm_n344);
	nand (gm_n1594, gm_n595, in_21, in_17, gm_n1593, gm_n373);
	nand (gm_n1595, gm_n1590, gm_n1589, gm_n1587, gm_n1594, gm_n1592);
	nand (gm_n1596, in_10, gm_n62, in_8, gm_n455, gm_n91);
	nor (gm_n1597, gm_n89, gm_n119, gm_n90, gm_n1596, gm_n531);
	nand (gm_n1598, gm_n281, gm_n79, in_15, gm_n998, gm_n449);
	nor (gm_n1599, gm_n72, in_20, gm_n56, gm_n1598);
	or (gm_n1600, gm_n430, in_13, gm_n62, gm_n988, gm_n480);
	nor (gm_n1601, gm_n121, in_21, in_17, gm_n1600, gm_n620);
	nor (gm_n1602, gm_n1597, gm_n1595, gm_n1585, gm_n1601, gm_n1599);
	or (gm_n1603, gm_n158, in_16, in_12, gm_n180, gm_n152);
	nor (gm_n1604, gm_n912, gm_n72, in_20, gm_n1603);
	nor (gm_n1605, gm_n93, in_6, gm_n97, gm_n238, gm_n94);
	nand (gm_n1606, gm_n90, in_10, in_9, gm_n1605, gm_n1011);
	nor (gm_n1607, gm_n246, gm_n211, in_18, gm_n1606);
	or (gm_n1608, gm_n147, in_10, gm_n62, gm_n462, gm_n430);
	nor (gm_n1609, gm_n211, gm_n119, in_14, gm_n1608, gm_n437);
	nor (gm_n1610, gm_n1609, gm_n1607, gm_n1604);
	and (gm_n1611, gm_n1067, gm_n291, gm_n94);
	nand (gm_n1612, gm_n90, gm_n78, gm_n62, gm_n1611, gm_n713);
	nor (gm_n1613, gm_n841, gm_n824, in_18, gm_n1612);
	not (gm_n1614, gm_n271);
	and (gm_n1615, gm_n124, gm_n97, gm_n108, gm_n169, in_7);
	nand (gm_n1616, gm_n1614, gm_n60, in_11, gm_n1615, gm_n449);
	nor (gm_n1617, gm_n72, in_20, gm_n56, gm_n1616, gm_n191);
	nand (gm_n1618, gm_n221, gm_n73, in_12, gm_n1451, gm_n222);
	nor (gm_n1619, gm_n58, in_21, in_20, gm_n1618);
	nor (gm_n1620, gm_n1619, gm_n1617, gm_n1613);
	nand (gm_n1621, gm_n1602, gm_n1582, gm_n1580, gm_n1620, gm_n1610);
	nor (gm_n1622, gm_n257, gm_n76, gm_n62, gm_n743, gm_n596);
	nand (gm_n1623, gm_n523, in_21, gm_n55, gm_n1622, gm_n254);
	nor (gm_n1624, gm_n1295, in_13, in_9, gm_n463, gm_n480);
	nand (gm_n1625, gm_n102, in_21, in_17, gm_n1624, gm_n523);
	nor (gm_n1626, gm_n274, in_16, in_12, gm_n1191, gm_n354);
	nand (gm_n1627, gm_n57, in_21, gm_n85, gm_n1626);
	nand (gm_n1628, gm_n1627, gm_n1625, gm_n1623);
	nor (gm_n1629, gm_n147, gm_n90, gm_n78, gm_n526, gm_n247);
	nand (gm_n1630, gm_n323, gm_n199, gm_n119, gm_n1629);
	nand (gm_n1631, gm_n93, gm_n124, in_5, gm_n519);
	nor (gm_n1632, in_10, in_9, gm_n94, gm_n1631, gm_n467);
	nand (gm_n1633, gm_n367, in_18, in_14, gm_n1632, gm_n436);
	nor (gm_n1634, gm_n358, in_13, gm_n62, gm_n359, gm_n596);
	nand (gm_n1635, gm_n327, gm_n72, in_17, gm_n1634, gm_n1076);
	nand (gm_n1636, gm_n1635, gm_n1633, gm_n1630);
	nor (gm_n1637, gm_n1621, gm_n1578, gm_n1577, gm_n1636, gm_n1628);
	nor (gm_n1638, gm_n274, gm_n141, gm_n94, gm_n643, gm_n572);
	nand (gm_n1639, gm_n55, gm_n73, in_15, gm_n1638);
	nor (gm_n1640, gm_n1639, gm_n374, in_21);
	or (gm_n1641, gm_n514, in_13, in_9, gm_n502, gm_n796);
	nor (gm_n1642, gm_n479, in_21, in_17, gm_n1641, gm_n313);
	nor (gm_n1643, gm_n406, in_13, gm_n62, gm_n988, gm_n596);
	and (gm_n1644, gm_n120, gm_n72, gm_n55, gm_n1643, gm_n122);
	nor (gm_n1645, gm_n1644, gm_n1642, gm_n1640);
	nand (gm_n1646, gm_n79, gm_n73, in_12, gm_n936, gm_n221);
	nor (gm_n1647, gm_n219, in_21, in_20, gm_n1646);
	or (gm_n1648, gm_n866, gm_n76, gm_n62, gm_n463, gm_n480);
	nor (gm_n1649, gm_n620, gm_n72, gm_n55, gm_n1648, gm_n662);
	or (gm_n1650, gm_n430, in_13, gm_n62, gm_n1583, gm_n480);
	nor (gm_n1651, gm_n103, in_21, gm_n55, gm_n1650, gm_n313);
	nor (gm_n1652, gm_n1651, gm_n1649, gm_n1647);
	nand (gm_n1653, gm_n1637, gm_n1575, gm_n1573, gm_n1652, gm_n1645);
	nor (gm_n1654, gm_n667, gm_n76, in_9, gm_n481, gm_n442);
	nand (gm_n1655, gm_n104, gm_n72, gm_n55, gm_n1654, gm_n373);
	nor (gm_n1656, gm_n263, gm_n74, in_15, gm_n1223, gm_n633);
	nand (gm_n1657, gm_n72, gm_n85, gm_n56, gm_n1656);
	nor (gm_n1658, in_13, gm_n62, in_8, gm_n939, gm_n431);
	nand (gm_n1659, gm_n174, in_21, in_17, gm_n1658, gm_n595);
	nand (gm_n1660, gm_n1659, gm_n1657, gm_n1655);
	or (gm_n1661, gm_n228, gm_n195, gm_n94);
	nor (gm_n1662, gm_n90, in_10, gm_n62, gm_n1661, gm_n369);
	nand (gm_n1663, gm_n323, gm_n164, in_18, gm_n1662);
	or (gm_n1664, gm_n194, gm_n67, gm_n94);
	nor (gm_n1665, in_14, in_10, gm_n62, gm_n1664, gm_n369);
	nand (gm_n1666, gm_n164, gm_n131, in_18, gm_n1665);
	nor (gm_n1667, gm_n155, in_16, in_12, gm_n1661, gm_n276);
	nand (gm_n1668, gm_n57, in_21, in_20, gm_n1667);
	nand (gm_n1669, gm_n1668, gm_n1666, gm_n1663);
	nor (gm_n1670, gm_n1653, gm_n1571, gm_n1568, gm_n1669, gm_n1660);
	or (gm_n1671, gm_n202, gm_n67, gm_n94);
	or (gm_n1672, in_14, in_10, in_9, gm_n1671, gm_n92);
	nor (gm_n1673, gm_n368, gm_n167, in_18, gm_n1672);
	or (gm_n1674, gm_n375, gm_n76, in_9, gm_n1542, gm_n480);
	nor (gm_n1675, gm_n388, in_21, gm_n55, gm_n1674);
	nor (gm_n1676, gm_n90, gm_n78, in_9, gm_n1246, gm_n807);
	and (gm_n1677, gm_n166, gm_n129, in_18, gm_n1676);
	nor (gm_n1678, gm_n1677, gm_n1675, gm_n1673);
	or (gm_n1679, gm_n147, gm_n78, in_9, gm_n1125);
	nor (gm_n1680, gm_n105, gm_n72, gm_n55, gm_n1679, gm_n620);
	or (gm_n1681, gm_n92, in_14, gm_n78, gm_n208, gm_n95);
	nor (gm_n1682, gm_n244, gm_n212, in_18, gm_n1681);
	or (gm_n1683, gm_n133, gm_n90, gm_n78, gm_n389, gm_n287);
	nor (gm_n1684, gm_n437, gm_n244, in_18, gm_n1683);
	nor (gm_n1685, gm_n1684, gm_n1682, gm_n1680);
	nand (gm_n1686, gm_n1670, gm_n1566, gm_n1564, gm_n1685, gm_n1678);
	nor (gm_n1687, gm_n430, in_13, gm_n62, gm_n743, gm_n431);
	nand (gm_n1688, gm_n339, gm_n72, in_17, gm_n1687, gm_n373);
	nand (gm_n1689, gm_n93, in_6, gm_n97, gm_n80, gm_n94);
	nor (gm_n1690, gm_n115, in_16, in_12, gm_n1689, gm_n385);
	nand (gm_n1691, gm_n138, in_21, in_20, gm_n1690);
	and (gm_n1692, gm_n454, gm_n81);
	and (gm_n1693, gm_n733, in_12, gm_n94, gm_n1692, gm_n264);
	nand (gm_n1694, gm_n72, in_20, in_16, gm_n1693, gm_n179);
	nand (gm_n1695, gm_n1694, gm_n1691, gm_n1688);
	and (gm_n1696, gm_n1614, gm_n60, gm_n63, gm_n1120, gm_n1398);
	nand (gm_n1697, gm_n72, gm_n85, gm_n56, gm_n1696, gm_n394);
	or (gm_n1698, gm_n234, gm_n194, gm_n94);
	nor (gm_n1699, in_14, gm_n76, gm_n59, gm_n1698, gm_n190);
	nand (gm_n1700, gm_n129, gm_n88, gm_n119, gm_n1699);
	nor (gm_n1701, gm_n271, gm_n60, in_11, gm_n643, gm_n282);
	nand (gm_n1702, in_21, gm_n85, gm_n56, gm_n1701, gm_n448);
	nand (gm_n1703, gm_n1702, gm_n1700, gm_n1697);
	nor (gm_n1704, gm_n1686, gm_n1562, gm_n1560, gm_n1703, gm_n1695);
	or (gm_n1705, gm_n818, gm_n76, in_9, gm_n502, gm_n358);
	nor (gm_n1706, gm_n103, in_21, in_17, gm_n1705, gm_n328);
	or (gm_n1707, gm_n431, gm_n76, in_9, gm_n503, gm_n443);
	nor (gm_n1708, gm_n479, gm_n72, gm_n55, gm_n1707, gm_n256);
	nor (gm_n1709, gm_n625, gm_n228, in_8);
	nand (gm_n1710, gm_n64, gm_n73, in_12, gm_n1709, gm_n949);
	nor (gm_n1711, gm_n496, in_21, gm_n85, gm_n1710);
	nor (gm_n1712, gm_n1711, gm_n1708, gm_n1706);
	and (gm_n1713, in_7, in_6, gm_n97, gm_n80, gm_n94);
	and (gm_n1714, gm_n1713, gm_n545, gm_n79);
	and (gm_n1715, gm_n806, gm_n164, gm_n119, gm_n1714);
	or (gm_n1716, gm_n223, gm_n68, gm_n94);
	or (gm_n1717, gm_n90, in_10, in_9, gm_n1716, gm_n467);
	nor (gm_n1718, gm_n841, gm_n165, gm_n119, gm_n1717);
	nand (gm_n1719, in_7, in_6, gm_n97, gm_n546, in_8);
	or (gm_n1720, gm_n114, in_16, gm_n59, gm_n1719, gm_n297);
	nor (gm_n1721, gm_n496, gm_n72, gm_n85, gm_n1720);
	nor (gm_n1722, gm_n1721, gm_n1718, gm_n1715);
	nand (gm_n1723, gm_n1704, gm_n1558, gm_n1556, gm_n1722, gm_n1712);
	nor (gm_n1724, gm_n358, in_13, gm_n62, gm_n344, gm_n866);
	nand (gm_n1725, gm_n102, in_21, in_17, gm_n1724, gm_n595);
	and (gm_n1726, gm_n335, in_14, in_10, gm_n793, gm_n1158);
	nand (gm_n1727, gm_n131, gm_n129, gm_n119, gm_n1726);
	nor (gm_n1728, gm_n406, in_13, in_9, gm_n481, gm_n443);
	nand (gm_n1729, gm_n523, gm_n72, gm_n55, gm_n1728, gm_n206);
	nand (gm_n1730, gm_n1729, gm_n1727, gm_n1725);
	or (gm_n1731, gm_n625, gm_n572, gm_n94);
	nor (gm_n1732, in_14, gm_n78, gm_n62, gm_n1731, gm_n369);
	nand (gm_n1733, gm_n245, gm_n164, gm_n119, gm_n1732);
	and (gm_n1734, gm_n76, in_9, gm_n94, gm_n1263, gm_n788);
	nand (gm_n1735, gm_n206, in_21, in_17, gm_n1734, gm_n1076);
	nor (gm_n1736, gm_n92, in_14, gm_n78, gm_n414, gm_n95);
	nand (gm_n1737, gm_n200, gm_n146, in_18, gm_n1736);
	nand (gm_n1738, gm_n1737, gm_n1735, gm_n1733);
	nor (gm_n1739, gm_n1723, gm_n1554, gm_n1552, gm_n1738, gm_n1730);
	nand (gm_n1740, gm_n281, gm_n143, gm_n60, gm_n1161, gm_n869);
	nor (gm_n1741, in_21, in_20, gm_n56, gm_n1740);
	nand (gm_n1742, gm_n90, gm_n78, gm_n62, gm_n884, gm_n713);
	nor (gm_n1743, gm_n244, gm_n841, in_18, gm_n1742);
	nand (gm_n1744, gm_n77, gm_n73, gm_n59, gm_n870, gm_n143);
	nor (gm_n1745, gm_n912, in_21, gm_n85, gm_n1744);
	nor (gm_n1746, gm_n1745, gm_n1743, gm_n1741);
	or (gm_n1747, gm_n313, gm_n208, in_13, gm_n438, gm_n406);
	nor (gm_n1748, gm_n312, in_21, in_17, gm_n1747);
	or (gm_n1749, gm_n297, gm_n59, in_8, gm_n417, gm_n319);
	nor (gm_n1750, gm_n72, in_20, gm_n73, gm_n1749, gm_n496);
	or (gm_n1751, gm_n202, gm_n195, gm_n94);
	nor (gm_n1752, gm_n220, gm_n155, in_12, gm_n1751);
	and (gm_n1753, in_21, gm_n85, in_19, gm_n1752, gm_n268);
	nor (gm_n1754, gm_n1753, gm_n1750, gm_n1748);
	nand (gm_n1755, gm_n1739, gm_n1550, gm_n1548, gm_n1754, gm_n1746);
	and (gm_n1756, gm_n64, in_12, in_8, gm_n455, gm_n733);
	nand (gm_n1757, in_21, in_20, in_16, gm_n1756, gm_n697);
	nor (gm_n1758, gm_n238, gm_n194, gm_n94);
	and (gm_n1759, gm_n233, gm_n75, gm_n60, gm_n1758, gm_n869);
	nand (gm_n1760, in_21, in_20, in_19, gm_n1759);
	and (gm_n1761, gm_n78, in_9, gm_n94, gm_n1496, gm_n1158);
	nand (gm_n1762, gm_n367, gm_n119, in_14, gm_n1761, gm_n436);
	nand (gm_n1763, gm_n1762, gm_n1760, gm_n1757);
	nor (gm_n1764, gm_n358, in_13, gm_n62, gm_n743, gm_n443);
	nand (gm_n1765, gm_n311, gm_n72, gm_n55, gm_n1764, gm_n595);
	nor (gm_n1766, gm_n148, gm_n99, gm_n76, gm_n442, gm_n375);
	nand (gm_n1767, gm_n206, gm_n72, in_17, gm_n1766);
	nor (gm_n1768, gm_n796, gm_n76, in_9, gm_n463, gm_n480);
	nand (gm_n1769, gm_n255, in_21, gm_n55, gm_n1768, gm_n327);
	nand (gm_n1770, gm_n1769, gm_n1767, gm_n1765);
	nor (gm_n1771, gm_n1755, gm_n1546, gm_n1544, gm_n1770, gm_n1763);
	or (gm_n1772, gm_n259, in_14, gm_n78, gm_n438, gm_n807);
	nor (gm_n1773, gm_n244, gm_n841, in_18, gm_n1772);
	or (gm_n1774, gm_n609, in_13, in_9, gm_n432, gm_n358);
	nor (gm_n1775, gm_n184, gm_n72, in_17, gm_n1774, gm_n374);
	nand (gm_n1776, gm_n154, in_16, gm_n59, gm_n1605, gm_n949);
	nor (gm_n1777, gm_n139, in_21, gm_n85, gm_n1776);
	nor (gm_n1778, gm_n1777, gm_n1775, gm_n1773);
	or (gm_n1779, gm_n115, gm_n73, in_12, gm_n648, gm_n220);
	nor (gm_n1780, gm_n384, gm_n72, gm_n85, gm_n1779);
	or (gm_n1781, gm_n92, in_14, gm_n78, gm_n491, gm_n286);
	nor (gm_n1782, gm_n437, gm_n824, gm_n119, gm_n1781);
	or (gm_n1783, gm_n155, gm_n74, in_15, gm_n1125, gm_n290);
	nor (gm_n1784, gm_n72, gm_n85, gm_n56, gm_n1783);
	nor (gm_n1785, gm_n1784, gm_n1782, gm_n1780);
	nand (gm_n1786, gm_n1771, gm_n1541, gm_n1539, gm_n1785, gm_n1778);
	nor (gm_n1787, gm_n461, gm_n121, gm_n76, gm_n775, gm_n370);
	nand (gm_n1788, gm_n311, in_21, in_17, gm_n1787);
	or (gm_n1789, gm_n63, gm_n78, gm_n62, gm_n463, gm_n1295);
	nor (gm_n1790, gm_n393, in_19, in_15, gm_n1789, gm_n764);
	nand (gm_n1791, gm_n1790, gm_n72, in_20);
	nor (gm_n1792, gm_n168, gm_n155, gm_n60, gm_n632, gm_n447);
	nand (gm_n1793, in_21, in_20, gm_n56, gm_n1792);
	nand (gm_n1794, gm_n1793, gm_n1791, gm_n1788);
	nand (gm_n1795, gm_n131, gm_n86, gm_n119, gm_n1020);
	nor (gm_n1796, gm_n818, gm_n76, in_9, gm_n463, gm_n442);
	nand (gm_n1797, gm_n104, in_21, gm_n55, gm_n1796, gm_n327);
	nor (gm_n1798, gm_n406, in_13, in_9, gm_n503, gm_n443);
	nand (gm_n1799, gm_n255, gm_n72, gm_n55, gm_n1798, gm_n373);
	nand (gm_n1800, gm_n1799, gm_n1797, gm_n1795);
	nor (gm_n1801, gm_n1786, gm_n1537, gm_n1535, gm_n1800, gm_n1794);
	or (gm_n1802, gm_n257, in_13, in_9, gm_n502, gm_n866);
	nor (gm_n1803, gm_n374, gm_n72, gm_n55, gm_n1802, gm_n375);
	or (gm_n1804, gm_n213, in_16, gm_n59, gm_n1125, gm_n220);
	nor (gm_n1805, gm_n262, in_21, gm_n85, gm_n1804);
	or (gm_n1806, gm_n430, gm_n76, in_9, gm_n621, gm_n442);
	nor (gm_n1807, gm_n388, in_21, gm_n55, gm_n1806, gm_n328);
	nor (gm_n1808, gm_n1807, gm_n1805, gm_n1803);
	nand (gm_n1809, gm_n64, gm_n73, in_12, gm_n586, gm_n77);
	nor (gm_n1810, gm_n219, gm_n72, gm_n85, gm_n1809);
	or (gm_n1811, gm_n359, in_13, gm_n62, gm_n502, gm_n442);
	nor (gm_n1812, gm_n183, in_21, in_17, gm_n1811, gm_n256);
	or (gm_n1813, gm_n147, gm_n90, in_10, gm_n389, gm_n349);
	nor (gm_n1814, gm_n246, gm_n244, in_18, gm_n1813);
	nor (gm_n1815, gm_n1814, gm_n1812, gm_n1810);
	nand (gm_n1816, gm_n1801, gm_n1533, gm_n1530, gm_n1815, gm_n1808);
	nor (gm_n1817, gm_n259, gm_n90, in_10, gm_n491, gm_n467);
	nand (gm_n1818, gm_n367, gm_n131, gm_n119, gm_n1817);
	nor (gm_n1819, gm_n133, in_14, in_10, gm_n349, gm_n208);
	nand (gm_n1820, gm_n88, gm_n86, in_18, gm_n1819);
	nor (gm_n1821, gm_n818, in_13, gm_n62, gm_n430, gm_n358);
	nand (gm_n1822, gm_n254, in_21, gm_n55, gm_n1821, gm_n255);
	nand (gm_n1823, gm_n1822, gm_n1820, gm_n1818);
	or (gm_n1824, gm_n93, in_6, gm_n97, gm_n215, in_8);
	nor (gm_n1825, gm_n90, in_10, gm_n62, gm_n1824, gm_n147);
	nand (gm_n1826, gm_n806, gm_n129, gm_n119, gm_n1825);
	nor (gm_n1827, in_14, gm_n78, in_9, gm_n399, gm_n362);
	nand (gm_n1828, gm_n166, gm_n86, in_18, gm_n1827);
	and (gm_n1829, gm_n449, in_15, gm_n63, gm_n1120, gm_n555);
	nand (gm_n1830, in_21, gm_n85, gm_n56, gm_n1829, gm_n281);
	nand (gm_n1831, gm_n1830, gm_n1828, gm_n1826);
	nor (gm_n1832, gm_n1816, gm_n1528, gm_n1526, gm_n1831, gm_n1823);
	nor (gm_n1833, gm_n90, gm_n76, in_12, gm_n1208, gm_n213);
	and (gm_n1834, gm_n146, gm_n88, in_18, gm_n1833);
	or (gm_n1835, gm_n461, gm_n76, gm_n62, gm_n503, gm_n344);
	nor (gm_n1836, gm_n105, in_21, gm_n55, gm_n1835, gm_n374);
	nand (gm_n1837, gm_n519, gm_n81, gm_n94);
	or (gm_n1838, gm_n90, in_10, gm_n62, gm_n1837, gm_n369);
	nor (gm_n1839, gm_n368, gm_n841, gm_n119, gm_n1838);
	nor (gm_n1840, gm_n1839, gm_n1836, gm_n1834);
	nor (gm_n1841, gm_n277, gm_n68, in_8);
	nand (gm_n1842, gm_n79, gm_n73, in_12, gm_n1841, gm_n275);
	nor (gm_n1843, gm_n781, gm_n72, in_20, gm_n1842);
	or (gm_n1844, gm_n148, gm_n90, gm_n78, gm_n526, gm_n362);
	nor (gm_n1845, gm_n211, gm_n89, gm_n119, gm_n1844);
	or (gm_n1846, gm_n133, in_14, gm_n78, gm_n438, gm_n208);
	nor (gm_n1847, gm_n437, gm_n244, gm_n119, gm_n1846);
	nor (gm_n1848, gm_n1847, gm_n1845, gm_n1843);
	nand (gm_n1849, gm_n1832, gm_n1523, gm_n1521, gm_n1848, gm_n1840);
	and (gm_n1850, gm_n1144, gm_n60, gm_n63, gm_n580, gm_n422);
	nand (gm_n1851, gm_n72, in_20, gm_n56, gm_n1850, gm_n281);
	nor (gm_n1852, gm_n667, gm_n76, gm_n62, gm_n345, gm_n257);
	nand (gm_n1853, gm_n120, gm_n72, gm_n55, gm_n1852, gm_n122);
	nor (gm_n1854, in_14, in_10, gm_n62, gm_n1284, gm_n92);
	nand (gm_n1855, gm_n146, gm_n131, gm_n119, gm_n1854);
	nand (gm_n1856, gm_n1855, gm_n1853, gm_n1851);
	nor (gm_n1857, gm_n609, gm_n76, in_9, gm_n743, gm_n480);
	nand (gm_n1858, gm_n122, gm_n72, gm_n55, gm_n1857, gm_n174);
	nand (gm_n1859, gm_n93, in_6, in_5, gm_n454, gm_n94);
	nor (gm_n1860, gm_n90, in_13, in_12, gm_n1859, gm_n263);
	nand (gm_n1861, gm_n806, gm_n129, in_18, gm_n1860);
	nor (gm_n1862, gm_n95, gm_n90, gm_n78, gm_n208, gm_n147);
	nand (gm_n1863, gm_n806, gm_n164, gm_n119, gm_n1862);
	nand (gm_n1864, gm_n1863, gm_n1861, gm_n1858);
	nor (gm_n1865, gm_n1849, gm_n1518, gm_n1516, gm_n1864, gm_n1856);
	nand (gm_n1866, gm_n1101, gm_n154, in_15, gm_n545, gm_n487);
	nor (gm_n1867, gm_n72, in_20, gm_n56, gm_n1866);
	nand (gm_n1868, gm_n90, in_10, in_9, gm_n1392, gm_n91);
	nor (gm_n1869, gm_n437, gm_n824, in_18, gm_n1868);
	nand (gm_n1870, gm_n79, gm_n73, gm_n59, gm_n1198, gm_n949);
	nor (gm_n1871, gm_n219, gm_n72, in_20, gm_n1870);
	nor (gm_n1872, gm_n1871, gm_n1869, gm_n1867);
	nand (gm_n1873, gm_n64, gm_n73, gm_n59, gm_n535, gm_n571);
	nor (gm_n1874, gm_n219, gm_n72, in_20, gm_n1873);
	nand (gm_n1875, gm_n61, in_16, in_12, gm_n672, gm_n143);
	nor (gm_n1876, gm_n58, gm_n72, gm_n85, gm_n1875);
	nand (gm_n1877, gm_n93, in_6, gm_n97, gm_n80, in_8);
	or (gm_n1878, gm_n115, in_16, in_12, gm_n1877, gm_n354);
	nor (gm_n1879, gm_n496, in_21, gm_n85, gm_n1878);
	nor (gm_n1880, gm_n1879, gm_n1876, gm_n1874);
	nand (gm_n1881, gm_n1865, gm_n1513, gm_n1511, gm_n1880, gm_n1872);
	nor (gm_n1882, gm_n406, gm_n76, gm_n62, gm_n621, gm_n443);
	nand (gm_n1883, gm_n206, gm_n72, in_17, gm_n1882, gm_n1076);
	nand (gm_n1884, in_7, gm_n124, gm_n97, gm_n134, in_8);
	nor (gm_n1885, gm_n514, gm_n76, gm_n62, gm_n1884, gm_n313);
	nand (gm_n1886, gm_n120, gm_n72, gm_n55, gm_n1885);
	nor (gm_n1887, gm_n282, gm_n60, gm_n63, gm_n764, gm_n283);
	nand (gm_n1888, in_21, in_20, in_19, gm_n1887, gm_n268);
	nand (gm_n1889, gm_n1888, gm_n1886, gm_n1883);
	or (gm_n1890, gm_n358, in_13, gm_n62, gm_n988, gm_n502);
	nor (gm_n1891, gm_n103, in_21, gm_n55, gm_n1890, gm_n256);
	nor (out_3, gm_n1889, gm_n1881, gm_n1509, gm_n1891);
	or (gm_n1893, gm_n247, gm_n90, in_10, gm_n389, gm_n362);
	nor (gm_n1894, gm_n531, gm_n167, in_18, gm_n1893);
	nand (gm_n1895, in_14, gm_n78, in_9, gm_n1416, gm_n532);
	nor (gm_n1896, gm_n167, gm_n130, in_18, gm_n1895);
	nor (gm_n1897, gm_n442, in_13, in_9, gm_n1132, gm_n463);
	nand (gm_n1898, gm_n104, in_21, gm_n55, gm_n1897, gm_n311);
	nor (gm_n1899, gm_n240, gm_n92, in_14, gm_n270);
	nand (gm_n1900, gm_n436, gm_n199, in_18, gm_n1899);
	or (gm_n1901, gm_n480, in_13, in_9, gm_n1583, gm_n463);
	nor (gm_n1902, gm_n103, in_21, gm_n55, gm_n1901, gm_n375);
	nand (gm_n1903, gm_n214, gm_n59, gm_n94, gm_n949, gm_n1379);
	nor (gm_n1904, in_21, gm_n85, in_16, gm_n1903, gm_n139);
	nand (gm_n1905, gm_n174, in_21, in_17, gm_n852, gm_n523);
	or (gm_n1906, gm_n572, gm_n67, gm_n94);
	or (gm_n1907, gm_n213, in_13, gm_n59, gm_n1906);
	or (gm_n1908, gm_n184, in_21, gm_n55, gm_n1907, gm_n620);
	nand (gm_n1909, gm_n77, gm_n73, in_12, gm_n838, gm_n222);
	nor (gm_n1910, gm_n139, gm_n72, gm_n85, gm_n1909);
	or (gm_n1911, gm_n155, in_16, gm_n59, gm_n1689, gm_n319);
	nor (gm_n1912, gm_n781, in_21, in_20, gm_n1911);
	nor (gm_n1913, gm_n358, in_13, gm_n62, gm_n345, gm_n667);
	nand (gm_n1914, gm_n104, gm_n72, in_17, gm_n1913, gm_n174);
	and (gm_n1915, gm_n316, in_13, in_9, gm_n1049, gm_n788);
	nand (gm_n1916, gm_n206, gm_n72, gm_n55, gm_n1915, gm_n405);
	nand (gm_n1917, gm_n171, in_15, in_11, gm_n869, gm_n756);
	nor (gm_n1918, in_21, gm_n85, in_19, gm_n1917, gm_n393);
	nand (gm_n1919, gm_n340, gm_n523, in_13, gm_n829, gm_n1345);
	nor (gm_n1920, gm_n103, in_21, gm_n55, gm_n1919);
	nor (gm_n1921, gm_n344, in_13, gm_n62, gm_n503, gm_n442);
	nand (gm_n1922, gm_n206, in_21, gm_n55, gm_n1921, gm_n339);
	or (gm_n1923, gm_n93, in_6, gm_n97, gm_n223, gm_n94);
	nor (gm_n1924, gm_n297, gm_n76, gm_n59, gm_n1923);
	nand (gm_n1925, gm_n523, in_21, in_17, gm_n1924, gm_n373);
	or (gm_n1926, in_13, gm_n62, gm_n94, gm_n981, gm_n442);
	nor (gm_n1927, gm_n103, in_21, in_17, gm_n1926, gm_n375);
	not (gm_n1928, gm_n605);
	and (gm_n1929, in_6, gm_n97, gm_n108, gm_n169, gm_n93);
	nand (gm_n1930, gm_n449, gm_n60, gm_n63, gm_n1929, gm_n1928);
	nor (gm_n1931, gm_n72, in_20, in_19, gm_n1930, gm_n393);
	nor (gm_n1932, gm_n263, in_13, in_12, gm_n292);
	nand (gm_n1933, gm_n311, in_21, in_17, gm_n1932, gm_n339);
	nor (gm_n1934, gm_n121, in_13, gm_n59, gm_n515, gm_n155);
	nand (gm_n1935, gm_n102, in_21, gm_n55, gm_n1934);
	or (gm_n1936, gm_n370, gm_n286, gm_n76, gm_n442);
	nor (gm_n1937, gm_n105, gm_n72, in_17, gm_n1936, gm_n441);
	nand (gm_n1938, gm_n61, gm_n59, gm_n94, gm_n69, gm_n64);
	nor (gm_n1939, in_21, gm_n85, in_16, gm_n1938, gm_n912);
	nor (gm_n1940, gm_n213, gm_n73, in_12, gm_n499, gm_n319);
	nand (gm_n1941, gm_n383, gm_n72, in_20, gm_n1940);
	nor (gm_n1942, gm_n78, in_9, in_8);
	and (gm_n1943, gm_n245, gm_n91, gm_n90, gm_n1942, gm_n756);
	nand (gm_n1944, gm_n1943, gm_n367, in_18);
	or (gm_n1945, gm_n1295, gm_n78, in_9, gm_n344, gm_n807);
	nor (gm_n1946, gm_n87, in_18, in_14, gm_n1945, gm_n89);
	nor (gm_n1947, gm_n141, gm_n68, in_8);
	nand (gm_n1948, gm_n61, gm_n73, gm_n59, gm_n1947, gm_n233);
	nor (gm_n1949, gm_n384, gm_n72, in_20, gm_n1948);
	nor (gm_n1950, gm_n514, in_13, in_9, gm_n1132, gm_n463);
	nand (gm_n1951, gm_n523, in_21, gm_n55, gm_n1950, gm_n206);
	nor (gm_n1952, gm_n430, gm_n76, gm_n62, gm_n1583, gm_n406);
	nand (gm_n1953, gm_n102, in_21, in_17, gm_n1952, gm_n523);
	or (gm_n1954, gm_n609, in_13, gm_n62, gm_n988, gm_n442);
	nor (gm_n1955, gm_n184, gm_n72, gm_n55, gm_n1954, gm_n620);
	nor (gm_n1956, gm_n103, in_21, in_17, gm_n1063, gm_n313);
	nor (gm_n1957, gm_n431, in_13, in_9, gm_n621, gm_n596);
	nand (gm_n1958, gm_n122, in_21, in_17, gm_n1957, gm_n327);
	and (gm_n1959, gm_n264, gm_n75, in_15, gm_n1605, gm_n545);
	nand (gm_n1960, gm_n72, gm_n85, in_19, gm_n1959);
	or (gm_n1961, gm_n359, gm_n76, in_9, gm_n502, gm_n442);
	nor (gm_n1962, gm_n105, in_21, gm_n55, gm_n1961, gm_n374);
	nand (gm_n1963, gm_n122, gm_n76, gm_n62, gm_n880, gm_n788);
	nor (gm_n1964, gm_n374, gm_n72, in_17, gm_n1963);
	nand (gm_n1965, gm_n93, in_6, gm_n97, gm_n546, in_8);
	nor (gm_n1966, gm_n760, gm_n297, gm_n60, gm_n1965);
	nand (gm_n1967, in_21, in_20, gm_n56, gm_n1966, gm_n281);
	nor (gm_n1968, gm_n431, gm_n76, gm_n62, gm_n621, gm_n502);
	nand (gm_n1969, gm_n122, in_21, gm_n55, gm_n1968, gm_n254);
	nor (gm_n1970, gm_n277, gm_n194, in_8);
	nand (gm_n1971, gm_n448, gm_n214, gm_n60, gm_n1970, gm_n1398);
	nor (gm_n1972, in_21, gm_n85, gm_n56, gm_n1971);
	nor (gm_n1973, gm_n358, in_13, in_9, gm_n503, gm_n430);
	nand (gm_n1974, gm_n254, gm_n72, gm_n55, gm_n1973, gm_n405);
	and (gm_n1975, gm_n110, gm_n76, gm_n62, gm_n1049, gm_n579);
	nand (gm_n1976, gm_n206, in_21, gm_n55, gm_n1975, gm_n255);
	nand (gm_n1977, gm_n1976, gm_n1974);
	and (gm_n1978, gm_n1067, gm_n304, in_8);
	nand (gm_n1979, gm_n106, gm_n76, in_9, gm_n1978);
	nor (gm_n1980, gm_n441, in_21, gm_n55, gm_n1979, gm_n375);
	nor (gm_n1981, gm_n103, in_21, gm_n55, gm_n1540, gm_n256);
	nand (gm_n1982, gm_n335, in_14, gm_n78, gm_n793, gm_n1011);
	nor (gm_n1983, gm_n244, gm_n841, gm_n119, gm_n1982);
	nor (gm_n1984, gm_n1980, gm_n1977, gm_n1972, gm_n1983, gm_n1981);
	or (gm_n1985, gm_n358, in_13, in_9, gm_n481, gm_n430);
	nor (gm_n1986, gm_n121, gm_n72, in_17, gm_n1985, gm_n620);
	or (gm_n1987, gm_n95, in_14, in_10, gm_n467, gm_n208);
	nor (gm_n1988, gm_n212, gm_n165, in_18, gm_n1987);
	not (gm_n1989, gm_n323);
	nor (gm_n1990, gm_n1989, gm_n130, in_18, gm_n784);
	nor (gm_n1991, gm_n1990, gm_n1988, gm_n1986);
	nand (gm_n1992, gm_n264, gm_n75, gm_n60, gm_n870, gm_n449);
	nor (gm_n1993, in_21, gm_n85, gm_n56, gm_n1992);
	nand (gm_n1994, gm_n143, gm_n73, in_12, gm_n1947, gm_n221);
	nor (gm_n1995, gm_n139, gm_n72, gm_n85, gm_n1994);
	nand (gm_n1996, in_14, in_10, gm_n62, gm_n825, gm_n91);
	nor (gm_n1997, gm_n437, gm_n824, gm_n119, gm_n1996);
	nor (gm_n1998, gm_n1997, gm_n1995, gm_n1993);
	nand (gm_n1999, gm_n1984, gm_n1969, gm_n1967, gm_n1998, gm_n1991);
	nor (gm_n2000, gm_n514, in_13, gm_n62, gm_n743, gm_n609);
	nand (gm_n2001, gm_n523, gm_n72, gm_n55, gm_n2000, gm_n254);
	nand (gm_n2002, in_7, in_6, gm_n97, gm_n546, gm_n94);
	nor (gm_n2003, in_14, gm_n78, in_9, gm_n2002, gm_n92);
	nand (gm_n2004, gm_n164, gm_n131, gm_n119, gm_n2003);
	nor (gm_n2005, gm_n269, gm_n115, in_15, gm_n855, gm_n290);
	nand (gm_n2006, in_21, in_20, in_19, gm_n2005);
	nand (gm_n2007, gm_n2006, gm_n2004, gm_n2001);
	nand (gm_n2008, gm_n93, in_6, gm_n97, gm_n519, gm_n94);
	nor (gm_n2009, in_14, gm_n78, in_9, gm_n2008, gm_n147);
	nand (gm_n2010, gm_n166, gm_n164, gm_n119, gm_n2009);
	nor (gm_n2011, in_14, in_10, in_9, gm_n1716, gm_n362);
	nand (gm_n2012, gm_n367, gm_n323, gm_n119, gm_n2011);
	nor (gm_n2013, gm_n141, gm_n68, in_8, gm_n643, gm_n213);
	nand (gm_n2014, gm_n348, gm_n166, gm_n119, gm_n2013);
	nand (gm_n2015, gm_n2014, gm_n2012, gm_n2010);
	nor (gm_n2016, gm_n1999, gm_n1964, gm_n1962, gm_n2015, gm_n2007);
	not (gm_n2017, gm_n1942);
	or (gm_n2018, gm_n764, in_15, in_11, gm_n2017, gm_n770);
	nor (gm_n2019, in_21, in_20, in_19, gm_n2018, gm_n447);
	or (gm_n2020, gm_n369, in_14, in_10, gm_n438, gm_n389);
	nor (gm_n2021, gm_n246, gm_n211, in_18, gm_n2020);
	or (gm_n2022, gm_n406, gm_n76, gm_n62, gm_n502, gm_n432);
	nor (gm_n2023, gm_n479, in_21, in_17, gm_n2022, gm_n256);
	nor (gm_n2024, gm_n2023, gm_n2021, gm_n2019);
	or (gm_n2025, gm_n480, gm_n76, gm_n62, gm_n1583, gm_n443);
	nor (gm_n2026, gm_n479, in_21, in_17, gm_n2025, gm_n313);
	or (gm_n2027, gm_n293, gm_n155, in_15, gm_n887, gm_n633);
	nor (gm_n2028, in_21, gm_n85, gm_n56, gm_n2027);
	nand (gm_n2029, gm_n454, gm_n304, in_8);
	or (gm_n2030, gm_n190, gm_n73, in_12, gm_n2029, gm_n354);
	nor (gm_n2031, gm_n384, in_21, in_20, gm_n2030);
	nor (gm_n2032, gm_n2031, gm_n2028, gm_n2026);
	nand (gm_n2033, gm_n2016, gm_n1960, gm_n1958, gm_n2032, gm_n2024);
	nor (gm_n2034, gm_n95, in_14, in_10, gm_n526, gm_n369);
	nand (gm_n2035, gm_n199, gm_n131, in_18, gm_n2034);
	nor (gm_n2036, gm_n148, in_14, in_10, gm_n589, gm_n467);
	nand (gm_n2037, gm_n245, gm_n86, gm_n119, gm_n2036);
	nand (gm_n2038, in_7, in_6, gm_n97, gm_n519, gm_n94);
	nor (gm_n2039, gm_n227, gm_n73, gm_n59, gm_n2038, gm_n158);
	nand (gm_n2040, gm_n495, in_21, in_20, gm_n2039);
	nand (gm_n2041, gm_n2040, gm_n2037, gm_n2035);
	and (gm_n2042, gm_n185, gm_n1157, gm_n76, gm_n722, gm_n339);
	nand (gm_n2043, gm_n327, gm_n72, in_17, gm_n2042);
	nor (gm_n2044, gm_n461, gm_n76, gm_n62, gm_n463, gm_n359);
	nand (gm_n2045, gm_n102, gm_n72, in_17, gm_n2044, gm_n595);
	nand (gm_n2046, gm_n199, gm_n131, gm_n119, gm_n1699);
	nand (gm_n2047, gm_n2046, gm_n2045, gm_n2043);
	nor (gm_n2048, gm_n2033, gm_n1956, gm_n1955, gm_n2047, gm_n2041);
	or (gm_n2049, gm_n95, in_14, gm_n78, gm_n248, gm_n207);
	nor (gm_n2050, gm_n1989, gm_n165, gm_n119, gm_n2049);
	or (gm_n2051, gm_n309, gm_n56, in_15, gm_n633, gm_n447);
	nor (gm_n2052, gm_n2051, in_21, in_20);
	or (gm_n2053, gm_n430, in_13, in_9, gm_n442, gm_n796);
	nor (gm_n2054, gm_n121, gm_n72, gm_n55, gm_n2053, gm_n388);
	nor (gm_n2055, gm_n2054, gm_n2052, gm_n2050);
	nand (gm_n2056, gm_n555, in_15, in_11, gm_n869, gm_n576);
	nor (gm_n2057, in_21, gm_n85, in_19, gm_n2056, gm_n1331);
	nand (gm_n2058, gm_n154, in_16, in_12, gm_n1605, gm_n949);
	nor (gm_n2059, gm_n384, in_21, in_20, gm_n2058);
	or (gm_n2060, gm_n93, in_6, gm_n97, gm_n238, in_8);
	or (gm_n2061, gm_n227, in_16, gm_n59, gm_n2060, gm_n213);
	nor (gm_n2062, gm_n496, in_21, in_20, gm_n2061);
	nor (gm_n2063, gm_n2062, gm_n2059, gm_n2057);
	nand (gm_n2064, gm_n2048, gm_n1953, gm_n1951, gm_n2063, gm_n2055);
	nor (gm_n2065, gm_n93, in_6, gm_n97, gm_n201, in_8);
	and (gm_n2066, gm_n379, gm_n233, gm_n60, gm_n2065, gm_n449);
	nand (gm_n2067, gm_n72, in_20, in_19, gm_n2066);
	nor (gm_n2068, gm_n344, gm_n76, gm_n62, gm_n1132, gm_n442);
	nand (gm_n2069, gm_n405, in_21, in_17, gm_n2068, gm_n327);
	nor (gm_n2070, gm_n93, in_6, gm_n97, gm_n215, gm_n94);
	and (gm_n2071, gm_n61, in_16, in_12, gm_n2070, gm_n233);
	nand (gm_n2072, gm_n383, in_21, gm_n85, gm_n2071);
	nand (gm_n2073, gm_n2072, gm_n2069, gm_n2067);
	and (gm_n2074, gm_n124, in_5, in_4, gm_n175, in_7);
	and (gm_n2075, gm_n449, in_15, gm_n63, gm_n2074, gm_n555);
	nand (gm_n2076, gm_n72, in_20, in_19, gm_n2075, gm_n486);
	nand (gm_n2077, gm_n93, gm_n124, in_5, gm_n519, gm_n94);
	nor (gm_n2078, gm_n369, gm_n78, in_9, gm_n2077);
	nand (gm_n2079, gm_n104, in_21, gm_n55, gm_n2078, gm_n206);
	or (gm_n2080, gm_n223, gm_n68, in_8);
	nor (gm_n2081, gm_n213, gm_n73, in_12, gm_n2080, gm_n276);
	nand (gm_n2082, gm_n383, gm_n72, gm_n85, gm_n2081);
	nand (gm_n2083, gm_n2082, gm_n2079, gm_n2076);
	nor (gm_n2084, gm_n2064, gm_n1949, gm_n1946, gm_n2083, gm_n2073);
	or (gm_n2085, gm_n442, in_13, gm_n62, gm_n502, gm_n481);
	nor (gm_n2086, gm_n313, gm_n72, in_17, gm_n2085, gm_n620);
	or (gm_n2087, gm_n406, in_13, in_9, gm_n443, gm_n432);
	nor (gm_n2088, gm_n184, gm_n72, gm_n55, gm_n2087, gm_n388);
	or (gm_n2089, gm_n667, in_13, gm_n62, gm_n621, gm_n461);
	nor (gm_n2090, gm_n620, in_21, gm_n55, gm_n2089, gm_n375);
	nor (gm_n2091, gm_n2090, gm_n2088, gm_n2086);
	nand (gm_n2092, gm_n192, gm_n60, gm_n63, gm_n1120, gm_n555);
	nor (gm_n2093, gm_n72, in_20, in_19, gm_n2092, gm_n293);
	or (gm_n2094, gm_n213, in_13, gm_n59, gm_n1223);
	nor (gm_n2095, gm_n103, in_21, in_17, gm_n2094, gm_n662);
	nor (gm_n2096, gm_n215, gm_n68, in_8);
	nand (gm_n2097, gm_n275, gm_n233, gm_n59, gm_n2096);
	nor (gm_n2098, gm_n72, gm_n85, gm_n56, gm_n2097, gm_n447);
	nor (gm_n2099, gm_n2098, gm_n2095, gm_n2093);
	nand (gm_n2100, gm_n2084, gm_n1944, gm_n1941, gm_n2099, gm_n2091);
	and (gm_n2101, gm_n449, gm_n60, gm_n63, gm_n601, gm_n555);
	nand (gm_n2102, in_21, gm_n85, in_19, gm_n2101, gm_n448);
	nor (gm_n2103, gm_n220, gm_n191, in_12, gm_n765, gm_n263);
	nand (gm_n2104, in_21, in_20, in_19, gm_n2103);
	and (gm_n2105, gm_n1345, gm_n255, in_13, gm_n829, gm_n402);
	nand (gm_n2106, gm_n311, in_21, in_17, gm_n2105);
	nand (gm_n2107, gm_n2106, gm_n2104, gm_n2102);
	and (gm_n2108, gm_n61, in_16, gm_n59, gm_n1970, gm_n143);
	nand (gm_n2109, gm_n697, in_21, gm_n85, gm_n2108);
	nor (gm_n2110, gm_n115, gm_n73, gm_n59, gm_n468, gm_n220);
	nand (gm_n2111, gm_n113, gm_n72, in_20, gm_n2110);
	nor (gm_n2112, gm_n220, gm_n73, gm_n59, gm_n1923, gm_n263);
	nand (gm_n2113, gm_n138, in_21, in_20, gm_n2112);
	nand (gm_n2114, gm_n2113, gm_n2111, gm_n2109);
	nor (gm_n2115, gm_n2100, gm_n1939, gm_n1937, gm_n2114, gm_n2107);
	or (gm_n2116, gm_n609, gm_n76, gm_n62, gm_n1583, gm_n461);
	nor (gm_n2117, gm_n121, in_21, gm_n55, gm_n2116, gm_n479);
	or (gm_n2118, gm_n344, gm_n76, in_9, gm_n481, gm_n442);
	nor (gm_n2119, gm_n662, in_21, gm_n55, gm_n2118, gm_n374);
	or (gm_n2120, gm_n213, gm_n73, gm_n59, gm_n1751, gm_n385);
	nor (gm_n2121, gm_n496, gm_n72, in_20, gm_n2120);
	nor (gm_n2122, gm_n2121, gm_n2119, gm_n2117);
	or (gm_n2123, gm_n90, gm_n78, gm_n62, gm_n562, gm_n467);
	nor (gm_n2124, gm_n246, gm_n165, gm_n119, gm_n2123);
	nand (gm_n2125, gm_n802, gm_n81, in_8);
	or (gm_n2126, gm_n633, gm_n297, in_15, gm_n2125);
	nor (gm_n2127, gm_n72, in_20, gm_n56, gm_n2126, gm_n393);
	nand (gm_n2128, gm_n422, gm_n214, in_15, gm_n1970, gm_n448);
	nor (gm_n2129, gm_n72, gm_n85, gm_n56, gm_n2128);
	nor (gm_n2130, gm_n2129, gm_n2127, gm_n2124);
	nand (gm_n2131, gm_n2115, gm_n1935, gm_n1933, gm_n2130, gm_n2122);
	nor (gm_n2132, gm_n263, gm_n168, gm_n60, gm_n2029, gm_n393);
	nand (gm_n2133, gm_n72, in_20, gm_n56, gm_n2132);
	nor (gm_n2134, in_14, in_13, in_12, gm_n1859, gm_n190);
	nand (gm_n2135, gm_n348, gm_n88, gm_n119, gm_n2134);
	nor (gm_n2136, gm_n257, in_13, gm_n62, gm_n503, gm_n596);
	nand (gm_n2137, gm_n523, in_21, gm_n55, gm_n2136, gm_n254);
	nand (gm_n2138, gm_n2137, gm_n2135, gm_n2133);
	nor (gm_n2139, gm_n193, gm_n297, gm_n60, gm_n1191, gm_n447);
	nand (gm_n2140, gm_n72, gm_n85, gm_n56, gm_n2139);
	nor (gm_n2141, gm_n95, gm_n90, gm_n78, gm_n389, gm_n207);
	nand (gm_n2142, gm_n367, gm_n806, gm_n119, gm_n2141);
	nor (gm_n2143, gm_n155, gm_n73, gm_n59, gm_n654, gm_n385);
	nand (gm_n2144, gm_n697, in_21, in_20, gm_n2143);
	nand (gm_n2145, gm_n2144, gm_n2142, gm_n2140);
	nor (gm_n2146, gm_n2131, gm_n1931, gm_n1927, gm_n2145, gm_n2138);
	and (gm_n2147, gm_n264, gm_n76, gm_n59, gm_n1095);
	and (gm_n2148, gm_n523, in_21, gm_n55, gm_n2147, gm_n327);
	or (gm_n2149, gm_n609, in_13, gm_n62, gm_n1583, gm_n442);
	nor (gm_n2150, gm_n103, gm_n72, in_17, gm_n2149, gm_n313);
	nand (gm_n2151, in_10, gm_n62, in_8, gm_n714, gm_n532);
	nor (gm_n2152, gm_n87, in_18, in_14, gm_n2151, gm_n132);
	nor (gm_n2153, gm_n2152, gm_n2150, gm_n2148);
	or (gm_n2154, gm_n290, gm_n274, gm_n60, gm_n1324, gm_n393);
	nor (gm_n2155, gm_n72, gm_n85, gm_n56, gm_n2154);
	nor (gm_n2156, gm_n388, in_21, gm_n55, gm_n317, gm_n313);
	or (gm_n2157, gm_n362, in_14, gm_n78, gm_n526, gm_n438);
	nor (gm_n2158, gm_n244, gm_n132, gm_n119, gm_n2157);
	nor (gm_n2159, gm_n2158, gm_n2156, gm_n2155);
	nand (gm_n2160, gm_n2146, gm_n1925, gm_n1922, gm_n2159, gm_n2153);
	nor (gm_n2161, gm_n90, in_10, in_9, gm_n799, gm_n133);
	nand (gm_n2162, gm_n367, gm_n166, gm_n119, gm_n2161);
	nor (gm_n2163, gm_n328, gm_n76, in_9, gm_n1481, gm_n406);
	nand (gm_n2164, gm_n174, gm_n72, gm_n55, gm_n2163);
	nor (gm_n2165, gm_n406, gm_n76, gm_n62, gm_n359, gm_n344);
	nand (gm_n2166, gm_n311, in_21, in_17, gm_n2165, gm_n595);
	nand (gm_n2167, gm_n2166, gm_n2164, gm_n2162);
	nor (gm_n2168, gm_n430, gm_n76, in_9, gm_n597, gm_n431);
	nand (gm_n2169, gm_n311, gm_n72, in_17, gm_n2168, gm_n339);
	and (gm_n2170, gm_n1144, in_15, in_11, gm_n1615, gm_n449);
	nand (gm_n2171, gm_n72, in_20, gm_n56, gm_n2170, gm_n448);
	nor (gm_n2172, gm_n671, gm_n194, in_8);
	and (gm_n2173, gm_n143, gm_n73, in_12, gm_n2172, gm_n275);
	nand (gm_n2174, gm_n179, gm_n72, gm_n85, gm_n2173);
	nand (gm_n2175, gm_n2174, gm_n2171, gm_n2169);
	nor (gm_n2176, gm_n2160, gm_n1920, gm_n1918, gm_n2175, gm_n2167);
	or (gm_n2177, gm_n115, in_16, gm_n59, gm_n1751, gm_n319);
	nor (gm_n2178, gm_n139, gm_n72, in_20, gm_n2177);
	or (gm_n2179, gm_n667, gm_n76, in_9, gm_n257, gm_n796);
	nor (gm_n2180, gm_n662, gm_n72, in_17, gm_n2179, gm_n374);
	or (gm_n2181, gm_n609, in_13, in_9, gm_n345, gm_n461);
	nor (gm_n2182, gm_n183, in_21, gm_n55, gm_n2181, gm_n256);
	nor (gm_n2183, gm_n2182, gm_n2180, gm_n2178);
	nand (gm_n2184, gm_n532, in_14, gm_n78, gm_n793, gm_n721);
	nor (gm_n2185, gm_n132, gm_n130, gm_n119, gm_n2184);
	nand (gm_n2186, gm_n555, gm_n192, gm_n63, gm_n1615);
	nor (gm_n2187, gm_n1989, gm_n824, gm_n119, gm_n2186);
	nand (gm_n2188, gm_n61, gm_n73, gm_n59, gm_n82, gm_n79);
	nor (gm_n2189, gm_n139, gm_n72, gm_n85, gm_n2188);
	nor (gm_n2190, gm_n2189, gm_n2187, gm_n2185);
	nand (gm_n2191, gm_n2176, gm_n1916, gm_n1914, gm_n2190, gm_n2183);
	nand (gm_n2192, in_2, in_1, in_0);
	nor (gm_n2193, in_5, gm_n108, in_3, gm_n2192, gm_n124);
	and (gm_n2194, gm_n2193, gm_n90, gm_n78, gm_n490, gm_n532);
	nand (gm_n2195, gm_n436, gm_n129, in_18, gm_n2194);
	nor (gm_n2196, gm_n461, gm_n76, gm_n62, gm_n345, gm_n596);
	nand (gm_n2197, gm_n102, gm_n72, in_17, gm_n2196, gm_n255);
	nand (gm_n2198, gm_n519, gm_n304, in_8);
	nor (gm_n2199, gm_n115, gm_n73, in_12, gm_n2198, gm_n276);
	nand (gm_n2200, gm_n179, gm_n72, gm_n85, gm_n2199);
	nand (gm_n2201, gm_n2200, gm_n2197, gm_n2195);
	and (gm_n2202, gm_n187, in_13, in_9, gm_n341, gm_n314);
	nand (gm_n2203, gm_n174, gm_n72, in_17, gm_n2202, gm_n339);
	and (gm_n2204, gm_n143, in_16, in_12, gm_n1456, gm_n221);
	nand (gm_n2205, gm_n138, gm_n72, gm_n85, gm_n2204);
	nor (gm_n2206, gm_n297, gm_n76, gm_n59, gm_n515);
	nand (gm_n2207, gm_n122, in_21, in_17, gm_n2206, gm_n206);
	nand (gm_n2208, gm_n2207, gm_n2205, gm_n2203);
	nor (gm_n2209, gm_n2191, gm_n1912, gm_n1910, gm_n2208, gm_n2201);
	nand (gm_n2210, gm_n104, gm_n76, in_9, gm_n1978, gm_n402);
	nor (gm_n2211, gm_n479, in_21, in_17, gm_n2210);
	nand (gm_n2212, gm_n314, gm_n104, gm_n76, gm_n829, gm_n1345);
	nor (gm_n2213, gm_n103, in_21, gm_n55, gm_n2212);
	nor (gm_n2214, gm_n105, gm_n72, gm_n55, gm_n1979, gm_n312);
	nor (gm_n2215, gm_n2214, gm_n2213, gm_n2211);
	or (gm_n2216, gm_n290, gm_n158, gm_n60, gm_n1689, gm_n447);
	nor (gm_n2217, in_21, in_20, gm_n56, gm_n2216);
	nor (gm_n2218, gm_n277, gm_n202, gm_n94);
	nand (gm_n2219, gm_n77, gm_n73, gm_n59, gm_n2218, gm_n233);
	nor (gm_n2220, gm_n262, gm_n72, in_20, gm_n2219);
	or (gm_n2221, gm_n228, gm_n201, in_8);
	or (gm_n2222, gm_n114, gm_n73, in_12, gm_n2221, gm_n274);
	nor (gm_n2223, gm_n384, in_21, gm_n85, gm_n2222);
	nor (gm_n2224, gm_n2223, gm_n2220, gm_n2217);
	nand (gm_n2225, gm_n2209, gm_n1908, gm_n1905, gm_n2224, gm_n2215);
	nor (gm_n2226, gm_n263, gm_n74, in_15, gm_n1519, gm_n764);
	nand (gm_n2227, gm_n72, in_20, in_19, gm_n2226);
	nor (gm_n2228, gm_n609, in_13, gm_n62, gm_n743, gm_n257);
	nand (gm_n2229, gm_n254, gm_n72, in_17, gm_n2228, gm_n339);
	and (gm_n2230, gm_n93, in_6, gm_n97, gm_n454, gm_n94);
	and (gm_n2231, gm_n233, gm_n73, in_12, gm_n2230, gm_n733);
	nand (gm_n2232, gm_n113, in_21, gm_n85, gm_n2231);
	nand (gm_n2233, gm_n2232, gm_n2229, gm_n2227);
	not (gm_n2234, gm_n502);
	and (gm_n2235, gm_n126, in_13, in_9, gm_n2234, gm_n314);
	nand (gm_n2236, gm_n122, in_21, gm_n55, gm_n2235, gm_n311);
	or (gm_n2237, in_7, in_6, in_5, gm_n671);
	nor (gm_n2238, in_13, in_9, gm_n94, gm_n2237, gm_n257);
	nand (gm_n2239, gm_n102, gm_n72, gm_n55, gm_n2238, gm_n104);
	nor (gm_n2240, gm_n541, gm_n168, in_11, gm_n842);
	nand (gm_n2241, gm_n199, gm_n88, in_18, gm_n2240);
	nand (gm_n2242, gm_n2241, gm_n2239, gm_n2236);
	nor (gm_n2243, gm_n2225, gm_n1904, gm_n1902, gm_n2242, gm_n2233);
	or (gm_n2244, gm_n671, gm_n228, in_8);
	or (gm_n2245, gm_n290, gm_n213, in_15, gm_n2244, gm_n293);
	nor (gm_n2246, in_21, in_20, in_19, gm_n2245);
	or (gm_n2247, gm_n227, in_16, gm_n59, gm_n657, gm_n263);
	nor (gm_n2248, gm_n781, in_21, in_20, gm_n2247);
	or (gm_n2249, gm_n430, in_13, in_9, gm_n743, gm_n480);
	nor (gm_n2250, gm_n312, gm_n72, gm_n55, gm_n2249, gm_n375);
	nor (gm_n2251, gm_n2250, gm_n2248, gm_n2246);
	nand (gm_n2252, gm_n170, in_15, in_11, gm_n602, gm_n422);
	nor (gm_n2253, in_21, in_20, gm_n56, gm_n2252, gm_n191);
	or (gm_n2254, gm_n667, in_13, in_9, gm_n597, gm_n480);
	nor (gm_n2255, gm_n441, in_21, in_17, gm_n2254, gm_n256);
	nand (gm_n2256, gm_n93, in_6, in_5, gm_n519, gm_n94);
	or (gm_n2257, gm_n328, in_13, in_9, gm_n2256, gm_n480);
	nor (gm_n2258, gm_n479, in_21, in_17, gm_n2257);
	nor (gm_n2259, gm_n2258, gm_n2255, gm_n2253);
	nand (gm_n2260, gm_n2243, gm_n1900, gm_n1898, gm_n2259, gm_n2251);
	and (gm_n2261, in_10, in_9, in_8, gm_n532, gm_n69);
	nand (gm_n2262, gm_n245, in_18, in_14, gm_n2261, gm_n348);
	nor (gm_n2263, gm_n274, gm_n74, gm_n60, gm_n2002, gm_n764);
	nand (gm_n2264, gm_n72, gm_n85, in_19, gm_n2263);
	nor (gm_n2265, gm_n514, in_13, in_9, gm_n988, gm_n596);
	nand (gm_n2266, gm_n122, gm_n72, gm_n55, gm_n2265, gm_n327);
	nand (gm_n2267, gm_n2266, gm_n2264, gm_n2262);
	nor (gm_n2268, gm_n90, in_13, gm_n59, gm_n855, gm_n263);
	nand (gm_n2269, gm_n200, gm_n129, gm_n119, gm_n2268);
	nor (gm_n2270, gm_n485, gm_n190, gm_n60, gm_n764, gm_n499);
	nand (gm_n2271, in_21, in_20, gm_n56, gm_n2270);
	nor (gm_n2272, gm_n95, in_14, gm_n78, gm_n369, gm_n350);
	nand (gm_n2273, gm_n323, gm_n164, gm_n119, gm_n2272);
	nand (gm_n2274, gm_n2273, gm_n2271, gm_n2269);
	nor (out_4, gm_n2260, gm_n1896, gm_n1894, gm_n2274, gm_n2267);
	nor (gm_n2276, gm_n202, gm_n141, in_8);
	nand (gm_n2277, gm_n90, in_10, in_9, gm_n2276, gm_n334);
	nor (gm_n2278, gm_n244, gm_n89, gm_n119, gm_n2277);
	nor (gm_n2279, gm_n76, gm_n62, in_8, gm_n417, gm_n406);
	nand (gm_n2280, gm_n311, gm_n72, gm_n55, gm_n2279, gm_n405);
	or (gm_n2281, gm_n92, gm_n90, in_10, gm_n491, gm_n350);
	nor (gm_n2282, gm_n368, gm_n212, in_18, gm_n2281);
	nor (gm_n2283, gm_n671, gm_n202, in_8);
	nand (gm_n2284, gm_n379, gm_n79, in_15, gm_n2283, gm_n449);
	nor (gm_n2285, in_21, gm_n85, gm_n56, gm_n2284);
	nor (gm_n2286, gm_n247, gm_n208, gm_n78, gm_n467);
	nand (gm_n2287, gm_n523, in_21, gm_n55, gm_n2286, gm_n206);
	nor (gm_n2288, gm_n461, gm_n121, in_13, gm_n350, gm_n287);
	nand (gm_n2289, gm_n373, gm_n72, gm_n55, gm_n2288);
	nand (gm_n2290, gm_n422, gm_n214, in_15, gm_n1531, gm_n486);
	nor (gm_n2291, gm_n72, gm_n85, in_19, gm_n2290);
	nand (gm_n2292, gm_n142, gm_n73, gm_n59, gm_n303, gm_n264);
	nor (gm_n2293, gm_n139, in_21, gm_n85, gm_n2292);
	nor (gm_n2294, gm_n406, in_13, gm_n62, gm_n481, gm_n463);
	nand (gm_n2295, gm_n311, gm_n72, in_17, gm_n2294, gm_n405);
	nor (gm_n2296, in_14, gm_n78, in_9, gm_n499, gm_n133);
	nand (gm_n2297, gm_n436, gm_n199, in_18, gm_n2296);
	nand (gm_n2298, gm_n392, gm_n143, gm_n60, gm_n486, gm_n411);
	nor (gm_n2299, in_21, in_20, gm_n56, gm_n2298);
	nand (gm_n2300, gm_n77, in_16, gm_n59, gm_n1416, gm_n264);
	nor (gm_n2301, gm_n496, in_21, gm_n85, gm_n2300);
	and (gm_n2302, gm_n90, gm_n78, gm_n62, gm_n1524, gm_n624);
	nand (gm_n2303, gm_n436, gm_n129, in_18, gm_n2302);
	nor (gm_n2304, gm_n155, gm_n73, in_12, gm_n385, gm_n180);
	nand (gm_n2305, gm_n383, in_21, gm_n85, gm_n2304);
	or (gm_n2306, gm_n485, gm_n263, in_15, gm_n760, gm_n654);
	nor (gm_n2307, in_21, in_20, gm_n56, gm_n2306);
	or (gm_n2308, gm_n667, gm_n76, gm_n62, gm_n480, gm_n796);
	nor (gm_n2309, gm_n183, gm_n72, gm_n55, gm_n2308, gm_n184);
	nor (gm_n2310, gm_n207, gm_n977, in_14, gm_n572, gm_n215);
	nand (gm_n2311, gm_n367, gm_n166, gm_n119, gm_n2310);
	nor (gm_n2312, gm_n92, in_14, in_10, gm_n259, gm_n148);
	nand (gm_n2313, gm_n243, gm_n131, in_18, gm_n2312);
	or (gm_n2314, gm_n430, gm_n76, gm_n62, gm_n743, gm_n480);
	nor (gm_n2315, gm_n121, gm_n72, gm_n55, gm_n2314, gm_n374);
	and (gm_n2316, gm_n255, in_21, gm_n55, gm_n2078, gm_n327);
	nor (gm_n2317, gm_n344, in_13, in_9, gm_n988, gm_n480);
	nand (gm_n2318, gm_n254, gm_n72, in_17, gm_n2317, gm_n339);
	nor (gm_n2319, gm_n514, gm_n76, in_9, gm_n1132, gm_n344);
	nand (gm_n2320, gm_n311, in_21, in_17, gm_n2319, gm_n339);
	or (gm_n2321, gm_n514, in_13, in_9, gm_n1132, gm_n443);
	nor (gm_n2322, gm_n105, in_21, in_17, gm_n2321, gm_n312);
	nand (gm_n2323, gm_n187, in_13, gm_n62, gm_n402, gm_n341);
	nor (gm_n2324, gm_n441, in_21, in_17, gm_n2323, gm_n662);
	and (gm_n2325, gm_n125, gm_n76, gm_n62, gm_n402, gm_n126);
	nand (gm_n2326, gm_n102, gm_n72, gm_n55, gm_n2325, gm_n255);
	nor (gm_n2327, gm_n514, gm_n76, in_9, gm_n463, gm_n866);
	nand (gm_n2328, gm_n311, in_21, gm_n55, gm_n2327, gm_n1076);
	nand (gm_n2329, gm_n1101, gm_n79, gm_n60, gm_n869, gm_n547);
	nor (gm_n2330, gm_n72, gm_n85, in_19, gm_n2329);
	nand (gm_n2331, gm_n214, gm_n73, gm_n59, gm_n547, gm_n949);
	nor (gm_n2332, gm_n781, in_21, gm_n85, gm_n2331);
	or (gm_n2333, gm_n223, gm_n194, in_8);
	nor (gm_n2334, in_14, gm_n78, in_9, gm_n2333, gm_n207);
	nand (gm_n2335, gm_n164, gm_n131, in_18, gm_n2334);
	nor (gm_n2336, gm_n152, in_16, gm_n59, gm_n932, gm_n155);
	nand (gm_n2337, gm_n138, in_21, gm_n85, gm_n2336);
	or (gm_n2338, in_14, gm_n78, in_9, gm_n648, gm_n207);
	nor (gm_n2339, gm_n824, gm_n167, gm_n119, gm_n2338);
	or (gm_n2340, gm_n93, in_6, gm_n97, gm_n67, in_8);
	or (gm_n2341, gm_n90, gm_n78, in_9, gm_n2340, gm_n147);
	nor (gm_n2342, gm_n132, gm_n87, gm_n119, gm_n2341);
	nor (gm_n2343, gm_n90, in_10, gm_n62, gm_n1176, gm_n133);
	nand (gm_n2344, gm_n323, gm_n129, gm_n119, gm_n2343);
	nand (gm_n2345, gm_n436, gm_n348, gm_n119, gm_n655);
	and (gm_n2346, gm_n802, gm_n291, gm_n94);
	nand (gm_n2347, gm_n104, in_13, gm_n62, gm_n2346, gm_n788);
	nor (gm_n2348, gm_n103, in_21, gm_n55, gm_n2347);
	nand (gm_n2349, gm_n755, gm_n60, in_11, gm_n756, gm_n422);
	nor (gm_n2350, gm_n72, in_20, gm_n56, gm_n2349, gm_n447);
	and (gm_n2351, gm_n90, in_13, gm_n59, gm_n216, gm_n143);
	nand (gm_n2352, gm_n348, gm_n166, gm_n119, gm_n2351);
	nor (gm_n2353, gm_n297, gm_n74, gm_n60, gm_n887, gm_n193);
	nand (gm_n2354, gm_n72, gm_n85, gm_n56, gm_n2353);
	nor (gm_n2355, gm_n147, gm_n90, in_10, gm_n376, gm_n287);
	nand (gm_n2356, gm_n436, gm_n129, gm_n119, gm_n2355);
	or (gm_n2357, gm_n194, gm_n67, in_8);
	nor (gm_n2358, gm_n155, gm_n73, in_12, gm_n2357, gm_n220);
	nand (gm_n2359, gm_n383, gm_n72, gm_n85, gm_n2358);
	nor (gm_n2360, gm_n257, gm_n76, gm_n62, gm_n1132, gm_n463);
	nand (gm_n2361, gm_n339, gm_n72, in_17, gm_n2360, gm_n373);
	nand (gm_n2362, gm_n2356, gm_n2354, gm_n2352, gm_n2361, gm_n2359);
	nor (gm_n2363, gm_n133, in_14, in_10, gm_n247, gm_n208);
	nand (gm_n2364, gm_n323, gm_n129, gm_n119, gm_n2363);
	nor (gm_n2365, gm_n269, gm_n115, in_15, gm_n799, gm_n633);
	nand (gm_n2366, gm_n72, in_20, in_19, gm_n2365);
	nor (gm_n2367, gm_n274, in_16, gm_n59, gm_n2244, gm_n276);
	nand (gm_n2368, gm_n113, in_21, in_20, gm_n2367);
	nand (gm_n2369, gm_n2368, gm_n2366, gm_n2364);
	nor (gm_n2370, gm_n909, gm_n133, in_14, gm_n240, gm_n212);
	nand (gm_n2371, gm_n2370, gm_n199, in_18);
	nor (gm_n2372, gm_n158, gm_n59, in_8, gm_n354, gm_n161);
	nand (gm_n2373, gm_n72, gm_n85, gm_n56, gm_n2372, gm_n486);
	nor (gm_n2374, gm_n514, gm_n76, gm_n62, gm_n502, gm_n462);
	nand (gm_n2375, gm_n311, in_21, in_17, gm_n2374, gm_n595);
	nand (gm_n2376, gm_n2375, gm_n2373, gm_n2371);
	nor (gm_n2377, gm_n2362, gm_n2350, gm_n2348, gm_n2376, gm_n2369);
	nand (gm_n2378, gm_n123, in_13, in_9, gm_n316, gm_n186);
	nor (gm_n2379, gm_n388, gm_n72, in_17, gm_n2378, gm_n256);
	or (gm_n2380, gm_n286, gm_n121, in_13, gm_n438, gm_n480);
	nor (gm_n2381, gm_n103, in_21, in_17, gm_n2380);
	or (gm_n2382, gm_n358, in_13, in_9, gm_n345, gm_n344);
	nor (gm_n2383, gm_n105, gm_n72, gm_n55, gm_n2382, gm_n183);
	nor (gm_n2384, gm_n2383, gm_n2381, gm_n2379);
	or (gm_n2385, gm_n358, gm_n76, gm_n62, gm_n462, gm_n667);
	nor (gm_n2386, gm_n441, gm_n72, in_17, gm_n2385, gm_n662);
	or (gm_n2387, gm_n149, gm_n90, in_10, gm_n362, gm_n349);
	nor (gm_n2388, gm_n244, gm_n212, in_18, gm_n2387);
	or (gm_n2389, gm_n430, in_13, gm_n62, gm_n503, gm_n442);
	nor (gm_n2390, gm_n183, gm_n72, gm_n55, gm_n2389, gm_n375);
	nor (gm_n2391, gm_n2390, gm_n2388, gm_n2386);
	nand (gm_n2392, gm_n2377, gm_n2345, gm_n2344, gm_n2391, gm_n2384);
	and (gm_n2393, in_14, in_10, in_9, gm_n2065, gm_n600);
	nand (gm_n2394, gm_n367, gm_n88, in_18, gm_n2393);
	nor (gm_n2395, gm_n461, in_13, in_9, gm_n503, gm_n430);
	nand (gm_n2396, gm_n122, in_21, in_17, gm_n2395, gm_n206);
	nor (gm_n2397, gm_n114, gm_n73, in_12, gm_n1016, gm_n274);
	nand (gm_n2398, gm_n383, gm_n72, gm_n85, gm_n2397);
	nand (gm_n2399, gm_n2398, gm_n2396, gm_n2394);
	nor (gm_n2400, gm_n263, in_16, in_12, gm_n1319, gm_n385);
	nand (gm_n2401, gm_n697, gm_n72, in_20, gm_n2400);
	or (gm_n2402, gm_n671, gm_n194, gm_n94);
	nor (gm_n2403, in_14, in_10, gm_n62, gm_n2402, gm_n92);
	nand (gm_n2404, gm_n166, gm_n129, gm_n119, gm_n2403);
	nor (gm_n2405, gm_n227, gm_n73, in_12, gm_n520, gm_n297);
	nand (gm_n2406, gm_n495, in_21, gm_n85, gm_n2405);
	nand (gm_n2407, gm_n2406, gm_n2404, gm_n2401);
	nor (gm_n2408, gm_n2392, gm_n2342, gm_n2339, gm_n2407, gm_n2399);
	nand (gm_n2409, gm_n143, in_16, gm_n59, gm_n1427, gm_n303);
	nor (gm_n2410, gm_n496, gm_n72, gm_n85, gm_n2409);
	or (gm_n2411, gm_n263, gm_n59, in_8, gm_n508, gm_n276);
	nor (gm_n2412, in_21, in_20, gm_n73, gm_n2411, gm_n58);
	nand (gm_n2413, gm_n143, gm_n73, in_12, gm_n1456, gm_n949);
	nor (gm_n2414, gm_n496, in_21, gm_n85, gm_n2413);
	nor (gm_n2415, gm_n2414, gm_n2412, gm_n2410);
	nor (gm_n2416, gm_n228, gm_n223, in_8);
	nand (gm_n2417, gm_n64, in_16, in_12, gm_n2416, gm_n77);
	nor (gm_n2418, gm_n262, gm_n72, in_20, gm_n2417);
	or (gm_n2419, gm_n158, gm_n73, in_12, gm_n552, gm_n276);
	nor (gm_n2420, gm_n912, in_21, in_20, gm_n2419);
	nand (gm_n2421, in_7, in_6, in_5, gm_n546, gm_n94);
	or (gm_n2422, gm_n152, gm_n73, in_12, gm_n2421, gm_n263);
	nor (gm_n2423, gm_n781, in_21, in_20, gm_n2422);
	nor (gm_n2424, gm_n2423, gm_n2420, gm_n2418);
	nand (gm_n2425, gm_n2408, gm_n2337, gm_n2335, gm_n2424, gm_n2415);
	and (gm_n2426, gm_n123, gm_n76, in_9, gm_n1427);
	nand (gm_n2427, gm_n102, in_21, gm_n55, gm_n2426, gm_n405);
	and (gm_n2428, in_14, in_10, in_9, gm_n998, gm_n624);
	nand (gm_n2429, gm_n436, gm_n146, gm_n119, gm_n2428);
	and (gm_n2430, in_14, gm_n78, gm_n62, gm_n1095, gm_n600);
	nand (gm_n2431, gm_n243, gm_n200, in_18, gm_n2430);
	nand (gm_n2432, gm_n2431, gm_n2429, gm_n2427);
	nor (gm_n2433, gm_n114, gm_n73, gm_n59, gm_n1324, gm_n155);
	nand (gm_n2434, gm_n697, in_21, gm_n85, gm_n2433);
	or (gm_n2435, gm_n193, gm_n194, gm_n63, gm_n271, gm_n238);
	nor (gm_n2436, in_21, gm_n56, gm_n60, gm_n2435, gm_n447);
	nand (gm_n2437, gm_n2436, in_20);
	nor (gm_n2438, gm_n190, in_16, in_12, gm_n765, gm_n227);
	nand (gm_n2439, gm_n57, in_21, gm_n85, gm_n2438);
	nand (gm_n2440, gm_n2439, gm_n2437, gm_n2434);
	nor (gm_n2441, gm_n2425, gm_n2332, gm_n2330, gm_n2440, gm_n2432);
	and (gm_n2442, gm_n102, in_21, gm_n55, gm_n2136, gm_n595);
	nor (gm_n2443, gm_n93, in_6, in_5, gm_n671, in_8);
	nand (gm_n2444, gm_n222, gm_n484, gm_n60, gm_n2443, gm_n486);
	nor (gm_n2445, in_21, in_20, in_19, gm_n2444);
	nand (gm_n2446, gm_n90, gm_n78, gm_n62, gm_n2218, gm_n713);
	nor (gm_n2447, gm_n212, gm_n165, gm_n119, gm_n2446);
	nor (gm_n2448, gm_n2447, gm_n2445, gm_n2442);
	nand (gm_n2449, gm_n110, gm_n76, gm_n62, gm_n579, gm_n186);
	nor (gm_n2450, gm_n256, gm_n72, gm_n55, gm_n2449, gm_n620);
	or (gm_n2451, gm_n159, gm_n60, in_11, gm_n981, gm_n980);
	nor (gm_n2452, gm_n72, gm_n85, in_19, gm_n2451, gm_n1331);
	or (gm_n2453, gm_n287, gm_n90, gm_n78, gm_n526, gm_n369);
	nor (gm_n2454, gm_n531, gm_n1989, gm_n119, gm_n2453);
	nor (gm_n2455, gm_n2454, gm_n2452, gm_n2450);
	nand (gm_n2456, gm_n2441, gm_n2328, gm_n2326, gm_n2455, gm_n2448);
	nor (gm_n2457, gm_n152, in_16, gm_n59, gm_n2421, gm_n274);
	nand (gm_n2458, gm_n697, gm_n72, gm_n85, gm_n2457);
	nor (gm_n2459, gm_n114, gm_n73, in_12, gm_n230, gm_n274);
	nand (gm_n2460, gm_n57, gm_n72, in_20, gm_n2459);
	nor (gm_n2461, gm_n149, gm_n358, gm_n76, gm_n438, gm_n313);
	nand (gm_n2462, gm_n120, gm_n72, gm_n55, gm_n2461);
	nand (gm_n2463, gm_n2462, gm_n2460, gm_n2458);
	nor (gm_n2464, gm_n227, gm_n73, gm_n59, gm_n1484, gm_n158);
	nand (gm_n2465, gm_n296, in_21, in_20, gm_n2464);
	and (gm_n2466, gm_n268, gm_n143, in_15, gm_n636, gm_n422);
	nand (gm_n2467, in_21, in_20, in_19, gm_n2466);
	and (gm_n2468, gm_n1157, in_14, in_10, gm_n829, gm_n1011);
	nand (gm_n2469, gm_n367, gm_n806, gm_n119, gm_n2468);
	nand (gm_n2470, gm_n2469, gm_n2467, gm_n2465);
	nor (gm_n2471, gm_n2456, gm_n2324, gm_n2322, gm_n2470, gm_n2463);
	nand (gm_n2472, gm_n264, gm_n73, in_12, gm_n2065, gm_n571);
	nor (gm_n2473, gm_n139, in_21, gm_n85, gm_n2472);
	or (gm_n2474, gm_n93, in_6, gm_n97, gm_n671, gm_n94);
	or (gm_n2475, gm_n461, in_13, in_9, gm_n2474, gm_n662);
	nor (gm_n2476, gm_n441, gm_n72, in_17, gm_n2475);
	nand (gm_n2477, gm_n221, in_16, gm_n59, gm_n991, gm_n264);
	nor (gm_n2478, gm_n781, gm_n72, in_20, gm_n2477);
	nor (gm_n2479, gm_n2478, gm_n2476, gm_n2473);
	or (gm_n2480, gm_n193, gm_n60, gm_n63, gm_n1382, gm_n541);
	nor (gm_n2481, in_21, gm_n85, gm_n56, gm_n2480, gm_n393);
	nand (gm_n2482, gm_n402, gm_n335, gm_n76, gm_n722);
	nor (gm_n2483, gm_n121, gm_n72, in_17, gm_n2482, gm_n388);
	or (gm_n2484, gm_n256, gm_n99, in_13, gm_n442, gm_n438);
	nor (gm_n2485, gm_n441, in_21, in_17, gm_n2484);
	nor (gm_n2486, gm_n2485, gm_n2483, gm_n2481);
	nand (gm_n2487, gm_n2471, gm_n2320, gm_n2318, gm_n2486, gm_n2479);
	nor (gm_n2488, gm_n95, in_14, gm_n78, gm_n526, gm_n147);
	nand (gm_n2489, gm_n436, gm_n199, gm_n119, gm_n2488);
	nor (gm_n2490, in_14, gm_n78, gm_n62, gm_n1689, gm_n147);
	nand (gm_n2491, gm_n129, gm_n88, in_18, gm_n2490);
	and (gm_n2492, gm_n532, gm_n90, in_10, gm_n335, gm_n333);
	nand (gm_n2493, gm_n131, gm_n86, in_18, gm_n2492);
	nand (gm_n2494, gm_n2493, gm_n2491, gm_n2489);
	nor (gm_n2495, gm_n514, in_13, gm_n62, gm_n502, gm_n345);
	nand (gm_n2496, gm_n174, in_21, in_17, gm_n2495, gm_n1076);
	and (gm_n2497, gm_n93, gm_n124, in_5, gm_n426, gm_n94);
	and (gm_n2498, gm_n61, in_16, gm_n59, gm_n2497, gm_n222);
	nand (gm_n2499, gm_n383, gm_n72, gm_n85, gm_n2498);
	nor (gm_n2500, gm_n220, gm_n73, gm_n59, gm_n399, gm_n274);
	nand (gm_n2501, gm_n383, in_21, in_20, gm_n2500);
	nand (gm_n2502, gm_n2501, gm_n2499, gm_n2496);
	nor (gm_n2503, gm_n2487, gm_n2316, gm_n2315, gm_n2502, gm_n2494);
	or (gm_n2504, in_13, in_9, in_8, gm_n842, gm_n406);
	nor (gm_n2505, gm_n103, gm_n72, in_17, gm_n2504, gm_n328);
	or (gm_n2506, gm_n796, in_13, gm_n62, gm_n502, gm_n480);
	nor (gm_n2507, gm_n103, in_21, gm_n55, gm_n2506, gm_n121);
	or (gm_n2508, gm_n121, gm_n76, in_12, gm_n835, gm_n274);
	nor (gm_n2509, gm_n620, gm_n72, gm_n55, gm_n2508);
	nor (gm_n2510, gm_n2509, gm_n2507, gm_n2505);
	nand (gm_n2511, gm_n90, in_10, in_9, gm_n626, gm_n713);
	nor (gm_n2512, gm_n841, gm_n824, gm_n119, gm_n2511);
	or (gm_n2513, gm_n115, in_16, in_12, gm_n385, gm_n135);
	nor (gm_n2514, gm_n384, gm_n72, in_20, gm_n2513);
	nand (gm_n2515, gm_n222, gm_n75, in_15, gm_n1095, gm_n1398);
	nor (gm_n2516, in_21, in_20, gm_n56, gm_n2515);
	nor (gm_n2517, gm_n2516, gm_n2514, gm_n2512);
	nand (gm_n2518, gm_n2503, gm_n2313, gm_n2311, gm_n2517, gm_n2510);
	nor (gm_n2519, gm_n480, gm_n76, gm_n62, gm_n988, gm_n502);
	nand (gm_n2520, gm_n174, in_21, in_17, gm_n2519, gm_n523);
	nor (gm_n2521, gm_n148, gm_n90, in_10, gm_n414, gm_n369);
	nand (gm_n2522, gm_n88, gm_n86, gm_n119, gm_n2521);
	nor (gm_n2523, gm_n92, in_14, gm_n78, gm_n389, gm_n370);
	nand (gm_n2524, gm_n348, gm_n245, in_18, gm_n2523);
	nand (gm_n2525, gm_n2524, gm_n2522, gm_n2520);
	or (gm_n2526, in_11, gm_n78, in_9, gm_n988, gm_n609);
	nor (gm_n2527, gm_n393, in_19, in_15, gm_n2526, gm_n633);
	nand (gm_n2528, gm_n2527, in_21, gm_n85);
	nor (gm_n2529, gm_n155, gm_n76, gm_n59, gm_n458);
	nand (gm_n2530, gm_n104, in_21, gm_n55, gm_n2529, gm_n327);
	nor (gm_n2531, gm_n1295, in_13, in_9, gm_n463, gm_n461);
	nand (gm_n2532, gm_n120, gm_n72, in_17, gm_n2531, gm_n523);
	nand (gm_n2533, gm_n2532, gm_n2530, gm_n2528);
	nor (gm_n2534, gm_n2518, gm_n2309, gm_n2307, gm_n2533, gm_n2525);
	nand (gm_n2535, gm_n265, gm_n154, in_15, gm_n1398, gm_n1101);
	nor (gm_n2536, in_21, gm_n85, in_19, gm_n2535);
	or (gm_n2537, gm_n141, gm_n194, in_14, gm_n605, gm_n807);
	nor (gm_n2538, gm_n437, gm_n244, gm_n119, gm_n2537);
	or (gm_n2539, gm_n190, gm_n73, in_12, gm_n152, gm_n116);
	nor (gm_n2540, gm_n384, gm_n72, gm_n85, gm_n2539);
	nor (gm_n2541, gm_n2540, gm_n2538, gm_n2536);
	nor (gm_n2542, gm_n349, in_11, gm_n78, gm_n526);
	nand (gm_n2543, gm_n281, in_19, gm_n60, gm_n2542, gm_n422);
	nor (gm_n2544, gm_n2543, in_21, in_20);
	or (gm_n2545, gm_n406, in_13, in_9, gm_n743, gm_n596);
	nor (gm_n2546, gm_n312, gm_n72, in_17, gm_n2545, gm_n313);
	and (gm_n2547, gm_n93, gm_n124, in_5, gm_n454, gm_n94);
	nand (gm_n2548, gm_n61, in_16, in_12, gm_n2547, gm_n222);
	nor (gm_n2549, gm_n139, in_21, in_20, gm_n2548);
	nor (gm_n2550, gm_n2549, gm_n2546, gm_n2544);
	nand (gm_n2551, gm_n2534, gm_n2305, gm_n2303, gm_n2550, gm_n2541);
	and (gm_n2552, gm_n214, gm_n73, gm_n59, gm_n1095, gm_n303);
	nand (gm_n2553, gm_n57, gm_n72, in_20, gm_n2552);
	nand (gm_n2554, gm_n104, gm_n72, gm_n55, gm_n2147, gm_n174);
	nor (gm_n2555, gm_n278, gm_n190, in_15, gm_n760, gm_n1331);
	nand (gm_n2556, gm_n72, gm_n85, in_19, gm_n2555);
	nand (gm_n2557, gm_n2556, gm_n2554, gm_n2553);
	nor (gm_n2558, gm_n148, gm_n90, in_10, gm_n389, gm_n362);
	nand (gm_n2559, gm_n166, gm_n164, in_18, gm_n2558);
	nor (gm_n2560, gm_n667, gm_n76, in_9, gm_n503, gm_n461);
	nand (gm_n2561, gm_n174, in_21, in_17, gm_n2560, gm_n1076);
	nand (gm_n2562, gm_n222, gm_n76, gm_n59, gm_n2218);
	or (gm_n2563, gm_n620, gm_n72, gm_n55, gm_n2562, gm_n662);
	nand (gm_n2564, gm_n2563, gm_n2561, gm_n2559);
	nor (gm_n2565, gm_n2551, gm_n2301, gm_n2299, gm_n2564, gm_n2557);
	or (gm_n2566, gm_n227, in_16, gm_n59, gm_n2357, gm_n213);
	nor (gm_n2567, gm_n139, gm_n72, in_20, gm_n2566);
	or (gm_n2568, gm_n480, in_13, in_9, gm_n1583, gm_n443);
	nor (gm_n2569, gm_n312, in_21, gm_n55, gm_n2568, gm_n375);
	or (gm_n2570, gm_n431, in_13, in_9, gm_n988, gm_n502);
	nor (gm_n2571, gm_n103, gm_n72, gm_n55, gm_n2570, gm_n375);
	nor (gm_n2572, gm_n2571, gm_n2569, gm_n2567);
	nor (gm_n2573, gm_n238, gm_n202, in_8);
	nand (gm_n2574, in_14, gm_n78, gm_n62, gm_n2573, gm_n600);
	nor (gm_n2575, gm_n1989, gm_n824, gm_n119, gm_n2574);
	nor (gm_n2576, gm_n121, gm_n72, gm_n55, gm_n1979, gm_n479);
	nand (gm_n2577, gm_n143, gm_n60, gm_n94, gm_n455, gm_n422);
	nor (gm_n2578, gm_n72, gm_n85, gm_n56, gm_n2577, gm_n393);
	nor (gm_n2579, gm_n2578, gm_n2576, gm_n2575);
	nand (gm_n2580, gm_n2565, gm_n2297, gm_n2295, gm_n2579, gm_n2572);
	nor (gm_n2581, gm_n248, gm_n90, in_10, gm_n491, gm_n369);
	nand (gm_n2582, gm_n200, gm_n129, gm_n119, gm_n2581);
	and (gm_n2583, gm_n90, gm_n78, gm_n62, gm_n2218, gm_n334);
	nand (gm_n2584, gm_n146, gm_n88, gm_n119, gm_n2583);
	nand (gm_n2585, gm_n104, gm_n72, gm_n55, gm_n1565, gm_n373);
	nand (gm_n2586, gm_n2585, gm_n2584, gm_n2582);
	nor (gm_n2587, gm_n115, gm_n74, in_15, gm_n180, gm_n159);
	nand (gm_n2588, gm_n72, in_20, in_19, gm_n2587);
	or (gm_n2589, gm_n277, gm_n228, gm_n94);
	nor (gm_n2590, gm_n115, in_16, in_12, gm_n2589, gm_n152);
	nand (gm_n2591, gm_n296, gm_n72, in_20, gm_n2590);
	nor (gm_n2592, gm_n514, in_13, gm_n62, gm_n1583, gm_n463);
	nand (gm_n2593, gm_n174, gm_n72, in_17, gm_n2592, gm_n595);
	nand (gm_n2594, gm_n2593, gm_n2591, gm_n2588);
	nor (gm_n2595, gm_n2580, gm_n2293, gm_n2291, gm_n2594, gm_n2586);
	or (gm_n2596, gm_n358, gm_n76, in_9, gm_n597, gm_n344);
	nor (gm_n2597, gm_n256, gm_n72, gm_n55, gm_n2596, gm_n620);
	or (gm_n2598, gm_n431, in_13, gm_n62, gm_n502, gm_n481);
	nor (gm_n2599, gm_n256, in_21, in_17, gm_n2598, gm_n312);
	nand (gm_n2600, gm_n79, in_16, in_12, gm_n884, gm_n221);
	nor (gm_n2601, gm_n912, in_21, in_20, gm_n2600);
	nor (gm_n2602, gm_n2601, gm_n2599, gm_n2597);
	or (gm_n2603, gm_n247, in_14, in_10, gm_n362, gm_n350);
	nor (gm_n2604, gm_n1989, gm_n211, gm_n119, gm_n2603);
	and (gm_n2605, in_7, in_6, in_5, gm_n426, in_8);
	nand (gm_n2606, gm_n64, in_16, gm_n59, gm_n2605, gm_n221);
	nor (gm_n2607, gm_n139, in_21, in_20, gm_n2606);
	and (gm_n2608, gm_n519, gm_n81, in_8);
	nand (gm_n2609, gm_n222, gm_n221, in_12, gm_n2608, gm_n394);
	nor (gm_n2610, in_21, gm_n85, in_19, gm_n2609);
	nor (gm_n2611, gm_n2610, gm_n2607, gm_n2604);
	nand (gm_n2612, gm_n2595, gm_n2289, gm_n2287, gm_n2611, gm_n2602);
	nor (gm_n2613, gm_n227, in_16, in_12, gm_n1125, gm_n274);
	nand (gm_n2614, gm_n383, gm_n72, gm_n85, gm_n2613);
	nor (gm_n2615, gm_n263, gm_n159, gm_n60, gm_n1751, gm_n293);
	nand (gm_n2616, gm_n72, in_20, in_19, gm_n2615);
	nor (gm_n2617, in_14, gm_n78, gm_n62, gm_n1731, gm_n133);
	nand (gm_n2618, gm_n323, gm_n164, gm_n119, gm_n2617);
	nand (gm_n2619, gm_n2618, gm_n2616, gm_n2614);
	nor (gm_n2620, gm_n115, in_16, in_12, gm_n468, gm_n319);
	nand (gm_n2621, gm_n113, in_21, gm_n85, gm_n2620);
	nor (gm_n2622, gm_n168, gm_n158, gm_n60, gm_n1514, gm_n393);
	nand (gm_n2623, in_21, in_20, in_19, gm_n2622);
	nor (gm_n2624, gm_n671, gm_n572, in_8);
	and (gm_n2625, gm_n733, in_16, gm_n59, gm_n2624, gm_n214);
	nand (gm_n2626, gm_n495, gm_n72, gm_n85, gm_n2625);
	nand (gm_n2627, gm_n2626, gm_n2623, gm_n2621);
	nor (gm_n2628, gm_n2612, gm_n2285, gm_n2282, gm_n2627, gm_n2619);
	nor (gm_n2629, gm_n99, in_14, in_10, gm_n467, gm_n349);
	nand (gm_n2630, gm_n436, gm_n199, in_18, gm_n2629);
	nor (gm_n2631, gm_n92, gm_n90, gm_n78, gm_n389, gm_n287);
	nand (gm_n2632, gm_n199, gm_n88, gm_n119, gm_n2631);
	and (gm_n2633, gm_n422, gm_n143, in_15, gm_n612, gm_n448);
	nand (gm_n2634, in_21, gm_n85, in_19, gm_n2633);
	nand (gm_n2635, gm_n2630, gm_n2628, gm_n2280, gm_n2634, gm_n2632);
	nor (gm_n2636, gm_n406, in_13, in_9, gm_n743, gm_n443);
	nand (gm_n2637, gm_n254, in_21, in_17, gm_n2636, gm_n339);
	and (gm_n2638, gm_n214, gm_n73, gm_n59, gm_n235, gm_n221);
	nand (gm_n2639, gm_n697, gm_n72, in_20, gm_n2638);
	nor (gm_n2640, in_10, gm_n62, gm_n94, gm_n761, gm_n467);
	nand (gm_n2641, gm_n243, in_18, gm_n90, gm_n2640, gm_n245);
	nand (gm_n2642, gm_n2641, gm_n2639, gm_n2637);
	or (gm_n2643, gm_n208, gm_n184, gm_n76, gm_n491, gm_n406);
	nor (gm_n2644, gm_n374, in_21, gm_n55, gm_n2643);
	nor (out_5, gm_n2642, gm_n2635, gm_n2278, gm_n2644);
	and (gm_n2646, gm_n305, gm_n291, gm_n94);
	nand (gm_n2647, gm_n90, gm_n78, in_9, gm_n2646, gm_n532);
	nor (gm_n2648, gm_n437, gm_n87, in_18, gm_n2647);
	nor (gm_n2649, gm_n153, gm_n190, in_15, gm_n760, gm_n269);
	nand (gm_n2650, in_21, gm_n85, gm_n56, gm_n2649);
	or (gm_n2651, gm_n406, in_13, in_9, gm_n502, gm_n462);
	nor (gm_n2652, gm_n103, gm_n72, gm_n55, gm_n2651, gm_n328);
	nand (gm_n2653, gm_n392, gm_n154, gm_n60, gm_n1359, gm_n1101);
	nor (gm_n2654, in_21, in_20, gm_n56, gm_n2653);
	nor (gm_n2655, gm_n596, in_13, in_9, gm_n481, gm_n442);
	nand (gm_n2656, gm_n174, gm_n72, gm_n55, gm_n2655, gm_n255);
	nor (gm_n2657, gm_n152, gm_n73, gm_n59, gm_n675, gm_n213);
	nand (gm_n2658, gm_n113, in_21, gm_n85, gm_n2657);
	or (gm_n2659, gm_n430, gm_n76, gm_n62, gm_n442, gm_n359);
	nor (gm_n2660, gm_n105, in_21, gm_n55, gm_n2659, gm_n479);
	nand (gm_n2661, gm_n264, gm_n76, in_12, gm_n734);
	nor (gm_n2662, gm_n183, gm_n72, gm_n55, gm_n2661, gm_n121);
	nor (gm_n2663, gm_n431, gm_n76, gm_n62, gm_n515);
	nand (gm_n2664, gm_n327, gm_n72, gm_n55, gm_n2663, gm_n1076);
	nor (gm_n2665, gm_n93, in_6, gm_n97, gm_n229, in_8);
	and (gm_n2666, gm_n61, in_16, in_12, gm_n2665, gm_n154);
	nand (gm_n2667, gm_n697, gm_n72, gm_n85, gm_n2666);
	nand (gm_n2668, gm_n334, gm_n90, in_10, gm_n793, gm_n1345);
	nor (gm_n2669, gm_n841, gm_n130, in_18, gm_n2668);
	not (gm_n2670, gm_n287);
	nand (gm_n2671, gm_n2670, gm_n122, gm_n76, gm_n829, gm_n788);
	nor (gm_n2672, gm_n479, in_21, in_17, gm_n2671);
	and (gm_n2673, gm_n379, gm_n64, gm_n60, gm_n1392, gm_n545);
	nand (gm_n2674, gm_n72, in_20, in_19, gm_n2673);
	nor (gm_n2675, gm_n239, gm_n60, in_11, gm_n633, gm_n240);
	nand (gm_n2676, gm_n72, in_20, in_19, gm_n2675, gm_n486);
	or (gm_n2677, gm_n461, gm_n76, gm_n62, gm_n359, gm_n596);
	nor (gm_n2678, gm_n441, in_21, gm_n55, gm_n2677, gm_n184);
	or (gm_n2679, gm_n514, in_13, in_9, gm_n345, gm_n596);
	nor (gm_n2680, gm_n184, gm_n72, gm_n55, gm_n2679, gm_n479);
	and (gm_n2681, gm_n233, gm_n76, gm_n59, gm_n1569);
	nand (gm_n2682, gm_n104, gm_n72, gm_n55, gm_n2681, gm_n254);
	and (gm_n2683, gm_n519, gm_n304, gm_n94);
	and (gm_n2684, gm_n523, in_13, in_9, gm_n2683, gm_n402);
	nand (gm_n2685, gm_n120, in_21, in_17, gm_n2684);
	or (gm_n2686, gm_n90, gm_n78, gm_n62, gm_n832, gm_n362);
	nor (gm_n2687, gm_n437, gm_n244, in_18, gm_n2686);
	or (gm_n2688, in_10, in_9, in_8, gm_n939, gm_n133);
	nor (gm_n2689, gm_n841, in_18, in_14, gm_n2688, gm_n368);
	nand (gm_n2690, in_7, in_6, gm_n97, gm_n80);
	nor (gm_n2691, gm_n240, in_15, gm_n63, gm_n2690, gm_n633);
	nand (gm_n2692, in_21, gm_n85, in_19, gm_n2691, gm_n394);
	nor (gm_n2693, gm_n95, in_14, in_10, gm_n807, gm_n286);
	nand (gm_n2694, gm_n245, gm_n164, gm_n119, gm_n2693);
	nand (gm_n2695, gm_n126, gm_n76, gm_n62, gm_n1049, gm_n314);
	nor (gm_n2696, gm_n121, in_21, in_17, gm_n2695, gm_n441);
	or (gm_n2697, gm_n215, gm_n194, gm_n94);
	or (gm_n2698, gm_n358, gm_n76, in_9, gm_n2697, gm_n184);
	nor (gm_n2699, gm_n441, gm_n72, gm_n55, gm_n2698);
	nor (gm_n2700, gm_n149, in_14, gm_n78, gm_n349, gm_n807);
	nand (gm_n2701, gm_n348, gm_n131, in_18, gm_n2700);
	nor (gm_n2702, in_14, gm_n78, gm_n62, gm_n207, gm_n203);
	nand (gm_n2703, gm_n166, gm_n129, gm_n119, gm_n2702);
	nand (gm_n2704, gm_n64, gm_n73, gm_n59, gm_n1524, gm_n733);
	nor (gm_n2705, gm_n219, in_21, in_20, gm_n2704);
	nand (gm_n2706, gm_n733, gm_n73, gm_n59, gm_n950, gm_n214);
	nor (gm_n2707, gm_n58, gm_n72, gm_n85, gm_n2706);
	and (gm_n2708, in_10, in_9, gm_n94, gm_n176, gm_n91);
	nand (gm_n2709, gm_n164, in_18, in_14, gm_n2708, gm_n245);
	nor (gm_n2710, gm_n643, in_15, in_11, gm_n1382, gm_n541);
	nand (gm_n2711, in_21, in_20, gm_n56, gm_n2710, gm_n1101);
	nor (gm_n2712, gm_n93, in_6, in_5, gm_n671, gm_n94);
	nand (gm_n2713, gm_n214, gm_n192, in_15, gm_n2712, gm_n394);
	nor (gm_n2714, gm_n72, in_20, in_19, gm_n2713);
	nand (gm_n2715, gm_n214, gm_n76, in_12, gm_n2547, gm_n1076);
	nor (gm_n2716, gm_n441, in_21, in_17, gm_n2715);
	nor (gm_n2717, gm_n240, gm_n68, in_14, gm_n671, gm_n467);
	nand (gm_n2718, gm_n367, gm_n323, in_18, gm_n2717);
	nor (gm_n2719, gm_n93, in_6, in_5, gm_n141);
	and (gm_n2720, in_13, gm_n62, gm_n94, gm_n402, gm_n2719);
	nand (gm_n2721, gm_n120, in_21, in_17, gm_n2720, gm_n405);
	or (gm_n2722, gm_n263, gm_n73, in_12, gm_n520, gm_n319);
	nor (gm_n2723, gm_n912, gm_n72, in_20, gm_n2722);
	or (gm_n2724, gm_n354, gm_n115, gm_n59, gm_n2080);
	nor (gm_n2725, in_21, in_20, in_19, gm_n2724, gm_n1331);
	nand (gm_n2726, gm_n102, gm_n72, gm_n55, gm_n1485, gm_n122);
	nor (gm_n2727, gm_n572, gm_n234, in_8);
	and (gm_n2728, in_14, in_10, gm_n62, gm_n2727, gm_n624);
	nand (gm_n2729, gm_n131, gm_n86, in_18, gm_n2728);
	nand (gm_n2730, in_7, in_6, gm_n97, gm_n426, in_8);
	nor (gm_n2731, gm_n297, in_16, gm_n59, gm_n2730, gm_n220);
	nand (gm_n2732, gm_n495, in_21, in_20, gm_n2731);
	nor (gm_n2733, gm_n184, gm_n358, gm_n76, gm_n526, gm_n491);
	nand (gm_n2734, gm_n174, gm_n72, in_17, gm_n2733);
	nor (gm_n2735, gm_n643, gm_n60, gm_n63, gm_n1382, gm_n541);
	nand (gm_n2736, gm_n72, gm_n85, in_19, gm_n2735, gm_n281);
	nand (gm_n2737, gm_n2732, gm_n2729, gm_n2726, gm_n2736, gm_n2734);
	nor (gm_n2738, gm_n461, in_13, in_9, gm_n705, gm_n256);
	nand (gm_n2739, gm_n102, in_21, gm_n55, gm_n2738);
	nor (gm_n2740, gm_n430, gm_n76, in_9, gm_n1132, gm_n257);
	nand (gm_n2741, gm_n104, gm_n72, in_17, gm_n2740, gm_n254);
	nor (gm_n2742, gm_n414, gm_n313, in_13, gm_n491, gm_n442);
	nand (gm_n2743, gm_n311, in_21, gm_n55, gm_n2742);
	nand (gm_n2744, gm_n2743, gm_n2741, gm_n2739);
	nor (gm_n2745, gm_n514, gm_n76, gm_n62, gm_n502, gm_n359);
	nand (gm_n2746, gm_n102, in_21, gm_n55, gm_n2745, gm_n104);
	nor (gm_n2747, gm_n609, in_13, in_9, gm_n480, gm_n359);
	nand (gm_n2748, gm_n206, in_21, in_17, gm_n2747, gm_n255);
	and (gm_n2749, gm_n126, gm_n76, gm_n62, gm_n1049, gm_n402);
	nand (gm_n2750, gm_n595, in_21, gm_n55, gm_n2749, gm_n373);
	nand (gm_n2751, gm_n2750, gm_n2748, gm_n2746);
	nor (gm_n2752, gm_n2737, gm_n2725, gm_n2723, gm_n2751, gm_n2744);
	or (gm_n2753, gm_n461, in_13, in_9, gm_n621, gm_n443);
	nor (gm_n2754, gm_n312, gm_n72, gm_n55, gm_n2753, gm_n375);
	nor (gm_n2755, gm_n190, gm_n59, in_8, gm_n572, gm_n223);
	nand (gm_n2756, gm_n733, in_20, gm_n73, gm_n2755, gm_n179);
	nor (gm_n2757, gm_n2756, in_21);
	or (gm_n2758, gm_n76, gm_n59, in_11, gm_n1382, gm_n541);
	nor (gm_n2759, gm_n312, gm_n72, in_17, gm_n2758, gm_n662);
	nor (gm_n2760, gm_n2759, gm_n2757, gm_n2754);
	or (gm_n2761, gm_n609, in_13, in_9, gm_n345, gm_n257);
	nor (gm_n2762, gm_n105, in_21, in_17, gm_n2761, gm_n388);
	or (gm_n2763, gm_n430, in_13, in_9, gm_n743, gm_n442);
	nor (gm_n2764, gm_n313, in_21, in_17, gm_n2763, gm_n374);
	or (gm_n2765, gm_n133, in_14, gm_n78, gm_n526, gm_n247);
	nor (gm_n2766, gm_n531, gm_n167, gm_n119, gm_n2765);
	nor (gm_n2767, gm_n2766, gm_n2764, gm_n2762);
	nand (gm_n2768, gm_n2752, gm_n2721, gm_n2718, gm_n2767, gm_n2760);
	or (gm_n2769, in_7, in_6, in_5, gm_n238);
	nor (gm_n2770, gm_n158, in_12, gm_n94, gm_n2769, gm_n354);
	nand (gm_n2771, gm_n72, in_20, in_16, gm_n2770, gm_n296);
	nor (gm_n2772, gm_n430, in_13, in_9, gm_n621, gm_n480);
	nand (gm_n2773, gm_n523, gm_n72, gm_n55, gm_n2772, gm_n327);
	nor (gm_n2774, gm_n191, gm_n190, gm_n60, gm_n2357, gm_n633);
	nand (gm_n2775, gm_n72, gm_n85, gm_n56, gm_n2774);
	nand (gm_n2776, gm_n2775, gm_n2773, gm_n2771);
	nor (gm_n2777, in_13, in_12, in_11, gm_n770, gm_n271);
	nand (gm_n2778, gm_n255, in_21, in_17, gm_n2777, gm_n327);
	nor (gm_n2779, gm_n286, in_14, gm_n78, gm_n467, gm_n349);
	nand (gm_n2780, gm_n129, gm_n88, gm_n119, gm_n2779);
	nand (gm_n2781, gm_n348, gm_n166, in_18, gm_n1362);
	nand (gm_n2782, gm_n2781, gm_n2780, gm_n2778);
	nor (gm_n2783, gm_n2768, gm_n2716, gm_n2714, gm_n2782, gm_n2776);
	nand (gm_n2784, gm_n484, gm_n233, in_15, gm_n547, gm_n281);
	nor (gm_n2785, in_21, in_20, in_19, gm_n2784);
	nand (gm_n2786, gm_n61, gm_n73, gm_n59, gm_n235, gm_n233);
	nor (gm_n2787, gm_n496, gm_n72, in_20, gm_n2786);
	nand (gm_n2788, gm_n79, in_16, in_12, gm_n2646, gm_n571);
	nor (gm_n2789, gm_n58, gm_n72, gm_n85, gm_n2788);
	nor (gm_n2790, gm_n2789, gm_n2787, gm_n2785);
	nand (gm_n2791, gm_n90, gm_n78, in_9, gm_n1531, gm_n624);
	nor (gm_n2792, gm_n212, gm_n87, in_18, gm_n2791);
	or (gm_n2793, gm_n1331, gm_n213, in_15, gm_n2244, gm_n764);
	nor (gm_n2794, in_21, gm_n85, in_19, gm_n2793);
	nand (gm_n2795, gm_n555, in_15, in_11, gm_n1398, gm_n601);
	nor (gm_n2796, in_21, gm_n85, gm_n56, gm_n2795, gm_n1331);
	nor (gm_n2797, gm_n2796, gm_n2794, gm_n2792);
	nand (gm_n2798, gm_n2783, gm_n2711, gm_n2709, gm_n2797, gm_n2790);
	nor (gm_n2799, gm_n147, in_14, gm_n78, gm_n589, gm_n148);
	nand (gm_n2800, gm_n436, gm_n146, in_18, gm_n2799);
	nor (gm_n2801, gm_n667, gm_n76, gm_n62, gm_n621, gm_n257);
	nand (gm_n2802, gm_n174, in_21, in_17, gm_n2801, gm_n1076);
	nor (gm_n2803, gm_n297, gm_n73, gm_n59, gm_n1751, gm_n276);
	nand (gm_n2804, gm_n296, in_21, in_20, gm_n2803);
	nand (gm_n2805, gm_n2804, gm_n2802, gm_n2800);
	and (gm_n2806, gm_n107, gm_n76, gm_n62, gm_n126, gm_n123);
	nand (gm_n2807, gm_n206, gm_n72, in_17, gm_n2806, gm_n595);
	nor (gm_n2808, gm_n369, in_14, gm_n78, gm_n389, gm_n370);
	nand (gm_n2809, gm_n245, gm_n86, gm_n119, gm_n2808);
	nor (gm_n2810, gm_n257, in_13, in_9, gm_n462, gm_n344);
	nand (gm_n2811, gm_n174, gm_n72, in_17, gm_n2810, gm_n595);
	nand (gm_n2812, gm_n2811, gm_n2809, gm_n2807);
	nor (gm_n2813, gm_n2798, gm_n2707, gm_n2705, gm_n2812, gm_n2805);
	nand (gm_n2814, gm_n268, gm_n79, gm_n60, gm_n1758, gm_n1398);
	nor (gm_n2815, gm_n72, gm_n85, gm_n56, gm_n2814);
	or (gm_n2816, gm_n78, in_9, in_8, gm_n981, gm_n147);
	nor (gm_n2817, gm_n244, in_18, in_14, gm_n2816, gm_n246);
	or (gm_n2818, gm_n274, in_16, gm_n59, gm_n1719, gm_n319);
	nor (gm_n2819, gm_n912, in_21, gm_n85, gm_n2818);
	nor (gm_n2820, gm_n2819, gm_n2817, gm_n2815);
	nand (gm_n2821, gm_n107, gm_n78, in_9, gm_n600, gm_n126);
	nor (gm_n2822, gm_n165, gm_n119, gm_n90, gm_n2821, gm_n1989);
	nand (gm_n2823, gm_n454, gm_n291, gm_n94);
	or (gm_n2824, gm_n114, gm_n73, gm_n59, gm_n2823, gm_n213);
	nor (gm_n2825, gm_n139, gm_n72, in_20, gm_n2824);
	or (gm_n2826, gm_n572, gm_n201, in_8);
	or (gm_n2827, gm_n152, gm_n73, gm_n59, gm_n2826, gm_n213);
	nor (gm_n2828, gm_n781, gm_n72, in_20, gm_n2827);
	nor (gm_n2829, gm_n2828, gm_n2825, gm_n2822);
	nand (gm_n2830, gm_n2813, gm_n2703, gm_n2701, gm_n2829, gm_n2820);
	and (gm_n2831, gm_n281, gm_n64, gm_n60, gm_n962, gm_n422);
	nand (gm_n2832, gm_n72, gm_n85, in_19, gm_n2831);
	and (gm_n2833, gm_n394, gm_n222, gm_n60, gm_n2096, gm_n545);
	nand (gm_n2834, in_21, in_20, gm_n56, gm_n2833);
	and (gm_n2835, gm_n106, gm_n76, gm_n62, gm_n2346, gm_n122);
	nand (gm_n2836, gm_n311, in_21, gm_n55, gm_n2835);
	nand (gm_n2837, gm_n2836, gm_n2834, gm_n2832);
	and (gm_n2838, gm_n76, in_12, in_8, gm_n455, gm_n64);
	nand (gm_n2839, gm_n206, in_21, in_17, gm_n2838, gm_n255);
	nor (gm_n2840, gm_n667, gm_n76, gm_n62, gm_n1132, gm_n406);
	nand (gm_n2841, gm_n254, gm_n72, in_17, gm_n2840, gm_n255);
	nor (gm_n2842, gm_n92, gm_n90, gm_n78, gm_n589, gm_n438);
	nand (gm_n2843, gm_n164, gm_n88, in_18, gm_n2842);
	nand (gm_n2844, gm_n2843, gm_n2841, gm_n2839);
	nor (gm_n2845, gm_n2830, gm_n2699, gm_n2696, gm_n2844, gm_n2837);
	nand (gm_n2846, in_14, in_10, in_9, gm_n2065, gm_n1011);
	nor (gm_n2847, gm_n437, gm_n165, gm_n119, gm_n2846);
	or (gm_n2848, gm_n133, gm_n90, gm_n78, gm_n370, gm_n259);
	nor (gm_n2849, gm_n368, gm_n246, gm_n119, gm_n2848);
	or (gm_n2850, gm_n514, gm_n76, in_9, gm_n621, gm_n430);
	nor (gm_n2851, gm_n388, gm_n72, gm_n55, gm_n2850, gm_n328);
	nor (gm_n2852, gm_n2851, gm_n2849, gm_n2847);
	or (gm_n2853, gm_n609, gm_n76, gm_n62, gm_n462, gm_n461);
	nor (gm_n2854, gm_n312, gm_n72, in_17, gm_n2853, gm_n313);
	or (gm_n2855, gm_n442, gm_n76, in_9, gm_n502, gm_n462);
	nor (gm_n2856, gm_n620, in_21, in_17, gm_n2855, gm_n375);
	nor (gm_n2857, gm_n437, gm_n130, gm_n119, gm_n2186);
	nor (gm_n2858, gm_n2857, gm_n2856, gm_n2854);
	nand (gm_n2859, gm_n2845, gm_n2694, gm_n2692, gm_n2858, gm_n2852);
	and (gm_n2860, gm_n93, in_6, in_5, gm_n80, gm_n94);
	and (gm_n2861, gm_n233, gm_n76, gm_n59, gm_n2860);
	nand (gm_n2862, gm_n174, gm_n72, in_17, gm_n2861, gm_n255);
	nand (gm_n2863, gm_n254, gm_n72, gm_n55, gm_n1482, gm_n1076);
	nor (gm_n2864, gm_n431, in_13, in_9, gm_n621, gm_n502);
	nand (gm_n2865, gm_n311, in_21, gm_n55, gm_n2864, gm_n339);
	nand (gm_n2866, gm_n2865, gm_n2863, gm_n2862);
	and (gm_n2867, gm_n222, gm_n192, gm_n60, gm_n2172, gm_n1101);
	nand (gm_n2868, gm_n72, in_20, in_19, gm_n2867);
	and (gm_n2869, gm_n214, gm_n76, gm_n59, gm_n1456);
	nand (gm_n2870, gm_n311, gm_n72, gm_n55, gm_n2869, gm_n595);
	and (gm_n2871, gm_n264, in_16, gm_n59, gm_n1531, gm_n303);
	nand (gm_n2872, gm_n296, in_21, in_20, gm_n2871);
	nand (gm_n2873, gm_n2872, gm_n2870, gm_n2868);
	nor (gm_n2874, gm_n2859, gm_n2689, gm_n2687, gm_n2873, gm_n2866);
	or (gm_n2875, gm_n328, gm_n257, in_13, gm_n589, gm_n349);
	nor (gm_n2876, gm_n103, in_21, in_17, gm_n2875);
	or (gm_n2877, gm_n155, gm_n73, in_12, gm_n1661, gm_n385);
	nor (gm_n2878, gm_n262, in_21, gm_n85, gm_n2877);
	nor (gm_n2879, gm_n93, in_6, in_5, gm_n201, gm_n94);
	nand (gm_n2880, gm_n143, in_16, gm_n59, gm_n2879, gm_n949);
	nor (gm_n2881, gm_n58, in_21, gm_n85, gm_n2880);
	nor (gm_n2882, gm_n2881, gm_n2878, gm_n2876);
	or (gm_n2883, gm_n609, in_13, in_9, gm_n359, gm_n257);
	nor (gm_n2884, gm_n105, gm_n72, in_17, gm_n2883, gm_n388);
	nor (gm_n2885, gm_n671, gm_n572, gm_n94);
	nand (gm_n2886, gm_n733, in_16, gm_n59, gm_n2885, gm_n222);
	nor (gm_n2887, gm_n781, gm_n72, gm_n85, gm_n2886);
	or (gm_n2888, gm_n220, gm_n73, in_12, gm_n855, gm_n263);
	nor (gm_n2889, gm_n781, in_21, gm_n85, gm_n2888);
	nor (gm_n2890, gm_n2889, gm_n2887, gm_n2884);
	nand (gm_n2891, gm_n2874, gm_n2685, gm_n2682, gm_n2890, gm_n2882);
	and (gm_n2892, gm_n143, in_16, gm_n59, gm_n1135, gm_n303);
	nand (gm_n2893, gm_n296, in_21, gm_n85, gm_n2892);
	and (gm_n2894, gm_n484, gm_n154, gm_n60, gm_n2065, gm_n268);
	nand (gm_n2895, in_21, gm_n85, gm_n56, gm_n2894);
	and (gm_n2896, gm_n264, gm_n73, in_12, gm_n547, gm_n571);
	nand (gm_n2897, gm_n495, gm_n72, gm_n85, gm_n2896);
	nand (gm_n2898, gm_n2897, gm_n2895, gm_n2893);
	and (gm_n2899, gm_n90, gm_n78, gm_n62, gm_n1611, gm_n624);
	nand (gm_n2900, gm_n348, gm_n323, gm_n119, gm_n2899);
	nor (gm_n2901, gm_n213, gm_n73, gm_n59, gm_n632, gm_n220);
	nand (gm_n2902, gm_n57, in_21, gm_n85, gm_n2901);
	nor (gm_n2903, gm_n78, in_9, in_8, gm_n270, gm_n147);
	nand (gm_n2904, gm_n146, gm_n119, gm_n90, gm_n2903, gm_n323);
	nand (gm_n2905, gm_n2904, gm_n2902, gm_n2900);
	nor (gm_n2906, gm_n2891, gm_n2680, gm_n2678, gm_n2905, gm_n2898);
	nand (gm_n2907, gm_n2670, gm_n106, gm_n76, gm_n829, gm_n595);
	nor (gm_n2908, gm_n441, in_21, gm_n55, gm_n2907);
	or (gm_n2909, gm_n358, in_13, in_9, gm_n503, gm_n667);
	nor (gm_n2910, gm_n184, in_21, in_17, gm_n2909, gm_n479);
	or (gm_n2911, in_14, gm_n78, in_9, gm_n399, gm_n207);
	nor (gm_n2912, gm_n437, gm_n165, gm_n119, gm_n2911);
	nor (gm_n2913, gm_n2912, gm_n2910, gm_n2908);
	nor (gm_n2914, gm_n369, gm_n78, gm_n62, gm_n2198);
	and (gm_n2915, gm_n174, gm_n72, gm_n55, gm_n2914, gm_n405);
	nor (gm_n2916, gm_n229, gm_n194, in_8);
	nand (gm_n2917, gm_n394, gm_n154, gm_n60, gm_n1398, gm_n2916);
	nor (gm_n2918, gm_n72, gm_n85, in_19, gm_n2917);
	nand (gm_n2919, gm_n2719, in_15, gm_n63, gm_n422, gm_n171);
	nor (gm_n2920, gm_n72, gm_n85, in_19, gm_n2919, gm_n74);
	nor (gm_n2921, gm_n2920, gm_n2918, gm_n2915);
	nand (gm_n2922, gm_n2906, gm_n2676, gm_n2674, gm_n2921, gm_n2913);
	nor (gm_n2923, gm_n190, in_16, gm_n59, gm_n815, gm_n354);
	nand (gm_n2924, gm_n383, in_21, in_20, gm_n2923);
	nor (gm_n2925, gm_n213, in_16, in_12, gm_n2697, gm_n276);
	nand (gm_n2926, gm_n383, gm_n72, gm_n85, gm_n2925);
	or (gm_n2927, in_11, gm_n78, in_9, gm_n1583, gm_n430);
	nor (gm_n2928, gm_n191, gm_n56, gm_n60, gm_n2927, gm_n633);
	nand (gm_n2929, gm_n2928, in_21, gm_n85);
	nand (gm_n2930, gm_n2929, gm_n2926, gm_n2924);
	nand (gm_n2931, gm_n1067, gm_n81, gm_n94);
	nor (gm_n2932, gm_n115, gm_n73, in_12, gm_n2931, gm_n276);
	nand (gm_n2933, gm_n138, gm_n72, in_20, gm_n2932);
	nor (gm_n2934, gm_n350, gm_n514, in_13, gm_n370);
	nand (gm_n2935, gm_n104, in_21, in_17, gm_n2934, gm_n206);
	nor (gm_n2936, gm_n609, in_13, in_9, gm_n432, gm_n461);
	nand (gm_n2937, gm_n311, gm_n72, in_17, gm_n2936, gm_n595);
	nand (gm_n2938, gm_n2937, gm_n2935, gm_n2933);
	nor (gm_n2939, gm_n2922, gm_n2672, gm_n2669, gm_n2938, gm_n2930);
	nor (gm_n2940, gm_n114, gm_n73, in_12, gm_n2125, gm_n274);
	and (gm_n2941, gm_n495, gm_n72, in_20, gm_n2940);
	nor (gm_n2942, in_7, in_6, in_5, gm_n141, in_8);
	nand (gm_n2943, gm_n123, in_13, gm_n62, gm_n2942, gm_n595);
	nor (gm_n2944, gm_n441, gm_n72, gm_n55, gm_n2943);
	or (gm_n2945, gm_n168, gm_n297, gm_n60, gm_n2125, gm_n1331);
	nor (gm_n2946, gm_n72, in_20, in_19, gm_n2945);
	nor (gm_n2947, gm_n2946, gm_n2944, gm_n2941);
	and (gm_n2948, gm_n254, gm_n72, gm_n55, gm_n1209, gm_n1076);
	nor (gm_n2949, gm_n93, in_6, in_5, gm_n229, in_8);
	nand (gm_n2950, gm_n448, gm_n79, gm_n60, gm_n2949, gm_n1398);
	nor (gm_n2951, gm_n72, in_20, in_19, gm_n2950);
	nand (gm_n2952, in_10, in_9, gm_n94, gm_n176, gm_n624);
	nor (gm_n2953, gm_n211, in_18, gm_n90, gm_n2952, gm_n841);
	nor (gm_n2954, gm_n2953, gm_n2951, gm_n2948);
	nand (gm_n2955, gm_n2939, gm_n2667, gm_n2664, gm_n2954, gm_n2947);
	or (gm_n2956, gm_n572, gm_n141, gm_n94);
	nor (gm_n2957, gm_n190, gm_n73, gm_n59, gm_n2956, gm_n385);
	nand (gm_n2958, gm_n57, in_21, in_20, gm_n2957);
	nor (gm_n2959, gm_n431, gm_n76, in_9, gm_n502, gm_n432);
	nand (gm_n2960, gm_n311, in_21, in_17, gm_n2959, gm_n595);
	nand (gm_n2961, gm_n102, in_21, gm_n55, gm_n1034, gm_n595);
	nand (gm_n2962, gm_n2961, gm_n2960, gm_n2958);
	nand (gm_n2963, gm_n93, in_6, in_5, gm_n454, in_8);
	nor (gm_n2964, in_14, gm_n78, in_9, gm_n2963, gm_n467);
	nand (gm_n2965, gm_n245, gm_n164, gm_n119, gm_n2964);
	nor (gm_n2966, gm_n667, in_13, in_9, gm_n988, gm_n431);
	nand (gm_n2967, gm_n254, gm_n72, gm_n55, gm_n2966, gm_n405);
	nor (gm_n2968, gm_n257, gm_n76, in_9, gm_n1132, gm_n344);
	nand (gm_n2969, gm_n174, gm_n72, in_17, gm_n2968, gm_n405);
	nand (gm_n2970, gm_n2969, gm_n2967, gm_n2965);
	nor (gm_n2971, gm_n2955, gm_n2662, gm_n2660, gm_n2970, gm_n2962);
	nand (gm_n2972, gm_n405, gm_n76, gm_n62, gm_n1709, gm_n340);
	nor (gm_n2973, gm_n103, gm_n72, gm_n55, gm_n2972);
	nand (gm_n2974, gm_n1928, in_15, gm_n63, gm_n1929, gm_n869);
	nor (gm_n2975, in_21, gm_n85, gm_n56, gm_n2974, gm_n191);
	nand (gm_n2976, gm_n79, in_16, gm_n59, gm_n1012, gm_n303);
	nor (gm_n2977, gm_n219, in_21, in_20, gm_n2976);
	nor (gm_n2978, gm_n2977, gm_n2975, gm_n2973);
	nor (gm_n2979, gm_n981, gm_n283, in_11);
	and (gm_n2980, gm_n131, gm_n129, gm_n119, gm_n2979, gm_n449);
	or (gm_n2981, gm_n442, in_13, in_9, gm_n597, gm_n443);
	nor (gm_n2982, gm_n388, gm_n72, in_17, gm_n2981, gm_n662);
	or (gm_n2983, gm_n514, in_13, in_9, gm_n597, gm_n596);
	nor (gm_n2984, gm_n121, gm_n72, in_17, gm_n2983, gm_n479);
	nor (gm_n2985, gm_n2984, gm_n2982, gm_n2980);
	nand (gm_n2986, gm_n2971, gm_n2658, gm_n2656, gm_n2985, gm_n2978);
	and (gm_n2987, gm_n106, gm_n76, gm_n62, gm_n1049, gm_n316);
	nand (gm_n2988, gm_n373, gm_n72, gm_n55, gm_n2987, gm_n1076);
	and (gm_n2989, gm_n186, gm_n76, in_9, gm_n402, gm_n316);
	nand (gm_n2990, gm_n327, gm_n72, in_17, gm_n2989, gm_n339);
	nor (gm_n2991, gm_n240, in_15, gm_n63, gm_n2690, gm_n290);
	nand (gm_n2992, gm_n72, gm_n85, gm_n56, gm_n2991, gm_n379);
	nand (gm_n2993, gm_n2992, gm_n2990, gm_n2988);
	nor (gm_n2994, gm_n667, gm_n76, in_9, gm_n503, gm_n406);
	nand (gm_n2995, gm_n206, in_21, gm_n55, gm_n2994, gm_n405);
	nor (gm_n2996, gm_n344, in_13, in_9, gm_n1132, gm_n442);
	nand (gm_n2997, gm_n120, gm_n72, gm_n55, gm_n2996, gm_n523);
	nor (gm_n2998, gm_n152, in_16, in_12, gm_n730, gm_n155);
	nand (gm_n2999, gm_n113, gm_n72, in_20, gm_n2998);
	nand (gm_n3000, gm_n2999, gm_n2997, gm_n2995);
	nor (gm_n3001, gm_n2986, gm_n2654, gm_n2652, gm_n3000, gm_n2993);
	nor (gm_n3002, gm_n406, gm_n76, gm_n62, gm_n463, gm_n359);
	nand (gm_n3003, gm_n104, gm_n72, in_17, gm_n3002, gm_n327);
	nor (gm_n3004, gm_n114, gm_n73, gm_n59, gm_n887, gm_n274);
	nand (gm_n3005, gm_n495, gm_n72, gm_n85, gm_n3004);
	nand (gm_n3006, gm_n93, in_6, in_5, gm_n546, in_8);
	nor (gm_n3007, gm_n293, gm_n297, in_15, gm_n3006, gm_n760);
	nand (gm_n3008, gm_n72, gm_n85, in_19, gm_n3007);
	nand (gm_n3009, gm_n3003, gm_n3001, gm_n2650, gm_n3008, gm_n3005);
	nor (gm_n3010, gm_n152, gm_n73, in_12, gm_n1837, gm_n274);
	nand (gm_n3011, gm_n296, gm_n72, gm_n85, gm_n3010);
	nor (gm_n3012, gm_n114, in_16, gm_n59, gm_n2421, gm_n190);
	nand (gm_n3013, gm_n296, in_21, in_20, gm_n3012);
	nor (gm_n3014, in_14, gm_n78, in_9, gm_n2333, gm_n369);
	nand (gm_n3015, gm_n243, gm_n131, in_18, gm_n3014);
	nand (gm_n3016, gm_n3015, gm_n3013, gm_n3011);
	or (gm_n3017, gm_n344, in_10, gm_n62, gm_n597, gm_n369);
	nor (gm_n3018, gm_n89, in_18, gm_n90, gm_n3017, gm_n211);
	nor (out_6, gm_n3016, gm_n3009, gm_n2648, gm_n3018);
	or (gm_n3020, gm_n148, gm_n90, gm_n78, gm_n207, gm_n149);
	nor (gm_n3021, gm_n130, gm_n89, in_18, gm_n3020);
	and (gm_n3022, gm_n192, gm_n64, gm_n60, gm_n870, gm_n281);
	nand (gm_n3023, in_21, in_20, in_19, gm_n3022);
	nand (gm_n3024, gm_n733, in_16, gm_n59, gm_n1179, gm_n154);
	nor (gm_n3025, gm_n219, gm_n72, gm_n85, gm_n3024);
	nand (gm_n3026, gm_n245, gm_n91, gm_n90, gm_n602, gm_n601);
	nor (gm_n3027, gm_n3026, gm_n531, in_18);
	nor (gm_n3028, gm_n207, in_14, in_10, gm_n589, gm_n370);
	nand (gm_n3029, gm_n367, gm_n88, gm_n119, gm_n3028);
	nor (gm_n3030, in_14, in_10, gm_n62, gm_n807, gm_n320);
	nand (gm_n3031, gm_n200, gm_n199, in_18, gm_n3030);
	nand (gm_n3032, in_13, in_9, gm_n94, gm_n556, gm_n106);
	nor (gm_n3033, gm_n105, gm_n72, in_17, gm_n3032, gm_n388);
	or (gm_n3034, gm_n190, in_16, gm_n59, gm_n1923, gm_n385);
	nor (gm_n3035, gm_n139, in_21, gm_n85, gm_n3034);
	nor (gm_n3036, gm_n263, in_16, in_12, gm_n2421, gm_n319);
	nand (gm_n3037, gm_n113, in_21, gm_n85, gm_n3036);
	nor (gm_n3038, gm_n90, gm_n78, gm_n62, gm_n203, gm_n92);
	nand (gm_n3039, gm_n199, gm_n131, gm_n119, gm_n3038);
	and (gm_n3040, gm_n806, gm_n86, gm_n119, gm_n1819);
	nor (gm_n3041, gm_n234, gm_n194, gm_n94);
	nand (gm_n3042, gm_n222, in_16, gm_n59, gm_n3041, gm_n275);
	nor (gm_n3043, gm_n384, in_21, gm_n85, gm_n3042);
	and (gm_n3044, gm_n221, gm_n73, in_12, gm_n264, gm_n224);
	nand (gm_n3045, gm_n138, gm_n72, in_20, gm_n3044);
	nor (gm_n3046, gm_n90, gm_n78, gm_n62, gm_n3006, gm_n369);
	nand (gm_n3047, gm_n348, gm_n323, in_18, gm_n3046);
	nand (gm_n3048, gm_n192, gm_n60, in_11, gm_n602, gm_n556);
	nor (gm_n3049, gm_n72, gm_n85, gm_n56, gm_n3048, gm_n293);
	or (gm_n3050, gm_n345, in_13, gm_n62, gm_n502, gm_n442);
	nor (gm_n3051, gm_n183, in_21, in_17, gm_n3050, gm_n328);
	or (gm_n3052, gm_n228, gm_n223, gm_n94);
	nor (gm_n3053, gm_n3052, gm_n274, gm_n60, gm_n633, gm_n269);
	nand (gm_n3054, gm_n72, in_20, gm_n56, gm_n3053);
	and (gm_n3055, gm_n77, gm_n73, in_12, gm_n612, gm_n233);
	nand (gm_n3056, gm_n495, gm_n72, in_20, gm_n3055);
	or (gm_n3057, gm_n344, gm_n76, gm_n62, gm_n432, gm_n480);
	nor (gm_n3058, gm_n103, gm_n72, gm_n55, gm_n3057, gm_n105);
	or (gm_n3059, gm_n461, in_13, gm_n62, gm_n503, gm_n344);
	nor (gm_n3060, gm_n103, gm_n72, gm_n55, gm_n3059, gm_n328);
	nor (gm_n3061, gm_n358, in_13, in_9, gm_n463, gm_n432);
	nand (gm_n3062, gm_n595, in_21, in_17, gm_n3061, gm_n373);
	and (gm_n3063, gm_n1067, gm_n81, in_8);
	and (gm_n3064, gm_n90, in_10, in_9, gm_n3063, gm_n532);
	nand (gm_n3065, gm_n166, gm_n146, gm_n119, gm_n3064);
	nand (gm_n3066, gm_n123, in_13, gm_n62, gm_n962);
	nor (gm_n3067, gm_n105, gm_n72, in_17, gm_n3066, gm_n441);
	or (gm_n3068, gm_n105, in_13, in_9, gm_n1542, gm_n406);
	nor (gm_n3069, gm_n374, in_21, in_17, gm_n3068);
	nor (gm_n3070, gm_n667, gm_n76, gm_n62, gm_n621, gm_n431);
	nand (gm_n3071, gm_n102, gm_n72, in_17, gm_n3070, gm_n523);
	nor (gm_n3072, gm_n369, gm_n90, gm_n78, gm_n775, gm_n491);
	nand (gm_n3073, gm_n436, gm_n164, in_18, gm_n3072);
	nand (gm_n3074, gm_n422, gm_n233, in_15, gm_n2416, gm_n394);
	nor (gm_n3075, gm_n72, gm_n85, gm_n56, gm_n3074);
	or (gm_n3076, gm_n290, gm_n155, gm_n60, gm_n695, gm_n393);
	nor (gm_n3077, gm_n72, gm_n85, gm_n56, gm_n3076);
	nor (gm_n3078, gm_n667, in_13, in_9, gm_n481, gm_n406);
	nand (gm_n3079, gm_n523, in_21, in_17, gm_n3078, gm_n373);
	nor (gm_n3080, gm_n168, gm_n60, gm_n94, gm_n508, gm_n213);
	nand (gm_n3081, in_21, in_20, gm_n56, gm_n3080, gm_n281);
	or (gm_n3082, gm_n248, in_14, gm_n78, gm_n467, gm_n438);
	nor (gm_n3083, gm_n368, gm_n89, gm_n119, gm_n3082);
	nand (gm_n3084, gm_n1101, gm_n143, in_15, gm_n1758, gm_n869);
	nor (gm_n3085, in_21, gm_n85, in_19, gm_n3084);
	nor (gm_n3086, gm_n667, in_13, in_9, gm_n481, gm_n257);
	nand (gm_n3087, gm_n104, in_21, in_17, gm_n3086, gm_n174);
	nor (gm_n3088, gm_n274, in_16, in_12, gm_n695, gm_n385);
	nand (gm_n3089, gm_n113, gm_n72, gm_n85, gm_n3088);
	nand (gm_n3090, in_10, in_9, in_8, gm_n624, gm_n69);
	nor (gm_n3091, gm_n132, gm_n119, in_14, gm_n3090, gm_n368);
	or (gm_n3092, gm_n213, gm_n73, gm_n59, gm_n2333, gm_n385);
	nor (gm_n3093, gm_n219, in_21, in_20, gm_n3092);
	nor (gm_n3094, gm_n99, gm_n90, gm_n78, gm_n362, gm_n287);
	nand (gm_n3095, gm_n436, gm_n348, gm_n119, gm_n3094);
	nand (gm_n3096, gm_n93, gm_n124, in_5, gm_n454, in_8);
	nor (gm_n3097, gm_n121, gm_n76, gm_n62, gm_n3096, gm_n480);
	nand (gm_n3098, gm_n311, in_21, in_17, gm_n3097);
	nand (gm_n3099, gm_n305, gm_n81, gm_n94);
	nor (gm_n3100, gm_n263, in_16, in_12, gm_n3099, gm_n276);
	nand (gm_n3101, gm_n113, in_21, gm_n85, gm_n3100);
	nor (gm_n3102, gm_n213, in_16, gm_n59, gm_n2826, gm_n354);
	nand (gm_n3103, gm_n383, in_21, in_20, gm_n3102);
	nor (gm_n3104, gm_n370, gm_n90, gm_n78, gm_n467, gm_n389);
	nand (gm_n3105, gm_n243, gm_n88, gm_n119, gm_n3104);
	nand (gm_n3106, gm_n3101, gm_n3098, gm_n3095, gm_n3105, gm_n3103);
	nor (gm_n3107, gm_n114, in_16, in_12, gm_n2963, gm_n274);
	nand (gm_n3108, gm_n113, gm_n72, gm_n85, gm_n3107);
	nor (gm_n3109, gm_n362, gm_n78, in_9, gm_n2402);
	nand (gm_n3110, gm_n102, gm_n72, in_17, gm_n3109, gm_n1076);
	nor (gm_n3111, gm_n149, gm_n514, in_13, gm_n438, gm_n328);
	nand (gm_n3112, gm_n311, gm_n72, in_17, gm_n3111);
	nand (gm_n3113, gm_n3112, gm_n3110, gm_n3108);
	nor (gm_n3114, gm_n213, in_16, gm_n59, gm_n1542, gm_n385);
	nand (gm_n3115, gm_n138, in_21, gm_n85, gm_n3114);
	nor (gm_n3116, gm_n115, gm_n73, gm_n59, gm_n152, gm_n116);
	nand (gm_n3117, gm_n138, in_21, in_20, gm_n3116);
	nor (gm_n3118, gm_n263, gm_n168, in_15, gm_n293, gm_n278);
	nand (gm_n3119, in_21, gm_n85, in_19, gm_n3118);
	nand (gm_n3120, gm_n3119, gm_n3117, gm_n3115);
	nor (gm_n3121, gm_n3106, gm_n3093, gm_n3091, gm_n3120, gm_n3113);
	nand (gm_n3122, gm_n90, in_10, gm_n62, gm_n2727, gm_n532);
	nor (gm_n3123, gm_n211, gm_n89, gm_n119, gm_n3122);
	nand (gm_n3124, gm_n222, gm_n392, in_15, gm_n1095, gm_n268);
	nor (gm_n3125, gm_n72, gm_n85, gm_n56, gm_n3124);
	nand (gm_n3126, gm_n448, gm_n214, in_15, gm_n1569, gm_n545);
	nor (gm_n3127, gm_n72, gm_n85, gm_n56, gm_n3126);
	nor (gm_n3128, gm_n3127, gm_n3125, gm_n3123);
	nand (gm_n3129, gm_n61, in_16, gm_n59, gm_n2885, gm_n222);
	nor (gm_n3130, gm_n384, in_21, in_20, gm_n3129);
	nand (gm_n3131, gm_n106, gm_n76, in_9, gm_n1012, gm_n255);
	nor (gm_n3132, gm_n312, gm_n72, gm_n55, gm_n3131);
	or (gm_n3133, gm_n115, in_16, gm_n59, gm_n2002, gm_n354);
	nor (gm_n3134, gm_n58, in_21, gm_n85, gm_n3133);
	nor (gm_n3135, gm_n3134, gm_n3132, gm_n3130);
	nand (gm_n3136, gm_n3121, gm_n3089, gm_n3087, gm_n3135, gm_n3128);
	nor (gm_n3137, gm_n92, in_14, in_10, gm_n438, gm_n99);
	nand (gm_n3138, gm_n131, gm_n86, gm_n119, gm_n3137);
	nor (gm_n3139, gm_n190, in_13, in_12, gm_n1150);
	nand (gm_n3140, gm_n102, in_21, gm_n55, gm_n3139, gm_n405);
	and (gm_n3141, in_10, gm_n62, in_8, gm_n601, gm_n600);
	nand (gm_n3142, gm_n199, in_18, in_14, gm_n3141, gm_n200);
	nand (gm_n3143, gm_n3142, gm_n3140, gm_n3138);
	nor (gm_n3144, gm_n257, gm_n76, gm_n62, gm_n597, gm_n463);
	nand (gm_n3145, gm_n255, in_21, gm_n55, gm_n3144, gm_n373);
	nor (gm_n3146, gm_n76, in_9, gm_n94, gm_n2237, gm_n461);
	nand (gm_n3147, gm_n174, in_21, in_17, gm_n3146, gm_n405);
	nor (gm_n3148, gm_n95, in_14, gm_n78, gm_n807, gm_n149);
	nand (gm_n3149, gm_n200, gm_n129, gm_n119, gm_n3148);
	nand (gm_n3150, gm_n3149, gm_n3147, gm_n3145);
	nor (gm_n3151, gm_n3136, gm_n3085, gm_n3083, gm_n3150, gm_n3143);
	nand (gm_n3152, gm_n392, in_15, in_11, gm_n756, gm_n171);
	nor (gm_n3153, gm_n72, in_20, gm_n56, gm_n3152, gm_n485);
	or (gm_n3154, gm_n818, in_13, in_9, gm_n344, gm_n358);
	nor (gm_n3155, gm_n313, gm_n72, in_17, gm_n3154, gm_n374);
	nand (gm_n3156, gm_n79, in_16, in_12, gm_n953, gm_n221);
	nor (gm_n3157, gm_n912, in_21, in_20, gm_n3156);
	nor (gm_n3158, gm_n3157, gm_n3155, gm_n3153);
	or (gm_n3159, gm_n155, gm_n73, gm_n59, gm_n1906, gm_n319);
	nor (gm_n3160, gm_n58, in_21, in_20, gm_n3159);
	nor (gm_n3161, gm_n105, gm_n72, gm_n55, gm_n646, gm_n388);
	or (gm_n3162, gm_n196, gm_n73, gm_n59, gm_n220, gm_n213);
	nor (gm_n3163, gm_n912, gm_n72, in_20, gm_n3162);
	nor (gm_n3164, gm_n3163, gm_n3161, gm_n3160);
	nand (gm_n3165, gm_n3151, gm_n3081, gm_n3079, gm_n3164, gm_n3158);
	nor (gm_n3166, gm_n257, gm_n76, gm_n62, gm_n502, gm_n481);
	nand (gm_n3167, gm_n120, gm_n72, gm_n55, gm_n3166, gm_n405);
	nor (gm_n3168, gm_n362, in_14, gm_n78, gm_n376, gm_n370);
	nand (gm_n3169, gm_n806, gm_n199, in_18, gm_n3168);
	nor (gm_n3170, gm_n269, gm_n263, in_15, gm_n1170, gm_n764);
	nand (gm_n3171, in_21, in_20, in_19, gm_n3170);
	nand (gm_n3172, gm_n3171, gm_n3169, gm_n3167);
	nor (gm_n3173, gm_n514, gm_n76, gm_n62, gm_n597, gm_n463);
	nand (gm_n3174, gm_n174, in_21, gm_n55, gm_n3173, gm_n523);
	nor (gm_n3175, gm_n287, gm_n358, gm_n76, gm_n350, gm_n662);
	nand (gm_n3176, gm_n174, gm_n72, gm_n55, gm_n3175);
	nor (gm_n3177, gm_n147, in_14, in_10, gm_n438, gm_n389);
	nand (gm_n3178, gm_n436, gm_n146, in_18, gm_n3177);
	nand (gm_n3179, gm_n3178, gm_n3176, gm_n3174);
	nor (gm_n3180, gm_n3165, gm_n3077, gm_n3075, gm_n3179, gm_n3172);
	nand (gm_n3181, gm_n106, gm_n76, gm_n62, gm_n2712, gm_n255);
	nor (gm_n3182, gm_n312, in_21, gm_n55, gm_n3181);
	or (gm_n3183, gm_n442, gm_n76, in_9, gm_n597, gm_n502);
	nor (gm_n3184, gm_n103, in_21, in_17, gm_n3183, gm_n105);
	or (gm_n3185, gm_n95, gm_n90, in_10, gm_n248, gm_n147);
	nor (gm_n3186, gm_n368, gm_n167, gm_n119, gm_n3185);
	nor (gm_n3187, gm_n3186, gm_n3184, gm_n3182);
	nor (gm_n3188, gm_n1639, gm_n312, in_21);
	nand (gm_n3189, gm_n171, gm_n60, in_11, gm_n1929, gm_n449);
	nor (gm_n3190, gm_n72, in_20, gm_n56, gm_n3189, gm_n191);
	or (gm_n3191, gm_n133, in_14, gm_n78, gm_n349, gm_n208);
	nor (gm_n3192, gm_n437, gm_n368, in_18, gm_n3191);
	nor (gm_n3193, gm_n3192, gm_n3190, gm_n3188);
	nand (gm_n3194, gm_n3180, gm_n3073, gm_n3071, gm_n3193, gm_n3187);
	nor (gm_n3195, gm_n393, gm_n158, gm_n60, gm_n760, gm_n515);
	nand (gm_n3196, gm_n72, gm_n85, in_19, gm_n3195);
	nor (gm_n3197, gm_n349, gm_n248, gm_n76, gm_n480, gm_n375);
	nand (gm_n3198, gm_n206, gm_n72, gm_n55, gm_n3197);
	nor (gm_n3199, gm_n92, gm_n90, in_10, gm_n247, gm_n208);
	nand (gm_n3200, gm_n806, gm_n86, gm_n119, gm_n3199);
	nand (gm_n3201, gm_n3200, gm_n3198, gm_n3196);
	and (gm_n3202, gm_n64, in_16, gm_n59, gm_n586, gm_n77);
	nand (gm_n3203, gm_n138, in_21, in_20, gm_n3202);
	and (gm_n3204, gm_n392, gm_n64, gm_n60, gm_n427, gm_n1101);
	nand (gm_n3205, in_21, in_20, gm_n56, gm_n3204);
	and (gm_n3206, gm_n392, gm_n56, gm_n60, gm_n1068, gm_n394);
	nand (gm_n3207, gm_n3206, gm_n72, gm_n85);
	nand (gm_n3208, gm_n3207, gm_n3205, gm_n3203);
	nor (gm_n3209, gm_n3194, gm_n3069, gm_n3067, gm_n3208, gm_n3201);
	or (gm_n3210, gm_n328, gm_n286, gm_n76, gm_n438, gm_n406);
	nor (gm_n3211, gm_n374, gm_n72, in_17, gm_n3210);
	nand (gm_n3212, gm_n600, gm_n90, in_10, gm_n333, gm_n995);
	nor (gm_n3213, gm_n212, gm_n824, gm_n119, gm_n3212);
	nand (gm_n3214, gm_n1076, in_13, in_9, gm_n1012, gm_n402);
	nor (gm_n3215, gm_n388, gm_n72, gm_n55, gm_n3214);
	nor (gm_n3216, gm_n3215, gm_n3213, gm_n3211);
	and (gm_n3217, gm_n206, gm_n72, in_17, gm_n567, gm_n339);
	or (gm_n3218, gm_n344, in_10, gm_n62, gm_n467, gm_n462);
	nor (gm_n3219, gm_n132, in_18, gm_n90, gm_n3218, gm_n244);
	nand (gm_n3220, gm_n233, in_16, in_12, gm_n1198, gm_n733);
	nor (gm_n3221, gm_n219, in_21, gm_n85, gm_n3220);
	nor (gm_n3222, gm_n3221, gm_n3219, gm_n3217);
	nand (gm_n3223, gm_n3209, gm_n3065, gm_n3062, gm_n3222, gm_n3216);
	nor (gm_n3224, gm_n135, gm_n158, gm_n60, gm_n293, gm_n159);
	nand (gm_n3225, gm_n72, in_20, in_19, gm_n3224);
	nand (gm_n3226, gm_n245, gm_n146, in_18, gm_n2310);
	nor (gm_n3227, in_14, gm_n78, in_9, gm_n467, gm_n153);
	nand (gm_n3228, gm_n245, gm_n129, in_18, gm_n3227);
	nand (gm_n3229, gm_n3228, gm_n3226, gm_n3225);
	nor (gm_n3230, gm_n208, in_14, gm_n78, gm_n362, gm_n349);
	nand (gm_n3231, gm_n200, gm_n146, in_18, gm_n3230);
	nor (gm_n3232, gm_n116, gm_n76, in_12, gm_n213);
	nand (gm_n3233, gm_n254, gm_n72, in_17, gm_n3232, gm_n339);
	nor (gm_n3234, gm_n514, in_13, gm_n62, gm_n345, gm_n430);
	nand (gm_n3235, gm_n206, in_21, in_17, gm_n3234, gm_n1076);
	nand (gm_n3236, gm_n3235, gm_n3233, gm_n3231);
	nor (gm_n3237, gm_n3223, gm_n3060, gm_n3058, gm_n3236, gm_n3229);
	or (gm_n3238, gm_n105, in_13, in_9, gm_n1150, gm_n431);
	nor (gm_n3239, gm_n479, gm_n72, in_17, gm_n3238);
	nand (gm_n3240, gm_n224, gm_n64, gm_n60, gm_n545, gm_n486);
	nor (gm_n3241, gm_n72, gm_n85, in_19, gm_n3240);
	or (gm_n3242, gm_n114, gm_n73, gm_n59, gm_n520, gm_n263);
	nor (gm_n3243, gm_n912, gm_n72, in_20, gm_n3242);
	nor (gm_n3244, gm_n3243, gm_n3241, gm_n3239);
	nand (gm_n3245, in_14, in_10, in_9, gm_n2276, gm_n713);
	nor (gm_n3246, gm_n841, gm_n211, in_18, gm_n3245);
	nand (gm_n3247, gm_n555, gm_n60, in_11, gm_n1398, gm_n556);
	nor (gm_n3248, gm_n72, gm_n85, in_19, gm_n3247, gm_n293);
	nand (gm_n3249, gm_n154, in_16, in_12, gm_n3041, gm_n571);
	nor (gm_n3250, gm_n384, gm_n72, in_20, gm_n3249);
	nor (gm_n3251, gm_n3250, gm_n3248, gm_n3246);
	nand (gm_n3252, gm_n3237, gm_n3056, gm_n3054, gm_n3251, gm_n3244);
	nor (gm_n3253, gm_n115, in_16, gm_n59, gm_n385, gm_n153);
	nand (gm_n3254, gm_n57, in_21, gm_n85, gm_n3253);
	nor (gm_n3255, gm_n213, gm_n73, gm_n59, gm_n2956, gm_n220);
	nand (gm_n3256, gm_n296, in_21, gm_n85, gm_n3255);
	nor (gm_n3257, gm_n207, gm_n909, in_14, gm_n605);
	nand (gm_n3258, gm_n348, gm_n88, in_18, gm_n3257);
	nand (gm_n3259, gm_n3258, gm_n3256, gm_n3254);
	nor (gm_n3260, gm_n190, in_16, gm_n59, gm_n354, gm_n324);
	nand (gm_n3261, gm_n138, in_21, in_20, gm_n3260);
	nand (gm_n3262, gm_n351, gm_n348, in_18, gm_n436);
	nor (gm_n3263, gm_n95, gm_n90, gm_n78, gm_n526, gm_n467);
	nand (gm_n3264, gm_n166, gm_n164, in_18, gm_n3263);
	nand (gm_n3265, gm_n3264, gm_n3262, gm_n3261);
	nor (gm_n3266, gm_n3252, gm_n3051, gm_n3049, gm_n3265, gm_n3259);
	nand (gm_n3267, gm_n192, gm_n154, in_15, gm_n1427, gm_n281);
	nor (gm_n3268, gm_n72, gm_n85, gm_n56, gm_n3267);
	nand (gm_n3269, gm_n579, gm_n76, gm_n62, gm_n471, gm_n405);
	nor (gm_n3270, gm_n441, in_21, in_17, gm_n3269);
	nand (gm_n3271, gm_n523, in_13, gm_n62, gm_n788, gm_n306);
	nor (gm_n3272, gm_n312, in_21, gm_n55, gm_n3271);
	nor (gm_n3273, gm_n3272, gm_n3270, gm_n3268);
	and (gm_n3274, in_21, gm_n85, gm_n56, gm_n448, gm_n83);
	nand (gm_n3275, in_10, in_9, gm_n94, gm_n1120, gm_n1011);
	nor (gm_n3276, gm_n87, in_18, gm_n90, gm_n3275, gm_n132);
	nand (gm_n3277, gm_n392, gm_n143, in_15, gm_n2624, gm_n448);
	nor (gm_n3278, gm_n72, gm_n85, gm_n56, gm_n3277);
	nor (gm_n3279, gm_n3278, gm_n3276, gm_n3274);
	nand (gm_n3280, gm_n3266, gm_n3047, gm_n3045, gm_n3279, gm_n3273);
	nor (gm_n3281, gm_n293, gm_n297, gm_n60, gm_n760, gm_n515);
	nand (gm_n3282, in_21, gm_n85, gm_n56, gm_n3281);
	nor (gm_n3283, gm_n274, in_16, in_12, gm_n1125, gm_n354);
	nand (gm_n3284, gm_n179, in_21, in_20, gm_n3283);
	nor (gm_n3285, gm_n133, in_14, gm_n78, gm_n247, gm_n149);
	nand (gm_n3286, gm_n166, gm_n164, gm_n119, gm_n3285);
	nand (gm_n3287, gm_n3286, gm_n3284, gm_n3282);
	nor (gm_n3288, gm_n114, gm_n73, gm_n59, gm_n3099, gm_n158);
	nand (gm_n3289, gm_n383, gm_n72, in_20, gm_n3288);
	nor (gm_n3290, gm_n190, gm_n73, gm_n59, gm_n1191, gm_n385);
	nand (gm_n3291, gm_n383, gm_n72, gm_n85, gm_n3290);
	and (gm_n3292, gm_n1157, gm_n90, in_10, gm_n829, gm_n600);
	nand (gm_n3293, gm_n348, gm_n245, gm_n119, gm_n3292);
	nand (gm_n3294, gm_n3293, gm_n3291, gm_n3289);
	nor (gm_n3295, gm_n3280, gm_n3043, gm_n3040, gm_n3294, gm_n3287);
	or (gm_n3296, gm_n155, gm_n74, gm_n60, gm_n1319, gm_n159);
	nor (gm_n3297, in_21, in_20, gm_n56, gm_n3296);
	or (gm_n3298, gm_n609, in_13, in_9, gm_n462, gm_n406);
	nor (gm_n3299, gm_n105, in_21, gm_n55, gm_n3298, gm_n479);
	or (gm_n3300, gm_n430, gm_n76, in_9, gm_n462, gm_n442);
	nor (gm_n3301, gm_n121, gm_n72, in_17, gm_n3300, gm_n312);
	nor (gm_n3302, gm_n3301, gm_n3299, gm_n3297);
	nand (gm_n3303, gm_n110, in_13, in_9, gm_n1049, gm_n314);
	nor (gm_n3304, gm_n441, in_21, in_17, gm_n3303, gm_n662);
	nand (gm_n3305, gm_n78, gm_n62, gm_n94, gm_n1263, gm_n532);
	nor (gm_n3306, gm_n211, in_18, gm_n90, gm_n3305, gm_n167);
	or (gm_n3307, gm_n207, in_10, gm_n62, gm_n1664, gm_n375);
	nor (gm_n3308, gm_n441, in_21, in_17, gm_n3307);
	nor (gm_n3309, gm_n3308, gm_n3306, gm_n3304);
	nand (gm_n3310, gm_n3295, gm_n3039, gm_n3037, gm_n3309, gm_n3302);
	nor (gm_n3311, gm_n297, in_16, in_12, gm_n319, gm_n230);
	nand (gm_n3312, gm_n138, gm_n72, gm_n85, gm_n3311);
	nor (gm_n3313, gm_n133, in_10, gm_n62, gm_n462, gm_n430);
	nand (gm_n3314, gm_n131, in_18, gm_n90, gm_n3313, gm_n367);
	or (gm_n3315, gm_n228, gm_n141, gm_n94);
	nor (gm_n3316, gm_n227, gm_n73, in_12, gm_n3315, gm_n158);
	nand (gm_n3317, gm_n296, in_21, gm_n85, gm_n3316);
	nand (gm_n3318, gm_n3317, gm_n3314, gm_n3312);
	nand (gm_n3319, gm_n243, gm_n200, gm_n119, gm_n2979, gm_n449);
	nand (gm_n3320, gm_n327, gm_n72, gm_n55, gm_n3175);
	and (gm_n3321, gm_n154, in_16, gm_n59, gm_n1179, gm_n949);
	nand (gm_n3322, gm_n495, in_21, in_20, gm_n3321);
	nand (gm_n3323, gm_n3322, gm_n3320, gm_n3319);
	nor (gm_n3324, gm_n3310, gm_n3035, gm_n3033, gm_n3323, gm_n3318);
	nand (gm_n3325, gm_n123, gm_n76, gm_n62, gm_n186, gm_n126);
	nor (gm_n3326, gm_n184, gm_n72, gm_n55, gm_n3325, gm_n312);
	nand (gm_n3327, gm_n122, in_13, gm_n62, gm_n880, gm_n340);
	nor (gm_n3328, gm_n479, in_21, gm_n55, gm_n3327);
	or (gm_n3329, gm_n406, gm_n76, in_9, gm_n462, gm_n443);
	nor (gm_n3330, gm_n388, gm_n72, in_17, gm_n3329, gm_n375);
	nor (gm_n3331, gm_n3330, gm_n3328, gm_n3326);
	nand (gm_n3332, gm_n78, gm_n62, in_8, gm_n2074, gm_n334);
	nor (gm_n3333, gm_n132, gm_n119, gm_n90, gm_n3332, gm_n824);
	or (gm_n3334, gm_n514, gm_n76, gm_n62, gm_n621, gm_n502);
	nor (gm_n3335, gm_n313, gm_n72, gm_n55, gm_n3334, gm_n374);
	nand (gm_n3336, gm_n602, gm_n624, gm_n90, gm_n756);
	nor (gm_n3337, gm_n212, gm_n824, in_18, gm_n3336);
	nor (gm_n3338, gm_n3337, gm_n3335, gm_n3333);
	nand (gm_n3339, gm_n3324, gm_n3031, gm_n3029, gm_n3338, gm_n3331);
	or (gm_n3340, gm_n262, in_21, in_20, gm_n1646);
	nor (gm_n3341, gm_n442, gm_n76, gm_n62, gm_n502, gm_n481);
	nand (gm_n3342, gm_n339, in_21, in_17, gm_n3341, gm_n373);
	nor (gm_n3343, gm_n60, gm_n90, gm_n76, t_2, in_16);
	nand (gm_n3344, gm_n697, in_21, in_20, gm_n3343);
	nand (gm_n3345, gm_n3344, gm_n3342, gm_n3340);
	and (gm_n3346, gm_n77, in_16, gm_n59, gm_n2283, gm_n143);
	nand (gm_n3347, gm_n57, in_21, gm_n85, gm_n3346);
	and (gm_n3348, gm_n214, gm_n59, gm_n94, gm_n1379, gm_n221);
	nand (gm_n3349, in_21, in_20, in_16, gm_n3348, gm_n179);
	and (gm_n3350, gm_n64, in_16, in_12, gm_n2860, gm_n733);
	nand (gm_n3351, gm_n697, in_21, gm_n85, gm_n3350);
	nand (gm_n3352, gm_n3351, gm_n3349, gm_n3347);
	nor (gm_n3353, gm_n3339, gm_n3027, gm_n3025, gm_n3352, gm_n3345);
	nor (gm_n3354, gm_n287, gm_n90, in_10, gm_n775, gm_n467);
	nand (gm_n3355, gm_n367, gm_n245, in_18, gm_n3354);
	or (gm_n3356, gm_n461, in_13, in_9, gm_n597, gm_n344);
	or (gm_n3357, gm_n103, in_21, in_17, gm_n3356, gm_n328);
	and (gm_n3358, in_14, in_10, in_9, gm_n880, gm_n91);
	nand (gm_n3359, gm_n146, gm_n88, gm_n119, gm_n3358);
	nand (gm_n3360, gm_n3355, gm_n3353, gm_n3023, gm_n3359, gm_n3357);
	nor (gm_n3361, gm_n256, gm_n208, gm_n76, gm_n438, gm_n406);
	nand (gm_n3362, gm_n254, gm_n72, in_17, gm_n3361);
	nor (gm_n3363, gm_n609, gm_n76, gm_n62, gm_n597, gm_n406);
	nand (gm_n3364, gm_n254, in_21, in_17, gm_n3363, gm_n595);
	and (gm_n3365, gm_n61, in_16, gm_n59, gm_n423, gm_n64);
	nand (gm_n3366, gm_n296, gm_n72, in_20, gm_n3365);
	nand (gm_n3367, gm_n3366, gm_n3364, gm_n3362);
	nor (gm_n3368, gm_n93, in_6, gm_n97, gm_n141, gm_n94);
	nand (gm_n3369, gm_n281, gm_n233, gm_n60, gm_n3368, gm_n545);
	nor (gm_n3370, in_21, gm_n85, in_19, gm_n3369);
	nor (out_7, gm_n3367, gm_n3360, gm_n3021, gm_n3370);
	nand (gm_n3372, gm_n79, in_16, gm_n59, gm_n2547, gm_n949);
	nor (gm_n3373, gm_n384, in_21, gm_n85, gm_n3372);
	nand (gm_n3374, gm_n422, gm_n264, in_15, gm_n2172, gm_n1101);
	nor (gm_n3375, gm_n72, in_20, in_19, gm_n3374);
	and (gm_n3376, gm_n75, in_19, in_15, gm_n2542, gm_n545);
	nand (gm_n3377, gm_n3376, in_21, gm_n85);
	nor (gm_n3378, gm_n596, in_13, in_9, gm_n597, gm_n480);
	nand (gm_n3379, gm_n174, in_21, in_17, gm_n3378, gm_n1076);
	or (gm_n3380, gm_n227, gm_n73, in_12, gm_n230, gm_n158);
	nor (gm_n3381, gm_n384, in_21, in_20, gm_n3380);
	or (gm_n3382, gm_n93, in_6, gm_n97, gm_n229, gm_n94);
	or (gm_n3383, gm_n293, gm_n190, in_15, gm_n3382, gm_n643);
	nor (gm_n3384, gm_n72, gm_n85, in_19, gm_n3383);
	nor (gm_n3385, gm_n168, gm_n115, gm_n60, gm_n1698, gm_n269);
	nand (gm_n3386, in_21, in_20, gm_n56, gm_n3385);
	and (gm_n3387, gm_n1144, gm_n60, gm_n63, gm_n580, gm_n545);
	nand (gm_n3388, in_21, gm_n85, gm_n56, gm_n3387, gm_n268);
	and (gm_n3389, gm_n1011, in_10, in_9, gm_n1446);
	and (gm_n3390, gm_n254, gm_n72, gm_n55, gm_n3389, gm_n595);
	or (gm_n3391, gm_n431, gm_n76, in_9, gm_n481, gm_n443);
	nor (gm_n3392, gm_n184, in_21, in_17, gm_n3391, gm_n620);
	nor (gm_n3393, gm_n358, gm_n76, gm_n62, gm_n988, gm_n430);
	nand (gm_n3394, gm_n254, in_21, gm_n55, gm_n3393, gm_n405);
	and (gm_n3395, gm_n733, gm_n73, in_12, gm_n2065, gm_n264);
	nand (gm_n3396, gm_n383, in_21, gm_n85, gm_n3395);
	or (gm_n3397, gm_n447, gm_n115, gm_n60, gm_n760, gm_n552);
	nor (gm_n3398, in_21, in_20, in_19, gm_n3397);
	and (gm_n3399, gm_n122, in_21, in_17, gm_n2987, gm_n174);
	nor (gm_n3400, gm_n263, in_16, gm_n59, gm_n1203, gm_n319);
	nand (gm_n3401, gm_n383, in_21, in_20, gm_n3400);
	nand (gm_n3402, gm_n454, gm_n291, in_8);
	nor (gm_n3403, gm_n313, gm_n76, gm_n62, gm_n3402, gm_n480);
	nand (gm_n3404, gm_n254, in_21, gm_n55, gm_n3403);
	nand (gm_n3405, gm_n214, gm_n379, in_15, gm_n449, gm_n265);
	nor (gm_n3406, in_21, gm_n85, gm_n56, gm_n3405);
	nand (gm_n3407, gm_n233, gm_n73, gm_n59, gm_n870, gm_n221);
	nor (gm_n3408, gm_n912, gm_n72, in_20, gm_n3407);
	or (gm_n3409, gm_n312, in_21, gm_n55, gm_n2149, gm_n313);
	nor (gm_n3410, gm_n796, gm_n76, gm_n62, gm_n480, gm_n344);
	nand (gm_n3411, gm_n311, gm_n72, gm_n55, gm_n3410, gm_n595);
	and (gm_n3412, in_14, gm_n76, gm_n59, gm_n1071, gm_n64);
	and (gm_n3413, gm_n200, gm_n146, gm_n119, gm_n3412);
	or (gm_n3414, gm_n158, gm_n74, in_15, gm_n764, gm_n135);
	nor (gm_n3415, gm_n72, gm_n85, gm_n56, gm_n3414);
	nand (gm_n3416, gm_n296, gm_n72, in_20, gm_n1940);
	and (gm_n3417, gm_n214, gm_n192, gm_n60, gm_n1947, gm_n394);
	nand (gm_n3418, gm_n72, gm_n85, gm_n56, gm_n3417);
	nand (gm_n3419, gm_n186, gm_n76, in_9, gm_n340, gm_n187);
	nor (gm_n3420, gm_n121, gm_n72, gm_n55, gm_n3419, gm_n620);
	and (gm_n3421, gm_n174, gm_n72, gm_n55, gm_n1376, gm_n405);
	nand (gm_n3422, gm_n131, gm_n129, in_18, gm_n2899);
	nor (gm_n3423, gm_n115, gm_n73, in_12, gm_n385, gm_n292);
	nand (gm_n3424, gm_n138, gm_n72, in_20, gm_n3423);
	nand (gm_n3425, gm_n392, in_15, gm_n63, gm_n601, gm_n555);
	nor (gm_n3426, in_21, gm_n85, gm_n56, gm_n3425, gm_n485);
	nor (gm_n3427, gm_n72, gm_n85, gm_n56, gm_n1402, gm_n485);
	and (gm_n3428, gm_n64, gm_n73, in_12, gm_n1147, gm_n303);
	nand (gm_n3429, gm_n57, in_21, in_20, gm_n3428);
	nor (gm_n3430, gm_n480, in_13, in_9, gm_n481, gm_n463);
	nand (gm_n3431, gm_n327, gm_n72, gm_n55, gm_n3430, gm_n595);
	or (gm_n3432, gm_n270, gm_n60, in_11, gm_n643, gm_n283);
	nor (gm_n3433, gm_n72, in_20, gm_n56, gm_n3432, gm_n393);
	or (gm_n3434, gm_n190, in_16, gm_n59, gm_n1719, gm_n385);
	nor (gm_n3435, gm_n496, gm_n72, in_20, gm_n3434);
	and (gm_n3436, gm_n79, gm_n73, in_12, gm_n2172, gm_n221);
	nand (gm_n3437, gm_n383, in_21, gm_n85, gm_n3436);
	nor (gm_n3438, gm_n159, gm_n60, gm_n63, gm_n2690, gm_n240);
	nand (gm_n3439, gm_n72, gm_n85, in_19, gm_n3438, gm_n1101);
	or (gm_n3440, in_7, in_6, in_5, gm_n223, in_8);
	nor (gm_n3441, gm_n760, gm_n155, in_15, gm_n3440);
	and (gm_n3442, in_21, in_20, gm_n56, gm_n3441, gm_n1101);
	or (gm_n3443, gm_n430, gm_n76, gm_n62, gm_n1583, gm_n431);
	or (gm_n3444, gm_n103, gm_n72, in_17, gm_n3443, gm_n184);
	nor (gm_n3445, gm_n514, gm_n76, gm_n62, gm_n481, gm_n596);
	nand (gm_n3446, gm_n405, in_21, in_17, gm_n3445, gm_n327);
	nor (gm_n3447, gm_n667, gm_n76, in_9, gm_n481, gm_n461);
	nand (gm_n3448, gm_n174, in_21, in_17, gm_n3447, gm_n1076);
	nor (gm_n3449, gm_n271, gm_n60, gm_n63, gm_n770, gm_n764);
	nand (gm_n3450, gm_n72, in_20, gm_n56, gm_n3449, gm_n268);
	nor (gm_n3451, gm_n190, gm_n73, in_12, gm_n835, gm_n319);
	nand (gm_n3452, gm_n179, in_21, gm_n85, gm_n3451);
	nand (gm_n3453, gm_n3448, gm_n3446, gm_n3444, gm_n3452, gm_n3450);
	and (gm_n3454, gm_n305, gm_n81, in_8);
	nand (gm_n3455, gm_n90, gm_n78, gm_n62, gm_n3454, gm_n600);
	nor (gm_n3456, gm_n1989, gm_n211, in_18, gm_n3455);
	or (gm_n3457, gm_n406, gm_n76, in_9, gm_n743, gm_n463);
	nor (gm_n3458, gm_n312, gm_n72, gm_n55, gm_n3457, gm_n313);
	or (gm_n3459, gm_n344, gm_n76, gm_n62, gm_n480, gm_n359);
	nor (gm_n3460, gm_n103, gm_n72, gm_n55, gm_n3459, gm_n256);
	nor (gm_n3461, gm_n3456, gm_n3453, gm_n3442, gm_n3460, gm_n3458);
	or (gm_n3462, gm_n406, in_13, gm_n62, gm_n463, gm_n359);
	nor (gm_n3463, gm_n121, in_21, in_17, gm_n3462, gm_n620);
	or (gm_n3464, gm_n115, in_13, in_12, gm_n1223);
	nor (gm_n3465, gm_n184, in_21, in_17, gm_n3464, gm_n374);
	nand (gm_n3466, in_14, in_10, in_9, gm_n1158, gm_n2916);
	nor (gm_n3467, gm_n841, gm_n211, in_18, gm_n3466);
	nor (gm_n3468, gm_n3467, gm_n3465, gm_n3463);
	or (gm_n3469, gm_n240, gm_n68, in_14, gm_n671, gm_n369);
	nor (gm_n3470, gm_n368, gm_n132, in_18, gm_n3469);
	nand (gm_n3471, in_14, gm_n78, gm_n62, gm_n838, gm_n600);
	nor (gm_n3472, gm_n368, gm_n132, in_18, gm_n3471);
	or (gm_n3473, in_14, in_10, in_9, gm_n2244, gm_n133);
	nor (gm_n3474, gm_n531, gm_n89, gm_n119, gm_n3473);
	nor (gm_n3475, gm_n3474, gm_n3472, gm_n3470);
	nand (gm_n3476, gm_n3461, gm_n3439, gm_n3437, gm_n3475, gm_n3468);
	or (gm_n3477, gm_n183, gm_n72, in_17, gm_n1901, gm_n375);
	nand (gm_n3478, gm_n339, in_21, in_17, gm_n1643, gm_n373);
	nor (gm_n3479, gm_n609, in_13, gm_n62, gm_n621, gm_n480);
	nand (gm_n3480, gm_n120, gm_n72, in_17, gm_n3479, gm_n523);
	nand (gm_n3481, gm_n3480, gm_n3478, gm_n3477);
	nor (gm_n3482, in_13, gm_n62, gm_n94, gm_n431, gm_n161);
	nand (gm_n3483, gm_n104, gm_n72, in_17, gm_n3482, gm_n327);
	nor (gm_n3484, gm_n461, gm_n76, in_9, gm_n344, gm_n796);
	nand (gm_n3485, gm_n311, gm_n72, in_17, gm_n3484, gm_n595);
	nor (gm_n3486, gm_n461, gm_n76, in_9, gm_n1583, gm_n502);
	nand (gm_n3487, gm_n102, in_21, in_17, gm_n3486, gm_n122);
	nand (gm_n3488, gm_n3487, gm_n3485, gm_n3483);
	nor (gm_n3489, gm_n3476, gm_n3435, gm_n3433, gm_n3488, gm_n3481);
	nand (gm_n3490, gm_n90, gm_n78, in_9, gm_n1446, gm_n713);
	nor (gm_n3491, gm_n246, gm_n130, in_18, gm_n3490);
	or (gm_n3492, gm_n247, in_14, in_10, gm_n369, gm_n350);
	nor (gm_n3493, gm_n167, gm_n87, gm_n119, gm_n3492);
	or (gm_n3494, gm_n667, in_13, in_9, gm_n462, gm_n461);
	nor (gm_n3495, gm_n183, in_21, in_17, gm_n3494, gm_n121);
	nor (gm_n3496, gm_n3495, gm_n3493, gm_n3491);
	or (gm_n3497, gm_n393, gm_n297, gm_n60, gm_n3440, gm_n633);
	nor (gm_n3498, gm_n72, gm_n85, gm_n56, gm_n3497);
	nand (gm_n3499, gm_n422, gm_n143, in_15, gm_n678, gm_n448);
	nor (gm_n3500, gm_n72, in_20, gm_n56, gm_n3499);
	nand (gm_n3501, gm_n91, gm_n78, gm_n62, gm_n2605);
	nor (gm_n3502, gm_n184, gm_n72, gm_n55, gm_n3501, gm_n374);
	nor (gm_n3503, gm_n3502, gm_n3500, gm_n3498);
	nand (gm_n3504, gm_n3489, gm_n3431, gm_n3429, gm_n3503, gm_n3496);
	nor (gm_n3505, gm_n807, in_14, in_10, gm_n389, gm_n349);
	nand (gm_n3506, gm_n164, gm_n88, gm_n119, gm_n3505);
	and (gm_n3507, gm_n143, in_16, gm_n59, gm_n1970, gm_n221);
	nand (gm_n3508, gm_n296, gm_n72, gm_n85, gm_n3507);
	nor (gm_n3509, gm_n282, gm_n60, in_11, gm_n633, gm_n283);
	nand (gm_n3510, in_21, gm_n85, gm_n56, gm_n3509, gm_n379);
	nand (gm_n3511, gm_n3510, gm_n3508, gm_n3506);
	nor (gm_n3512, in_14, gm_n78, in_9, gm_n2340, gm_n133);
	nand (gm_n3513, gm_n245, gm_n199, gm_n119, gm_n3512);
	nor (gm_n3514, gm_n148, in_14, in_10, gm_n259, gm_n207);
	nand (gm_n3515, gm_n806, gm_n146, in_18, gm_n3514);
	nor (gm_n3516, gm_n90, in_10, gm_n62, gm_n1406, gm_n362);
	nand (gm_n3517, gm_n436, gm_n146, gm_n119, gm_n3516);
	nand (gm_n3518, gm_n3517, gm_n3515, gm_n3513);
	nor (gm_n3519, gm_n3504, gm_n3427, gm_n3426, gm_n3518, gm_n3511);
	nand (gm_n3520, gm_n143, in_16, in_12, gm_n586, gm_n571);
	nor (gm_n3521, gm_n262, in_21, in_20, gm_n3520);
	nor (gm_n3522, gm_n276, gm_n190, gm_n59, gm_n860);
	and (gm_n3523, in_21, in_20, in_19, gm_n3522, gm_n379);
	nand (gm_n3524, gm_n123, in_13, in_9, gm_n2949);
	nor (gm_n3525, gm_n388, gm_n72, gm_n55, gm_n3524, gm_n662);
	nor (gm_n3526, gm_n3525, gm_n3523, gm_n3521);
	or (gm_n3527, in_14, in_10, in_9, gm_n657, gm_n92);
	nor (gm_n3528, gm_n824, gm_n89, gm_n119, gm_n3527);
	or (gm_n3529, gm_n152, in_16, gm_n59, gm_n2589, gm_n263);
	nor (gm_n3530, gm_n781, in_21, in_20, gm_n3529);
	nand (gm_n3531, gm_n79, gm_n73, in_12, gm_n678, gm_n303);
	nor (gm_n3532, gm_n58, gm_n72, in_20, gm_n3531);
	nor (gm_n3533, gm_n3532, gm_n3530, gm_n3528);
	nand (gm_n3534, gm_n3519, gm_n3424, gm_n3422, gm_n3533, gm_n3526);
	nor (gm_n3535, gm_n1295, in_13, gm_n62, gm_n344, gm_n461);
	nand (gm_n3536, gm_n104, gm_n72, in_17, gm_n3535, gm_n120);
	and (gm_n3537, gm_n233, in_16, gm_n59, gm_n1392, gm_n221);
	nand (gm_n3538, gm_n138, in_21, in_20, gm_n3537);
	nor (gm_n3539, gm_n105, gm_n76, gm_n62, gm_n442, gm_n298);
	nand (gm_n3540, gm_n373, gm_n72, in_17, gm_n3539);
	nand (gm_n3541, gm_n3540, gm_n3538, gm_n3536);
	and (gm_n3542, gm_n192, gm_n154, gm_n60, gm_n1135, gm_n448);
	nand (gm_n3543, in_21, gm_n85, in_19, gm_n3542);
	nor (gm_n3544, gm_n90, in_10, in_9, gm_n1406, gm_n369);
	nand (gm_n3545, gm_n367, gm_n166, gm_n119, gm_n3544);
	nor (gm_n3546, gm_n207, gm_n121, gm_n78, gm_n491, gm_n248);
	nand (gm_n3547, gm_n206, gm_n72, in_17, gm_n3546);
	nand (gm_n3548, gm_n3547, gm_n3545, gm_n3543);
	nor (gm_n3549, gm_n3534, gm_n3421, gm_n3420, gm_n3548, gm_n3541);
	or (gm_n3550, gm_n114, gm_n73, gm_n59, gm_n263, gm_n230);
	nor (gm_n3551, gm_n496, in_21, gm_n85, gm_n3550);
	or (gm_n3552, gm_n90, in_10, gm_n62, gm_n1824, gm_n467);
	nor (gm_n3553, gm_n841, gm_n824, in_18, gm_n3552);
	nand (gm_n3554, gm_n143, gm_n73, gm_n59, gm_n969, gm_n221);
	nor (gm_n3555, gm_n262, in_21, in_20, gm_n3554);
	nor (gm_n3556, gm_n3555, gm_n3553, gm_n3551);
	nand (gm_n3557, gm_n79, gm_n73, in_12, gm_n2497, gm_n303);
	nor (gm_n3558, gm_n58, in_21, in_20, gm_n3557);
	or (gm_n3559, gm_n99, in_14, in_10, gm_n467, gm_n370);
	nor (gm_n3560, gm_n531, gm_n212, gm_n119, gm_n3559);
	or (gm_n3561, gm_n609, gm_n76, in_9, gm_n1132, gm_n480);
	nor (gm_n3562, gm_n103, in_21, gm_n55, gm_n3561, gm_n121);
	nor (gm_n3563, gm_n3562, gm_n3560, gm_n3558);
	nand (gm_n3564, gm_n3549, gm_n3418, gm_n3416, gm_n3563, gm_n3556);
	nor (gm_n3565, gm_n227, gm_n73, in_12, gm_n835, gm_n213);
	nand (gm_n3566, gm_n138, in_21, in_20, gm_n3565);
	nor (gm_n3567, gm_n78, gm_n62, gm_n94, gm_n417, gm_n207);
	nand (gm_n3568, gm_n164, gm_n119, in_14, gm_n3567, gm_n166);
	nor (gm_n3569, gm_n442, gm_n76, gm_n62, gm_n988, gm_n502);
	nand (gm_n3570, gm_n405, gm_n72, gm_n55, gm_n3569, gm_n327);
	nand (gm_n3571, gm_n3570, gm_n3568, gm_n3566);
	nor (gm_n3572, gm_n344, in_13, in_9, gm_n480, gm_n345);
	nand (gm_n3573, gm_n595, in_21, in_17, gm_n3572, gm_n373);
	and (gm_n3574, gm_n484, in_15, gm_n63, gm_n756, gm_n755);
	nand (gm_n3575, in_21, gm_n85, gm_n56, gm_n3574, gm_n394);
	nor (gm_n3576, gm_n90, gm_n78, gm_n62, gm_n2008, gm_n133);
	nand (gm_n3577, gm_n245, gm_n146, gm_n119, gm_n3576);
	nand (gm_n3578, gm_n3577, gm_n3575, gm_n3573);
	nor (gm_n3579, gm_n3564, gm_n3415, gm_n3413, gm_n3578, gm_n3571);
	nand (gm_n3580, gm_n76, gm_n62, gm_n94, gm_n402, gm_n2719);
	nor (gm_n3581, gm_n441, in_21, in_17, gm_n3580, gm_n313);
	or (gm_n3582, gm_n609, gm_n76, in_9, gm_n345, gm_n431);
	nor (gm_n3583, gm_n103, in_21, in_17, gm_n3582, gm_n313);
	nand (gm_n3584, gm_n110, gm_n76, gm_n62, gm_n402, gm_n341);
	nor (gm_n3585, gm_n183, in_21, in_17, gm_n3584, gm_n375);
	nor (gm_n3586, gm_n3585, gm_n3583, gm_n3581);
	and (gm_n3587, gm_n1067, gm_n291, in_8);
	and (gm_n3588, gm_n713, gm_n78, gm_n62, gm_n3587);
	and (gm_n3589, gm_n405, gm_n72, in_17, gm_n3588, gm_n373);
	or (gm_n3590, gm_n358, gm_n76, gm_n62, gm_n481, gm_n596);
	nor (gm_n3591, gm_n183, in_21, in_17, gm_n3590, gm_n328);
	or (gm_n3592, gm_n274, gm_n193, gm_n60, gm_n632, gm_n485);
	nor (gm_n3593, gm_n72, gm_n85, in_19, gm_n3592);
	nor (gm_n3594, gm_n3593, gm_n3591, gm_n3589);
	nand (gm_n3595, gm_n3579, gm_n3411, gm_n3409, gm_n3594, gm_n3586);
	nor (gm_n3596, gm_n213, in_16, gm_n59, gm_n2060, gm_n319);
	nand (gm_n3597, gm_n697, in_21, gm_n85, gm_n3596);
	and (gm_n3598, gm_n90, gm_n78, gm_n62, gm_n1451, gm_n624);
	nand (gm_n3599, gm_n199, gm_n88, gm_n119, gm_n3598);
	nor (gm_n3600, gm_n297, gm_n73, in_12, gm_n1484, gm_n276);
	nand (gm_n3601, gm_n138, in_21, gm_n85, gm_n3600);
	nand (gm_n3602, gm_n3601, gm_n3599, gm_n3597);
	nor (gm_n3603, gm_n191, gm_n297, gm_n60, gm_n3382, gm_n760);
	nand (gm_n3604, gm_n72, gm_n85, in_19, gm_n3603);
	nor (gm_n3605, gm_n514, gm_n76, gm_n62, gm_n3402, gm_n184);
	nand (gm_n3606, gm_n102, gm_n72, in_17, gm_n3605);
	nor (gm_n3607, gm_n358, gm_n76, in_9, gm_n502, gm_n462);
	nand (gm_n3608, gm_n122, in_21, in_17, gm_n3607, gm_n311);
	nand (gm_n3609, gm_n3608, gm_n3606, gm_n3604);
	nor (gm_n3610, gm_n3595, gm_n3408, gm_n3406, gm_n3609, gm_n3602);
	nand (gm_n3611, gm_n126, gm_n76, in_9, gm_n341, gm_n185);
	nor (gm_n3612, gm_n620, gm_n72, in_17, gm_n3611, gm_n328);
	or (gm_n3613, gm_n115, gm_n73, in_12, gm_n1223, gm_n152);
	nor (gm_n3614, gm_n496, in_21, gm_n85, gm_n3613);
	nand (gm_n3615, gm_n484, gm_n60, in_11, gm_n714, gm_n1144);
	nor (gm_n3616, gm_n72, gm_n85, in_19, gm_n3615, gm_n447);
	nor (gm_n3617, gm_n3616, gm_n3614, gm_n3612);
	nand (gm_n3618, gm_n110, in_13, gm_n62, gm_n402, gm_n341);
	nor (gm_n3619, gm_n388, in_21, in_17, gm_n3618, gm_n375);
	nor (gm_n3620, gm_n312, gm_n72, gm_n55, gm_n1532);
	nand (gm_n3621, gm_n76, gm_n59, in_11, gm_n756, gm_n602);
	nor (gm_n3622, gm_n211, gm_n119, gm_n90, gm_n3621, gm_n246);
	nor (gm_n3623, gm_n3622, gm_n3620, gm_n3619);
	nand (gm_n3624, gm_n3610, gm_n3404, gm_n3401, gm_n3623, gm_n3617);
	nor (gm_n3625, gm_n572, gm_n215, gm_n977);
	and (gm_n3626, gm_n268, in_15, in_11, gm_n3625, gm_n545);
	nand (gm_n3627, gm_n72, gm_n85, gm_n56, gm_n3626);
	and (gm_n3628, gm_n600, gm_n170, in_14, gm_n1942);
	nand (gm_n3629, gm_n806, gm_n129, gm_n119, gm_n3628);
	nor (gm_n3630, gm_n430, in_13, gm_n62, gm_n442, gm_n345);
	nand (gm_n3631, gm_n255, gm_n72, in_17, gm_n3630, gm_n373);
	nand (gm_n3632, gm_n3631, gm_n3629, gm_n3627);
	nand (gm_n3633, gm_n93, in_6, gm_n97, gm_n426, gm_n94);
	nor (gm_n3634, gm_n263, in_16, gm_n59, gm_n3633, gm_n354);
	nand (gm_n3635, gm_n383, in_21, in_20, gm_n3634);
	nor (gm_n3636, gm_n514, gm_n76, gm_n62, gm_n345, gm_n667);
	nand (gm_n3637, gm_n523, in_21, in_17, gm_n3636, gm_n373);
	nand (gm_n3638, gm_n546, gm_n81, in_8);
	nor (gm_n3639, gm_n227, gm_n73, gm_n59, gm_n3638, gm_n155);
	nand (gm_n3640, gm_n138, in_21, gm_n85, gm_n3639);
	nand (gm_n3641, gm_n3640, gm_n3637, gm_n3635);
	nor (gm_n3642, gm_n3624, gm_n3399, gm_n3398, gm_n3641, gm_n3632);
	or (gm_n3643, gm_n442, gm_n76, gm_n62, gm_n1132, gm_n443);
	nor (gm_n3644, gm_n479, in_21, gm_n55, gm_n3643, gm_n375);
	nand (gm_n3645, gm_n90, in_10, gm_n62, gm_n626, gm_n600);
	nor (gm_n3646, gm_n212, gm_n130, in_18, gm_n3645);
	or (gm_n3647, gm_n442, gm_n76, in_9, gm_n988, gm_n463);
	nor (gm_n3648, gm_n312, gm_n72, in_17, gm_n3647, gm_n313);
	nor (gm_n3649, gm_n3648, gm_n3646, gm_n3644);
	or (gm_n3650, gm_n406, in_13, in_9, gm_n481, gm_n596);
	nor (gm_n3651, gm_n103, in_21, gm_n55, gm_n3650, gm_n375);
	or (gm_n3652, in_14, gm_n78, gm_n62, gm_n2474, gm_n133);
	nor (gm_n3653, gm_n246, gm_n87, gm_n119, gm_n3652);
	or (gm_n3654, gm_n514, in_13, in_9, gm_n481, gm_n667);
	nor (gm_n3655, gm_n312, gm_n72, in_17, gm_n3654, gm_n662);
	nor (gm_n3656, gm_n3655, gm_n3653, gm_n3651);
	nand (gm_n3657, gm_n3642, gm_n3396, gm_n3394, gm_n3656, gm_n3649);
	nand (gm_n3658, in_21, in_20, in_19, gm_n613, gm_n448);
	nand (gm_n3659, gm_n348, gm_n806, gm_n119, gm_n1833);
	nand (gm_n3660, in_7, gm_n124, gm_n97, gm_n80, in_8);
	nor (gm_n3661, gm_n152, in_16, in_12, gm_n3660, gm_n274);
	nand (gm_n3662, gm_n495, in_21, gm_n85, gm_n3661);
	nand (gm_n3663, gm_n3662, gm_n3659, gm_n3658);
	nor (gm_n3664, gm_n358, gm_n76, gm_n62, gm_n988, gm_n502);
	nand (gm_n3665, gm_n104, gm_n72, in_17, gm_n3664, gm_n327);
	nor (gm_n3666, in_14, in_10, in_9, gm_n2421, gm_n807);
	nand (gm_n3667, gm_n245, gm_n164, gm_n119, gm_n3666);
	nor (gm_n3668, gm_n227, gm_n73, in_12, gm_n180, gm_n155);
	nand (gm_n3669, gm_n57, gm_n72, gm_n85, gm_n3668);
	nand (gm_n3670, gm_n3669, gm_n3667, gm_n3665);
	nor (gm_n3671, gm_n3657, gm_n3392, gm_n3390, gm_n3670, gm_n3663);
	nand (gm_n3672, gm_n110, gm_n76, in_9, gm_n341, gm_n185);
	nor (gm_n3673, gm_n183, gm_n72, gm_n55, gm_n3672, gm_n662);
	nand (gm_n3674, gm_n2719, in_15, gm_n63, gm_n1398, gm_n171);
	nor (gm_n3675, gm_n72, gm_n85, gm_n56, gm_n3674, gm_n191);
	nand (gm_n3676, gm_n245, gm_n600, gm_n90, gm_n1120, gm_n602);
	nor (gm_n3677, gm_n3676, gm_n165, in_18);
	nor (gm_n3678, gm_n3677, gm_n3675, gm_n3673);
	and (gm_n3679, gm_n93, in_6, in_5, gm_n426, gm_n94);
	nand (gm_n3680, gm_n214, in_16, in_12, gm_n3679, gm_n275);
	nor (gm_n3681, gm_n781, gm_n72, in_20, gm_n3680);
	or (gm_n3682, gm_n257, gm_n76, in_9, gm_n1583, gm_n463);
	nor (gm_n3683, gm_n103, in_21, in_17, gm_n3682, gm_n184);
	nand (gm_n3684, in_13, gm_n62, in_8, gm_n580, gm_n402);
	nor (gm_n3685, gm_n388, gm_n72, gm_n55, gm_n3684, gm_n313);
	nor (gm_n3686, gm_n3685, gm_n3683, gm_n3681);
	nand (gm_n3687, gm_n3671, gm_n3388, gm_n3386, gm_n3686, gm_n3678);
	and (gm_n3688, gm_n214, gm_n61, gm_n59, gm_n734);
	nand (gm_n3689, gm_n72, in_20, in_19, gm_n3688, gm_n268);
	nor (gm_n3690, gm_n667, in_13, gm_n62, gm_n1132, gm_n480);
	nand (gm_n3691, gm_n102, in_21, gm_n55, gm_n3690, gm_n339);
	nor (gm_n3692, gm_n467, in_14, in_10, gm_n589, gm_n491);
	nand (gm_n3693, gm_n348, gm_n200, gm_n119, gm_n3692);
	nand (gm_n3694, gm_n3693, gm_n3691, gm_n3689);
	nor (gm_n3695, gm_n1331, gm_n213, in_15, gm_n2589, gm_n643);
	nand (gm_n3696, in_21, gm_n85, in_19, gm_n3695);
	nor (gm_n3697, gm_n213, in_16, in_12, gm_n2080, gm_n354);
	nand (gm_n3698, gm_n57, gm_n72, in_20, gm_n3697);
	and (gm_n3699, gm_n221, gm_n73, gm_n59, gm_n1456, gm_n264);
	nand (gm_n3700, gm_n113, in_21, gm_n85, gm_n3699);
	nand (gm_n3701, gm_n3700, gm_n3698, gm_n3696);
	nor (gm_n3702, gm_n3687, gm_n3384, gm_n3381, gm_n3701, gm_n3694);
	or (gm_n3703, gm_n609, gm_n76, gm_n62, gm_n1132, gm_n406);
	nor (gm_n3704, gm_n183, gm_n72, in_17, gm_n3703, gm_n313);
	or (gm_n3705, gm_n99, in_14, in_10, gm_n491, gm_n362);
	nor (gm_n3706, gm_n368, gm_n167, in_18, gm_n3705);
	nor (gm_n3707, gm_n183, gm_n72, in_17, gm_n2449, gm_n184);
	nor (gm_n3708, gm_n3707, gm_n3706, gm_n3704);
	nand (gm_n3709, gm_n61, in_16, gm_n59, gm_n1012, gm_n264);
	nor (gm_n3710, gm_n219, gm_n72, in_20, gm_n3709);
	or (gm_n3711, gm_n514, in_13, gm_n62, gm_n1583, gm_n502);
	nor (gm_n3712, gm_n184, gm_n72, in_17, gm_n3711, gm_n312);
	or (gm_n3713, gm_n148, in_14, gm_n78, gm_n775, gm_n467);
	nor (gm_n3714, gm_n841, gm_n87, in_18, gm_n3713);
	nor (gm_n3715, gm_n3714, gm_n3712, gm_n3710);
	nand (gm_n3716, gm_n3702, gm_n3379, gm_n3377, gm_n3715, gm_n3708);
	nor (gm_n3717, gm_n147, gm_n67, gm_n90, gm_n2017, gm_n572);
	nand (gm_n3718, gm_n348, gm_n88, gm_n119, gm_n3717);
	nor (gm_n3719, gm_n257, in_13, gm_n62, gm_n597, gm_n596);
	nand (gm_n3720, gm_n255, gm_n72, gm_n55, gm_n3719, gm_n373);
	or (gm_n3721, gm_n93, in_6, in_5, gm_n215, in_8);
	nor (gm_n3722, gm_n227, gm_n73, in_12, gm_n3721, gm_n263);
	nand (gm_n3723, gm_n57, in_21, in_20, gm_n3722);
	nand (gm_n3724, gm_n3723, gm_n3720, gm_n3718);
	nor (out_8, gm_n3716, gm_n3375, gm_n3373, gm_n3724);
	or (gm_n3726, gm_n442, in_13, in_9, gm_n621, gm_n443);
	nor (gm_n3727, gm_n105, gm_n72, in_17, gm_n3726, gm_n183);
	nor (gm_n3728, gm_n609, gm_n76, in_9, gm_n1583, gm_n461);
	nand (gm_n3729, gm_n523, gm_n72, gm_n55, gm_n3728, gm_n311);
	nor (gm_n3730, gm_n95, in_14, in_10, gm_n807, gm_n259);
	nand (gm_n3731, gm_n199, gm_n166, gm_n119, gm_n3730);
	nand (gm_n3732, in_14, gm_n78, gm_n62, gm_n803, gm_n334);
	nor (gm_n3733, gm_n824, gm_n89, gm_n119, gm_n3732);
	nor (gm_n3734, gm_n293, gm_n263, gm_n60, gm_n1751, gm_n760);
	nand (gm_n3735, gm_n72, in_20, gm_n56, gm_n3734);
	nor (gm_n3736, gm_n274, gm_n74, in_15, gm_n821, gm_n290);
	nand (gm_n3737, in_21, in_20, in_19, gm_n3736);
	nand (gm_n3738, in_10, gm_n62, in_8, gm_n756, gm_n624);
	nor (gm_n3739, gm_n167, gm_n119, gm_n90, gm_n3738, gm_n368);
	or (gm_n3740, gm_n430, gm_n76, in_9, gm_n481, gm_n406);
	nor (gm_n3741, gm_n312, gm_n72, gm_n55, gm_n3740, gm_n328);
	nor (gm_n3742, gm_n213, in_16, gm_n59, gm_n1664, gm_n319);
	nand (gm_n3743, gm_n57, gm_n72, in_20, gm_n3742);
	nor (gm_n3744, gm_n194, gm_n92, in_14, gm_n240, gm_n141);
	nand (gm_n3745, gm_n436, gm_n146, in_18, gm_n3744);
	or (gm_n3746, gm_n514, in_13, in_9, gm_n1132, gm_n667);
	nor (gm_n3747, gm_n183, in_21, gm_n55, gm_n3746, gm_n256);
	or (gm_n3748, gm_n431, gm_n99, in_13, gm_n370, gm_n662);
	nor (gm_n3749, gm_n479, in_21, in_17, gm_n3748);
	nor (gm_n3750, gm_n78, gm_n62, gm_n94, gm_n417, gm_n362);
	nand (gm_n3751, gm_n200, in_18, gm_n90, gm_n3750, gm_n243);
	nor (gm_n3752, gm_n269, gm_n56, in_15, gm_n2927, gm_n290);
	nand (gm_n3753, gm_n3752, gm_n72, gm_n85);
	or (gm_n3754, gm_n671, gm_n68);
	nor (gm_n3755, gm_n290, gm_n60, gm_n63, gm_n3754, gm_n605);
	nand (gm_n3756, in_21, in_20, in_19, gm_n3755, gm_n75);
	and (gm_n3757, gm_n154, gm_n73, in_12, gm_n2497, gm_n949);
	nand (gm_n3758, gm_n113, in_21, in_20, gm_n3757);
	nand (gm_n3759, gm_n3753, gm_n3751, t_4, gm_n3758, gm_n3756);
	and (gm_n3760, gm_n79, gm_n73, gm_n59, gm_n2547, gm_n733);
	nand (gm_n3761, gm_n138, gm_n72, gm_n85, gm_n3760);
	nor (gm_n3762, gm_n866, in_13, gm_n62, gm_n463, gm_n406);
	nand (gm_n3763, gm_n102, gm_n72, gm_n55, gm_n3762, gm_n595);
	nor (gm_n3764, gm_n514, gm_n76, in_9, gm_n481, gm_n430);
	nand (gm_n3765, gm_n120, gm_n72, in_17, gm_n3764, gm_n339);
	nand (gm_n3766, gm_n3765, gm_n3763, gm_n3761);
	nor (gm_n3767, gm_n90, in_10, gm_n62, gm_n3660, gm_n92);
	nand (gm_n3768, gm_n348, gm_n323, gm_n119, gm_n3767);
	nand (gm_n3769, gm_n304, gm_n59, gm_n94, gm_n546, gm_n264);
	nor (gm_n3770, gm_n139, in_20, gm_n73, gm_n3769, gm_n319);
	nand (gm_n3771, gm_n3770, in_21);
	nor (gm_n3772, gm_n430, in_13, gm_n62, gm_n359, gm_n406);
	nand (gm_n3773, gm_n104, gm_n72, gm_n55, gm_n3772, gm_n254);
	nand (gm_n3774, gm_n3773, gm_n3771, gm_n3768);
	nor (gm_n3775, gm_n3759, gm_n3749, gm_n3747, gm_n3774, gm_n3766);
	nor (gm_n3776, gm_n620, in_21, in_17, gm_n584, gm_n375);
	or (gm_n3777, gm_n158, gm_n74, in_15, gm_n515, gm_n290);
	nor (gm_n3778, gm_n72, gm_n85, in_19, gm_n3777);
	nand (gm_n3779, gm_n316, gm_n76, in_9, gm_n1049, gm_n402);
	nor (gm_n3780, gm_n441, gm_n72, gm_n55, gm_n3779, gm_n184);
	nor (gm_n3781, gm_n3780, gm_n3778, gm_n3776);
	or (gm_n3782, gm_n286, gm_n90, gm_n78, gm_n491, gm_n369);
	nor (gm_n3783, gm_n167, gm_n87, gm_n119, gm_n3782);
	or (gm_n3784, gm_n257, in_13, gm_n62, gm_n1132, gm_n344);
	nor (gm_n3785, gm_n105, gm_n72, in_17, gm_n3784, gm_n183);
	not (gm_n3786, gm_n722);
	or (gm_n3787, gm_n92, gm_n90, gm_n78, gm_n3786, gm_n287);
	nor (gm_n3788, gm_n824, gm_n89, in_18, gm_n3787);
	nor (gm_n3789, gm_n3788, gm_n3785, gm_n3783);
	nand (gm_n3790, gm_n3775, gm_n3745, gm_n3743, gm_n3789, gm_n3781);
	nor (gm_n3791, gm_n313, gm_n76, gm_n62, gm_n2340, gm_n480);
	nand (gm_n3792, gm_n120, gm_n72, gm_n55, gm_n3791);
	nor (gm_n3793, in_14, gm_n78, in_9, gm_n2008, gm_n807);
	nand (gm_n3794, gm_n348, gm_n200, in_18, gm_n3793);
	nor (gm_n3795, gm_n431, in_13, gm_n62, gm_n345, gm_n344);
	nand (gm_n3796, gm_n311, in_21, in_17, gm_n3795, gm_n595);
	nand (gm_n3797, gm_n3796, gm_n3794, gm_n3792);
	nand (gm_n3798, gm_n104, in_21, gm_n55, gm_n2206, gm_n254);
	nor (gm_n3799, gm_n90, in_10, gm_n62, gm_n1906, gm_n92);
	nand (gm_n3800, gm_n245, gm_n243, gm_n119, gm_n3799);
	nand (gm_n3801, gm_n323, gm_n199, in_18, gm_n1055);
	nand (gm_n3802, gm_n3801, gm_n3800, gm_n3798);
	nor (gm_n3803, gm_n3790, gm_n3741, gm_n3739, gm_n3802, gm_n3797);
	or (gm_n3804, gm_n207, in_14, in_10, gm_n526, gm_n287);
	nor (gm_n3805, gm_n1989, gm_n130, gm_n119, gm_n3804);
	nand (gm_n3806, gm_n107, gm_n76, gm_n62, gm_n788, gm_n316);
	nor (gm_n3807, gm_n312, gm_n72, gm_n55, gm_n3806, gm_n328);
	and (gm_n3808, in_21, in_20, in_19, gm_n735, gm_n394);
	nor (gm_n3809, gm_n3808, gm_n3807, gm_n3805);
	or (gm_n3810, gm_n155, gm_n73, gm_n59, gm_n2357, gm_n354);
	nor (gm_n3811, gm_n58, gm_n72, in_20, gm_n3810);
	nor (gm_n3812, gm_n467, gm_n78, gm_n62, gm_n1689);
	and (gm_n3813, gm_n122, gm_n72, gm_n55, gm_n3812, gm_n174);
	or (gm_n3814, gm_n667, in_13, gm_n62, gm_n480, gm_n345);
	nor (gm_n3815, gm_n388, gm_n72, in_17, gm_n3814, gm_n328);
	nor (gm_n3816, gm_n3815, gm_n3813, gm_n3811);
	nand (gm_n3817, gm_n3803, gm_n3737, gm_n3735, gm_n3816, gm_n3809);
	and (gm_n3818, gm_n426, gm_n81);
	nand (gm_n3819, gm_n192, in_15, in_11, gm_n3818, gm_n1942);
	nor (gm_n3820, in_21, in_20, in_19, gm_n3819, gm_n485);
	or (gm_n3821, gm_n271, in_15, gm_n63, gm_n770, gm_n633);
	nor (gm_n3822, gm_n72, in_20, in_19, gm_n3821, gm_n393);
	or (gm_n3823, gm_n406, gm_n76, gm_n62, gm_n621, gm_n596);
	nor (gm_n3824, gm_n121, gm_n72, gm_n55, gm_n3823, gm_n312);
	nor (gm_n3825, gm_n3820, gm_n3817, gm_n3733, gm_n3824, gm_n3822);
	nand (gm_n3826, gm_n143, gm_n75, gm_n60, gm_n2276, gm_n545);
	nor (gm_n3827, gm_n72, in_20, gm_n56, gm_n3826);
	or (gm_n3828, gm_n227, gm_n73, in_12, gm_n849, gm_n213);
	nor (gm_n3829, gm_n912, in_21, gm_n85, gm_n3828);
	or (gm_n3830, gm_n193, gm_n155, in_15, gm_n648, gm_n447);
	nor (gm_n3831, gm_n72, gm_n85, gm_n56, gm_n3830);
	nor (gm_n3832, gm_n3831, gm_n3829, gm_n3827);
	nand (gm_n3833, gm_n394, gm_n79, in_15, gm_n1398, gm_n423);
	nor (gm_n3834, in_21, in_20, in_19, gm_n3833);
	or (gm_n3835, gm_n227, gm_n73, in_12, gm_n1542, gm_n115);
	nor (gm_n3836, gm_n58, gm_n72, in_20, gm_n3835);
	or (gm_n3837, gm_n90, gm_n78, gm_n62, gm_n654, gm_n92);
	nor (gm_n3838, gm_n246, gm_n87, gm_n119, gm_n3837);
	nor (gm_n3839, gm_n3838, gm_n3836, gm_n3834);
	nand (gm_n3840, gm_n3825, gm_n3731, gm_n3729, gm_n3839, gm_n3832);
	nor (gm_n3841, in_14, in_10, in_9, gm_n657, gm_n467);
	nand (gm_n3842, gm_n806, gm_n199, in_18, gm_n3841);
	nand (gm_n3843, gm_n199, gm_n88, in_18, gm_n2351);
	and (gm_n3844, gm_n125, gm_n76, in_9, gm_n340, gm_n126);
	nand (gm_n3845, gm_n373, gm_n72, gm_n55, gm_n3844, gm_n1076);
	nand (gm_n3846, gm_n3845, gm_n3843, gm_n3842);
	nand (gm_n3847, gm_n61, gm_n73, in_12, gm_n998, gm_n264);
	nor (gm_n3848, gm_n384, in_21, in_20, gm_n3847);
	nor (out_9, gm_n3846, gm_n3840, gm_n3727, gm_n3848);
	or (gm_n3850, gm_n362, gm_n90, gm_n78, gm_n438, gm_n389);
	nor (gm_n3851, gm_n1989, gm_n211, in_18, gm_n3850);
	and (gm_n3852, gm_n449, gm_n60, in_11, gm_n1120, gm_n1928);
	nand (gm_n3853, in_21, gm_n85, in_19, gm_n3852, gm_n394);
	nand (gm_n3854, gm_n76, in_9, gm_n94, gm_n2074, gm_n185);
	nor (gm_n3855, gm_n388, gm_n72, in_17, gm_n3854, gm_n328);
	and (gm_n3856, gm_n106, in_13, gm_n62, gm_n187, gm_n186);
	and (gm_n3857, gm_n122, gm_n72, in_17, gm_n3856, gm_n327);
	nor (gm_n3858, gm_n344, in_13, in_9, gm_n442, gm_n432);
	nand (gm_n3859, gm_n327, gm_n72, gm_n55, gm_n3858, gm_n595);
	nor (gm_n3860, in_10, gm_n62, gm_n94, gm_n467, gm_n417);
	nand (gm_n3861, gm_n131, in_18, gm_n90, gm_n3860, gm_n348);
	nand (gm_n3862, gm_n154, in_16, gm_n59, gm_n586, gm_n303);
	nor (gm_n3863, gm_n781, in_21, in_20, gm_n3862);
	nand (gm_n3864, in_14, gm_n78, in_9, gm_n1011, gm_n446);
	nor (gm_n3865, gm_n531, gm_n212, in_18, gm_n3864);
	nor (gm_n3866, gm_n297, in_16, in_12, gm_n520, gm_n354);
	nand (gm_n3867, gm_n383, in_21, in_20, gm_n3866);
	nor (gm_n3868, gm_n190, gm_n73, in_12, gm_n3638, gm_n319);
	nand (gm_n3869, gm_n138, in_21, gm_n85, gm_n3868);
	nand (gm_n3870, gm_n222, in_16, gm_n59, gm_n3041, gm_n303);
	nor (gm_n3871, gm_n58, gm_n72, gm_n85, gm_n3870);
	nand (gm_n3872, gm_n122, gm_n76, in_9, gm_n1611, gm_n579);
	nor (gm_n3873, gm_n374, gm_n72, in_17, gm_n3872);
	nor (gm_n3874, gm_n290, gm_n60, gm_n63, gm_n770, gm_n605);
	nand (gm_n3875, in_21, gm_n85, in_19, gm_n3874, gm_n75);
	nor (gm_n3876, gm_n572, gm_n141, in_8);
	nand (gm_n3877, gm_n154, in_16, gm_n59, gm_n3876, gm_n221);
	or (gm_n3878, gm_n781, gm_n72, in_20, gm_n3877);
	and (gm_n3879, gm_n102, in_21, in_17, gm_n2663, gm_n255);
	or (gm_n3880, gm_n155, gm_n73, in_12, gm_n3315, gm_n319);
	nor (gm_n3881, gm_n139, in_21, in_20, gm_n3880);
	and (gm_n3882, gm_n233, in_16, gm_n59, gm_n275, gm_n235);
	nand (gm_n3883, gm_n138, gm_n72, gm_n85, gm_n3882);
	nor (gm_n3884, gm_n193, gm_n190, in_15, gm_n2357, gm_n269);
	nand (gm_n3885, gm_n72, gm_n85, gm_n56, gm_n3884);
	nor (gm_n3886, gm_n93, in_6, in_5, gm_n238, gm_n94);
	nand (gm_n3887, gm_n192, gm_n75, in_15, gm_n3886, gm_n214);
	nor (gm_n3888, in_21, gm_n85, gm_n56, gm_n3887);
	or (gm_n3889, gm_n191, gm_n155, gm_n60, gm_n2008, gm_n193);
	nor (gm_n3890, in_21, gm_n85, gm_n56, gm_n3889);
	nor (gm_n3891, gm_n430, in_13, gm_n62, gm_n743, gm_n480);
	nand (gm_n3892, gm_n120, gm_n72, gm_n55, gm_n3891, gm_n339);
	nor (gm_n3893, gm_n447, gm_n213, in_15, gm_n1319, gm_n633);
	nand (gm_n3894, gm_n72, in_20, in_19, gm_n3893);
	nor (gm_n3895, gm_n389, gm_n207, in_10, gm_n491);
	and (gm_n3896, gm_n104, gm_n72, in_17, gm_n3895, gm_n327);
	and (gm_n3897, gm_n334, gm_n171, gm_n81, gm_n426);
	and (gm_n3898, gm_n206, in_21, in_17, gm_n3897, gm_n1076);
	nor (gm_n3899, gm_n293, gm_n155, gm_n60, gm_n2008, gm_n643);
	nand (gm_n3900, gm_n72, in_20, gm_n56, gm_n3899);
	nor (gm_n3901, gm_n158, gm_n74, in_15, gm_n760, gm_n116);
	nand (gm_n3902, gm_n72, in_20, gm_n56, gm_n3901);
	or (gm_n3903, gm_n442, in_13, gm_n62, gm_n621, gm_n502);
	nor (gm_n3904, gm_n103, gm_n72, in_17, gm_n3903, gm_n105);
	nand (gm_n3905, gm_n222, gm_n379, in_15, gm_n2172, gm_n449);
	nor (gm_n3906, gm_n72, gm_n85, gm_n56, gm_n3905);
	nor (gm_n3907, gm_n207, gm_n167, in_14, gm_n981, gm_n271);
	nand (gm_n3908, gm_n3907, gm_n199, gm_n119);
	nor (gm_n3909, in_14, gm_n78, in_9, gm_n1006, gm_n467);
	nand (gm_n3910, gm_n806, gm_n129, in_18, gm_n3909);
	or (gm_n3911, gm_n977, gm_n60, gm_n63, gm_n770, gm_n193);
	nor (gm_n3912, in_21, gm_n85, in_19, gm_n3911, gm_n191);
	or (gm_n3913, gm_n207, gm_n167, gm_n90, gm_n770, gm_n240);
	nor (gm_n3914, gm_n3913, gm_n211, gm_n119);
	nor (gm_n3915, gm_n274, in_16, in_12, gm_n354, gm_n251);
	nand (gm_n3916, gm_n296, gm_n72, gm_n85, gm_n3915);
	and (gm_n3917, gm_n316, in_13, in_9, gm_n402, gm_n341);
	nand (gm_n3918, gm_n523, in_21, gm_n55, gm_n3917, gm_n327);
	nand (gm_n3919, gm_n143, in_16, gm_n59, gm_n3041, gm_n275);
	nor (gm_n3920, gm_n384, gm_n72, gm_n85, gm_n3919);
	nand (gm_n3921, gm_n154, in_16, gm_n59, gm_n571, gm_n446);
	nor (gm_n3922, gm_n781, gm_n72, in_20, gm_n3921);
	nor (gm_n3923, gm_n158, in_16, in_12, gm_n815, gm_n152);
	nand (gm_n3924, gm_n113, gm_n72, in_20, gm_n3923);
	nor (gm_n3925, gm_n431, gm_n76, gm_n62, gm_n503, gm_n502);
	nand (gm_n3926, gm_n122, in_21, gm_n55, gm_n3925, gm_n373);
	nor (gm_n3927, gm_n596, in_13, gm_n62, gm_n621, gm_n480);
	nand (gm_n3928, gm_n102, gm_n72, in_17, gm_n3927, gm_n405);
	nand (gm_n3929, gm_n519, gm_n291, gm_n94);
	nor (gm_n3930, gm_n227, gm_n73, in_12, gm_n3929, gm_n213);
	nand (gm_n3931, gm_n138, in_21, in_20, gm_n3930);
	nor (gm_n3932, in_14, in_10, gm_n62, gm_n2697, gm_n807);
	nand (gm_n3933, gm_n200, gm_n164, in_18, gm_n3932);
	nand (gm_n3934, gm_n3928, gm_n3926, gm_n3924, gm_n3933, gm_n3931);
	nor (gm_n3935, gm_n297, gm_n73, in_12, gm_n1689, gm_n319);
	nand (gm_n3936, gm_n138, in_21, in_20, gm_n3935);
	and (gm_n3937, gm_n233, in_16, gm_n59, gm_n962, gm_n275);
	nand (gm_n3938, gm_n57, gm_n72, gm_n85, gm_n3937);
	nor (gm_n3939, gm_n114, in_16, in_12, gm_n278, gm_n213);
	nand (gm_n3940, gm_n296, gm_n72, gm_n85, gm_n3939);
	nand (gm_n3941, gm_n3940, gm_n3938, gm_n3936);
	nor (gm_n3942, gm_n227, in_16, gm_n59, gm_n552, gm_n297);
	nand (gm_n3943, gm_n179, in_21, in_20, gm_n3942);
	nor (gm_n3944, gm_n133, in_14, in_10, gm_n526, gm_n370);
	nand (gm_n3945, gm_n200, gm_n146, in_18, gm_n3944);
	and (gm_n3946, gm_n107, in_10, gm_n62, gm_n600, gm_n110);
	nand (gm_n3947, gm_n129, in_18, gm_n90, gm_n3946, gm_n131);
	nand (gm_n3948, gm_n3947, gm_n3945, gm_n3943);
	nor (gm_n3949, gm_n3934, gm_n3922, gm_n3920, gm_n3948, gm_n3941);
	nand (gm_n3950, gm_n154, in_16, in_12, gm_n2276, gm_n221);
	nor (gm_n3951, gm_n219, in_21, gm_n85, gm_n3950);
	or (gm_n3952, gm_n358, gm_n76, gm_n62, gm_n345, gm_n596);
	nor (gm_n3953, gm_n121, gm_n72, in_17, gm_n3952, gm_n620);
	nand (gm_n3954, gm_n187, in_13, in_9, gm_n341, gm_n579);
	nor (gm_n3955, gm_n620, in_21, gm_n55, gm_n3954, gm_n375);
	nor (gm_n3956, gm_n3955, gm_n3953, gm_n3951);
	nand (gm_n3957, gm_n143, in_13, gm_n59, gm_n778);
	nor (gm_n3958, gm_n441, in_21, gm_n55, gm_n3957, gm_n662);
	nand (gm_n3959, gm_n523, in_13, in_9, gm_n2346, gm_n185);
	nor (gm_n3960, gm_n479, in_21, gm_n55, gm_n3959);
	nand (gm_n3961, gm_n76, in_9, gm_n94, gm_n576, gm_n579);
	nor (gm_n3962, gm_n312, gm_n72, in_17, gm_n3961, gm_n328);
	nor (gm_n3963, gm_n3962, gm_n3960, gm_n3958);
	nand (gm_n3964, gm_n3949, gm_n3918, gm_n3916, gm_n3963, gm_n3956);
	nor (gm_n3965, gm_n74, in_19, gm_n60, gm_n2526, gm_n159);
	nand (gm_n3966, gm_n3965, gm_n72, gm_n85);
	and (gm_n3967, gm_n61, in_16, in_12, gm_n1071, gm_n154);
	nand (gm_n3968, gm_n113, gm_n72, in_20, gm_n3967);
	nor (gm_n3969, gm_n159, gm_n60, gm_n63, gm_n761, gm_n283);
	nand (gm_n3970, in_21, gm_n85, in_19, gm_n3969, gm_n448);
	nand (gm_n3971, gm_n3970, gm_n3968, gm_n3966);
	and (gm_n3972, gm_n214, gm_n73, in_12, gm_n636, gm_n303);
	nand (gm_n3973, gm_n383, in_21, gm_n85, gm_n3972);
	nor (gm_n3974, gm_n818, in_13, gm_n62, gm_n463, gm_n431);
	nand (gm_n3975, gm_n104, gm_n72, in_17, gm_n3974, gm_n254);
	nor (gm_n3976, gm_n190, gm_n73, in_12, gm_n2221, gm_n385);
	nand (gm_n3977, gm_n138, gm_n72, gm_n85, gm_n3976);
	nand (gm_n3978, gm_n3977, gm_n3975, gm_n3973);
	nor (gm_n3979, gm_n3964, gm_n3914, gm_n3912, gm_n3978, gm_n3971);
	nand (gm_n3980, gm_n233, gm_n73, gm_n59, gm_n3454, gm_n221);
	nor (gm_n3981, gm_n384, gm_n72, gm_n85, gm_n3980);
	nor (gm_n3982, gm_n531, gm_n132, in_18, gm_n439);
	or (gm_n3983, gm_n431, in_13, in_9, gm_n1132, gm_n344);
	nor (gm_n3984, gm_n105, gm_n72, in_17, gm_n3983, gm_n479);
	nor (gm_n3985, gm_n3984, gm_n3982, gm_n3981);
	nand (gm_n3986, gm_n233, gm_n73, gm_n59, gm_n936, gm_n221);
	nor (gm_n3987, gm_n384, gm_n72, gm_n85, gm_n3986);
	or (gm_n3988, gm_n159, in_15, in_11, gm_n761, gm_n605);
	nor (gm_n3989, in_21, gm_n85, in_19, gm_n3988, gm_n191);
	nand (gm_n3990, gm_n79, in_16, in_12, gm_n1451, gm_n303);
	nor (gm_n3991, gm_n58, gm_n72, gm_n85, gm_n3990);
	nor (gm_n3992, gm_n3991, gm_n3989, gm_n3987);
	nand (gm_n3993, gm_n3979, gm_n3910, gm_n3908, gm_n3992, gm_n3985);
	nor (gm_n3994, gm_n190, in_16, gm_n59, gm_n1173, gm_n385);
	nand (gm_n3995, gm_n138, in_21, gm_n85, gm_n3994);
	nor (gm_n3996, gm_n430, in_13, gm_n62, gm_n621, gm_n431);
	nand (gm_n3997, gm_n120, in_21, gm_n55, gm_n3996, gm_n122);
	nor (gm_n3998, gm_n430, in_13, in_9, gm_n432, gm_n406);
	nand (gm_n3999, gm_n405, in_21, gm_n55, gm_n3998, gm_n327);
	nand (gm_n4000, gm_n3999, gm_n3997, gm_n3995);
	nor (gm_n4001, gm_n358, in_13, in_9, gm_n988, gm_n502);
	nand (gm_n4002, gm_n523, gm_n72, in_17, gm_n4001, gm_n373);
	and (gm_n4003, gm_n334, in_14, gm_n78, gm_n829, gm_n721);
	nand (gm_n4004, gm_n243, gm_n166, gm_n119, gm_n4003);
	nor (gm_n4005, gm_n430, in_13, gm_n62, gm_n743, gm_n406);
	nand (gm_n4006, gm_n104, gm_n72, gm_n55, gm_n4005, gm_n120);
	nand (gm_n4007, gm_n4006, gm_n4004, gm_n4002);
	nor (gm_n4008, gm_n3993, gm_n3906, gm_n3904, gm_n4007, gm_n4000);
	or (gm_n4009, gm_n609, in_13, gm_n62, gm_n1132, gm_n257);
	nor (gm_n4010, gm_n103, in_21, in_17, gm_n4009, gm_n256);
	and (gm_n4011, in_7, in_6, in_5, gm_n134, gm_n94);
	nand (gm_n4012, gm_n90, gm_n78, gm_n62, gm_n4011, gm_n91);
	nor (gm_n4013, gm_n368, gm_n167, in_18, gm_n4012);
	nand (gm_n4014, gm_n170, in_15, in_11, gm_n869, gm_n602);
	nor (gm_n4015, in_21, in_20, gm_n56, gm_n4014, gm_n393);
	nor (gm_n4016, gm_n4015, gm_n4013, gm_n4010);
	or (gm_n4017, gm_n461, gm_n76, in_9, gm_n481, gm_n463);
	nor (gm_n4018, gm_n441, in_21, in_17, gm_n4017, gm_n662);
	nand (gm_n4019, gm_n392, gm_n233, gm_n60, gm_n2860, gm_n268);
	nor (gm_n4020, in_21, in_20, in_19, gm_n4019);
	or (gm_n4021, gm_n95, gm_n90, in_10, gm_n526, gm_n807);
	nor (gm_n4022, gm_n244, gm_n212, gm_n119, gm_n4021);
	nor (gm_n4023, gm_n4022, gm_n4020, gm_n4018);
	nand (gm_n4024, gm_n4008, gm_n3902, gm_n3900, gm_n4023, gm_n4016);
	nor (gm_n4025, gm_n362, gm_n283, in_14, gm_n842);
	nand (gm_n4026, gm_n323, gm_n164, in_18, gm_n4025);
	nor (gm_n4027, gm_n190, in_16, in_12, gm_n468, gm_n276);
	nand (gm_n4028, gm_n57, in_21, in_20, gm_n4027);
	and (gm_n4029, gm_n143, in_16, in_12, gm_n875, gm_n733);
	nand (gm_n4030, gm_n138, gm_n72, gm_n85, gm_n4029);
	nand (gm_n4031, gm_n4030, gm_n4028, gm_n4026);
	nor (gm_n4032, gm_n263, gm_n191, gm_n60, gm_n1170, gm_n290);
	nand (gm_n4033, gm_n72, in_20, gm_n56, gm_n4032);
	and (gm_n4034, gm_n555, in_15, gm_n63, gm_n1398, gm_n556);
	nand (gm_n4035, in_21, gm_n85, gm_n56, gm_n4034, gm_n486);
	nor (gm_n4036, gm_n406, gm_n76, in_9, gm_n502, gm_n359);
	nand (gm_n4037, gm_n122, in_21, in_17, gm_n4036, gm_n254);
	nand (gm_n4038, gm_n4037, gm_n4035, gm_n4033);
	nor (gm_n4039, gm_n4024, gm_n3898, gm_n3896, gm_n4038, gm_n4031);
	or (gm_n4040, gm_n461, gm_n76, gm_n62, gm_n2077, gm_n375);
	nor (gm_n4041, gm_n183, in_21, gm_n55, gm_n4040);
	or (gm_n4042, gm_n276, gm_n297, in_12, gm_n447, gm_n320);
	nor (gm_n4043, gm_n72, gm_n85, gm_n56, gm_n4042);
	nand (gm_n4044, gm_n314, gm_n76, in_9, gm_n803, gm_n339);
	nor (gm_n4045, gm_n441, in_21, gm_n55, gm_n4044);
	nor (gm_n4046, gm_n4045, gm_n4043, gm_n4041);
	nand (gm_n4047, gm_n90, in_10, gm_n62, gm_n2443, gm_n624);
	nor (gm_n4048, gm_n368, gm_n246, gm_n119, gm_n4047);
	nand (gm_n4049, in_14, in_10, in_9, gm_n1071, gm_n334);
	nor (gm_n4050, gm_n824, gm_n167, in_18, gm_n4049);
	nand (gm_n4051, in_13, in_9, gm_n94, gm_n1692, gm_n123);
	nor (gm_n4052, gm_n105, in_21, in_17, gm_n4051, gm_n620);
	nor (gm_n4053, gm_n4052, gm_n4050, gm_n4048);
	nand (gm_n4054, gm_n4039, gm_n3894, gm_n3892, gm_n4053, gm_n4046);
	nor (gm_n4055, gm_n133, gm_n90, gm_n78, gm_n350, gm_n148);
	nand (gm_n4056, gm_n806, gm_n199, in_18, gm_n4055);
	and (gm_n4057, gm_n61, in_16, gm_n59, gm_n535, gm_n222);
	nand (gm_n4058, gm_n495, in_21, gm_n85, gm_n4057);
	nor (gm_n4059, gm_n193, gm_n56, gm_n60, gm_n1789, gm_n485);
	nand (gm_n4060, gm_n4059, gm_n72, gm_n85);
	nand (gm_n4061, gm_n4060, gm_n4058, gm_n4056);
	nor (gm_n4062, gm_n406, in_13, in_9, gm_n743, gm_n344);
	nand (gm_n4063, gm_n122, gm_n72, in_17, gm_n4062, gm_n327);
	nor (gm_n4064, gm_n358, gm_n76, in_9, gm_n503, gm_n596);
	nand (gm_n4065, gm_n311, gm_n72, in_17, gm_n4064, gm_n339);
	nor (gm_n4066, gm_n92, gm_n78, in_9, gm_n344, gm_n1295);
	nand (gm_n4067, gm_n199, gm_n119, gm_n90, gm_n4066, gm_n245);
	nand (gm_n4068, gm_n4067, gm_n4065, gm_n4063);
	nor (gm_n4069, gm_n4054, gm_n3890, gm_n3888, gm_n4068, gm_n4061);
	nand (gm_n4070, gm_n1076, in_13, in_9, gm_n1186, gm_n402);
	nor (gm_n4071, gm_n441, in_21, in_17, gm_n4070);
	nand (gm_n4072, gm_n64, gm_n59, gm_n94, gm_n455, gm_n571);
	nor (gm_n4073, in_21, gm_n85, in_16, gm_n4072, gm_n384);
	nand (gm_n4074, gm_n122, in_13, in_9, gm_n586, gm_n314);
	nor (gm_n4075, gm_n183, gm_n72, in_17, gm_n4074);
	nor (gm_n4076, gm_n4075, gm_n4073, gm_n4071);
	and (gm_n4077, gm_n166, gm_n164, gm_n119, gm_n2134);
	nand (gm_n4078, gm_n126, in_13, gm_n62, gm_n341, gm_n340);
	nor (gm_n4079, gm_n183, gm_n72, in_17, gm_n4078, gm_n313);
	nand (gm_n4080, gm_n264, in_16, in_12, gm_n2646, gm_n949);
	nor (gm_n4081, gm_n219, in_21, in_20, gm_n4080);
	nor (gm_n4082, gm_n4081, gm_n4079, gm_n4077);
	nand (gm_n4083, gm_n4069, gm_n3885, gm_n3883, gm_n4082, gm_n4076);
	nor (gm_n4084, gm_n115, in_16, in_12, gm_n1052, gm_n220);
	nand (gm_n4085, gm_n495, gm_n72, gm_n85, gm_n4084);
	and (gm_n4086, in_13, in_9, gm_n94, gm_n756, gm_n402);
	nand (gm_n4087, gm_n104, in_21, in_17, gm_n4086, gm_n206);
	nand (gm_n4088, in_7, in_6, in_5, gm_n134, in_8);
	nor (gm_n4089, gm_n158, in_16, gm_n59, gm_n4088, gm_n220);
	nand (gm_n4090, gm_n383, gm_n72, gm_n85, gm_n4089);
	nand (gm_n4091, gm_n4090, gm_n4087, gm_n4085);
	nor (gm_n4092, gm_n114, in_16, in_12, gm_n230, gm_n158);
	nand (gm_n4093, gm_n113, in_21, gm_n85, gm_n4092);
	nor (gm_n4094, gm_n406, gm_n76, in_9, gm_n621, gm_n443);
	nand (gm_n4095, gm_n405, in_21, in_17, gm_n4094, gm_n327);
	nor (gm_n4096, gm_n152, gm_n59, gm_n94, gm_n2769, gm_n274);
	nand (gm_n4097, in_21, in_20, gm_n73, gm_n4096, gm_n697);
	nand (gm_n4098, gm_n4097, gm_n4095, gm_n4093);
	nor (gm_n4099, gm_n4083, gm_n3881, gm_n3879, gm_n4098, gm_n4091);
	nand (gm_n4100, gm_n233, in_16, gm_n59, gm_n1970, gm_n303);
	nor (gm_n4101, gm_n219, gm_n72, gm_n85, gm_n4100);
	or (gm_n4102, gm_n461, gm_n76, gm_n62, gm_n1132, gm_n430);
	nor (gm_n4103, gm_n183, in_21, in_17, gm_n4102, gm_n184);
	nand (gm_n4104, gm_n64, in_13, in_12, gm_n547);
	nor (gm_n4105, gm_n441, in_21, in_17, gm_n4104, gm_n184);
	nor (gm_n4106, gm_n4105, gm_n4103, gm_n4101);
	or (gm_n4107, gm_n609, gm_n76, gm_n62, gm_n462, gm_n431);
	nor (gm_n4108, gm_n121, in_21, in_17, gm_n4107, gm_n441);
	nand (gm_n4109, gm_n222, gm_n192, gm_n60, gm_n2096, gm_n486);
	nor (gm_n4110, in_21, in_20, gm_n56, gm_n4109);
	or (gm_n4111, gm_n213, gm_n191, gm_n60, gm_n1170, gm_n290);
	nor (gm_n4112, gm_n72, in_20, gm_n56, gm_n4111);
	nor (gm_n4113, gm_n4112, gm_n4110, gm_n4108);
	nand (gm_n4114, gm_n4099, gm_n3878, gm_n3875, gm_n4113, gm_n4106);
	nor (gm_n4115, in_14, gm_n78, in_9, gm_n2002, gm_n207);
	nand (gm_n4116, gm_n245, gm_n86, in_18, gm_n4115);
	nor (gm_n4117, gm_n358, in_13, in_9, gm_n503, gm_n443);
	nand (gm_n4118, gm_n102, in_21, in_17, gm_n4117, gm_n339);
	nor (gm_n4119, gm_n362, gm_n90, in_10, gm_n589, gm_n370);
	nand (gm_n4120, gm_n245, gm_n164, gm_n119, gm_n4119);
	nand (gm_n4121, gm_n4120, gm_n4118, gm_n4116);
	nor (gm_n4122, gm_n358, in_13, gm_n62, gm_n1583, gm_n344);
	nand (gm_n4123, gm_n254, in_21, in_17, gm_n4122, gm_n1076);
	or (gm_n4124, in_21, in_20, in_19, gm_n2724, gm_n269);
	nor (gm_n4125, gm_n667, in_13, gm_n62, gm_n597, gm_n442);
	nand (gm_n4126, gm_n595, gm_n72, in_17, gm_n4125, gm_n373);
	nand (gm_n4127, gm_n4126, gm_n4124, gm_n4123);
	nor (gm_n4128, gm_n4114, gm_n3873, gm_n3871, gm_n4127, gm_n4121);
	or (gm_n4129, gm_n1295, gm_n76, gm_n62, gm_n344, gm_n257);
	nor (gm_n4130, gm_n374, gm_n72, gm_n55, gm_n4129, gm_n375);
	or (gm_n4131, gm_n227, gm_n73, in_12, gm_n1475, gm_n297);
	nor (gm_n4132, gm_n219, in_21, in_20, gm_n4131);
	or (gm_n4133, gm_n358, in_13, in_9, gm_n1583, gm_n463);
	nor (gm_n4134, gm_n121, in_21, gm_n55, gm_n4133, gm_n479);
	nor (gm_n4135, gm_n4134, gm_n4132, gm_n4130);
	nand (gm_n4136, in_14, gm_n78, gm_n62, gm_n2608, gm_n600);
	nor (gm_n4137, gm_n212, gm_n130, in_18, gm_n4136);
	or (gm_n4138, gm_n191, gm_n190, gm_n60, gm_n562, gm_n643);
	nor (gm_n4139, in_21, in_20, in_19, gm_n4138);
	or (gm_n4140, in_13, gm_n62, in_8, gm_n442, gm_n909);
	nor (gm_n4141, gm_n121, in_21, in_17, gm_n4140, gm_n374);
	nor (gm_n4142, gm_n4141, gm_n4139, gm_n4137);
	nand (gm_n4143, gm_n4128, gm_n3869, gm_n3867, gm_n4142, gm_n4135);
	nor (gm_n4144, gm_n667, gm_n76, gm_n62, gm_n1132, gm_n461);
	nand (gm_n4145, gm_n174, in_21, in_17, gm_n4144, gm_n1076);
	and (gm_n4146, gm_n61, in_16, in_12, gm_n884, gm_n79);
	nand (gm_n4147, gm_n383, gm_n72, gm_n85, gm_n4146);
	nor (gm_n4148, gm_n818, in_13, in_9, gm_n344, gm_n461);
	nand (gm_n4149, gm_n104, in_21, gm_n55, gm_n4148, gm_n120);
	nand (gm_n4150, gm_n4149, gm_n4147, gm_n4145);
	nor (gm_n4151, gm_n297, in_16, in_12, gm_n324, gm_n385);
	nand (gm_n4152, gm_n138, gm_n72, gm_n85, gm_n4151);
	nor (gm_n4153, gm_n514, in_13, gm_n62, gm_n743, gm_n344);
	nand (gm_n4154, gm_n311, in_21, in_17, gm_n4153, gm_n339);
	and (gm_n4155, gm_n61, gm_n73, in_12, gm_n1001, gm_n64);
	nand (gm_n4156, gm_n383, gm_n72, gm_n85, gm_n4155);
	nand (gm_n4157, gm_n4156, gm_n4154, gm_n4152);
	nor (gm_n4158, gm_n4143, gm_n3865, gm_n3863, gm_n4157, gm_n4150);
	nand (gm_n4159, gm_n1158, gm_n90, gm_n78, gm_n722, gm_n490);
	nor (gm_n4160, gm_n824, gm_n167, gm_n119, gm_n4159);
	and (gm_n4161, gm_n523, in_21, gm_n55, gm_n1249, gm_n311);
	nand (gm_n4162, gm_n122, gm_n76, gm_n62, gm_n2942, gm_n788);
	nor (gm_n4163, gm_n620, in_21, gm_n55, gm_n4162);
	nor (gm_n4164, gm_n4163, gm_n4161, gm_n4160);
	nand (gm_n4165, gm_n61, in_16, in_12, gm_n685, gm_n154);
	nor (gm_n4166, gm_n262, in_21, in_20, gm_n4165);
	nand (gm_n4167, gm_n264, gm_n75, in_15, gm_n1427, gm_n449);
	nor (gm_n4168, gm_n72, in_20, in_19, gm_n4167);
	or (gm_n4169, gm_n114, in_12, in_8, gm_n417, gm_n297);
	nor (gm_n4170, gm_n72, gm_n85, in_16, gm_n4169, gm_n262);
	nor (gm_n4171, gm_n4170, gm_n4168, gm_n4166);
	nand (gm_n4172, gm_n4158, gm_n3861, gm_n3859, gm_n4171, gm_n4164);
	nor (gm_n4173, gm_n358, gm_n76, in_9, gm_n1132, gm_n667);
	nand (gm_n4174, gm_n104, in_21, gm_n55, gm_n4173, gm_n174);
	nor (gm_n4175, gm_n358, gm_n76, in_9, gm_n1583, gm_n596);
	nand (gm_n4176, gm_n102, gm_n72, gm_n55, gm_n4175, gm_n122);
	and (gm_n4177, gm_n64, in_13, in_12, gm_n998);
	nand (gm_n4178, gm_n523, in_21, gm_n55, gm_n4177, gm_n254);
	nand (gm_n4179, gm_n4178, gm_n4176, gm_n4174);
	nor (gm_n4180, gm_n514, gm_n76, in_9, gm_n1583, gm_n463);
	nand (gm_n4181, gm_n327, in_21, in_17, gm_n4180, gm_n339);
	nor (gm_n4182, gm_n248, gm_n90, in_10, gm_n438, gm_n369);
	nand (gm_n4183, gm_n348, gm_n806, gm_n119, gm_n4182);
	and (gm_n4184, gm_n484, gm_n60, in_11, gm_n576, gm_n555);
	nand (gm_n4185, gm_n72, in_20, gm_n56, gm_n4184, gm_n75);
	nand (gm_n4186, gm_n4185, gm_n4183, gm_n4181);
	nor (gm_n4187, gm_n4172, gm_n3857, gm_n3855, gm_n4186, gm_n4179);
	nor (gm_n4188, gm_n90, gm_n78, gm_n62, gm_n1475, gm_n147);
	nand (gm_n4189, gm_n243, gm_n166, gm_n119, gm_n4188);
	and (gm_n4190, in_14, in_10, gm_n62, gm_n2624, gm_n91);
	nand (gm_n4191, gm_n348, gm_n88, gm_n119, gm_n4190);
	and (gm_n4192, in_13, gm_n62, gm_n94, gm_n601, gm_n314);
	nand (gm_n4193, gm_n255, gm_n72, in_17, gm_n4192, gm_n373);
	nand (gm_n4194, gm_n4189, gm_n4187, gm_n3853, gm_n4193, gm_n4191);
	and (gm_n4195, in_14, in_10, in_9, gm_n2070, gm_n624);
	nand (gm_n4196, gm_n367, gm_n131, in_18, gm_n4195);
	nor (gm_n4197, gm_n95, in_14, gm_n78, gm_n133, gm_n99);
	nand (gm_n4198, gm_n323, gm_n243, gm_n119, gm_n4197);
	and (gm_n4199, gm_n106, gm_n828, gm_n76, gm_n793, gm_n595);
	nand (gm_n4200, gm_n206, in_21, gm_n55, gm_n4199);
	nand (gm_n4201, gm_n4200, gm_n4198, gm_n4196);
	nor (out_10, gm_n4194, gm_n3851, t_1, gm_n4201);
	nand (gm_n4203, gm_n523, gm_n76, gm_n62, gm_n2712, gm_n314);
	nor (gm_n4204, gm_n620, in_21, in_17, gm_n4203);
	nand (gm_n4205, gm_n102, gm_n72, gm_n55, gm_n1224, gm_n104);
	nand (gm_n4206, gm_n106, gm_n76, in_9, gm_n2346, gm_n523);
	nor (gm_n4207, gm_n374, gm_n72, gm_n55, gm_n4206);
	nand (gm_n4208, gm_n555, in_15, in_11, gm_n756, gm_n545);
	nor (gm_n4209, gm_n72, in_20, gm_n56, gm_n4208, gm_n191);
	nand (gm_n4210, gm_n102, in_21, in_17, gm_n3389, gm_n104);
	nor (gm_n4211, gm_n430, gm_n76, gm_n62, gm_n359, gm_n431);
	nand (gm_n4212, gm_n405, in_21, gm_n55, gm_n4211, gm_n373);
	or (gm_n4213, gm_n358, in_13, gm_n62, gm_n743, gm_n596);
	nor (gm_n4214, gm_n121, in_21, gm_n55, gm_n4213, gm_n479);
	or (gm_n4215, gm_n1331, gm_n158, gm_n60, gm_n1191, gm_n760);
	nor (gm_n4216, in_21, in_20, in_19, gm_n4215);
	nor (gm_n4217, in_14, gm_n78, in_9, gm_n1837, gm_n467);
	nand (gm_n4218, gm_n367, gm_n88, in_18, gm_n4217);
	nor (gm_n4219, gm_n263, in_16, in_12, gm_n821, gm_n276);
	nand (gm_n4220, gm_n138, gm_n72, gm_n85, gm_n4219);
	or (gm_n4221, gm_n90, in_10, gm_n62, gm_n1284, gm_n467);
	nor (gm_n4222, gm_n531, gm_n167, in_18, gm_n4221);
	or (gm_n4223, gm_n247, gm_n121, in_13, gm_n431, gm_n259);
	nor (gm_n4224, gm_n374, gm_n72, gm_n55, gm_n4223);
	and (gm_n4225, gm_n264, gm_n75, in_15, gm_n1427, gm_n422);
	nand (gm_n4226, gm_n72, gm_n85, in_19, gm_n4225);
	nor (gm_n4227, gm_n220, in_16, gm_n59, gm_n2333, gm_n274);
	nand (gm_n4228, gm_n383, gm_n72, gm_n85, gm_n4227);
	nand (gm_n4229, gm_n379, gm_n143, gm_n60, gm_n1398, gm_n547);
	nor (gm_n4230, in_21, in_20, in_19, gm_n4229);
	nand (gm_n4231, gm_n76, in_9, gm_n94, gm_n556, gm_n106);
	nor (gm_n4232, gm_n388, gm_n72, gm_n55, gm_n4231, gm_n256);
	nor (gm_n4233, gm_n461, in_13, in_9, gm_n675, gm_n328);
	nand (gm_n4234, gm_n373, in_21, gm_n55, gm_n4233);
	nor (gm_n4235, gm_n90, in_10, gm_n62, gm_n3099, gm_n362);
	nand (gm_n4236, gm_n323, gm_n86, in_18, gm_n4235);
	nand (gm_n4237, gm_n107, in_13, gm_n62, gm_n316, gm_n579);
	nor (gm_n4238, gm_n184, in_21, in_17, gm_n4237, gm_n620);
	nand (gm_n4239, gm_n104, gm_n76, in_9, gm_n1359, gm_n340);
	nor (gm_n4240, gm_n620, gm_n72, in_17, gm_n4239);
	nand (gm_n4241, gm_n104, in_21, gm_n55, gm_n3812, gm_n120);
	nor (gm_n4242, in_14, in_10, gm_n62, gm_n1906, gm_n207);
	nand (gm_n4243, gm_n348, gm_n88, gm_n119, gm_n4242);
	nand (gm_n4244, gm_n123, in_13, in_9, gm_n2283, gm_n405);
	nor (gm_n4245, gm_n388, in_21, gm_n55, gm_n4244);
	nor (gm_n4246, gm_n461, gm_n76, gm_n62, gm_n462, gm_n596);
	and (gm_n4247, gm_n120, gm_n72, gm_n55, gm_n4246, gm_n405);
	nor (gm_n4248, gm_n514, in_13, gm_n62, gm_n432, gm_n609);
	nand (gm_n4249, gm_n311, gm_n72, in_17, gm_n4248, gm_n1076);
	nand (gm_n4250, gm_n574, gm_n164);
	nand (gm_n4251, gm_n490, gm_n91, in_10, gm_n722);
	nor (gm_n4252, gm_n121, gm_n72, in_17, gm_n4251, gm_n441);
	or (gm_n4253, gm_n227, in_16, in_12, gm_n695, gm_n297);
	nor (gm_n4254, gm_n496, in_21, gm_n85, gm_n4253);
	nor (gm_n4255, gm_n431, in_13, in_9, gm_n743, gm_n463);
	nand (gm_n4256, gm_n523, in_21, in_17, gm_n4255, gm_n206);
	nor (gm_n4257, gm_n841, gm_n92, gm_n90, gm_n981, gm_n271);
	nand (gm_n4258, gm_n4257, gm_n164, gm_n119);
	or (gm_n4259, gm_n257, in_13, in_9, gm_n481, gm_n596);
	nor (gm_n4260, gm_n620, gm_n72, in_17, gm_n4259, gm_n375);
	nand (gm_n4261, gm_n64, gm_n73, gm_n59, gm_n1758, gm_n303);
	nor (gm_n4262, gm_n58, gm_n72, in_20, gm_n4261);
	and (gm_n4263, gm_n106, in_13, gm_n62, gm_n1076, gm_n235);
	nand (gm_n4264, gm_n373, gm_n72, in_17, gm_n4263);
	nor (gm_n4265, gm_n99, gm_n90, in_10, gm_n362, gm_n148);
	nand (gm_n4266, gm_n243, gm_n88, gm_n119, gm_n4265);
	nand (gm_n4267, gm_n448, gm_n154, in_15, gm_n1135, gm_n449);
	nor (gm_n4268, gm_n72, gm_n85, in_19, gm_n4267);
	or (gm_n4269, gm_n514, in_13, in_9, gm_n481, gm_n609);
	nor (gm_n4270, gm_n479, gm_n72, in_17, gm_n4269, gm_n375);
	nor (gm_n4271, gm_n667, gm_n76, gm_n62, gm_n462, gm_n442);
	nand (gm_n4272, gm_n255, in_21, gm_n55, gm_n4271, gm_n373);
	nor (gm_n4273, gm_n269, gm_n213, gm_n60, gm_n355, gm_n290);
	nand (gm_n4274, gm_n72, in_20, in_19, gm_n4273);
	nor (gm_n4275, gm_n667, in_13, in_9, gm_n988, gm_n442);
	nand (gm_n4276, gm_n174, gm_n72, gm_n55, gm_n4275, gm_n339);
	nor (gm_n4277, gm_n358, gm_n76, gm_n62, gm_n2077, gm_n256);
	nand (gm_n4278, gm_n373, in_21, gm_n55, gm_n4277);
	nand (gm_n4279, gm_n367, gm_n166, gm_n119, gm_n3412);
	nand (gm_n4280, gm_n4276, gm_n4274, gm_n4272, gm_n4279, gm_n4278);
	nor (gm_n4281, gm_n155, gm_n73, gm_n59, gm_n2340, gm_n385);
	nand (gm_n4282, gm_n57, gm_n72, gm_n85, gm_n4281);
	and (gm_n4283, in_10, in_9, in_8, gm_n714, gm_n624);
	nand (gm_n4284, gm_n146, gm_n119, in_14, gm_n4283, gm_n436);
	nor (gm_n4285, gm_n213, gm_n159, in_15, gm_n485, gm_n3052);
	nand (gm_n4286, gm_n72, gm_n85, gm_n56, gm_n4285);
	nand (gm_n4287, gm_n4286, gm_n4284, gm_n4282);
	nor (gm_n4288, gm_n605, in_15, gm_n63, gm_n3754, gm_n760);
	nand (gm_n4289, gm_n72, gm_n85, in_19, gm_n4288, gm_n486);
	or (gm_n4290, gm_n105, in_21, in_17, gm_n2321, gm_n620);
	nor (gm_n4291, gm_n190, in_16, gm_n59, gm_n648, gm_n152);
	nand (gm_n4292, gm_n296, gm_n72, gm_n85, gm_n4291);
	nand (gm_n4293, gm_n4292, gm_n4290, gm_n4289);
	nor (gm_n4294, gm_n4280, gm_n4270, gm_n4268, gm_n4293, gm_n4287);
	nand (gm_n4295, gm_n222, gm_n75, gm_n60, gm_n953, gm_n422);
	nor (gm_n4296, gm_n72, in_20, gm_n56, gm_n4295);
	nand (gm_n4297, gm_n64, in_16, gm_n59, gm_n586, gm_n949);
	nor (gm_n4298, gm_n219, gm_n72, in_20, gm_n4297);
	nand (gm_n4299, gm_n90, in_10, in_9, gm_n672, gm_n1158);
	nor (gm_n4300, gm_n368, gm_n212, gm_n119, gm_n4299);
	nor (gm_n4301, gm_n4300, gm_n4298, gm_n4296);
	nand (gm_n4302, gm_n995, in_14, in_10, gm_n793, gm_n1011);
	nor (gm_n4303, gm_n531, gm_n246, gm_n119, gm_n4302);
	nand (gm_n4304, gm_n61, gm_n73, gm_n59, gm_n487, gm_n143);
	nor (gm_n4305, gm_n384, gm_n72, in_20, gm_n4304);
	nand (gm_n4306, in_14, in_10, in_9, gm_n1392, gm_n600);
	nor (gm_n4307, gm_n437, gm_n87, in_18, gm_n4306);
	nor (gm_n4308, gm_n4307, gm_n4305, gm_n4303);
	nand (gm_n4309, gm_n4294, gm_n4266, gm_n4264, gm_n4308, gm_n4301);
	nor (gm_n4310, gm_n121, in_13, in_9, gm_n2697, gm_n431);
	nand (gm_n4311, gm_n206, gm_n72, in_17, gm_n4310);
	nor (gm_n4312, gm_n461, in_13, in_9, gm_n462, gm_n443);
	nand (gm_n4313, gm_n122, gm_n72, gm_n55, gm_n4312, gm_n311);
	nor (gm_n4314, gm_n257, gm_n76, gm_n62, gm_n988, gm_n596);
	nand (gm_n4315, gm_n311, gm_n72, in_17, gm_n4314, gm_n339);
	nand (gm_n4316, gm_n4315, gm_n4313, gm_n4311);
	and (gm_n4317, gm_n1144, gm_n60, gm_n63, gm_n714, gm_n545);
	nand (gm_n4318, gm_n72, in_20, in_19, gm_n4317, gm_n486);
	nor (gm_n4319, gm_n461, in_13, in_9, gm_n988, gm_n596);
	nand (gm_n4320, gm_n102, in_21, in_17, gm_n4319, gm_n1076);
	nor (gm_n4321, gm_n461, gm_n76, in_9, gm_n503, gm_n502);
	nand (gm_n4322, gm_n102, gm_n72, in_17, gm_n4321, gm_n122);
	nand (gm_n4323, gm_n4322, gm_n4320, gm_n4318);
	nor (gm_n4324, gm_n4309, gm_n4262, gm_n4260, gm_n4323, gm_n4316);
	or (gm_n4325, gm_n480, gm_n76, gm_n62, gm_n597, gm_n463);
	nor (gm_n4326, gm_n105, gm_n72, in_17, gm_n4325, gm_n441);
	nand (gm_n4327, gm_n77, gm_n73, in_12, gm_n1970, gm_n143);
	nor (gm_n4328, gm_n384, in_21, in_20, gm_n4327);
	or (gm_n4329, gm_n358, gm_n76, in_9, gm_n1583, gm_n502);
	nor (gm_n4330, gm_n441, gm_n72, in_17, gm_n4329, gm_n184);
	nor (gm_n4331, gm_n4330, gm_n4328, gm_n4326);
	or (gm_n4332, gm_n90, gm_n78, in_9, gm_n355, gm_n207);
	nor (gm_n4333, gm_n1989, gm_n87, in_18, gm_n4332);
	or (gm_n4334, gm_n259, in_14, gm_n78, gm_n491, gm_n807);
	nor (gm_n4335, gm_n244, gm_n212, gm_n119, gm_n4334);
	or (gm_n4336, gm_n155, gm_n74, gm_n60, gm_n2589, gm_n643);
	nor (gm_n4337, gm_n72, gm_n85, gm_n56, gm_n4336);
	nor (gm_n4338, gm_n4337, gm_n4335, gm_n4333);
	nand (gm_n4339, gm_n4324, gm_n4258, gm_n4256, gm_n4338, gm_n4331);
	nor (gm_n4340, gm_n596, gm_n76, in_9, gm_n462, gm_n480);
	nand (gm_n4341, gm_n102, in_21, in_17, gm_n4340, gm_n122);
	nor (gm_n4342, gm_n358, gm_n76, gm_n62, gm_n443, gm_n432);
	nand (gm_n4343, gm_n102, in_21, gm_n55, gm_n4342, gm_n339);
	and (gm_n4344, gm_n76, gm_n62, in_8, gm_n1263, gm_n579);
	nand (gm_n4345, gm_n523, in_21, in_17, gm_n4344, gm_n206);
	nand (gm_n4346, gm_n4345, gm_n4343, gm_n4341);
	nor (gm_n4347, gm_n114, in_16, in_12, gm_n730, gm_n155);
	nand (gm_n4348, gm_n383, gm_n72, in_20, gm_n4347);
	nor (gm_n4349, gm_n358, gm_n76, in_9, gm_n988, gm_n667);
	nand (gm_n4350, gm_n523, in_21, gm_n55, gm_n4349, gm_n206);
	nor (gm_n4351, gm_n78, gm_n62, in_8, gm_n508, gm_n807);
	nand (gm_n4352, gm_n86, in_18, gm_n90, gm_n4351, gm_n200);
	nand (gm_n4353, gm_n4352, gm_n4350, gm_n4348);
	nor (gm_n4354, gm_n4339, gm_n4254, gm_n4252, gm_n4353, gm_n4346);
	or (gm_n4355, gm_n667, in_13, gm_n62, gm_n462, gm_n480);
	nor (gm_n4356, gm_n183, in_21, gm_n55, gm_n4355, gm_n184);
	nand (gm_n4357, gm_n221, in_16, in_12, gm_n751, gm_n264);
	nor (gm_n4358, gm_n139, in_21, in_20, gm_n4357);
	or (gm_n4359, gm_n90, gm_n78, in_9, gm_n835, gm_n133);
	nor (gm_n4360, gm_n244, gm_n89, in_18, gm_n4359);
	nor (gm_n4361, gm_n4360, gm_n4358, gm_n4356);
	or (gm_n4362, gm_n313, gm_n76, in_9, gm_n675, gm_n406);
	nor (gm_n4363, gm_n103, in_21, in_17, gm_n4362);
	nand (gm_n4364, gm_n339, in_13, in_9, gm_n1186, gm_n340);
	nor (gm_n4365, gm_n388, in_21, in_17, gm_n4364);
	nand (gm_n4366, gm_n90, gm_n78, gm_n62, gm_n1501, gm_n600);
	nor (gm_n4367, gm_n531, gm_n212, in_18, gm_n4366);
	nor (gm_n4368, gm_n4367, gm_n4365, gm_n4363);
	nand (gm_n4369, gm_n4354, gm_n4250, gm_n4249, gm_n4368, gm_n4361);
	nor (gm_n4370, gm_n247, gm_n461, gm_n76, gm_n414, gm_n328);
	nand (gm_n4371, gm_n311, gm_n72, in_17, gm_n4370);
	nor (gm_n4372, gm_n220, gm_n73, in_12, gm_n1731, gm_n263);
	nand (gm_n4373, gm_n383, in_21, gm_n85, gm_n4372);
	nand (gm_n4374, gm_n523, gm_n72, in_17, gm_n3856, gm_n373);
	nand (gm_n4375, gm_n4374, gm_n4373, gm_n4371);
	and (gm_n4376, gm_n126, gm_n76, in_9, gm_n340, gm_n186);
	nand (gm_n4377, gm_n206, gm_n72, in_17, gm_n4376, gm_n595);
	nand (gm_n4378, gm_n122, in_21, gm_n55, gm_n3895, gm_n327);
	and (gm_n4379, gm_n90, gm_n78, gm_n62, gm_n3454, gm_n713);
	nand (gm_n4380, gm_n245, gm_n146, in_18, gm_n4379);
	nand (gm_n4381, gm_n4380, gm_n4378, gm_n4377);
	nor (gm_n4382, gm_n4369, gm_n4247, gm_n4245, gm_n4381, gm_n4375);
	nand (gm_n4383, gm_n214, gm_n73, in_12, gm_n2573, gm_n571);
	nor (gm_n4384, gm_n262, gm_n72, gm_n85, gm_n4383);
	nand (gm_n4385, gm_n78, gm_n62, gm_n94, gm_n1263, gm_n334);
	nor (gm_n4386, gm_n130, in_18, gm_n90, gm_n4385, gm_n132);
	or (gm_n4387, gm_n480, gm_n76, in_9, gm_n743, gm_n502);
	nor (gm_n4388, gm_n620, in_21, in_17, gm_n4387, gm_n662);
	nor (gm_n4389, gm_n4388, gm_n4386, gm_n4384);
	nand (gm_n4390, gm_n143, in_12, in_8, gm_n455, gm_n949);
	nor (gm_n4391, in_21, gm_n85, gm_n73, gm_n4390, gm_n912);
	or (gm_n4392, gm_n609, in_13, in_9, gm_n432, gm_n406);
	nor (gm_n4393, gm_n105, in_21, gm_n55, gm_n4392, gm_n312);
	or (gm_n4394, gm_n133, in_14, in_10, gm_n491, gm_n248);
	nor (gm_n4395, gm_n244, gm_n89, in_18, gm_n4394);
	nor (gm_n4396, gm_n4395, gm_n4393, gm_n4391);
	nand (gm_n4397, gm_n4382, gm_n4243, gm_n4241, gm_n4396, gm_n4389);
	nor (gm_n4398, gm_n168, gm_n60, gm_n63, gm_n842, gm_n240);
	nand (gm_n4399, gm_n72, in_20, gm_n56, gm_n4398, gm_n394);
	nor (gm_n4400, gm_n155, gm_n73, in_12, gm_n1246, gm_n319);
	nand (gm_n4401, gm_n697, gm_n72, in_20, gm_n4400);
	nor (gm_n4402, gm_n158, gm_n73, in_12, gm_n1884, gm_n220);
	nand (gm_n4403, gm_n138, in_21, in_20, gm_n4402);
	nand (gm_n4404, gm_n4403, gm_n4401, gm_n4399);
	nor (gm_n4405, gm_n274, gm_n193, in_15, gm_n705, gm_n447);
	nand (gm_n4406, gm_n72, in_20, in_19, gm_n4405);
	nor (gm_n4407, gm_n461, in_13, in_9, gm_n502, gm_n345);
	nand (gm_n4408, gm_n122, in_21, in_17, gm_n4407, gm_n311);
	nor (gm_n4409, gm_n158, gm_n74, gm_n60, gm_n849, gm_n643);
	nand (gm_n4410, in_21, in_20, gm_n56, gm_n4409);
	nand (gm_n4411, gm_n4410, gm_n4408, gm_n4406);
	nor (gm_n4412, gm_n4397, gm_n4240, gm_n4238, gm_n4411, gm_n4404);
	or (gm_n4413, gm_n121, gm_n99, gm_n76, gm_n442, gm_n349);
	nor (gm_n4414, gm_n103, in_21, in_17, gm_n4413);
	nand (gm_n4415, gm_n523, in_13, gm_n62, gm_n1030, gm_n579);
	nor (gm_n4416, gm_n183, gm_n72, in_17, gm_n4415);
	or (gm_n4417, gm_n90, in_10, in_9, gm_n3402, gm_n467);
	nor (gm_n4418, gm_n1989, gm_n87, in_18, gm_n4417);
	nor (gm_n4419, gm_n4418, gm_n4416, gm_n4414);
	or (gm_n4420, gm_n274, in_16, in_12, gm_n385, gm_n278);
	nor (gm_n4421, gm_n139, in_21, in_20, gm_n4420);
	nand (gm_n4422, gm_n571, gm_n233, gm_n59, gm_n1392);
	nor (gm_n4423, gm_n72, in_20, gm_n56, gm_n4422, gm_n269);
	nand (gm_n4424, gm_n402, gm_n76, in_9, gm_n1401);
	nor (gm_n4425, gm_n183, in_21, in_17, gm_n4424, gm_n662);
	nor (gm_n4426, gm_n4425, gm_n4423, gm_n4421);
	nand (gm_n4427, gm_n4412, gm_n4236, gm_n4234, gm_n4426, gm_n4419);
	nor (gm_n4428, gm_n190, gm_n73, gm_n59, gm_n2963, gm_n152);
	nand (gm_n4429, gm_n138, gm_n72, in_20, gm_n4428);
	nor (gm_n4430, gm_n344, in_13, in_9, gm_n442, gm_n359);
	nand (gm_n4431, gm_n120, gm_n72, gm_n55, gm_n4430, gm_n523);
	nor (gm_n4432, gm_n430, gm_n76, gm_n62, gm_n481, gm_n406);
	nand (gm_n4433, gm_n120, gm_n72, in_17, gm_n4432, gm_n339);
	nand (gm_n4434, gm_n4433, gm_n4431, gm_n4429);
	nand (gm_n4435, gm_n123, in_13, in_9, gm_n1401, gm_n595);
	or (gm_n4436, gm_n620, gm_n72, gm_n55, gm_n4435);
	nand (gm_n4437, gm_n305, gm_n304, in_8);
	nor (gm_n4438, gm_n297, in_16, gm_n59, gm_n4437, gm_n385);
	nand (gm_n4439, gm_n495, gm_n72, gm_n85, gm_n4438);
	nor (gm_n4440, gm_n461, in_13, gm_n62, gm_n481, gm_n463);
	nand (gm_n4441, gm_n120, gm_n72, gm_n55, gm_n4440, gm_n255);
	nand (gm_n4442, gm_n4441, gm_n4439, gm_n4436);
	nor (gm_n4443, gm_n4427, gm_n4232, gm_n4230, gm_n4442, gm_n4434);
	or (gm_n4444, gm_n227, in_16, gm_n59, gm_n3315, gm_n297);
	nor (gm_n4445, gm_n262, gm_n72, gm_n85, gm_n4444);
	nand (gm_n4446, gm_n214, in_16, in_12, gm_n875, gm_n221);
	nor (gm_n4447, gm_n912, gm_n72, gm_n85, gm_n4446);
	or (gm_n4448, gm_n514, in_13, in_9, gm_n597, gm_n443);
	nor (gm_n4449, gm_n105, gm_n72, in_17, gm_n4448, gm_n388);
	nor (gm_n4450, gm_n4449, gm_n4447, gm_n4445);
	nand (gm_n4451, gm_n233, in_16, in_12, gm_n2070, gm_n733);
	nor (gm_n4452, gm_n912, gm_n72, in_20, gm_n4451);
	nand (gm_n4453, gm_n125, in_13, in_9, gm_n316, gm_n185);
	nor (gm_n4454, gm_n374, in_21, in_17, gm_n4453, gm_n375);
	or (gm_n4455, in_14, in_10, gm_n62, gm_n1319, gm_n147);
	nor (gm_n4456, gm_n246, gm_n165, gm_n119, gm_n4455);
	nor (gm_n4457, gm_n4456, gm_n4454, gm_n4452);
	nand (gm_n4458, gm_n4443, gm_n4228, gm_n4226, gm_n4457, gm_n4450);
	nor (gm_n4459, gm_n263, in_16, in_12, gm_n552, gm_n354);
	nand (gm_n4460, gm_n179, gm_n72, gm_n85, gm_n4459);
	nor (gm_n4461, gm_n431, gm_n76, gm_n62, gm_n502, gm_n462);
	nand (gm_n4462, gm_n104, in_21, in_17, gm_n4461, gm_n174);
	nor (gm_n4463, gm_n114, gm_n73, in_12, gm_n2060, gm_n158);
	nand (gm_n4464, gm_n296, in_21, in_20, gm_n4463);
	nand (gm_n4465, gm_n4464, gm_n4462, gm_n4460);
	nor (gm_n4466, gm_n227, gm_n73, gm_n59, gm_n3929, gm_n297);
	nand (gm_n4467, gm_n296, gm_n72, gm_n85, gm_n4466);
	nor (gm_n4468, gm_n190, in_16, in_12, gm_n1519, gm_n152);
	nand (gm_n4469, gm_n383, gm_n72, in_20, gm_n4468);
	and (gm_n4470, gm_n264, in_16, in_12, gm_n2885, gm_n949);
	nand (gm_n4471, gm_n383, in_21, in_20, gm_n4470);
	nand (gm_n4472, gm_n4471, gm_n4469, gm_n4467);
	nor (gm_n4473, gm_n4458, gm_n4224, gm_n4222, gm_n4472, gm_n4465);
	nand (gm_n4474, gm_n61, gm_n73, in_12, gm_n487, gm_n79);
	nor (gm_n4475, gm_n496, gm_n72, gm_n85, gm_n4474);
	nor (gm_n4476, gm_n287, gm_n358, in_13, gm_n350);
	and (gm_n4477, gm_n122, in_21, in_17, gm_n4476, gm_n254);
	or (gm_n4478, gm_n256, gm_n461, gm_n76, gm_n589, gm_n349);
	nor (gm_n4479, gm_n479, gm_n72, gm_n55, gm_n4478);
	nor (gm_n4480, gm_n4479, gm_n4477, gm_n4475);
	or (gm_n4481, gm_n155, in_16, in_12, gm_n1324, gm_n276);
	nor (gm_n4482, gm_n781, gm_n72, in_20, gm_n4481);
	nand (gm_n4483, gm_n392, gm_n233, in_15, gm_n3368, gm_n394);
	nor (gm_n4484, gm_n72, in_20, in_19, gm_n4483);
	or (gm_n4485, gm_n257, in_13, gm_n62, gm_n502, gm_n359);
	nor (gm_n4486, gm_n441, gm_n72, in_17, gm_n4485, gm_n662);
	nor (gm_n4487, gm_n4486, gm_n4484, gm_n4482);
	nand (gm_n4488, gm_n4473, gm_n4220, gm_n4218, gm_n4487, gm_n4480);
	nor (gm_n4489, gm_n90, in_10, in_9, gm_n2402, gm_n207);
	nand (gm_n4490, gm_n243, gm_n166, gm_n119, gm_n4489);
	nand (gm_n4491, gm_n110, in_13, gm_n62, gm_n341, gm_n185);
	or (gm_n4492, gm_n183, gm_n72, gm_n55, gm_n4491, gm_n328);
	nor (gm_n4493, gm_n190, in_16, gm_n59, gm_n3006, gm_n227);
	nand (gm_n4494, gm_n113, gm_n72, in_20, gm_n4493);
	nand (gm_n4495, gm_n4494, gm_n4492, gm_n4490);
	nor (gm_n4496, gm_n514, in_13, gm_n62, gm_n596, gm_n818);
	nand (gm_n4497, gm_n254, in_21, in_17, gm_n4496, gm_n1076);
	nor (gm_n4498, gm_n274, gm_n193, gm_n60, gm_n1716, gm_n485);
	nand (gm_n4499, in_21, gm_n85, gm_n56, gm_n4498);
	nor (gm_n4500, gm_n442, gm_n76, gm_n62, gm_n621, gm_n502);
	nand (gm_n4501, gm_n327, in_21, gm_n55, gm_n4500, gm_n595);
	nand (gm_n4502, gm_n4501, gm_n4499, gm_n4497);
	nor (gm_n4503, gm_n4488, gm_n4216, gm_n4214, gm_n4502, gm_n4495);
	and (gm_n4504, gm_n523, gm_n72, in_17, gm_n3086, gm_n311);
	nand (gm_n4505, gm_n143, gm_n60, gm_n94, gm_n869, gm_n455);
	nor (gm_n4506, gm_n72, gm_n85, in_19, gm_n4505, gm_n447);
	nand (gm_n4507, gm_n595, in_13, gm_n62, gm_n875, gm_n402);
	nor (gm_n4508, gm_n312, gm_n72, in_17, gm_n4507);
	nor (gm_n4509, gm_n4508, gm_n4506, gm_n4504);
	or (gm_n4510, gm_n643, gm_n60, gm_n63, gm_n770, gm_n541);
	nor (gm_n4511, in_21, gm_n85, gm_n56, gm_n4510, gm_n269);
	nor (gm_n4512, gm_n202, gm_n115, gm_n94, gm_n223);
	nand (gm_n4513, gm_n392, gm_n56, in_15, gm_n4512, gm_n379);
	nor (gm_n4514, gm_n4513, in_21, gm_n85);
	or (gm_n4515, gm_n1331, gm_n213, in_15, gm_n633, gm_n399);
	nor (gm_n4516, in_21, gm_n85, in_19, gm_n4515);
	nor (gm_n4517, gm_n4516, gm_n4514, gm_n4511);
	nand (gm_n4518, gm_n4503, gm_n4212, gm_n4210, gm_n4517, gm_n4509);
	nor (gm_n4519, gm_n667, gm_n76, in_9, gm_n359, gm_n461);
	nand (gm_n4520, gm_n523, in_21, in_17, gm_n4519, gm_n311);
	nor (gm_n4521, gm_n514, in_13, gm_n62, gm_n808, gm_n184);
	nand (gm_n4522, gm_n311, in_21, in_17, gm_n4521);
	nor (gm_n4523, gm_n213, gm_n73, gm_n59, gm_n1324, gm_n354);
	nand (gm_n4524, gm_n296, in_21, in_20, gm_n4523);
	nand (gm_n4525, gm_n4524, gm_n4522, gm_n4520);
	nor (gm_n4526, gm_n662, in_13, in_9, gm_n3660, gm_n480);
	nand (gm_n4527, gm_n102, in_21, in_17, gm_n4526);
	nor (gm_n4528, gm_n168, gm_n60, in_11, gm_n2690, gm_n240);
	nand (gm_n4529, in_21, gm_n85, gm_n56, gm_n4528, gm_n268);
	nor (gm_n4530, gm_n76, gm_n62, gm_n94, gm_n981, gm_n442);
	nand (gm_n4531, gm_n104, gm_n72, in_17, gm_n4530, gm_n206);
	nand (gm_n4532, gm_n4531, gm_n4529, gm_n4527);
	nor (gm_n4533, gm_n4518, gm_n4209, gm_n4207, gm_n4532, gm_n4525);
	and (gm_n4534, gm_n61, in_16, gm_n59, gm_n1186, gm_n79);
	nand (gm_n4535, gm_n57, in_21, gm_n85, gm_n4534);
	nor (gm_n4536, gm_n514, in_13, in_9, gm_n743, gm_n344);
	nand (gm_n4537, gm_n206, in_21, gm_n55, gm_n4536, gm_n1076);
	nand (gm_n4538, gm_n311, in_21, gm_n55, gm_n2869, gm_n405);
	nand (gm_n4539, gm_n4535, gm_n4533, gm_n4205, gm_n4538, gm_n4537);
	and (gm_n4540, gm_n339, in_13, gm_n62, gm_n3679, gm_n402);
	nand (gm_n4541, gm_n311, gm_n72, gm_n55, gm_n4540);
	and (gm_n4542, gm_n64, gm_n73, in_12, gm_n1135, gm_n949);
	nand (gm_n4543, gm_n495, gm_n72, gm_n85, gm_n4542);
	nor (gm_n4544, gm_n158, gm_n73, gm_n59, gm_n1052, gm_n220);
	nand (gm_n4545, gm_n138, in_21, gm_n85, gm_n4544);
	nand (gm_n4546, gm_n4545, gm_n4543, gm_n4541);
	nand (gm_n4547, gm_n90, gm_n78, in_9, gm_n1841, gm_n1158);
	nor (gm_n4548, gm_n132, gm_n130, gm_n119, gm_n4547);
	nor (out_11, gm_n4546, gm_n4539, gm_n4204, gm_n4548);
	nand (gm_n4550, gm_n268, gm_n233, gm_n60, gm_n3041, gm_n1398);
	nor (gm_n4551, in_21, gm_n85, in_19, gm_n4550);
	nor (gm_n4552, gm_n90, in_10, gm_n62, gm_n399, gm_n207);
	nand (gm_n4553, gm_n436, gm_n243, in_18, gm_n4552);
	nand (gm_n4554, gm_n107, gm_n76, in_9, gm_n314, gm_n187);
	nor (gm_n4555, gm_n103, gm_n72, in_17, gm_n4554, gm_n375);
	nor (gm_n4556, gm_n184, in_21, gm_n55, gm_n1679, gm_n388);
	nor (gm_n4557, gm_n159, gm_n158, in_15, gm_n1519, gm_n269);
	nand (gm_n4558, in_21, gm_n85, gm_n56, gm_n4557);
	and (gm_n4559, gm_n1614, gm_n131, gm_n90, gm_n1120, gm_n713);
	nand (gm_n4560, gm_n4559, gm_n199, in_18);
	and (gm_n4561, gm_n60, gm_n90, in_13, t_7, gm_n73);
	and (gm_n4562, gm_n697, in_21, gm_n85, gm_n4561);
	or (gm_n4563, gm_n274, in_16, in_12, gm_n3382, gm_n385);
	nor (gm_n4564, gm_n912, in_21, gm_n85, gm_n4563);
	nor (gm_n4565, gm_n159, gm_n190, gm_n60, gm_n1751, gm_n293);
	nand (gm_n4566, gm_n72, in_20, gm_n56, gm_n4565);
	and (gm_n4567, gm_n222, in_16, in_12, gm_n1416, gm_n949);
	nand (gm_n4568, gm_n383, in_21, gm_n85, gm_n4567);
	or (gm_n4569, gm_n90, gm_n78, gm_n62, gm_n657, gm_n467);
	nor (gm_n4570, gm_n368, gm_n841, gm_n119, gm_n4569);
	or (gm_n4571, gm_n158, gm_n60, in_8, gm_n2690, gm_n168);
	nor (gm_n4572, gm_n72, gm_n85, in_19, gm_n4571, gm_n269);
	nor (gm_n4573, gm_n239, gm_n60, in_11, gm_n2017, gm_n643);
	nand (gm_n4574, gm_n72, in_20, in_19, gm_n4573, gm_n1101);
	and (gm_n4575, in_14, in_10, gm_n62, gm_n946, gm_n713);
	nand (gm_n4576, gm_n348, gm_n323, in_18, gm_n4575);
	or (gm_n4577, gm_n259, gm_n247, in_13, gm_n406);
	nor (gm_n4578, gm_n105, gm_n72, in_17, gm_n4577, gm_n183);
	and (gm_n4579, gm_n200, gm_n146, gm_n119, gm_n236);
	and (gm_n4580, gm_n233, gm_n73, gm_n59, gm_n1147, gm_n221);
	nand (gm_n4581, gm_n179, gm_n72, in_20, gm_n4580);
	nor (gm_n4582, gm_n190, in_16, gm_n59, gm_n2080, gm_n152);
	nand (gm_n4583, gm_n138, in_21, gm_n85, gm_n4582);
	or (gm_n4584, gm_n667, gm_n76, in_9, gm_n743, gm_n406);
	nor (gm_n4585, gm_n105, in_21, gm_n55, gm_n4584, gm_n620);
	nand (gm_n4586, gm_n323, gm_n171, in_14, gm_n3818, gm_n713);
	nor (gm_n4587, gm_n4586, gm_n165, gm_n119);
	nor (gm_n4588, gm_n259, gm_n247, gm_n76, gm_n431);
	nand (gm_n4589, gm_n104, gm_n72, in_17, gm_n4588, gm_n206);
	nor (gm_n4590, gm_n76, gm_n59, gm_n63, gm_n981, gm_n977);
	nand (gm_n4591, gm_n120, in_21, in_17, gm_n4590, gm_n255);
	nand (gm_n4592, in_14, in_10, in_9, gm_n1501, gm_n600);
	nor (gm_n4593, gm_n1989, gm_n165, in_18, gm_n4592);
	nand (gm_n4594, gm_n214, gm_n73, gm_n59, gm_n1841, gm_n303);
	nor (gm_n4595, gm_n912, gm_n72, gm_n85, gm_n4594);
	and (gm_n4596, gm_n90, in_10, in_9, gm_n991, gm_n1158);
	nand (gm_n4597, gm_n166, gm_n164, gm_n119, gm_n4596);
	and (gm_n4598, gm_n110, in_13, in_9, gm_n341, gm_n314);
	nand (gm_n4599, gm_n339, in_21, gm_n55, gm_n4598, gm_n373);
	nand (gm_n4600, gm_n828, in_14, gm_n78, gm_n829, gm_n1011);
	nor (gm_n4601, gm_n246, gm_n244, gm_n119, gm_n4600);
	nand (gm_n4602, gm_n339, gm_n76, in_9, gm_n1611, gm_n788);
	nor (gm_n4603, gm_n183, in_21, gm_n55, gm_n4602);
	nor (gm_n4604, gm_n115, gm_n73, gm_n59, gm_n765, gm_n276);
	nand (gm_n4605, gm_n113, in_21, gm_n85, gm_n4604);
	nor (gm_n4606, gm_n90, in_10, gm_n62, gm_n4088, gm_n369);
	nand (gm_n4607, gm_n436, gm_n199, gm_n119, gm_n4606);
	or (gm_n4608, gm_n514, in_13, gm_n62, gm_n1583, gm_n609);
	nor (gm_n4609, gm_n183, in_21, in_17, gm_n4608, gm_n313);
	nand (gm_n4610, gm_n143, in_16, gm_n59, gm_n685, gm_n303);
	nor (gm_n4611, gm_n262, in_21, in_20, gm_n4610);
	nor (gm_n4612, gm_n133, in_14, in_10, gm_n526, gm_n247);
	nand (gm_n4613, gm_n323, gm_n146, gm_n119, gm_n4612);
	not (gm_n4614, gm_n919);
	nor (gm_n4615, gm_n293, gm_n274, in_15, gm_n4614, gm_n760);
	nand (gm_n4616, gm_n72, gm_n85, in_19, gm_n4615);
	or (gm_n4617, gm_n227, in_16, gm_n59, gm_n2002, gm_n115);
	nor (gm_n4618, gm_n912, gm_n72, in_20, gm_n4617);
	or (gm_n4619, gm_n158, in_12, gm_n94, gm_n939, gm_n152);
	nor (gm_n4620, gm_n72, gm_n85, in_16, gm_n4619, gm_n262);
	nor (gm_n4621, gm_n190, in_16, in_12, gm_n1923, gm_n354);
	nand (gm_n4622, gm_n697, gm_n72, in_20, gm_n4621);
	nor (gm_n4623, gm_n95, gm_n90, gm_n78, gm_n362, gm_n259);
	nand (gm_n4624, gm_n200, gm_n86, in_18, gm_n4623);
	nor (gm_n4625, gm_n115, gm_n73, in_12, gm_n1052, gm_n385);
	nand (gm_n4626, gm_n57, gm_n72, gm_n85, gm_n4625);
	nor (gm_n4627, gm_n358, in_13, gm_n62, gm_n796, gm_n667);
	nand (gm_n4628, gm_n104, in_21, gm_n55, gm_n4627, gm_n120);
	nor (gm_n4629, gm_n213, in_16, in_12, gm_n632, gm_n385);
	nand (gm_n4630, gm_n57, in_21, in_20, gm_n4629);
	nand (gm_n4631, gm_n4626, gm_n4624, gm_n4622, gm_n4630, gm_n4628);
	nor (gm_n4632, gm_n358, in_13, gm_n62, gm_n4437, gm_n328);
	nand (gm_n4633, gm_n102, gm_n72, in_17, gm_n4632);
	nor (gm_n4634, gm_n213, in_16, gm_n59, gm_n815, gm_n220);
	nand (gm_n4635, gm_n495, in_21, gm_n85, gm_n4634);
	nor (gm_n4636, gm_n193, gm_n190, in_15, gm_n2244, gm_n269);
	nand (gm_n4637, in_21, in_20, in_19, gm_n4636);
	nand (gm_n4638, gm_n4637, gm_n4635, gm_n4633);
	nor (gm_n4639, gm_n147, gm_n90, in_10, gm_n438, gm_n414);
	nand (gm_n4640, gm_n436, gm_n348, in_18, gm_n4639);
	and (gm_n4641, gm_n77, gm_n73, gm_n59, gm_n1978, gm_n154);
	nand (gm_n4642, gm_n697, gm_n72, in_20, gm_n4641);
	and (gm_n4643, gm_n90, gm_n76, in_12, gm_n2860, gm_n222);
	nand (gm_n4644, gm_n243, gm_n88, gm_n119, gm_n4643);
	nand (gm_n4645, gm_n4644, gm_n4642, gm_n4640);
	nor (gm_n4646, gm_n4631, gm_n4620, gm_n4618, gm_n4645, gm_n4638);
	nand (gm_n4647, gm_n143, gm_n75, in_15, gm_n869, gm_n411);
	nor (gm_n4648, gm_n72, in_20, gm_n56, gm_n4647);
	or (gm_n4649, gm_n257, gm_n76, in_9, gm_n462, gm_n596);
	nor (gm_n4650, gm_n388, in_21, in_17, gm_n4649, gm_n662);
	or (gm_n4651, gm_n99, in_14, in_10, gm_n438, gm_n362);
	nor (gm_n4652, gm_n1989, gm_n165, in_18, gm_n4651);
	nor (gm_n4653, gm_n4652, gm_n4650, gm_n4648);
	nand (gm_n4654, gm_n76, in_9, gm_n94, gm_n579, gm_n170);
	nor (gm_n4655, gm_n103, in_21, gm_n55, gm_n4654, gm_n662);
	or (gm_n4656, gm_n133, in_14, in_10, gm_n370, gm_n259);
	nor (gm_n4657, gm_n244, gm_n841, gm_n119, gm_n4656);
	or (gm_n4658, gm_n257, in_13, gm_n62, gm_n432, gm_n344);
	nor (gm_n4659, gm_n479, in_21, in_17, gm_n4658, gm_n375);
	nor (gm_n4660, gm_n4659, gm_n4657, gm_n4655);
	nand (gm_n4661, gm_n4646, gm_n4616, gm_n4613, gm_n4660, gm_n4653);
	nor (gm_n4662, gm_n193, gm_n297, in_15, gm_n1965, gm_n485);
	nand (gm_n4663, gm_n72, gm_n85, gm_n56, gm_n4662);
	and (gm_n4664, gm_n90, gm_n78, gm_n62, gm_n4011, gm_n600);
	nand (gm_n4665, gm_n367, gm_n166, in_18, gm_n4664);
	nor (gm_n4666, gm_n393, gm_n56, gm_n60, gm_n760, gm_n590);
	nand (gm_n4667, gm_n4666, gm_n72, gm_n85);
	nand (gm_n4668, gm_n4667, gm_n4665, gm_n4663);
	nor (gm_n4669, gm_n431, gm_n76, in_9, gm_n359, gm_n344);
	nand (gm_n4670, gm_n102, gm_n72, in_17, gm_n4669, gm_n339);
	nor (gm_n4671, gm_n807, in_14, in_10, gm_n775, gm_n438);
	nand (gm_n4672, gm_n243, gm_n131, in_18, gm_n4671);
	nor (gm_n4673, gm_n251, gm_n213, gm_n60, gm_n764, gm_n269);
	nand (gm_n4674, gm_n72, gm_n85, in_19, gm_n4673);
	nand (gm_n4675, gm_n4674, gm_n4672, gm_n4670);
	nor (gm_n4676, gm_n4661, gm_n4611, gm_n4609, gm_n4675, gm_n4668);
	nand (gm_n4677, gm_n214, in_16, gm_n59, gm_n919, gm_n571);
	nor (gm_n4678, gm_n384, in_21, gm_n85, gm_n4677);
	or (gm_n4679, gm_n358, in_13, gm_n62, gm_n481, gm_n430);
	nor (gm_n4680, gm_n256, gm_n72, gm_n55, gm_n4679, gm_n374);
	nand (gm_n4681, gm_n76, in_9, gm_n94, gm_n1692, gm_n185);
	nor (gm_n4682, gm_n121, gm_n72, gm_n55, gm_n4681, gm_n388);
	nor (gm_n4683, gm_n4682, gm_n4680, gm_n4678);
	nand (gm_n4684, gm_n76, in_9, in_8, gm_n1929, gm_n314);
	nor (gm_n4685, gm_n184, in_21, in_17, gm_n4684, gm_n479);
	nor (gm_n4686, gm_n620, gm_n72, in_17, gm_n2758, gm_n328);
	or (gm_n4687, gm_n159, gm_n155, gm_n60, gm_n3440, gm_n191);
	nor (gm_n4688, in_21, in_20, gm_n56, gm_n4687);
	nor (gm_n4689, gm_n4688, gm_n4686, gm_n4685);
	nand (gm_n4690, gm_n4676, gm_n4607, gm_n4605, gm_n4689, gm_n4683);
	nor (gm_n4691, gm_n193, gm_n191, in_15, gm_n1319, gm_n213);
	nand (gm_n4692, gm_n72, gm_n85, in_19, gm_n4691);
	nand (gm_n4693, gm_n122, gm_n72, gm_n55, gm_n3139, gm_n174);
	nor (gm_n4694, gm_n213, in_16, in_12, gm_n2221, gm_n319);
	nand (gm_n4695, gm_n296, in_21, gm_n85, gm_n4694);
	nand (gm_n4696, gm_n4695, gm_n4693, gm_n4692);
	nor (gm_n4697, gm_n158, gm_n59, gm_n94, gm_n2769, gm_n152);
	nand (gm_n4698, in_21, in_20, in_16, gm_n4697, gm_n179);
	nor (gm_n4699, gm_n159, in_15, gm_n63, gm_n2017, gm_n770);
	nand (gm_n4700, gm_n72, in_20, in_19, gm_n4699, gm_n379);
	and (gm_n4701, gm_n123, in_13, in_9, gm_n1049, gm_n126);
	nand (gm_n4702, gm_n206, in_21, gm_n55, gm_n4701, gm_n255);
	nand (gm_n4703, gm_n4702, gm_n4700, gm_n4698);
	nor (gm_n4704, gm_n4690, gm_n4603, gm_n4601, gm_n4703, gm_n4696);
	nand (gm_n4705, gm_n61, gm_n73, gm_n59, gm_n919, gm_n64);
	nor (gm_n4706, gm_n384, in_21, in_20, gm_n4705);
	or (gm_n4707, gm_n609, gm_n76, gm_n62, gm_n743, gm_n442);
	nor (gm_n4708, gm_n662, gm_n72, gm_n55, gm_n4707, gm_n374);
	or (gm_n4709, gm_n393, gm_n115, gm_n60, gm_n2421, gm_n643);
	nor (gm_n4710, in_21, in_20, in_19, gm_n4709);
	nor (gm_n4711, gm_n4710, gm_n4708, gm_n4706);
	or (gm_n4712, gm_n121, gm_n76, gm_n62, gm_n1884, gm_n442);
	nor (gm_n4713, gm_n441, in_21, in_17, gm_n4712);
	or (gm_n4714, gm_n514, gm_n76, gm_n62, gm_n359, gm_n596);
	nor (gm_n4715, gm_n441, gm_n72, in_17, gm_n4714, gm_n662);
	or (gm_n4716, gm_n274, in_16, gm_n59, gm_n2080, gm_n354);
	nor (gm_n4717, gm_n781, in_21, gm_n85, gm_n4716);
	nor (gm_n4718, gm_n4717, gm_n4715, gm_n4713);
	nand (gm_n4719, gm_n4704, gm_n4599, gm_n4597, gm_n4718, gm_n4711);
	and (gm_n4720, gm_n392, gm_n64, gm_n60, gm_n1095, gm_n394);
	nand (gm_n4721, gm_n72, in_20, gm_n56, gm_n4720);
	nand (gm_n4722, gm_n120, gm_n72, gm_n55, gm_n2864, gm_n595);
	nor (gm_n4723, gm_n514, gm_n76, in_9, gm_n597, gm_n463);
	nand (gm_n4724, gm_n104, gm_n72, in_17, gm_n4723, gm_n174);
	nand (gm_n4725, gm_n4724, gm_n4722, gm_n4721);
	and (gm_n4726, gm_n186, in_13, in_9, gm_n340, gm_n316);
	nand (gm_n4727, gm_n102, in_21, gm_n55, gm_n4726, gm_n339);
	nor (gm_n4728, gm_n207, gm_n194, gm_n90, gm_n283, gm_n238);
	nand (gm_n4729, gm_n367, gm_n200, in_18, gm_n4728);
	nor (gm_n4730, gm_n263, in_16, in_12, gm_n695, gm_n354);
	nand (gm_n4731, gm_n138, in_21, in_20, gm_n4730);
	nand (gm_n4732, gm_n4731, gm_n4729, gm_n4727);
	nor (gm_n4733, gm_n4719, gm_n4595, gm_n4593, gm_n4732, gm_n4725);
	nand (gm_n4734, gm_n222, gm_n73, in_12, gm_n2646, gm_n571);
	nor (gm_n4735, gm_n262, gm_n72, in_20, gm_n4734);
	or (gm_n4736, gm_n207, gm_n90, gm_n78, gm_n438, gm_n350);
	nor (gm_n4737, gm_n89, gm_n87, in_18, gm_n4736);
	or (gm_n4738, gm_n430, in_13, in_9, gm_n503, gm_n431);
	nor (gm_n4739, gm_n479, gm_n72, in_17, gm_n4738, gm_n256);
	nor (gm_n4740, gm_n4739, gm_n4737, gm_n4735);
	or (gm_n4741, gm_n461, in_13, in_9, gm_n597, gm_n430);
	nor (gm_n4742, gm_n183, gm_n72, gm_n55, gm_n4741, gm_n184);
	and (gm_n4743, gm_n102, gm_n72, in_17, gm_n1924, gm_n1076);
	nand (gm_n4744, in_14, gm_n78, in_9, gm_n2497, gm_n1158);
	nor (gm_n4745, gm_n244, gm_n841, gm_n119, gm_n4744);
	nor (gm_n4746, gm_n4745, gm_n4743, gm_n4742);
	nand (gm_n4747, gm_n4733, gm_n4591, gm_n4589, gm_n4746, gm_n4740);
	nor (gm_n4748, gm_n491, gm_n92, in_10, gm_n775);
	nand (gm_n4749, gm_n102, in_21, gm_n55, gm_n4748, gm_n595);
	nand (gm_n4750, gm_n131, gm_n86, gm_n119, gm_n1055);
	nor (gm_n4751, gm_n148, gm_n90, gm_n78, gm_n362, gm_n259);
	nand (gm_n4752, gm_n245, gm_n243, gm_n119, gm_n4751);
	nand (gm_n4753, gm_n4752, gm_n4750, gm_n4749);
	and (gm_n4754, gm_n222, in_12, gm_n94, gm_n275, gm_n1379);
	nand (gm_n4755, in_21, gm_n85, gm_n73, gm_n4754, gm_n179);
	nor (gm_n4756, in_13, gm_n62, gm_n94, gm_n406, gm_n161);
	nand (gm_n4757, gm_n120, gm_n72, in_17, gm_n4756, gm_n255);
	nor (gm_n4758, gm_n430, gm_n76, gm_n62, gm_n432, gm_n257);
	nand (gm_n4759, gm_n122, gm_n72, gm_n55, gm_n4758, gm_n174);
	nand (gm_n4760, gm_n4759, gm_n4757, gm_n4755);
	nor (gm_n4761, gm_n4747, gm_n4587, gm_n4585, gm_n4760, gm_n4753);
	nand (gm_n4762, gm_n143, gm_n75, gm_n60, gm_n1416, gm_n392);
	nor (gm_n4763, in_21, in_20, gm_n56, gm_n4762);
	nand (gm_n4764, gm_n192, gm_n154, in_15, gm_n486, gm_n216);
	nor (gm_n4765, gm_n72, in_20, in_19, gm_n4764);
	or (gm_n4766, gm_n447, gm_n155, gm_n60, gm_n1319, gm_n633);
	nor (gm_n4767, in_21, in_20, in_19, gm_n4766);
	nor (gm_n4768, gm_n4767, gm_n4765, gm_n4763);
	or (gm_n4769, gm_n596, gm_n76, in_9, gm_n988, gm_n442);
	nor (gm_n4770, gm_n184, in_21, in_17, gm_n4769, gm_n388);
	nand (gm_n4771, in_14, in_10, gm_n62, gm_n3063, gm_n600);
	nor (gm_n4772, gm_n244, gm_n841, in_18, gm_n4771);
	nand (gm_n4773, gm_n125, in_13, gm_n62, gm_n340, gm_n126);
	nor (gm_n4774, gm_n620, in_21, gm_n55, gm_n4773, gm_n375);
	nor (gm_n4775, gm_n4774, gm_n4772, gm_n4770);
	nand (gm_n4776, gm_n4761, gm_n4583, gm_n4581, gm_n4775, gm_n4768);
	nor (gm_n4777, gm_n115, in_16, gm_n59, gm_n1191, gm_n354);
	nand (gm_n4778, gm_n383, gm_n72, gm_n85, gm_n4777);
	nor (gm_n4779, gm_n609, gm_n76, in_9, gm_n481, gm_n406);
	nand (gm_n4780, gm_n120, in_21, gm_n55, gm_n4779, gm_n1076);
	or (gm_n4781, gm_n388, in_21, in_17, gm_n3356, gm_n313);
	nand (gm_n4782, gm_n4781, gm_n4780, gm_n4778);
	nor (gm_n4783, gm_n193, gm_n155, gm_n60, gm_n821, gm_n1331);
	nand (gm_n4784, in_21, in_20, in_19, gm_n4783);
	nor (gm_n4785, gm_n514, gm_n76, in_9, gm_n463, gm_n432);
	nand (gm_n4786, gm_n254, in_21, gm_n55, gm_n4785, gm_n405);
	nor (gm_n4787, gm_n257, gm_n76, in_9, gm_n502, gm_n359);
	nand (gm_n4788, gm_n174, gm_n72, gm_n55, gm_n4787, gm_n339);
	nand (gm_n4789, gm_n4788, gm_n4786, gm_n4784);
	nor (gm_n4790, gm_n4776, gm_n4579, gm_n4578, gm_n4789, gm_n4782);
	and (gm_n4791, gm_n131, gm_n129, gm_n119, gm_n4643);
	nand (gm_n4792, gm_n448, gm_n154, in_15, gm_n2065, gm_n545);
	nor (gm_n4793, in_21, gm_n85, gm_n56, gm_n4792);
	or (gm_n4794, gm_n149, gm_n90, in_10, gm_n467, gm_n370);
	nor (gm_n4795, gm_n1989, gm_n130, gm_n119, gm_n4794);
	nor (gm_n4796, gm_n4795, gm_n4793, gm_n4791);
	and (gm_n4797, gm_n436, gm_n129, gm_n119, gm_n1499);
	or (gm_n4798, gm_n431, gm_n149, in_13, gm_n438);
	nor (gm_n4799, gm_n105, gm_n72, gm_n55, gm_n4798, gm_n388);
	or (gm_n4800, in_14, gm_n78, in_9, gm_n1475, gm_n362);
	nor (gm_n4801, gm_n167, gm_n87, in_18, gm_n4800);
	nor (gm_n4802, gm_n4801, gm_n4799, gm_n4797);
	nand (gm_n4803, gm_n4790, gm_n4576, gm_n4574, gm_n4802, gm_n4796);
	nor (gm_n4804, gm_n257, in_13, in_9, gm_n443, gm_n359);
	nand (gm_n4805, gm_n102, gm_n72, in_17, gm_n4804, gm_n1076);
	nor (gm_n4806, gm_n168, gm_n190, gm_n60, gm_n1150, gm_n485);
	nand (gm_n4807, in_21, gm_n85, gm_n56, gm_n4806);
	nor (gm_n4808, gm_n95, gm_n90, in_10, gm_n259, gm_n147);
	nand (gm_n4809, gm_n245, gm_n243, gm_n119, gm_n4808);
	nand (gm_n4810, gm_n4809, gm_n4807, gm_n4805);
	nor (gm_n4811, gm_n358, in_13, in_9, gm_n359, gm_n667);
	nand (gm_n4812, gm_n254, gm_n72, gm_n55, gm_n4811, gm_n255);
	nor (gm_n4813, gm_n193, gm_n158, in_15, gm_n849, gm_n1331);
	nand (gm_n4814, gm_n72, gm_n85, in_19, gm_n4813);
	and (gm_n4815, gm_n64, in_16, in_12, gm_n265, gm_n77);
	nand (gm_n4816, gm_n138, gm_n72, gm_n85, gm_n4815);
	nand (gm_n4817, gm_n4816, gm_n4814, gm_n4812);
	nor (gm_n4818, gm_n4803, gm_n4572, gm_n4570, gm_n4817, gm_n4810);
	and (gm_n4819, gm_n104, in_21, gm_n55, gm_n1341, gm_n174);
	or (gm_n4820, gm_n191, gm_n155, gm_n60, gm_n821, gm_n760);
	nor (gm_n4821, in_21, in_20, gm_n56, gm_n4820);
	nand (gm_n4822, gm_n90, gm_n78, gm_n62, gm_n946, gm_n91);
	nor (gm_n4823, gm_n167, gm_n87, in_18, gm_n4822);
	nor (gm_n4824, gm_n4823, gm_n4821, gm_n4819);
	or (gm_n4825, gm_n596, gm_n76, in_9, gm_n503, gm_n480);
	nor (gm_n4826, gm_n105, in_21, gm_n55, gm_n4825, gm_n312);
	or (gm_n4827, gm_n207, in_14, in_10, gm_n350, gm_n349);
	nor (gm_n4828, gm_n531, gm_n246, in_18, gm_n4827);
	or (gm_n4829, gm_n238, gm_n194, in_14, gm_n369, gm_n283);
	nor (gm_n4830, gm_n165, gm_n132, gm_n119, gm_n4829);
	nor (gm_n4831, gm_n4830, gm_n4828, gm_n4826);
	nand (gm_n4832, gm_n4818, gm_n4568, gm_n4566, gm_n4831, gm_n4824);
	nor (gm_n4833, gm_n158, in_16, gm_n59, gm_n1223, gm_n152);
	nand (gm_n4834, gm_n495, in_21, gm_n85, gm_n4833);
	nand (gm_n4835, gm_n79, in_13, in_12, gm_n547);
	or (gm_n4836, gm_n105, gm_n72, in_17, gm_n4835, gm_n312);
	nor (gm_n4837, gm_n297, gm_n73, gm_n59, gm_n1223, gm_n385);
	nand (gm_n4838, gm_n383, in_21, gm_n85, gm_n4837);
	nand (gm_n4839, gm_n4838, gm_n4836, gm_n4834);
	nor (gm_n4840, gm_n362, in_14, in_10, gm_n775, gm_n491);
	nand (gm_n4841, gm_n243, gm_n166, in_18, gm_n4840);
	nor (gm_n4842, gm_n190, gm_n73, gm_n59, gm_n2963, gm_n319);
	nand (gm_n4843, gm_n495, in_21, in_20, gm_n4842);
	and (gm_n4844, gm_n392, gm_n60, gm_n63, gm_n1615, gm_n602);
	nand (gm_n4845, gm_n72, in_20, gm_n56, gm_n4844, gm_n75);
	nand (gm_n4846, gm_n4845, gm_n4843, gm_n4841);
	nor (gm_n4847, gm_n4832, gm_n4564, gm_n4562, gm_n4846, gm_n4839);
	and (gm_n4848, gm_n523, in_21, gm_n55, gm_n1171, gm_n311);
	nand (gm_n4849, in_10, gm_n62, in_8, gm_n756, gm_n91);
	nor (gm_n4850, gm_n87, in_18, in_14, gm_n4849, gm_n841);
	or (gm_n4851, gm_n431, gm_n99, gm_n76, gm_n370, gm_n328);
	nor (gm_n4852, gm_n183, gm_n72, gm_n55, gm_n4851);
	nor (gm_n4853, gm_n4852, gm_n4850, gm_n4848);
	and (gm_n4854, gm_n104, gm_n72, in_17, gm_n2861, gm_n311);
	nand (gm_n4855, in_13, in_9, gm_n94, gm_n576, gm_n185);
	nor (gm_n4856, gm_n374, gm_n72, gm_n55, gm_n4855, gm_n375);
	or (gm_n4857, gm_n485, gm_n155, gm_n60, gm_n648, gm_n633);
	nor (gm_n4858, gm_n72, gm_n85, gm_n56, gm_n4857);
	nor (gm_n4859, gm_n4858, gm_n4856, gm_n4854);
	nand (gm_n4860, gm_n4847, gm_n4560, gm_n4558, gm_n4859, gm_n4853);
	nor (gm_n4861, gm_n667, in_13, gm_n62, gm_n597, gm_n461);
	nand (gm_n4862, gm_n327, gm_n72, gm_n55, gm_n4861, gm_n339);
	nor (gm_n4863, gm_n461, gm_n76, in_9, gm_n988, gm_n502);
	nand (gm_n4864, gm_n122, gm_n72, gm_n55, gm_n4863, gm_n373);
	nor (gm_n4865, gm_n667, in_13, in_9, gm_n743, gm_n257);
	nand (gm_n4866, gm_n122, gm_n72, gm_n55, gm_n4865, gm_n373);
	nand (gm_n4867, gm_n4866, gm_n4864, gm_n4862);
	nor (gm_n4868, gm_n345, gm_n76, gm_n62, gm_n502, gm_n442);
	nand (gm_n4869, gm_n523, in_21, gm_n55, gm_n4868, gm_n254);
	nand (gm_n4870, gm_n206, gm_n72, gm_n55, gm_n3061, gm_n1076);
	nor (gm_n4871, in_14, gm_n78, gm_n62, gm_n2008, gm_n92);
	nand (gm_n4872, gm_n243, gm_n166, gm_n119, gm_n4871);
	nand (gm_n4873, gm_n4872, gm_n4870, gm_n4869);
	nor (gm_n4874, gm_n4860, gm_n4556, gm_n4555, gm_n4873, gm_n4867);
	or (gm_n4875, gm_n103, gm_n72, gm_n55, gm_n1261, gm_n313);
	nor (gm_n4876, gm_n667, gm_n76, gm_n62, gm_n1583, gm_n406);
	nand (gm_n4877, gm_n104, gm_n72, gm_n55, gm_n4876, gm_n120);
	nor (gm_n4878, gm_n213, in_16, in_12, gm_n3099, gm_n319);
	nand (gm_n4879, gm_n138, gm_n72, gm_n85, gm_n4878);
	nand (gm_n4880, gm_n4875, gm_n4874, gm_n4553, gm_n4879, gm_n4877);
	and (gm_n4881, gm_n316, gm_n76, in_9, gm_n1049, gm_n340);
	nand (gm_n4882, gm_n174, gm_n72, in_17, gm_n4881, gm_n255);
	nor (gm_n4883, gm_n442, in_13, in_9, gm_n463, gm_n462);
	nand (gm_n4884, gm_n405, in_21, gm_n55, gm_n4883, gm_n327);
	nor (gm_n4885, gm_n90, in_10, gm_n62, gm_n1406, gm_n133);
	nand (gm_n4886, gm_n243, gm_n166, gm_n119, gm_n4885);
	nand (gm_n4887, gm_n4886, gm_n4884, gm_n4882);
	nand (gm_n4888, gm_n106, gm_n2193, in_13, gm_n995, gm_n523);
	nor (gm_n4889, gm_n620, in_21, in_17, gm_n4888);
	nor (out_12, gm_n4887, gm_n4880, gm_n4551, gm_n4889);
	or (gm_n4891, gm_n95, in_14, in_10, gm_n589, gm_n133);
	nor (gm_n4892, gm_n167, gm_n130, in_18, gm_n4891);
	nor (gm_n4893, gm_n1331, gm_n274, in_15, gm_n1173, gm_n643);
	nand (gm_n4894, in_21, gm_n85, in_19, gm_n4893);
	nand (gm_n4895, gm_n143, in_16, gm_n59, gm_n2070, gm_n949);
	nor (gm_n4896, gm_n496, in_21, gm_n85, gm_n4895);
	or (gm_n4897, gm_n227, gm_n73, gm_n59, gm_n2333, gm_n213);
	nor (gm_n4898, gm_n384, gm_n72, in_20, gm_n4897);
	and (gm_n4899, gm_n90, gm_n78, in_9, gm_n2712, gm_n1158);
	nand (gm_n4900, gm_n146, gm_n88, in_18, gm_n4899);
	and (gm_n4901, in_13, gm_n62, in_8, gm_n788, gm_n176);
	nand (gm_n4902, gm_n327, gm_n72, in_17, gm_n4901, gm_n595);
	or (gm_n4903, gm_n609, gm_n76, in_9, gm_n432, gm_n431);
	nor (gm_n4904, gm_n183, in_21, gm_n55, gm_n4903, gm_n121);
	nand (gm_n4905, gm_n107, in_10, gm_n62, gm_n532, gm_n110);
	nor (gm_n4906, gm_n87, in_18, in_14, gm_n4905, gm_n167);
	nor (gm_n4907, gm_n514, in_13, gm_n62, gm_n462, gm_n667);
	nand (gm_n4908, gm_n339, gm_n72, in_17, gm_n4907, gm_n373);
	nor (gm_n4909, gm_n152, gm_n73, gm_n59, gm_n1208, gm_n263);
	nand (gm_n4910, gm_n495, gm_n72, in_20, gm_n4909);
	nor (gm_n4911, gm_n479, gm_n72, gm_n55, gm_n4714, gm_n313);
	nor (gm_n4912, gm_n105, gm_n72, in_17, gm_n4104, gm_n620);
	nor (gm_n4913, gm_n297, gm_n74, in_15, gm_n760, gm_n562);
	nand (gm_n4914, in_21, gm_n85, in_19, gm_n4913);
	nor (gm_n4915, gm_n227, gm_n73, in_12, gm_n849, gm_n263);
	nand (gm_n4916, gm_n495, gm_n72, in_20, gm_n4915);
	or (gm_n4917, in_7, in_6, in_5, gm_n141, gm_n94);
	or (gm_n4918, gm_n159, gm_n74, gm_n60, gm_n4917, gm_n263);
	nor (gm_n4919, gm_n72, gm_n85, in_19, gm_n4918);
	or (gm_n4920, gm_n148, gm_n121, gm_n76, gm_n406, gm_n286);
	nor (gm_n4921, gm_n388, gm_n72, in_17, gm_n4920);
	and (gm_n4922, gm_n61, gm_n73, in_12, gm_n1501, gm_n264);
	nand (gm_n4923, gm_n296, in_21, in_20, gm_n4922);
	nor (gm_n4924, gm_n115, gm_n76, in_12, gm_n855);
	nand (gm_n4925, gm_n595, gm_n72, in_17, gm_n4924, gm_n373);
	and (gm_n4926, gm_n426, gm_n304, in_8);
	nand (gm_n4927, gm_n233, in_16, gm_n59, gm_n4926, gm_n221);
	nor (gm_n4928, gm_n912, gm_n72, in_20, gm_n4927);
	nand (gm_n4929, gm_n264, in_16, gm_n59, gm_n3368, gm_n949);
	nor (gm_n4930, gm_n912, in_21, gm_n85, gm_n4929);
	and (gm_n4931, gm_n110, gm_n76, in_9, gm_n314, gm_n186);
	nand (gm_n4932, gm_n122, gm_n72, in_17, gm_n4931, gm_n311);
	nor (gm_n4933, gm_n257, gm_n76, gm_n62, gm_n597, gm_n443);
	nand (gm_n4934, gm_n120, gm_n72, gm_n55, gm_n4933, gm_n405);
	or (gm_n4935, gm_n625, gm_n202, gm_n94);
	or (gm_n4936, gm_n114, gm_n73, in_12, gm_n4935, gm_n190);
	nor (gm_n4937, gm_n58, gm_n72, gm_n85, gm_n4936);
	and (gm_n4938, gm_n206, gm_n72, in_17, gm_n898, gm_n1076);
	nor (gm_n4939, gm_n148, gm_n90, gm_n78, gm_n589, gm_n362);
	nand (gm_n4940, gm_n806, gm_n129, in_18, gm_n4939);
	and (gm_n4941, gm_n392, in_15, in_11, gm_n1615, gm_n1144);
	nand (gm_n4942, gm_n72, gm_n85, gm_n56, gm_n4941, gm_n1101);
	nor (gm_n4943, gm_n467, in_10, gm_n62, gm_n1484);
	and (gm_n4944, gm_n523, gm_n72, gm_n55, gm_n4943, gm_n206);
	nand (gm_n4945, gm_n484, gm_n60, gm_n63, gm_n601, gm_n1614);
	nor (gm_n4946, in_21, gm_n85, gm_n56, gm_n4945, gm_n485);
	and (gm_n4947, gm_n126, gm_n76, in_9, gm_n341, gm_n579);
	nand (gm_n4948, gm_n120, in_21, gm_n55, gm_n4947, gm_n405);
	and (gm_n4949, gm_n171, gm_n60, gm_n63, gm_n449, gm_n176);
	nand (gm_n4950, gm_n72, in_20, gm_n56, gm_n4949, gm_n281);
	or (gm_n4951, gm_n184, in_13, in_12, gm_n705, gm_n274);
	nor (gm_n4952, gm_n441, in_21, gm_n55, gm_n4951);
	nand (gm_n4953, gm_n221, gm_n73, gm_n59, gm_n1970, gm_n222);
	nor (gm_n4954, gm_n139, gm_n72, in_20, gm_n4953);
	nor (gm_n4955, gm_n227, gm_n73, gm_n59, gm_n1689, gm_n115);
	nand (gm_n4956, gm_n138, in_21, gm_n85, gm_n4955);
	nor (gm_n4957, gm_n344, in_13, gm_n62, gm_n481, gm_n480);
	nand (gm_n4958, gm_n255, in_21, in_17, gm_n4957, gm_n327);
	or (gm_n4959, gm_n349, gm_n90, in_10, gm_n389, gm_n362);
	nor (gm_n4960, gm_n246, gm_n244, in_18, gm_n4959);
	or (gm_n4961, gm_n95, gm_n90, gm_n78, gm_n467, gm_n208);
	nor (gm_n4962, gm_n1989, gm_n130, gm_n119, gm_n4961);
	and (gm_n4963, gm_n545, gm_n60, gm_n63, gm_n602, gm_n576);
	nand (gm_n4964, in_21, gm_n85, gm_n56, gm_n4963, gm_n394);
	nor (gm_n4965, gm_n269, gm_n190, gm_n60, gm_n2244, gm_n764);
	nand (gm_n4966, gm_n72, in_20, in_19, gm_n4965);
	or (gm_n4967, gm_n572, gm_n201, gm_n94);
	nor (gm_n4968, gm_n190, gm_n73, in_12, gm_n4967, gm_n319);
	nand (gm_n4969, gm_n296, in_21, gm_n85, gm_n4968);
	nor (gm_n4970, gm_n274, in_16, gm_n59, gm_n1191, gm_n385);
	nand (gm_n4971, gm_n495, in_21, in_20, gm_n4970);
	nor (gm_n4972, gm_n213, gm_n73, in_12, gm_n2256, gm_n319);
	nand (gm_n4973, gm_n495, gm_n72, gm_n85, gm_n4972);
	nand (gm_n4974, gm_n4969, gm_n4966, gm_n4964, gm_n4973, gm_n4971);
	or (gm_n4975, gm_n228, gm_n201, gm_n94);
	nor (gm_n4976, gm_n213, gm_n73, in_12, gm_n4975, gm_n220);
	nand (gm_n4977, gm_n138, gm_n72, in_20, gm_n4976);
	nor (gm_n4978, in_13, gm_n62, in_8, gm_n939, gm_n257);
	nand (gm_n4979, gm_n311, gm_n72, in_17, gm_n4978, gm_n1076);
	nor (gm_n4980, gm_n76, in_12, in_11, gm_n271, gm_n270);
	nand (gm_n4981, gm_n174, gm_n72, gm_n55, gm_n4980, gm_n339);
	nand (gm_n4982, gm_n4981, gm_n4979, gm_n4977);
	nor (gm_n4983, gm_n461, gm_n76, gm_n62, gm_n597, gm_n443);
	nand (gm_n4984, gm_n373, gm_n72, in_17, gm_n4983, gm_n1076);
	nor (gm_n4985, gm_n168, gm_n158, gm_n60, gm_n1191, gm_n1331);
	nand (gm_n4986, in_21, in_20, in_19, gm_n4985);
	nor (gm_n4987, gm_n274, gm_n73, gm_n59, gm_n2730, gm_n385);
	nand (gm_n4988, gm_n495, in_21, in_20, gm_n4987);
	nand (gm_n4989, gm_n4988, gm_n4986, gm_n4984);
	nor (gm_n4990, gm_n4974, gm_n4962, gm_n4960, gm_n4989, gm_n4982);
	or (gm_n4991, gm_n461, in_13, in_9, gm_n1583, gm_n502);
	nor (gm_n4992, gm_n183, in_21, gm_n55, gm_n4991, gm_n313);
	or (gm_n4993, gm_n227, in_16, in_12, gm_n1191, gm_n274);
	nor (gm_n4994, gm_n139, gm_n72, gm_n85, gm_n4993);
	or (gm_n4995, gm_n92, in_14, in_10, gm_n286, gm_n95);
	nor (gm_n4996, gm_n211, gm_n89, gm_n119, gm_n4995);
	nor (gm_n4997, gm_n4996, gm_n4994, gm_n4992);
	nand (gm_n4998, gm_n214, in_13, in_12, gm_n2665, gm_n595);
	nor (gm_n4999, gm_n312, gm_n72, in_17, gm_n4998);
	nand (gm_n5000, gm_n61, in_16, in_12, gm_n612, gm_n64);
	nor (gm_n5001, gm_n219, in_21, in_20, gm_n5000);
	or (gm_n5002, gm_n344, in_13, in_9, gm_n481, gm_n442);
	nor (gm_n5003, gm_n184, in_21, in_17, gm_n5002, gm_n388);
	nor (gm_n5004, gm_n5003, gm_n5001, gm_n4999);
	nand (gm_n5005, gm_n4990, gm_n4958, gm_n4956, gm_n5004, gm_n4997);
	nor (gm_n5006, gm_n358, gm_n76, gm_n62, gm_n481, gm_n430);
	nand (gm_n5007, gm_n206, gm_n72, gm_n55, gm_n5006, gm_n405);
	nor (gm_n5008, gm_n274, gm_n73, in_12, gm_n2589, gm_n319);
	nand (gm_n5009, gm_n697, in_21, gm_n85, gm_n5008);
	nor (gm_n5010, gm_n161, in_12, gm_n94, gm_n319, gm_n263);
	nand (gm_n5011, gm_n72, gm_n85, in_16, gm_n5010, gm_n383);
	nand (gm_n5012, gm_n5011, gm_n5009, gm_n5007);
	and (gm_n5013, gm_n76, in_9, gm_n94, gm_n756, gm_n340);
	nand (gm_n5014, gm_n206, gm_n72, in_17, gm_n5013, gm_n405);
	nor (gm_n5015, gm_n430, in_13, gm_n62, gm_n597, gm_n257);
	nand (gm_n5016, gm_n523, gm_n72, in_17, gm_n5015, gm_n373);
	nor (gm_n5017, gm_n461, gm_n76, in_9, gm_n502, gm_n462);
	nand (gm_n5018, gm_n206, gm_n72, gm_n55, gm_n5017, gm_n595);
	nand (gm_n5019, gm_n5018, gm_n5016, gm_n5014);
	nor (gm_n5020, gm_n5005, gm_n4954, gm_n4952, gm_n5019, gm_n5012);
	or (gm_n5021, gm_n514, gm_n76, in_9, gm_n468, gm_n184);
	nor (gm_n5022, gm_n103, gm_n72, in_17, gm_n5021);
	nand (gm_n5023, gm_n78, gm_n62, gm_n94, gm_n1692, gm_n624);
	nor (gm_n5024, gm_n87, gm_n119, gm_n90, gm_n5023, gm_n437);
	or (gm_n5025, gm_n406, gm_n76, in_9, gm_n481, gm_n596);
	nor (gm_n5026, gm_n121, gm_n72, in_17, gm_n5025, gm_n388);
	nor (gm_n5027, gm_n5026, gm_n5024, gm_n5022);
	nand (gm_n5028, gm_n143, in_16, gm_n59, gm_n275, gm_n224);
	nor (gm_n5029, gm_n219, gm_n72, gm_n85, gm_n5028);
	nor (gm_n5030, gm_n620, in_21, gm_n55, gm_n3066, gm_n328);
	or (gm_n5031, gm_n208, gm_n461, gm_n76, gm_n491, gm_n328);
	nor (gm_n5032, gm_n620, in_21, gm_n55, gm_n5031);
	nor (gm_n5033, gm_n5032, gm_n5030, gm_n5029);
	nand (gm_n5034, gm_n5020, gm_n4950, gm_n4948, gm_n5033, gm_n5027);
	and (gm_n5035, gm_n64, in_16, in_12, gm_n1451, gm_n949);
	nand (gm_n5036, gm_n179, gm_n72, in_20, gm_n5035);
	nor (gm_n5037, in_14, in_10, gm_n62, gm_n1260, gm_n467);
	nand (gm_n5038, gm_n436, gm_n86, gm_n119, gm_n5037);
	and (gm_n5039, gm_n268, gm_n64, in_15, gm_n449, gm_n427);
	nand (gm_n5040, gm_n72, gm_n85, in_19, gm_n5039);
	nand (gm_n5041, gm_n5040, gm_n5038, gm_n5036);
	nor (gm_n5042, gm_n148, gm_n99, in_13, gm_n461, gm_n184);
	nand (gm_n5043, gm_n120, in_21, gm_n55, gm_n5042);
	and (gm_n5044, in_13, gm_n62, in_8, gm_n1263, gm_n314);
	nand (gm_n5045, gm_n174, gm_n72, in_17, gm_n5044, gm_n595);
	nor (gm_n5046, gm_n344, gm_n76, in_9, gm_n503, gm_n480);
	nand (gm_n5047, gm_n102, in_21, in_17, gm_n5046, gm_n122);
	nand (gm_n5048, gm_n5047, gm_n5045, gm_n5043);
	nor (gm_n5049, gm_n5034, gm_n4946, gm_n4944, gm_n5048, gm_n5041);
	or (gm_n5050, in_14, in_10, gm_n62, gm_n1016, gm_n467);
	nor (gm_n5051, gm_n1989, gm_n244, in_18, gm_n5050);
	or (gm_n5052, gm_n152, gm_n73, in_12, gm_n3929, gm_n263);
	nor (gm_n5053, gm_n912, gm_n72, gm_n85, gm_n5052);
	or (gm_n5054, gm_n358, gm_n76, gm_n62, gm_n432, gm_n667);
	nor (gm_n5055, gm_n121, in_21, in_17, gm_n5054, gm_n479);
	nor (gm_n5056, gm_n5055, gm_n5053, gm_n5051);
	or (gm_n5057, gm_n159, gm_n297, gm_n60, gm_n3006, gm_n485);
	nor (gm_n5058, in_21, in_20, in_19, gm_n5057);
	nand (gm_n5059, gm_n126, gm_n76, gm_n62, gm_n314, gm_n186);
	nor (gm_n5060, gm_n183, gm_n72, in_17, gm_n5059, gm_n256);
	or (gm_n5061, gm_n259, in_14, gm_n78, gm_n362, gm_n349);
	nor (gm_n5062, gm_n368, gm_n132, in_18, gm_n5061);
	nor (gm_n5063, gm_n5062, gm_n5060, gm_n5058);
	nand (gm_n5064, gm_n5049, gm_n4942, gm_n4940, gm_n5063, gm_n5056);
	nor (gm_n5065, gm_n514, gm_n76, in_9, gm_n1583, gm_n609);
	nand (gm_n5066, gm_n102, in_21, gm_n55, gm_n5065, gm_n255);
	nand (gm_n5067, gm_n255, gm_n72, in_17, gm_n3897, gm_n327);
	and (gm_n5068, gm_n233, gm_n73, in_12, gm_n626, gm_n949);
	nand (gm_n5069, gm_n179, in_21, in_20, gm_n5068);
	nand (gm_n5070, gm_n5069, gm_n5067, gm_n5066);
	and (gm_n5071, gm_n64, gm_n76, in_12, gm_n2416);
	nand (gm_n5072, gm_n254, gm_n72, in_17, gm_n5071, gm_n1076);
	nor (gm_n5073, gm_n148, in_14, in_10, gm_n589, gm_n362);
	nand (gm_n5074, gm_n245, gm_n129, in_18, gm_n5073);
	and (gm_n5075, gm_n281, gm_n222, in_15, gm_n2218, gm_n422);
	nand (gm_n5076, gm_n72, gm_n85, in_19, gm_n5075);
	nand (gm_n5077, gm_n5076, gm_n5074, gm_n5072);
	nor (gm_n5078, gm_n5064, gm_n4938, gm_n4937, gm_n5077, gm_n5070);
	nand (gm_n5079, gm_n126, gm_n76, gm_n62, gm_n341, gm_n579);
	nor (gm_n5080, gm_n388, in_21, gm_n55, gm_n5079, gm_n375);
	nand (gm_n5081, gm_n222, in_12, gm_n94, gm_n571, gm_n1379);
	nor (gm_n5082, in_21, gm_n85, in_16, gm_n5081, gm_n384);
	and (gm_n5083, gm_n254, gm_n72, gm_n55, gm_n3232, gm_n595);
	nor (gm_n5084, gm_n5083, gm_n5082, gm_n5080);
	or (gm_n5085, gm_n431, in_13, gm_n62, gm_n743, gm_n344);
	nor (gm_n5086, gm_n184, in_21, gm_n55, gm_n5085, gm_n374);
	or (gm_n5087, gm_n431, in_13, gm_n62, gm_n988, gm_n596);
	nor (gm_n5088, gm_n441, gm_n72, in_17, gm_n5087, gm_n375);
	or (gm_n5089, gm_n662, gm_n76, gm_n62, gm_n3315, gm_n406);
	nor (gm_n5090, gm_n183, gm_n72, in_17, gm_n5089);
	nor (gm_n5091, gm_n5090, gm_n5088, gm_n5086);
	nand (gm_n5092, gm_n5078, gm_n4934, gm_n4932, gm_n5091, gm_n5084);
	nand (gm_n5093, gm_n122, gm_n72, in_17, gm_n3070, gm_n206);
	nor (gm_n5094, gm_n344, in_13, gm_n62, gm_n503, gm_n480);
	nand (gm_n5095, gm_n104, in_21, gm_n55, gm_n5094, gm_n206);
	nor (gm_n5096, gm_n193, in_15, gm_n63, gm_n541, gm_n407);
	nand (gm_n5097, gm_n72, gm_n85, gm_n56, gm_n5096, gm_n379);
	nand (gm_n5098, gm_n5097, gm_n5095, gm_n5093);
	nor (gm_n5099, gm_n344, gm_n76, gm_n62, gm_n621, gm_n442);
	nand (gm_n5100, gm_n174, in_21, gm_n55, gm_n5099, gm_n595);
	nor (gm_n5101, gm_n514, in_13, gm_n62, gm_n1583, gm_n430);
	nand (gm_n5102, gm_n122, gm_n72, in_17, gm_n5101, gm_n373);
	nor (gm_n5103, gm_n148, in_14, gm_n78, gm_n362, gm_n208);
	nand (gm_n5104, gm_n245, gm_n86, in_18, gm_n5103);
	nand (gm_n5105, gm_n5104, gm_n5102, gm_n5100);
	nor (gm_n5106, gm_n5092, gm_n4930, gm_n4928, gm_n5105, gm_n5098);
	or (gm_n5107, gm_n147, in_14, in_10, gm_n414, gm_n370);
	nor (gm_n5108, gm_n1989, gm_n87, gm_n119, gm_n5107);
	nor (gm_n5109, gm_n167, gm_n87, gm_n119, gm_n1987);
	nor (gm_n5110, gm_n247, gm_n208, gm_n78, gm_n362);
	and (gm_n5111, gm_n523, gm_n72, gm_n55, gm_n5110, gm_n373);
	nor (gm_n5112, gm_n5111, gm_n5109, gm_n5108);
	nand (gm_n5113, gm_n484, gm_n60, gm_n94, gm_n455, gm_n264);
	nor (gm_n5114, in_21, gm_n85, gm_n56, gm_n5113, gm_n191);
	or (gm_n5115, gm_n248, gm_n358, gm_n76, gm_n349);
	nor (gm_n5116, gm_n105, gm_n72, gm_n55, gm_n5115, gm_n312);
	or (gm_n5117, gm_n431, in_13, gm_n62, gm_n503, gm_n443);
	nor (gm_n5118, gm_n183, in_21, in_17, gm_n5117, gm_n328);
	nor (gm_n5119, gm_n5118, gm_n5116, gm_n5114);
	nand (gm_n5120, gm_n5106, gm_n4925, gm_n4923, gm_n5119, gm_n5112);
	nor (gm_n5121, gm_n431, in_13, gm_n62, gm_n4437, gm_n328);
	nand (gm_n5122, gm_n174, in_21, gm_n55, gm_n5121);
	nand (gm_n5123, gm_n72, in_20, in_19, gm_n3522, gm_n281);
	nor (gm_n5124, gm_n358, in_13, in_9, gm_n743, gm_n667);
	nand (gm_n5125, gm_n120, gm_n72, in_17, gm_n5124, gm_n122);
	nand (gm_n5126, gm_n5125, gm_n5123, gm_n5122);
	and (gm_n5127, gm_n422, gm_n143, in_15, gm_n1531);
	nand (gm_n5128, in_21, gm_n85, gm_n56, gm_n5127, gm_n448);
	or (gm_n5129, gm_n105, in_21, gm_n55, gm_n3464, gm_n183);
	nor (gm_n5130, gm_n514, in_13, in_9, gm_n1583, gm_n463);
	nand (gm_n5131, gm_n120, in_21, in_17, gm_n5130, gm_n122);
	nand (gm_n5132, gm_n5131, gm_n5129, gm_n5128);
	nor (gm_n5133, gm_n5120, gm_n4921, gm_n4919, gm_n5132, gm_n5126);
	nor (gm_n5134, gm_n368, gm_n167, in_18, gm_n4656);
	or (gm_n5135, in_14, in_10, gm_n62, gm_n520, gm_n467);
	nor (gm_n5136, gm_n167, gm_n130, gm_n119, gm_n5135);
	or (gm_n5137, gm_n297, in_16, in_12, gm_n1514, gm_n152);
	nor (gm_n5138, gm_n781, gm_n72, gm_n85, gm_n5137);
	nor (gm_n5139, gm_n5138, gm_n5136, gm_n5134);
	or (gm_n5140, gm_n818, gm_n76, in_9, gm_n344, gm_n358);
	nor (gm_n5141, gm_n184, gm_n72, in_17, gm_n5140, gm_n374);
	or (gm_n5142, gm_n99, in_14, in_10, gm_n438, gm_n807);
	nor (gm_n5143, gm_n212, gm_n165, gm_n119, gm_n5142);
	or (gm_n5144, gm_n152, gm_n73, in_12, gm_n263, gm_n196);
	nor (gm_n5145, gm_n219, gm_n72, gm_n85, gm_n5144);
	nor (gm_n5146, gm_n5145, gm_n5143, gm_n5141);
	nand (gm_n5147, gm_n5133, gm_n4916, gm_n4914, gm_n5146, gm_n5139);
	nand (gm_n5148, gm_n102, gm_n72, gm_n55, gm_n2681, gm_n255);
	nand (gm_n5149, gm_n327, gm_n72, in_17, gm_n2749, gm_n1076);
	nand (gm_n5150, gm_n436, gm_n243, in_18, gm_n1629);
	nand (gm_n5151, gm_n5150, gm_n5149, gm_n5148);
	and (gm_n5152, gm_n802, gm_n304, in_8);
	and (gm_n5153, gm_n214, gm_n192, gm_n60, gm_n5152, gm_n486);
	nand (gm_n5154, in_21, gm_n85, in_19, gm_n5153);
	nor (gm_n5155, in_14, in_10, gm_n62, gm_n705, gm_n207);
	nand (gm_n5156, gm_n806, gm_n164, in_18, gm_n5155);
	nor (gm_n5157, gm_n461, in_13, in_9, gm_n988, gm_n502);
	nand (gm_n5158, gm_n595, gm_n72, in_17, gm_n5157, gm_n373);
	nand (gm_n5159, gm_n5158, gm_n5156, gm_n5154);
	nor (gm_n5160, gm_n5147, gm_n4912, gm_n4911, gm_n5159, gm_n5151);
	or (gm_n5161, gm_n190, gm_n73, gm_n59, gm_n1052, gm_n227);
	nor (gm_n5162, gm_n781, in_21, gm_n85, gm_n5161);
	nand (gm_n5163, gm_n123, gm_n76, in_9, gm_n2683, gm_n1076);
	nor (gm_n5164, gm_n479, in_21, gm_n55, gm_n5163);
	or (gm_n5165, gm_n152, in_12, in_8, gm_n1382, gm_n274);
	nor (gm_n5166, gm_n72, in_20, in_16, gm_n5165, gm_n219);
	nor (gm_n5167, gm_n5166, gm_n5164, gm_n5162);
	or (gm_n5168, gm_n393, gm_n297, in_15, gm_n1191, gm_n764);
	nor (gm_n5169, gm_n72, in_20, gm_n56, gm_n5168);
	or (gm_n5170, gm_n147, in_14, in_10, gm_n370, gm_n208);
	nor (gm_n5171, gm_n212, gm_n87, gm_n119, gm_n5170);
	nand (gm_n5172, gm_n523, gm_n76, gm_n62, gm_n2230, gm_n340);
	nor (gm_n5173, gm_n441, in_21, in_17, gm_n5172);
	nor (gm_n5174, gm_n5173, gm_n5171, gm_n5169);
	nand (gm_n5175, gm_n5160, gm_n4910, gm_n4908, gm_n5174, gm_n5167);
	nand (gm_n5176, gm_n166, gm_n164, gm_n119, gm_n2240);
	nor (gm_n5177, gm_n239, in_15, in_11, gm_n605, gm_n643);
	nand (gm_n5178, gm_n72, in_20, in_19, gm_n5177, gm_n486);
	nor (gm_n5179, gm_n461, gm_n76, in_9, gm_n462, gm_n344);
	nand (gm_n5180, gm_n254, gm_n72, in_17, gm_n5179, gm_n405);
	nand (gm_n5181, gm_n5180, gm_n5178, gm_n5176);
	nor (gm_n5182, gm_n461, in_13, in_9, gm_n743, gm_n502);
	nand (gm_n5183, gm_n255, gm_n72, in_17, gm_n5182, gm_n311);
	nor (gm_n5184, gm_n274, in_16, in_12, gm_n1260, gm_n385);
	nand (gm_n5185, gm_n57, gm_n72, gm_n85, gm_n5184);
	nor (gm_n5186, in_14, gm_n78, in_9, gm_n1698, gm_n807);
	nand (gm_n5187, gm_n806, gm_n164, in_18, gm_n5186);
	nand (gm_n5188, gm_n5187, gm_n5185, gm_n5183);
	nor (gm_n5189, gm_n5175, gm_n4906, gm_n4904, gm_n5188, gm_n5181);
	or (gm_n5190, gm_n431, gm_n76, gm_n62, gm_n502, gm_n432);
	nor (gm_n5191, gm_n183, gm_n72, gm_n55, gm_n5190, gm_n121);
	or (gm_n5192, gm_n155, in_16, in_12, gm_n1176, gm_n385);
	nor (gm_n5193, gm_n262, in_21, gm_n85, gm_n5192);
	nand (gm_n5194, gm_n392, gm_n75, in_15, gm_n751, gm_n222);
	nor (gm_n5195, in_21, in_20, gm_n56, gm_n5194);
	nor (gm_n5196, gm_n5195, gm_n5193, gm_n5191);
	or (gm_n5197, gm_n461, in_13, in_9, gm_n432, gm_n430);
	nor (gm_n5198, gm_n184, in_21, in_17, gm_n5197, gm_n388);
	or (gm_n5199, gm_n514, in_13, in_9, gm_n502, gm_n818);
	nor (gm_n5200, gm_n256, gm_n72, gm_n55, gm_n5199, gm_n620);
	nand (gm_n5201, gm_n339, in_13, in_9, gm_n3876, gm_n402);
	nor (gm_n5202, gm_n441, gm_n72, gm_n55, gm_n5201);
	nor (gm_n5203, gm_n5202, gm_n5200, gm_n5198);
	nand (gm_n5204, gm_n5189, gm_n4902, gm_n4900, gm_n5203, gm_n5196);
	and (gm_n5205, gm_n107, in_13, gm_n62, gm_n402, gm_n316);
	nand (gm_n5206, gm_n122, gm_n72, in_17, gm_n5205, gm_n206);
	nor (gm_n5207, gm_n442, gm_n76, in_9, gm_n1132, gm_n443);
	nand (gm_n5208, gm_n255, gm_n72, in_17, gm_n5207, gm_n311);
	and (gm_n5209, gm_n79, in_13, gm_n59, gm_n685);
	nand (gm_n5210, gm_n122, gm_n72, gm_n55, gm_n5209, gm_n254);
	nand (gm_n5211, gm_n5210, gm_n5208, gm_n5206);
	nor (gm_n5212, gm_n133, in_14, in_10, gm_n259, gm_n148);
	nand (gm_n5213, gm_n164, gm_n88, gm_n119, gm_n5212);
	nor (gm_n5214, gm_n158, gm_n74, gm_n60, gm_n1965, gm_n764);
	nand (gm_n5215, gm_n72, in_20, in_19, gm_n5214);
	and (gm_n5216, gm_n1011, in_14, in_10, gm_n722, gm_n490);
	nand (gm_n5217, gm_n245, gm_n86, in_18, gm_n5216);
	nand (gm_n5218, gm_n5217, gm_n5215, gm_n5213);
	nor (gm_n5219, gm_n5204, gm_n4898, gm_n4896, gm_n5218, gm_n5211);
	and (gm_n5220, gm_n142, in_16, gm_n59, gm_n275, gm_n154);
	nand (gm_n5221, gm_n113, gm_n72, gm_n85, gm_n5220);
	nand (gm_n5222, gm_n120, in_21, in_17, gm_n5110, gm_n1076);
	and (gm_n5223, gm_n392, in_15, in_11, gm_n1615, gm_n171);
	nand (gm_n5224, in_21, gm_n85, gm_n56, gm_n5223, gm_n75);
	nand (gm_n5225, gm_n5221, gm_n5219, gm_n4894, gm_n5224, gm_n5222);
	nor (gm_n5226, gm_n227, in_16, in_12, gm_n499, gm_n155);
	nand (gm_n5227, gm_n179, in_21, in_20, gm_n5226);
	and (gm_n5228, gm_n107, in_13, gm_n62, gm_n788, gm_n316);
	nand (gm_n5229, gm_n102, in_21, in_17, gm_n5228, gm_n405);
	nor (gm_n5230, gm_n1331, gm_n274, gm_n60, gm_n1519, gm_n760);
	nand (gm_n5231, in_21, gm_n85, gm_n56, gm_n5230);
	nand (gm_n5232, gm_n5231, gm_n5229, gm_n5227);
	and (gm_n5233, gm_n1067, gm_n171, gm_n304);
	nand (gm_n5234, gm_n394, in_15, in_11, gm_n5233, gm_n869);
	nor (gm_n5235, gm_n72, gm_n85, gm_n56, gm_n5234);
	nor (out_13, gm_n5232, gm_n5225, gm_n4892, gm_n5235);
	nand (gm_n5237, gm_n392, gm_n79, gm_n60, gm_n1095, gm_n1101);
	nor (gm_n5238, in_21, in_20, in_19, gm_n5237);
	nor (gm_n5239, gm_n290, gm_n274, gm_n60, gm_n2956, gm_n393);
	nand (gm_n5240, gm_n72, gm_n85, in_19, gm_n5239);
	and (gm_n5241, gm_n91, in_14, in_10, gm_n333, gm_n995);
	nand (gm_n5242, gm_n367, gm_n245, in_18, gm_n5241);
	nand (gm_n5243, gm_n316, in_13, gm_n62, gm_n402, gm_n341);
	nor (gm_n5244, gm_n184, gm_n72, in_17, gm_n5243, gm_n620);
	or (gm_n5245, gm_n159, gm_n155, in_15, gm_n324, gm_n293);
	nor (gm_n5246, gm_n72, in_20, gm_n56, gm_n5245);
	and (gm_n5247, gm_n110, in_13, gm_n62, gm_n1049, gm_n314);
	nand (gm_n5248, gm_n327, in_21, gm_n55, gm_n5247, gm_n339);
	nand (gm_n5249, gm_n255, in_21, gm_n55, gm_n4590, gm_n327);
	and (gm_n5250, gm_n102, in_21, in_17, gm_n412, gm_n104);
	or (gm_n5251, gm_n158, in_16, gm_n59, gm_n1906, gm_n276);
	nor (gm_n5252, gm_n781, in_21, in_20, gm_n5251);
	nor (gm_n5253, gm_n818, in_13, in_9, gm_n463, gm_n257);
	nand (gm_n5254, gm_n254, gm_n72, in_17, gm_n5253, gm_n595);
	nor (gm_n5255, gm_n667, in_13, in_9, gm_n597, gm_n442);
	nand (gm_n5256, gm_n255, gm_n72, in_17, gm_n5255, gm_n373);
	or (gm_n5257, gm_n115, in_16, in_12, gm_n849, gm_n152);
	nor (gm_n5258, gm_n912, gm_n72, gm_n85, gm_n5257);
	nor (gm_n5259, gm_n105, gm_n72, in_17, gm_n2661, gm_n441);
	nor (gm_n5260, gm_n193, gm_n115, gm_n60, gm_n2826, gm_n293);
	nand (gm_n5261, in_21, in_20, in_19, gm_n5260);
	nor (gm_n5262, gm_n208, gm_n90, gm_n78, gm_n349, gm_n807);
	nand (gm_n5263, gm_n243, gm_n88, in_18, gm_n5262);
	or (gm_n5264, in_14, gm_n78, in_9, gm_n1284, gm_n369);
	nor (gm_n5265, gm_n244, gm_n167, gm_n119, gm_n5264);
	nand (gm_n5266, gm_n79, gm_n73, in_12, gm_n2497, gm_n275);
	nor (gm_n5267, gm_n262, in_21, gm_n85, gm_n5266);
	and (gm_n5268, gm_n187, in_13, gm_n62, gm_n1049, gm_n579);
	nand (gm_n5269, gm_n595, gm_n72, gm_n55, gm_n5268, gm_n373);
	and (gm_n5270, gm_n171, gm_n60, gm_n63, gm_n1398, gm_n556);
	nand (gm_n5271, gm_n72, in_20, gm_n56, gm_n5270, gm_n486);
	or (gm_n5272, gm_n596, gm_n76, in_9, gm_n442, gm_n345);
	nor (gm_n5273, gm_n441, in_21, in_17, gm_n5272, gm_n375);
	or (gm_n5274, gm_n609, gm_n76, gm_n62, gm_n743, gm_n480);
	nor (gm_n5275, gm_n313, gm_n72, in_17, gm_n5274, gm_n374);
	nor (gm_n5276, gm_n269, gm_n274, gm_n60, gm_n1716, gm_n633);
	and (gm_n5277, in_21, gm_n85, gm_n56, gm_n5276);
	nor (gm_n5278, gm_n461, in_13, gm_n62, gm_n502, gm_n345);
	and (gm_n5279, gm_n405, gm_n72, gm_n55, gm_n5278, gm_n373);
	and (gm_n5280, gm_n90, gm_n76, gm_n59, gm_n936, gm_n233);
	and (gm_n5281, gm_n348, gm_n88, in_18, gm_n5280);
	nor (gm_n5282, gm_n115, gm_n74, in_15, gm_n2038, gm_n290);
	and (gm_n5283, gm_n72, gm_n85, gm_n56, gm_n5282);
	or (gm_n5284, gm_n5279, gm_n5277, t_3, gm_n5283, gm_n5281);
	nor (gm_n5285, gm_n461, gm_n76, gm_n62, gm_n1514, gm_n662);
	nand (gm_n5286, gm_n102, gm_n72, in_17, gm_n5285);
	nor (gm_n5287, gm_n406, gm_n247, in_13, gm_n414, gm_n375);
	nand (gm_n5288, gm_n254, gm_n72, in_17, gm_n5287);
	nor (gm_n5289, gm_n95, in_14, in_10, gm_n389, gm_n133);
	nand (gm_n5290, gm_n436, gm_n146, gm_n119, gm_n5289);
	nand (gm_n5291, gm_n5290, gm_n5288, gm_n5286);
	nand (gm_n5292, gm_n436, gm_n243, in_18, gm_n3148);
	nand (gm_n5293, gm_n102, gm_n72, gm_n55, gm_n2286, gm_n1076);
	nor (gm_n5294, gm_n90, in_13, gm_n59, gm_n1698, gm_n274);
	nand (gm_n5295, gm_n367, gm_n245, in_18, gm_n5294);
	nand (gm_n5296, gm_n5295, gm_n5293, gm_n5292);
	nor (gm_n5297, gm_n5284, gm_n5275, gm_n5273, gm_n5296, gm_n5291);
	nand (gm_n5298, gm_n264, in_16, in_12, gm_n3587, gm_n949);
	nor (gm_n5299, gm_n139, in_21, in_20, gm_n5298);
	nand (gm_n5300, gm_n486, gm_n154, gm_n60, gm_n1427, gm_n1398);
	nor (gm_n5301, gm_n72, in_20, gm_n56, gm_n5300);
	or (gm_n5302, gm_n147, in_14, in_10, gm_n247, gm_n149);
	nor (gm_n5303, gm_n368, gm_n1989, in_18, gm_n5302);
	nor (gm_n5304, gm_n5303, gm_n5301, gm_n5299);
	nand (gm_n5305, in_14, in_10, gm_n62, gm_n1392, gm_n1011);
	nor (gm_n5306, gm_n246, gm_n211, gm_n119, gm_n5305);
	nor (gm_n5307, gm_n93, in_6, gm_n97, gm_n141, in_8);
	nand (gm_n5308, gm_n214, gm_n73, in_12, gm_n5307, gm_n571);
	nor (gm_n5309, gm_n781, in_21, gm_n85, gm_n5308);
	or (gm_n5310, gm_n168, gm_n297, in_15, gm_n3440, gm_n393);
	nor (gm_n5311, gm_n72, in_20, in_19, gm_n5310);
	nor (gm_n5312, gm_n5311, gm_n5309, gm_n5306);
	nand (gm_n5313, gm_n5297, gm_n5271, gm_n5269, gm_n5312, gm_n5304);
	and (gm_n5314, gm_n107, in_13, gm_n62, gm_n340, gm_n126);
	nand (gm_n5315, gm_n523, gm_n72, in_17, gm_n5314, gm_n206);
	and (gm_n5316, gm_n75, in_15, in_11, gm_n5233, gm_n484);
	nand (gm_n5317, gm_n72, gm_n85, gm_n56, gm_n5316);
	nor (gm_n5318, gm_n95, in_14, gm_n78, gm_n807, gm_n99);
	nand (gm_n5319, gm_n806, gm_n199, gm_n119, gm_n5318);
	nand (gm_n5320, gm_n5319, gm_n5317, gm_n5315);
	nor (gm_n5321, gm_n290, gm_n263, gm_n60, gm_n3440, gm_n393);
	nand (gm_n5322, gm_n72, gm_n85, in_19, gm_n5321);
	nor (gm_n5323, gm_n370, gm_n90, gm_n78, gm_n467, gm_n376);
	nand (gm_n5324, gm_n166, gm_n146, gm_n119, gm_n5323);
	nor (gm_n5325, gm_n293, gm_n115, in_15, gm_n2826, gm_n764);
	nand (gm_n5326, gm_n72, in_20, gm_n56, gm_n5325);
	nand (gm_n5327, gm_n5326, gm_n5324, gm_n5322);
	nor (gm_n5328, gm_n5313, gm_n5267, gm_n5265, gm_n5327, gm_n5320);
	nand (gm_n5329, gm_n448, gm_n233, in_15, gm_n2624, gm_n1398);
	nor (gm_n5330, gm_n72, in_20, gm_n56, gm_n5329);
	or (gm_n5331, gm_n99, in_14, gm_n78, gm_n369, gm_n287);
	nor (gm_n5332, gm_n368, gm_n841, in_18, gm_n5331);
	nand (gm_n5333, gm_n484, gm_n60, in_11, gm_n580, gm_n1614);
	nor (gm_n5334, gm_n72, in_20, gm_n56, gm_n5333, gm_n1331);
	nor (gm_n5335, gm_n5334, gm_n5332, gm_n5330);
	or (gm_n5336, gm_n227, in_16, gm_n59, gm_n849, gm_n297);
	nor (gm_n5337, gm_n496, in_21, gm_n85, gm_n5336);
	or (gm_n5338, gm_n461, gm_n76, in_9, gm_n443, gm_n345);
	nor (gm_n5339, gm_n479, in_21, in_17, gm_n5338, gm_n256);
	or (gm_n5340, gm_n158, gm_n59, gm_n94, gm_n2769, gm_n385);
	nor (gm_n5341, in_21, gm_n85, gm_n73, gm_n5340, gm_n139);
	nor (gm_n5342, gm_n5341, gm_n5339, gm_n5337);
	nand (gm_n5343, gm_n5328, gm_n5263, gm_n5261, gm_n5342, gm_n5335);
	and (gm_n5344, gm_n600, in_14, in_10, gm_n829, gm_n490);
	nand (gm_n5345, gm_n348, gm_n166, in_18, gm_n5344);
	nor (gm_n5346, gm_n609, in_13, in_9, gm_n743, gm_n406);
	nand (gm_n5347, gm_n102, gm_n72, in_17, gm_n5346, gm_n122);
	nor (gm_n5348, gm_n99, gm_n90, gm_n78, gm_n287, gm_n147);
	nand (gm_n5349, gm_n131, gm_n129, in_18, gm_n5348);
	nand (gm_n5350, gm_n5349, gm_n5347, gm_n5345);
	nor (gm_n5351, gm_n514, gm_n76, in_9, gm_n443, gm_n359);
	nand (gm_n5352, gm_n311, gm_n72, in_17, gm_n5351, gm_n405);
	and (gm_n5353, gm_n233, gm_n73, gm_n59, gm_n950, gm_n571);
	nand (gm_n5354, gm_n113, gm_n72, gm_n85, gm_n5353);
	nor (gm_n5355, gm_n293, gm_n263, in_15, gm_n1671, gm_n760);
	nand (gm_n5356, in_21, gm_n85, in_19, gm_n5355);
	nand (gm_n5357, gm_n5356, gm_n5354, gm_n5352);
	nor (gm_n5358, gm_n5343, gm_n5259, gm_n5258, gm_n5357, gm_n5350);
	or (gm_n5359, gm_n152, gm_n73, gm_n59, gm_n2357, gm_n274);
	nor (gm_n5360, gm_n262, gm_n72, gm_n85, gm_n5359);
	nand (gm_n5361, gm_n264, gm_n392, gm_n60, gm_n1605, gm_n394);
	nor (gm_n5362, in_21, gm_n85, in_19, gm_n5361);
	or (gm_n5363, gm_n344, in_10, gm_n62, gm_n597, gm_n467);
	nor (gm_n5364, gm_n1989, in_18, in_14, gm_n5363, gm_n368);
	nor (gm_n5365, gm_n5364, gm_n5362, gm_n5360);
	or (gm_n5366, gm_n313, in_13, gm_n62, gm_n406, gm_n329);
	nor (gm_n5367, gm_n103, gm_n72, in_17, gm_n5366);
	or (gm_n5368, gm_n257, gm_n76, in_9, gm_n502, gm_n345);
	nor (gm_n5369, gm_n388, gm_n72, gm_n55, gm_n5368, gm_n375);
	or (gm_n5370, gm_n514, in_13, gm_n62, gm_n1132, gm_n344);
	nor (gm_n5371, gm_n388, gm_n72, gm_n55, gm_n5370, gm_n662);
	nor (gm_n5372, gm_n5371, gm_n5369, gm_n5367);
	nand (gm_n5373, gm_n5358, gm_n5256, gm_n5254, gm_n5372, gm_n5365);
	nor (gm_n5374, gm_n442, gm_n76, gm_n62, gm_n621, gm_n443);
	nand (gm_n5375, gm_n174, gm_n72, gm_n55, gm_n5374, gm_n523);
	nor (gm_n5376, gm_n227, gm_n73, in_12, gm_n4917, gm_n158);
	nand (gm_n5377, gm_n138, gm_n72, in_20, gm_n5376);
	nor (gm_n5378, gm_n114, gm_n73, gm_n59, gm_n1751, gm_n297);
	nand (gm_n5379, gm_n57, gm_n72, in_20, gm_n5378);
	nand (gm_n5380, gm_n5379, gm_n5377, gm_n5375);
	and (gm_n5381, gm_n222, in_16, gm_n59, gm_n870, gm_n949);
	nand (gm_n5382, gm_n138, in_21, in_20, gm_n5381);
	nor (gm_n5383, gm_n257, gm_n76, in_9, gm_n502, gm_n462);
	nand (gm_n5384, gm_n523, in_21, gm_n55, gm_n5383, gm_n311);
	nor (gm_n5385, gm_n190, in_16, gm_n59, gm_n2826, gm_n354);
	nand (gm_n5386, gm_n383, in_21, in_20, gm_n5385);
	nand (gm_n5387, gm_n5386, gm_n5384, gm_n5382);
	nor (gm_n5388, gm_n5373, gm_n5252, gm_n5250, gm_n5387, gm_n5380);
	nor (gm_n5389, in_21, gm_n85, gm_n56, gm_n951, gm_n269);
	or (gm_n5390, gm_n115, gm_n74, gm_n60, gm_n1170, gm_n193);
	nor (gm_n5391, in_21, in_20, gm_n56, gm_n5390);
	or (gm_n5392, gm_n286, gm_n90, in_10, gm_n491, gm_n362);
	nor (gm_n5393, gm_n824, gm_n89, gm_n119, gm_n5392);
	nor (gm_n5394, gm_n5393, gm_n5391, gm_n5389);
	or (gm_n5395, gm_n514, in_13, gm_n62, gm_n481, gm_n344);
	nor (gm_n5396, gm_n388, in_21, in_17, gm_n5395, gm_n256);
	nand (gm_n5397, in_14, gm_n78, gm_n62, gm_n1501, gm_n91);
	nor (gm_n5398, gm_n246, gm_n211, in_18, gm_n5397);
	nand (gm_n5399, gm_n76, in_9, gm_n94, gm_n2074, gm_n579);
	nor (gm_n5400, gm_n256, gm_n72, gm_n55, gm_n5399, gm_n620);
	nor (gm_n5401, gm_n5400, gm_n5398, gm_n5396);
	nand (gm_n5402, gm_n5388, gm_n5249, gm_n5248, gm_n5401, gm_n5394);
	nor (gm_n5403, gm_n667, in_13, gm_n62, gm_n743, gm_n480);
	nand (gm_n5404, gm_n120, gm_n72, in_17, gm_n5403, gm_n523);
	nor (gm_n5405, gm_n115, in_13, gm_n59, gm_n2125);
	nand (gm_n5406, gm_n122, in_21, gm_n55, gm_n5405, gm_n254);
	and (gm_n5407, gm_n91, in_14, in_10, gm_n335, gm_n333);
	nand (gm_n5408, gm_n245, gm_n86, gm_n119, gm_n5407);
	nand (gm_n5409, gm_n5408, gm_n5406, gm_n5404);
	nor (gm_n5410, gm_n193, in_15, in_11, gm_n981, gm_n605);
	nand (gm_n5411, gm_n72, gm_n85, gm_n56, gm_n5410, gm_n448);
	nor (gm_n5412, gm_n514, in_13, gm_n62, gm_n621, gm_n502);
	nand (gm_n5413, gm_n523, in_21, in_17, gm_n5412, gm_n254);
	nor (gm_n5414, gm_n159, gm_n158, in_15, gm_n1671, gm_n191);
	nand (gm_n5415, gm_n72, in_20, in_19, gm_n5414);
	nand (gm_n5416, gm_n5415, gm_n5413, gm_n5411);
	nor (gm_n5417, gm_n5402, gm_n5246, gm_n5244, gm_n5416, gm_n5409);
	nand (gm_n5418, gm_n123, gm_n76, gm_n62, gm_n1049, gm_n316);
	nor (gm_n5419, gm_n105, gm_n72, gm_n55, gm_n5418, gm_n183);
	nor (gm_n5420, gm_n72, in_20, gm_n56, gm_n2126, gm_n74);
	nand (gm_n5421, gm_n143, gm_n73, gm_n59, gm_n685, gm_n733);
	nor (gm_n5422, gm_n139, in_21, gm_n85, gm_n5421);
	nor (gm_n5423, gm_n5422, gm_n5420, gm_n5419);
	nor (gm_n5424, gm_n441, in_21, gm_n55, gm_n5087, gm_n313);
	or (gm_n5425, gm_n114, in_16, in_12, gm_n2060, gm_n213);
	nor (gm_n5426, gm_n139, in_21, in_20, gm_n5425);
	or (gm_n5427, gm_n344, gm_n76, in_9, gm_n462, gm_n480);
	nor (gm_n5428, gm_n103, gm_n72, gm_n55, gm_n5427, gm_n256);
	nor (gm_n5429, gm_n5428, gm_n5426, gm_n5424);
	nand (gm_n5430, gm_n5417, gm_n5242, gm_n5240, gm_n5429, gm_n5423);
	or (gm_n5431, gm_n184, in_21, gm_n55, gm_n4584, gm_n620);
	nor (gm_n5432, gm_n514, in_13, in_9, gm_n443, gm_n818);
	nand (gm_n5433, gm_n120, in_21, gm_n55, gm_n5432, gm_n595);
	nor (gm_n5434, gm_n147, in_14, in_10, gm_n208, gm_n148);
	nand (gm_n5435, gm_n436, gm_n164, in_18, gm_n5434);
	nand (gm_n5436, gm_n5435, gm_n5433, gm_n5431);
	nand (gm_n5437, gm_n1076, in_13, gm_n62, gm_n1709, gm_n788);
	nor (gm_n5438, gm_n620, in_21, gm_n55, gm_n5437);
	nor (out_14, gm_n5436, gm_n5430, gm_n5238, gm_n5438);
	nand (gm_n5440, gm_n233, gm_n73, in_12, gm_n612, gm_n949);
	nor (gm_n5441, gm_n781, gm_n72, gm_n85, gm_n5440);
	or (gm_n5442, gm_n193, gm_n190, in_15, gm_n932, gm_n293);
	nor (gm_n5443, gm_n72, in_20, gm_n56, gm_n5442);
	nor (gm_n5444, gm_n269, gm_n297, gm_n60, gm_n2221, gm_n764);
	nand (gm_n5445, gm_n72, in_20, in_19, gm_n5444);
	nand (gm_n5446, gm_n64, gm_n73, gm_n59, gm_n2885, gm_n733);
	nor (gm_n5447, gm_n781, in_21, in_20, gm_n5446);
	and (gm_n5448, gm_n245, gm_n243, in_18, gm_n1360);
	nor (gm_n5449, gm_n431, in_13, gm_n62, gm_n432, gm_n344);
	and (gm_n5450, gm_n405, in_21, gm_n55, gm_n5449, gm_n327);
	nor (gm_n5451, gm_n514, gm_n76, gm_n62, gm_n1583, gm_n463);
	and (gm_n5452, gm_n327, in_21, gm_n55, gm_n5451, gm_n339);
	or (gm_n5453, gm_n5448, gm_n5447, t_9, gm_n5452, gm_n5450);
	nand (gm_n5454, gm_n192, in_15, gm_n63, gm_n714, gm_n1614);
	nor (gm_n5455, in_21, in_20, in_19, gm_n5454, gm_n269);
	or (gm_n5456, in_14, in_10, gm_n62, gm_n2697, gm_n369);
	nor (gm_n5457, gm_n165, gm_n89, in_18, gm_n5456);
	or (gm_n5458, gm_n190, in_16, in_12, gm_n1923, gm_n152);
	nor (gm_n5459, gm_n58, gm_n72, gm_n85, gm_n5458);
	nor (gm_n5460, gm_n5457, gm_n5455, gm_n5453, gm_n5459);
	nor (gm_n5461, gm_n393, gm_n297, gm_n60, gm_n1923, gm_n643);
	nand (gm_n5462, in_21, in_20, gm_n56, gm_n5461);
	nor (gm_n5463, gm_n358, in_13, gm_n62, gm_n359, gm_n430);
	nand (gm_n5464, gm_n104, gm_n72, gm_n55, gm_n5463, gm_n311);
	nor (gm_n5465, gm_n596, in_13, gm_n62, gm_n743, gm_n480);
	nand (gm_n5466, gm_n206, gm_n72, in_17, gm_n5465, gm_n255);
	nand (gm_n5467, gm_n5462, gm_n5460, gm_n5445, gm_n5466, gm_n5464);
	nor (gm_n5468, gm_n485, gm_n158, gm_n60, gm_n1671, gm_n764);
	nand (gm_n5469, gm_n72, in_20, gm_n56, gm_n5468);
	nor (gm_n5470, gm_n158, in_16, gm_n59, gm_n1052, gm_n385);
	nand (gm_n5471, gm_n383, in_21, gm_n85, gm_n5470);
	and (gm_n5472, gm_n755, gm_n60, gm_n63, gm_n556, gm_n422);
	nand (gm_n5473, in_21, gm_n85, in_19, gm_n5472, gm_n448);
	nand (gm_n5474, gm_n5473, gm_n5471, gm_n5469);
	nand (gm_n5475, gm_n123, gm_n76, in_9, gm_n685, gm_n255);
	nor (gm_n5476, gm_n441, gm_n72, gm_n55, gm_n5475);
	nor (out_15, gm_n5467, gm_n5443, gm_n5441, gm_n5476, gm_n5474);
	nand (gm_n5478, in_14, gm_n78, gm_n62, gm_n1713, gm_n1011);
	nor (gm_n5479, gm_n211, gm_n89, in_18, gm_n5478);
	nor (gm_n5480, gm_n431, gm_n76, in_9, gm_n503, gm_n596);
	nand (gm_n5481, gm_n174, in_21, in_17, gm_n5480, gm_n339);
	nand (gm_n5482, gm_n154, in_16, in_12, gm_n1230, gm_n303);
	nor (gm_n5483, gm_n781, in_21, gm_n85, gm_n5482);
	or (gm_n5484, gm_n609, in_13, in_9, gm_n743, gm_n461);
	nor (gm_n5485, gm_n388, in_21, gm_n55, gm_n5484, gm_n662);
	nand (gm_n5486, gm_n243, gm_n131, in_18, gm_n5280);
	nor (gm_n5487, gm_n227, gm_n73, gm_n59, gm_n1719, gm_n274);
	nand (gm_n5488, gm_n495, in_21, gm_n85, gm_n5487);
	or (gm_n5489, gm_n114, gm_n73, in_12, gm_n399, gm_n274);
	nor (gm_n5490, gm_n139, in_21, gm_n85, gm_n5489);
	or (gm_n5491, gm_n393, gm_n213, in_15, gm_n1246, gm_n633);
	nor (gm_n5492, in_21, in_20, in_19, gm_n5491);
	nor (gm_n5493, gm_n358, gm_n76, gm_n62, gm_n503, gm_n596);
	nand (gm_n5494, gm_n174, gm_n72, in_17, gm_n5493, gm_n523);
	nor (gm_n5495, gm_n257, gm_n76, gm_n62, gm_n743, gm_n502);
	nand (gm_n5496, gm_n523, in_21, in_17, gm_n5495, gm_n206);
	or (gm_n5497, gm_n114, gm_n73, in_12, gm_n860, gm_n115);
	nor (gm_n5498, gm_n58, in_21, in_20, gm_n5497);
	or (gm_n5499, gm_n359, gm_n76, gm_n62, gm_n502, gm_n442);
	nor (gm_n5500, gm_n105, gm_n72, in_17, gm_n5499, gm_n374);
	nor (gm_n5501, gm_n227, gm_n73, gm_n59, gm_n520, gm_n263);
	nand (gm_n5502, gm_n113, gm_n72, gm_n85, gm_n5501);
	and (gm_n5503, gm_n221, in_16, in_12, gm_n1947, gm_n264);
	nand (gm_n5504, gm_n113, gm_n72, in_20, gm_n5503);
	and (gm_n5505, gm_n122, gm_n72, gm_n55, gm_n1687, gm_n254);
	nand (gm_n5506, gm_n545, gm_n60, gm_n63, gm_n1120, gm_n1942);
	nor (gm_n5507, in_21, in_20, gm_n56, gm_n5506, gm_n74);
	nand (gm_n5508, gm_n436, gm_n146, in_18, gm_n5294);
	nor (gm_n5509, gm_n461, gm_n76, in_9, gm_n621, gm_n430);
	nand (gm_n5510, gm_n255, in_21, in_17, gm_n5509, gm_n327);
	or (gm_n5511, gm_n115, gm_n73, gm_n59, gm_n835, gm_n385);
	nor (gm_n5512, gm_n139, gm_n72, in_20, gm_n5511);
	nand (gm_n5513, gm_n192, in_15, gm_n63, gm_n1120, gm_n1942);
	nor (gm_n5514, in_21, in_20, in_19, gm_n5513, gm_n1331);
	and (gm_n5515, gm_n448, gm_n222, gm_n60, gm_n2443, gm_n449);
	nand (gm_n5516, gm_n72, in_20, in_19, gm_n5515);
	nor (gm_n5517, gm_n263, in_16, in_12, gm_n1965, gm_n319);
	nand (gm_n5518, gm_n57, in_21, in_20, gm_n5517);
	or (gm_n5519, gm_n274, gm_n193, in_15, gm_n520, gm_n293);
	nor (gm_n5520, gm_n72, gm_n85, in_19, gm_n5519);
	nor (gm_n5521, gm_n90, in_10, in_9, gm_n3402, gm_n147);
	and (gm_n5522, gm_n243, gm_n88, in_18, gm_n5521);
	nor (gm_n5523, gm_n155, in_13, in_12, gm_n1751);
	nand (gm_n5524, gm_n120, in_21, gm_n55, gm_n5523, gm_n405);
	nor (gm_n5525, gm_n207, gm_n90, in_10, gm_n491, gm_n286);
	nand (gm_n5526, gm_n166, gm_n146, gm_n119, gm_n5525);
	nand (gm_n5527, gm_n448, gm_n222, gm_n60, gm_n953, gm_n545);
	nor (gm_n5528, gm_n72, in_20, in_19, gm_n5527);
	and (gm_n5529, gm_n348, gm_n131, in_18, gm_n2268);
	nor (gm_n5530, gm_n196, gm_n190, gm_n60, gm_n760, gm_n269);
	nand (gm_n5531, gm_n72, in_20, in_19, gm_n5530);
	nor (gm_n5532, gm_n406, in_13, in_9, gm_n503, gm_n502);
	nand (gm_n5533, gm_n102, in_21, gm_n55, gm_n5532, gm_n339);
	nand (gm_n5534, gm_n107, gm_n76, gm_n62, gm_n340, gm_n187);
	nor (gm_n5535, gm_n388, in_21, in_17, gm_n5534, gm_n328);
	nor (gm_n5536, gm_n479, gm_n72, in_17, gm_n2562, gm_n328);
	and (gm_n5537, gm_n523, gm_n2193, gm_n76, gm_n490, gm_n314);
	nand (gm_n5538, gm_n102, gm_n72, in_17, gm_n5537);
	nor (gm_n5539, gm_n292, gm_n213, in_15, gm_n633, gm_n447);
	nand (gm_n5540, gm_n72, gm_n85, in_19, gm_n5539);
	nand (gm_n5541, gm_n545, gm_n60, in_11, gm_n2074, gm_n1942);
	nor (gm_n5542, gm_n72, in_20, in_19, gm_n5541, gm_n447);
	or (gm_n5543, gm_n358, gm_n76, gm_n62, gm_n345, gm_n344);
	nor (gm_n5544, gm_n479, gm_n72, gm_n55, gm_n5543, gm_n662);
	nor (gm_n5545, gm_n159, gm_n60, in_11, gm_n271, gm_n270);
	nand (gm_n5546, in_21, gm_n85, gm_n56, gm_n5545, gm_n379);
	nand (gm_n5547, gm_n131, gm_n86, in_18, gm_n5521);
	nor (gm_n5548, gm_n485, gm_n263, in_15, gm_n3440, gm_n764);
	nand (gm_n5549, gm_n72, gm_n85, in_19, gm_n5548);
	nor (gm_n5550, gm_n115, gm_n73, in_12, gm_n1689, gm_n152);
	nand (gm_n5551, gm_n697, in_21, gm_n85, gm_n5550);
	or (gm_n5552, gm_n202, gm_n67, in_8, gm_n263);
	nor (gm_n5553, gm_n191, gm_n56, gm_n60, gm_n5552, gm_n643);
	nand (gm_n5554, gm_n5553, gm_n72, gm_n85);
	nand (gm_n5555, gm_n5549, gm_n5547, gm_n5546, gm_n5554, gm_n5551);
	and (gm_n5556, gm_n126, gm_n76, gm_n62, gm_n186, gm_n185);
	nand (gm_n5557, gm_n102, in_21, gm_n55, gm_n5556, gm_n122);
	nand (gm_n5558, gm_n174, gm_n72, in_17, gm_n2529, gm_n523);
	nand (gm_n5559, gm_n383, in_21, in_20, gm_n2940);
	nand (gm_n5560, gm_n5559, gm_n5558, gm_n5557);
	nand (gm_n5561, gm_n72, in_20, gm_n56, gm_n3441, gm_n268);
	nor (gm_n5562, in_14, gm_n78, in_9, gm_n2963, gm_n362);
	nand (gm_n5563, gm_n367, gm_n131, gm_n119, gm_n5562);
	nor (gm_n5564, gm_n155, in_16, gm_n59, gm_n3382, gm_n354);
	nand (gm_n5565, gm_n138, gm_n72, gm_n85, gm_n5564);
	nand (gm_n5566, gm_n5565, gm_n5563, gm_n5561);
	nor (gm_n5567, gm_n5555, gm_n5544, gm_n5542, gm_n5566, gm_n5560);
	nor (gm_n5568, gm_n121, gm_n72, in_17, gm_n3443, gm_n388);
	nand (gm_n5569, gm_n392, in_15, gm_n63, gm_n1615, gm_n1144);
	nor (gm_n5570, gm_n72, gm_n85, in_19, gm_n5569, gm_n393);
	or (gm_n5571, gm_n358, gm_n76, in_9, gm_n462, gm_n344);
	nor (gm_n5572, gm_n388, gm_n72, gm_n55, gm_n5571, gm_n256);
	nor (gm_n5573, gm_n5572, gm_n5570, gm_n5568);
	nand (gm_n5574, gm_n90, gm_n78, in_9, gm_n1446, gm_n1158);
	nor (gm_n5575, gm_n165, gm_n89, in_18, gm_n5574);
	nand (gm_n5576, gm_n2719, gm_n60, in_11, gm_n449, gm_n171);
	nor (gm_n5577, in_21, in_20, in_19, gm_n5576, gm_n293);
	or (gm_n5578, gm_n269, gm_n115, gm_n60, gm_n2038, gm_n760);
	nor (gm_n5579, in_21, gm_n85, gm_n56, gm_n5578);
	nor (gm_n5580, gm_n5579, gm_n5577, gm_n5575);
	nand (gm_n5581, gm_n5567, gm_n5540, gm_n5538, gm_n5580, gm_n5573);
	nor (gm_n5582, gm_n297, gm_n73, gm_n59, gm_n3315, gm_n354);
	nand (gm_n5583, gm_n138, in_21, in_20, gm_n5582);
	and (gm_n5584, gm_n214, gm_n73, gm_n59, gm_n2942, gm_n275);
	nand (gm_n5585, gm_n296, in_21, in_20, gm_n5584);
	nand (gm_n5586, gm_n311, gm_n72, gm_n55, gm_n4669, gm_n405);
	nand (gm_n5587, gm_n5586, gm_n5585, gm_n5583);
	nor (gm_n5588, gm_n344, in_13, in_9, gm_n1583, gm_n442);
	nand (gm_n5589, gm_n122, in_21, gm_n55, gm_n5588, gm_n254);
	nor (gm_n5590, gm_n667, in_13, in_9, gm_n462, gm_n480);
	nand (gm_n5591, gm_n174, gm_n72, in_17, gm_n5590, gm_n523);
	nor (gm_n5592, in_14, gm_n78, gm_n62, gm_n562, gm_n92);
	nand (gm_n5593, gm_n199, gm_n166, in_18, gm_n5592);
	nand (gm_n5594, gm_n5593, gm_n5591, gm_n5589);
	nor (gm_n5595, gm_n5581, gm_n5536, gm_n5535, gm_n5594, gm_n5587);
	or (gm_n5596, gm_n263, gm_n73, in_12, gm_n2125, gm_n276);
	nor (gm_n5597, gm_n384, gm_n72, in_20, gm_n5596);
	or (gm_n5598, gm_n247, gm_n90, gm_n78, gm_n376, gm_n369);
	nor (gm_n5599, gm_n212, gm_n87, gm_n119, gm_n5598);
	nor (gm_n5600, gm_n121, gm_n72, gm_n55, gm_n3356, gm_n441);
	nor (gm_n5601, gm_n5600, gm_n5599, gm_n5597);
	or (gm_n5602, gm_n297, in_16, gm_n59, gm_n3929, gm_n385);
	nor (gm_n5603, gm_n384, gm_n72, in_20, gm_n5602);
	nor (gm_n5604, gm_n374, gm_n72, gm_n55, gm_n1907, gm_n375);
	nor (gm_n5605, gm_n312, in_21, in_17, gm_n3524, gm_n328);
	nor (gm_n5606, gm_n5605, gm_n5604, gm_n5603);
	nand (gm_n5607, gm_n5595, gm_n5533, gm_n5531, gm_n5606, gm_n5601);
	and (gm_n5608, gm_n76, gm_n59, in_11, gm_n1942, gm_n176);
	nand (gm_n5609, gm_n86, in_18, gm_n90, gm_n5608, gm_n166);
	nor (gm_n5610, gm_n298, gm_n155, gm_n60, gm_n633, gm_n447);
	nand (gm_n5611, in_21, gm_n85, in_19, gm_n5610);
	nor (gm_n5612, gm_n414, gm_n406, gm_n76, gm_n491);
	nand (gm_n5613, gm_n102, gm_n72, gm_n55, gm_n5612, gm_n104);
	nand (gm_n5614, gm_n5613, gm_n5611, gm_n5609);
	nor (gm_n5615, gm_n147, in_14, in_10, gm_n376, gm_n148);
	nand (gm_n5616, gm_n367, gm_n806, gm_n119, gm_n5615);
	nor (gm_n5617, gm_n227, in_16, gm_n59, gm_n2221, gm_n158);
	nand (gm_n5618, gm_n495, gm_n72, in_20, gm_n5617);
	nor (gm_n5619, gm_n406, gm_n76, in_9, gm_n743, gm_n596);
	nand (gm_n5620, gm_n206, gm_n72, in_17, gm_n5619, gm_n1076);
	nand (gm_n5621, gm_n5620, gm_n5618, gm_n5616);
	nor (gm_n5622, gm_n5607, gm_n5529, gm_n5528, gm_n5621, gm_n5614);
	or (gm_n5623, gm_n977, gm_n60, gm_n63, gm_n760, gm_n270);
	nor (gm_n5624, in_21, in_20, gm_n56, gm_n5623, gm_n191);
	and (gm_n5625, gm_n327, in_21, in_17, gm_n610, gm_n339);
	or (gm_n5626, gm_n115, gm_n73, gm_n59, gm_n932, gm_n319);
	nor (gm_n5627, gm_n139, in_21, in_20, gm_n5626);
	nor (gm_n5628, gm_n5627, gm_n5625, gm_n5624);
	nand (gm_n5629, gm_n76, in_9, gm_n94, gm_n1263, gm_n123);
	nor (gm_n5630, gm_n479, gm_n72, gm_n55, gm_n5629, gm_n256);
	and (gm_n5631, gm_n138, in_21, gm_n85, gm_n4155);
	nand (gm_n5632, gm_n484, gm_n60, in_11, gm_n1120, gm_n1144);
	nor (gm_n5633, in_21, gm_n85, gm_n56, gm_n5632, gm_n393);
	nor (gm_n5634, gm_n5633, gm_n5631, gm_n5630);
	nand (gm_n5635, gm_n5622, gm_n5526, gm_n5524, gm_n5634, gm_n5628);
	nor (gm_n5636, gm_n115, gm_n73, in_12, gm_n3638, gm_n385);
	nand (gm_n5637, gm_n113, in_21, gm_n85, gm_n5636);
	nand (gm_n5638, gm_n206, gm_n72, in_17, gm_n2777, gm_n339);
	and (gm_n5639, gm_n126, in_13, in_9, gm_n402, gm_n341);
	nand (gm_n5640, gm_n122, gm_n72, in_17, gm_n5639, gm_n311);
	nand (gm_n5641, gm_n5640, gm_n5638, gm_n5637);
	nor (gm_n5642, gm_n438, in_14, in_10, gm_n526, gm_n467);
	nand (gm_n5643, gm_n245, gm_n164, gm_n119, gm_n5642);
	nor (gm_n5644, gm_n270, gm_n60, gm_n63, gm_n605, gm_n764);
	nand (gm_n5645, gm_n72, in_20, in_19, gm_n5644, gm_n486);
	nor (gm_n5646, gm_n238, gm_n228, gm_n977, gm_n807, gm_n313);
	nand (gm_n5647, gm_n254, gm_n72, gm_n55, gm_n5646);
	nand (gm_n5648, gm_n5647, gm_n5645, gm_n5643);
	nor (gm_n5649, gm_n5635, gm_n5522, gm_n5520, gm_n5648, gm_n5641);
	or (gm_n5650, gm_n370, in_14, in_10, gm_n467, gm_n414);
	nor (gm_n5651, gm_n165, gm_n89, in_18, gm_n5650);
	nand (gm_n5652, gm_n77, in_16, in_12, gm_n82, gm_n79);
	nor (gm_n5653, gm_n139, gm_n72, in_20, gm_n5652);
	nor (gm_n5654, gm_n183, gm_n72, in_17, gm_n876, gm_n313);
	nor (gm_n5655, gm_n5654, gm_n5653, gm_n5651);
	and (gm_n5656, gm_n255, gm_n72, in_17, gm_n5071, gm_n311);
	or (gm_n5657, gm_n148, in_14, in_10, gm_n376, gm_n807);
	nor (gm_n5658, gm_n531, gm_n212, gm_n119, gm_n5657);
	nand (gm_n5659, gm_n122, gm_n76, gm_n62, gm_n427, gm_n123);
	nor (gm_n5660, gm_n479, in_21, gm_n55, gm_n5659);
	nor (gm_n5661, gm_n5660, gm_n5658, gm_n5656);
	nand (gm_n5662, gm_n5649, gm_n5518, gm_n5516, gm_n5661, gm_n5655);
	nor (gm_n5663, gm_n190, gm_n73, in_12, gm_n1246, gm_n152);
	nand (gm_n5664, gm_n697, in_21, in_20, gm_n5663);
	nor (gm_n5665, gm_n155, gm_n73, in_12, gm_n808, gm_n319);
	nand (gm_n5666, gm_n138, in_21, gm_n85, gm_n5665);
	nor (gm_n5667, gm_n240, in_15, gm_n63, gm_n842, gm_n633);
	nand (gm_n5668, in_21, in_20, gm_n56, gm_n5667, gm_n268);
	nand (gm_n5669, gm_n5668, gm_n5666, gm_n5664);
	and (gm_n5670, gm_n126, gm_n76, in_9, gm_n788, gm_n186);
	nand (gm_n5671, gm_n174, gm_n72, gm_n55, gm_n5670, gm_n523);
	nor (gm_n5672, gm_n461, in_13, in_9, gm_n2198, gm_n375);
	nand (gm_n5673, gm_n327, gm_n72, gm_n55, gm_n5672);
	nor (gm_n5674, gm_n461, gm_n76, gm_n62, gm_n597, gm_n430);
	nand (gm_n5675, gm_n122, gm_n72, in_17, gm_n5674, gm_n206);
	nand (gm_n5676, gm_n5675, gm_n5673, gm_n5671);
	nor (gm_n5677, gm_n5662, gm_n5514, gm_n5512, gm_n5676, gm_n5669);
	nand (gm_n5678, gm_n394, gm_n143, in_15, gm_n1416, gm_n545);
	nor (gm_n5679, gm_n72, gm_n85, gm_n56, gm_n5678);
	or (gm_n5680, gm_n358, gm_n76, in_9, gm_n463, gm_n866);
	nor (gm_n5681, gm_n479, gm_n72, in_17, gm_n5680, gm_n328);
	nand (gm_n5682, gm_n602, gm_n91, gm_n90, gm_n1120);
	nor (gm_n5683, gm_n244, gm_n212, in_18, gm_n5682);
	nor (gm_n5684, gm_n5683, gm_n5681, gm_n5679);
	or (gm_n5685, gm_n148, gm_n99, in_13, gm_n442);
	nor (gm_n5686, gm_n103, in_21, gm_n55, gm_n5685, gm_n105);
	nand (gm_n5687, gm_n392, gm_n79, in_15, gm_n423, gm_n1101);
	nor (gm_n5688, in_21, in_20, in_19, gm_n5687);
	and (gm_n5689, gm_n122, in_21, gm_n55, gm_n5314, gm_n373);
	nor (gm_n5690, gm_n5689, gm_n5688, gm_n5686);
	nand (gm_n5691, gm_n5677, gm_n5510, gm_n5508, gm_n5690, gm_n5684);
	and (gm_n5692, gm_n64, in_16, gm_n59, gm_n5152, gm_n221);
	nand (gm_n5693, gm_n495, gm_n72, gm_n85, gm_n5692);
	and (gm_n5694, in_14, in_10, in_9, gm_n1501, gm_n532);
	nand (gm_n5695, gm_n323, gm_n164, gm_n119, gm_n5694);
	nor (gm_n5696, gm_n155, in_16, in_12, gm_n3315, gm_n220);
	nand (gm_n5697, gm_n138, gm_n72, in_20, gm_n5696);
	nand (gm_n5698, gm_n5697, gm_n5695, gm_n5693);
	nor (gm_n5699, gm_n213, in_15, gm_n94, gm_n764, gm_n508);
	nand (gm_n5700, in_21, gm_n85, gm_n56, gm_n5699, gm_n486);
	and (gm_n5701, gm_n449, gm_n60, gm_n63, gm_n1929, gm_n1942);
	nand (gm_n5702, gm_n72, in_20, gm_n56, gm_n5701, gm_n268);
	nor (gm_n5703, gm_n345, in_13, in_9, gm_n502, gm_n480);
	nand (gm_n5704, gm_n311, in_21, in_17, gm_n5703, gm_n405);
	nand (gm_n5705, gm_n5704, gm_n5702, gm_n5700);
	nor (gm_n5706, gm_n5691, gm_n5507, gm_n5505, gm_n5705, gm_n5698);
	or (gm_n5707, gm_n358, gm_n76, in_9, gm_n1583, gm_n463);
	nor (gm_n5708, gm_n441, gm_n72, in_17, gm_n5707, gm_n328);
	or (gm_n5709, gm_n274, in_16, gm_n59, gm_n2826, gm_n276);
	nor (gm_n5710, gm_n496, in_21, in_20, gm_n5709);
	or (gm_n5711, gm_n596, in_13, in_9, gm_n462, gm_n442);
	nor (gm_n5712, gm_n388, in_21, gm_n55, gm_n5711, gm_n313);
	nor (gm_n5713, gm_n5712, gm_n5710, gm_n5708);
	or (gm_n5714, gm_n207, in_14, gm_n78, gm_n370, gm_n208);
	nor (gm_n5715, gm_n89, gm_n87, gm_n119, gm_n5714);
	and (gm_n5716, gm_n233, in_13, gm_n59, gm_n142);
	and (gm_n5717, gm_n174, gm_n72, gm_n55, gm_n5716, gm_n255);
	nand (gm_n5718, gm_n828, gm_n90, gm_n78, gm_n829, gm_n624);
	nor (gm_n5719, gm_n841, gm_n87, gm_n119, gm_n5718);
	nor (gm_n5720, gm_n5719, gm_n5717, gm_n5715);
	nand (gm_n5721, gm_n5706, gm_n5504, gm_n5502, gm_n5720, gm_n5713);
	nor (gm_n5722, gm_n78, in_9, in_8, gm_n981, gm_n133);
	nand (gm_n5723, gm_n245, in_18, gm_n90, gm_n5722, gm_n367);
	nor (gm_n5724, in_10, in_9, gm_n94, gm_n1631, gm_n147);
	nand (gm_n5725, gm_n86, in_18, gm_n90, gm_n5724, gm_n806);
	nor (gm_n5726, gm_n609, gm_n76, in_9, gm_n481, gm_n461);
	nand (gm_n5727, gm_n120, in_21, gm_n55, gm_n5726, gm_n339);
	nand (gm_n5728, gm_n5727, gm_n5725, gm_n5723);
	nor (gm_n5729, gm_n155, in_16, gm_n59, gm_n1661, gm_n319);
	nand (gm_n5730, gm_n57, gm_n72, in_20, gm_n5729);
	nor (gm_n5731, gm_n133, in_14, in_10, gm_n287, gm_n149);
	nand (gm_n5732, gm_n436, gm_n146, gm_n119, gm_n5731);
	nor (gm_n5733, gm_n213, gm_n73, gm_n59, gm_n799, gm_n220);
	nand (gm_n5734, gm_n296, in_21, in_20, gm_n5733);
	nand (gm_n5735, gm_n5734, gm_n5732, gm_n5730);
	nor (gm_n5736, gm_n5721, gm_n5500, gm_n5498, gm_n5735, gm_n5728);
	or (gm_n5737, gm_n369, gm_n283, gm_n90, gm_n842);
	nor (gm_n5738, gm_n244, gm_n89, in_18, gm_n5737);
	nand (gm_n5739, gm_n264, gm_n60, gm_n94, gm_n1398, gm_n455);
	nor (gm_n5740, gm_n72, in_20, in_19, gm_n5739, gm_n293);
	or (gm_n5741, gm_n1331, gm_n115, in_15, gm_n2008, gm_n764);
	nor (gm_n5742, gm_n72, gm_n85, in_19, gm_n5741);
	nor (gm_n5743, gm_n5742, gm_n5740, gm_n5738);
	or (gm_n5744, gm_n358, gm_n76, in_9, gm_n443, gm_n345);
	nor (gm_n5745, gm_n184, in_21, gm_n55, gm_n5744, gm_n374);
	or (gm_n5746, gm_n430, in_13, gm_n62, gm_n442, gm_n432);
	nor (gm_n5747, gm_n105, gm_n72, in_17, gm_n5746, gm_n183);
	or (gm_n5748, gm_n362, gm_n841, gm_n90, gm_n1382, gm_n980);
	nor (gm_n5749, gm_n5748, gm_n87, gm_n119);
	nor (gm_n5750, gm_n5749, gm_n5747, gm_n5745);
	nand (gm_n5751, gm_n5736, gm_n5496, gm_n5494, gm_n5750, gm_n5743);
	nand (gm_n5752, gm_n174, gm_n72, gm_n55, gm_n4669, gm_n339);
	and (gm_n5753, gm_n64, in_16, in_12, gm_n3587, gm_n275);
	nand (gm_n5754, gm_n697, in_21, in_20, gm_n5753);
	nand (gm_n5755, gm_n102, in_21, in_17, gm_n4943, gm_n1076);
	nand (gm_n5756, gm_n5755, gm_n5754, gm_n5752);
	nor (gm_n5757, gm_n431, gm_n76, in_9, gm_n481, gm_n344);
	nand (gm_n5758, gm_n102, in_21, in_17, gm_n5757, gm_n122);
	nor (gm_n5759, gm_n114, gm_n73, gm_n59, gm_n2589, gm_n263);
	nand (gm_n5760, gm_n697, in_21, in_20, gm_n5759);
	nand (gm_n5761, gm_n129, t_5, in_18, gm_n806);
	nand (gm_n5762, gm_n5761, gm_n5760, gm_n5758);
	nor (gm_n5763, gm_n5751, gm_n5492, gm_n5490, gm_n5762, gm_n5756);
	nand (gm_n5764, gm_n91, gm_n90, in_10, gm_n793, gm_n1345);
	nor (gm_n5765, gm_n368, gm_n246, gm_n119, gm_n5764);
	or (gm_n5766, in_14, in_10, gm_n62, gm_n1319, gm_n207);
	nor (gm_n5767, gm_n368, gm_n841, gm_n119, gm_n5766);
	nand (gm_n5768, gm_n713, gm_n131, gm_n90, gm_n1928, gm_n601);
	nor (gm_n5769, gm_n5768, gm_n244, gm_n119);
	nor (gm_n5770, gm_n5769, gm_n5767, gm_n5765);
	or (gm_n5771, gm_n431, in_13, in_9, gm_n621, gm_n463);
	nor (gm_n5772, gm_n103, gm_n72, in_17, gm_n5771, gm_n256);
	nand (gm_n5773, gm_n222, gm_n192, in_15, gm_n875, gm_n486);
	nor (gm_n5774, in_21, gm_n85, gm_n56, gm_n5773);
	nand (gm_n5775, gm_n90, in_10, gm_n62, gm_n1524, gm_n334);
	nor (gm_n5776, gm_n368, gm_n89, in_18, gm_n5775);
	nor (gm_n5777, gm_n5776, gm_n5774, gm_n5772);
	nand (gm_n5778, gm_n5763, gm_n5488, gm_n5486, gm_n5777, gm_n5770);
	nor (gm_n5779, in_14, in_10, gm_n62, gm_n1484, gm_n362);
	nand (gm_n5780, gm_n245, gm_n243, gm_n119, gm_n5779);
	nor (gm_n5781, gm_n90, gm_n78, gm_n62, gm_n1475, gm_n133);
	nand (gm_n5782, gm_n243, gm_n806, in_18, gm_n5781);
	or (gm_n5783, gm_n184, gm_n72, gm_n55, gm_n3459, gm_n374);
	nand (gm_n5784, gm_n5783, gm_n5782, gm_n5780);
	nor (gm_n5785, gm_n430, gm_n76, in_9, gm_n345, gm_n431);
	nand (gm_n5786, gm_n255, in_21, gm_n55, gm_n5785, gm_n327);
	nor (gm_n5787, gm_n480, in_13, in_9, gm_n988, gm_n443);
	nand (gm_n5788, gm_n122, gm_n72, in_17, gm_n5787, gm_n206);
	and (gm_n5789, gm_n1144, in_15, in_11, gm_n1398, gm_n601);
	nand (gm_n5790, in_21, gm_n85, gm_n56, gm_n5789, gm_n486);
	nand (gm_n5791, gm_n5790, gm_n5788, gm_n5786);
	nor (gm_n5792, gm_n5778, gm_n5485, gm_n5483, gm_n5791, gm_n5784);
	nor (gm_n5793, gm_n514, gm_n76, gm_n62, gm_n597, gm_n443);
	nand (gm_n5794, gm_n255, in_21, gm_n55, gm_n5793, gm_n327);
	nor (gm_n5795, gm_n190, gm_n73, gm_n59, gm_n815, gm_n227);
	nand (gm_n5796, gm_n495, in_21, in_20, gm_n5795);
	and (gm_n5797, gm_n486, gm_n222, gm_n60, gm_n1841, gm_n545);
	nand (gm_n5798, in_21, in_20, in_19, gm_n5797);
	nand (gm_n5799, gm_n5794, gm_n5792, gm_n5481, gm_n5798, gm_n5796);
	and (gm_n5800, gm_n448, gm_n222, in_15, gm_n1161, gm_n869);
	nand (gm_n5801, gm_n72, in_20, in_19, gm_n5800);
	nor (gm_n5802, gm_n90, in_10, gm_n62, gm_n821, gm_n147);
	nand (gm_n5803, gm_n131, gm_n129, in_18, gm_n5802);
	nor (gm_n5804, gm_n662, gm_n247, gm_n76, gm_n414, gm_n406);
	nand (gm_n5805, gm_n327, gm_n72, in_17, gm_n5804);
	nand (gm_n5806, gm_n5805, gm_n5803, gm_n5801);
	or (gm_n5807, gm_n220, gm_n73, gm_n59, gm_n887, gm_n263);
	nor (gm_n5808, gm_n384, gm_n72, in_20, gm_n5807);
	nor (out_16, gm_n5806, gm_n5799, gm_n5479, gm_n5808);
	or (gm_n5810, gm_n461, gm_n76, gm_n62, gm_n597, gm_n463);
	nor (gm_n5811, gm_n256, gm_n72, in_17, gm_n5810, gm_n312);
	or (gm_n5812, gm_n620, gm_n72, in_17, gm_n2850, gm_n328);
	nor (gm_n5813, in_10, gm_n62, gm_n94, gm_n761, gm_n369);
	nand (gm_n5814, gm_n131, in_18, in_14, gm_n5813, gm_n367);
	or (gm_n5815, gm_n667, gm_n76, in_9, gm_n597, gm_n431);
	nor (gm_n5816, gm_n441, gm_n72, in_17, gm_n5815, gm_n184);
	or (gm_n5817, gm_n190, gm_n73, in_12, gm_n3638, gm_n276);
	nor (gm_n5818, gm_n912, gm_n72, gm_n85, gm_n5817);
	nor (gm_n5819, gm_n359, gm_n76, in_9, gm_n443, gm_n442);
	nand (gm_n5820, gm_n104, gm_n72, gm_n55, gm_n5819, gm_n254);
	and (gm_n5821, gm_n264, in_16, gm_n59, gm_n2860, gm_n303);
	nand (gm_n5822, gm_n179, in_21, in_20, gm_n5821);
	or (gm_n5823, gm_n168, gm_n155, in_15, gm_n860, gm_n447);
	nor (gm_n5824, gm_n72, gm_n85, gm_n56, gm_n5823);
	or (gm_n5825, gm_n431, gm_n76, in_9, gm_n1664, gm_n328);
	nor (gm_n5826, gm_n479, gm_n72, gm_n55, gm_n5825);
	and (gm_n5827, gm_n123, gm_n76, in_9, gm_n341, gm_n187);
	nand (gm_n5828, gm_n174, gm_n72, gm_n55, gm_n5827, gm_n1076);
	nor (gm_n5829, gm_n114, in_16, gm_n59, gm_n3440, gm_n190);
	nand (gm_n5830, gm_n697, gm_n72, gm_n85, gm_n5829);
	and (gm_n5831, gm_n323, t_5, in_18, gm_n348);
	nand (gm_n5832, gm_n122, gm_n76, in_9, gm_n2283, gm_n402);
	nor (gm_n5833, gm_n103, in_21, in_17, gm_n5832);
	nand (gm_n5834, gm_n311, in_21, gm_n55, gm_n5405, gm_n1076);
	nor (gm_n5835, in_13, in_9, in_8, gm_n2769, gm_n406);
	nand (gm_n5836, gm_n254, in_21, in_17, gm_n5835, gm_n405);
	nand (gm_n5837, gm_n61, gm_n73, gm_n59, gm_n2605, gm_n79);
	nor (gm_n5838, gm_n781, in_21, gm_n85, gm_n5837);
	nand (gm_n5839, gm_n486, gm_n143, in_15, gm_n1392, gm_n1398);
	nor (gm_n5840, in_21, gm_n85, in_19, gm_n5839);
	nand (gm_n5841, gm_n104, in_21, in_17, gm_n4748, gm_n120);
	and (gm_n5842, gm_n79, in_16, gm_n59, gm_n1611, gm_n949);
	nand (gm_n5843, gm_n296, in_21, in_20, gm_n5842);
	nor (gm_n5844, gm_n121, gm_n72, gm_n55, gm_n1936, gm_n312);
	nand (gm_n5845, gm_n91, in_14, gm_n78, gm_n793, gm_n490);
	nor (gm_n5846, gm_n246, gm_n244, gm_n119, gm_n5845);
	nor (gm_n5847, in_14, in_10, in_9, gm_n1406, gm_n467);
	nand (gm_n5848, gm_n348, gm_n323, in_18, gm_n5847);
	nor (gm_n5849, in_14, in_10, in_9, gm_n2956, gm_n133);
	nand (gm_n5850, gm_n367, gm_n131, gm_n119, gm_n5849);
	nand (gm_n5851, gm_n76, in_9, gm_n94, gm_n556, gm_n402);
	nor (gm_n5852, gm_n184, gm_n72, in_17, gm_n5851, gm_n312);
	nand (gm_n5853, gm_n394, gm_n222, in_15, gm_n1147, gm_n869);
	nor (gm_n5854, gm_n72, gm_n85, gm_n56, gm_n5853);
	nor (gm_n5855, gm_n153, in_16, gm_n59, gm_n319, gm_n155);
	nand (gm_n5856, gm_n113, in_21, gm_n85, gm_n5855);
	nor (gm_n5857, gm_n213, in_16, gm_n59, gm_n2002, gm_n354);
	nand (gm_n5858, gm_n495, in_21, gm_n85, gm_n5857);
	or (gm_n5859, gm_n90, in_10, in_9, gm_n832, gm_n807);
	nor (gm_n5860, gm_n531, gm_n1989, in_18, gm_n5859);
	nand (gm_n5861, gm_n143, in_13, gm_n59, gm_n919);
	nor (gm_n5862, gm_n662, in_21, gm_n55, gm_n5861, gm_n374);
	nor (gm_n5863, gm_n667, gm_n76, gm_n62, gm_n480, gm_n345);
	nand (gm_n5864, gm_n104, in_21, gm_n55, gm_n5863, gm_n120);
	and (gm_n5865, gm_n547, gm_n422, gm_n143);
	nand (gm_n5866, gm_n164, gm_n88, gm_n119, gm_n5865);
	nand (gm_n5867, gm_n79, gm_n59, gm_n94, gm_n1379, gm_n221);
	nor (gm_n5868, in_21, gm_n85, in_16, gm_n5867, gm_n384);
	nand (gm_n5869, gm_n123, gm_n76, gm_n62, gm_n126, gm_n125);
	nor (gm_n5870, gm_n184, in_21, gm_n55, gm_n5869, gm_n479);
	nand (gm_n5871, gm_n436, gm_n367, gm_n119, gm_n459);
	nor (gm_n5872, gm_n213, gm_n73, in_12, gm_n821, gm_n220);
	nand (gm_n5873, gm_n383, gm_n72, gm_n85, gm_n5872);
	nand (gm_n5874, gm_n143, gm_n75, in_15, gm_n2624, gm_n869);
	nor (gm_n5875, gm_n72, gm_n85, gm_n56, gm_n5874);
	nor (gm_n5876, gm_n193, in_15, in_11, gm_n842, gm_n283);
	nand (gm_n5877, gm_n72, gm_n85, gm_n56, gm_n5876, gm_n486);
	nor (gm_n5878, gm_n447, gm_n158, in_15, gm_n1016, gm_n643);
	nand (gm_n5879, in_21, gm_n85, gm_n56, gm_n5878);
	and (gm_n5880, gm_n123, gm_n2193, in_13, gm_n995, gm_n523);
	nand (gm_n5881, gm_n254, gm_n72, gm_n55, gm_n5880);
	nand (gm_n5882, gm_n5881, gm_n5879, gm_n5877);
	or (gm_n5883, gm_n147, gm_n90, gm_n78, gm_n414, gm_n287);
	nor (gm_n5884, gm_n531, gm_n89, gm_n119, gm_n5883);
	nor (gm_n5885, gm_n67, gm_n59, in_8, gm_n194, gm_n115);
	nand (gm_n5886, gm_n119, gm_n55, gm_n73, gm_n5885, gm_n571);
	nor (gm_n5887, gm_n5886, gm_n531);
	nand (gm_n5888, gm_n77, gm_n73, in_12, gm_n636, gm_n264);
	nor (gm_n5889, gm_n384, gm_n72, gm_n85, gm_n5888);
	nor (gm_n5890, gm_n5884, gm_n5882, gm_n5875, gm_n5889, gm_n5887);
	or (gm_n5891, gm_n431, in_13, in_9, gm_n1583, gm_n463);
	nor (gm_n5892, gm_n103, gm_n72, gm_n55, gm_n5891, gm_n256);
	nand (gm_n5893, gm_n394, gm_n64, in_15, gm_n962, gm_n449);
	nor (gm_n5894, gm_n72, in_20, in_19, gm_n5893);
	nor (gm_n5895, gm_n912, in_21, gm_n85, gm_n3877);
	nor (gm_n5896, gm_n5895, gm_n5894, gm_n5892);
	nand (gm_n5897, gm_n186, gm_n76, gm_n62, gm_n402, gm_n316);
	nor (gm_n5898, gm_n183, gm_n72, gm_n55, gm_n5897, gm_n256);
	or (gm_n5899, gm_n909, in_15, gm_n63, gm_n633, gm_n977);
	nor (gm_n5900, in_21, gm_n85, in_19, gm_n5899, gm_n1331);
	nor (gm_n5901, gm_n441, in_21, in_17, gm_n4835, gm_n184);
	nor (gm_n5902, gm_n5901, gm_n5900, gm_n5898);
	nand (gm_n5903, gm_n5890, gm_n5873, gm_n5871, gm_n5902, gm_n5896);
	nor (gm_n5904, gm_n114, gm_n73, in_12, gm_n3315, gm_n297);
	nand (gm_n5905, gm_n697, gm_n72, gm_n85, gm_n5904);
	nor (gm_n5906, gm_n514, gm_n76, in_9, gm_n1132, gm_n667);
	nand (gm_n5907, gm_n254, gm_n72, gm_n55, gm_n5906, gm_n255);
	nor (gm_n5908, gm_n90, in_10, gm_n62, gm_n4975, gm_n92);
	nand (gm_n5909, gm_n436, gm_n348, in_18, gm_n5908);
	nand (gm_n5910, gm_n5909, gm_n5907, gm_n5905);
	nor (gm_n5911, gm_n213, gm_n73, in_12, gm_n675, gm_n385);
	nand (gm_n5912, gm_n179, in_21, gm_n85, gm_n5911);
	nand (gm_n5913, gm_n102, in_21, in_17, gm_n986, gm_n1076);
	nor (gm_n5914, gm_n407, gm_n369, in_14, gm_n605);
	nand (gm_n5915, gm_n348, gm_n131, in_18, gm_n5914);
	nand (gm_n5916, gm_n5915, gm_n5913, gm_n5912);
	nor (gm_n5917, gm_n5903, gm_n5870, gm_n5868, gm_n5916, gm_n5910);
	nand (gm_n5918, gm_n264, gm_n73, in_12, gm_n2683, gm_n275);
	nor (gm_n5919, gm_n262, gm_n72, gm_n85, gm_n5918);
	nand (gm_n5920, gm_n110, in_13, in_9, gm_n1049, gm_n402);
	nor (gm_n5921, gm_n183, gm_n72, in_17, gm_n5920, gm_n256);
	nand (gm_n5922, gm_n90, in_10, gm_n62, gm_n1079, gm_n91);
	nor (gm_n5923, gm_n1989, gm_n211, in_18, gm_n5922);
	nor (gm_n5924, gm_n5923, gm_n5921, gm_n5919);
	nand (gm_n5925, in_14, in_10, in_9, gm_n1071, gm_n532);
	nor (gm_n5926, gm_n437, gm_n165, in_18, gm_n5925);
	or (gm_n5927, gm_n514, gm_n76, gm_n62, gm_n988, gm_n609);
	nor (gm_n5928, gm_n103, gm_n72, in_17, gm_n5927, gm_n328);
	nand (gm_n5929, gm_n78, gm_n62, in_8, gm_n1120, gm_n532);
	nor (gm_n5930, gm_n132, in_18, gm_n90, gm_n5929, gm_n211);
	nor (gm_n5931, gm_n5930, gm_n5928, gm_n5926);
	nand (gm_n5932, gm_n5917, gm_n5866, gm_n5864, gm_n5931, gm_n5924);
	nor (gm_n5933, gm_n90, in_10, gm_n62, gm_n2474, gm_n133);
	nand (gm_n5934, gm_n166, gm_n86, in_18, gm_n5933);
	nor (gm_n5935, gm_n485, gm_n213, gm_n60, gm_n633, gm_n520);
	nand (gm_n5936, gm_n72, gm_n85, gm_n56, gm_n5935);
	nor (gm_n5937, gm_n92, gm_n90, gm_n78, gm_n376, gm_n370);
	nand (gm_n5938, gm_n348, gm_n323, gm_n119, gm_n5937);
	nand (gm_n5939, gm_n5938, gm_n5936, gm_n5934);
	nor (gm_n5940, gm_n105, gm_n76, gm_n62, gm_n3721, gm_n431);
	nand (gm_n5941, gm_n254, in_21, gm_n55, gm_n5940);
	and (gm_n5942, gm_n422, gm_n60, gm_n63, gm_n2074, gm_n555);
	nand (gm_n5943, gm_n72, gm_n85, in_19, gm_n5942, gm_n394);
	nor (gm_n5944, gm_n447, gm_n115, gm_n60, gm_n1170, gm_n764);
	nand (gm_n5945, gm_n72, gm_n85, in_19, gm_n5944);
	nand (gm_n5946, gm_n5945, gm_n5943, gm_n5941);
	nor (gm_n5947, gm_n5932, gm_n5862, gm_n5860, gm_n5946, gm_n5939);
	nand (gm_n5948, gm_n143, gm_n73, in_12, gm_n825, gm_n221);
	nor (gm_n5949, gm_n219, in_21, gm_n85, gm_n5948);
	or (gm_n5950, gm_n358, in_13, in_9, gm_n743, gm_n344);
	nor (gm_n5951, gm_n479, gm_n72, gm_n55, gm_n5950, gm_n256);
	or (gm_n5952, gm_n95, in_14, gm_n78, gm_n350, gm_n147);
	nor (gm_n5953, gm_n437, gm_n87, in_18, gm_n5952);
	nor (gm_n5954, gm_n5953, gm_n5951, gm_n5949);
	nand (gm_n5955, gm_n64, gm_n73, in_12, gm_n1147, gm_n733);
	nor (gm_n5956, gm_n219, in_21, gm_n85, gm_n5955);
	nand (gm_n5957, gm_n79, gm_n75, gm_n60, gm_n1758, gm_n484);
	nor (gm_n5958, in_21, gm_n85, gm_n56, gm_n5957);
	nand (gm_n5959, gm_n64, in_16, gm_n59, gm_n4011, gm_n571);
	nor (gm_n5960, gm_n58, gm_n72, in_20, gm_n5959);
	nor (gm_n5961, gm_n5960, gm_n5958, gm_n5956);
	nand (gm_n5962, gm_n5947, gm_n5858, gm_n5856, gm_n5961, gm_n5954);
	nor (gm_n5963, in_14, gm_n78, gm_n62, gm_n832, gm_n467);
	nand (gm_n5964, gm_n199, gm_n131, in_18, gm_n5963);
	nor (gm_n5965, gm_n257, in_13, in_9, gm_n597, gm_n596);
	nand (gm_n5966, gm_n311, gm_n72, in_17, gm_n5965, gm_n595);
	and (gm_n5967, gm_n90, in_10, gm_n62, gm_n2624, gm_n334);
	nand (gm_n5968, gm_n131, gm_n86, gm_n119, gm_n5967);
	nand (gm_n5969, gm_n5968, gm_n5966, gm_n5964);
	and (gm_n5970, gm_n104, gm_n2193, in_13, gm_n490, gm_n402);
	nand (gm_n5971, gm_n120, gm_n72, in_17, gm_n5970);
	nand (gm_n5972, gm_n104, in_21, in_17, gm_n2317, gm_n327);
	and (gm_n5973, gm_n392, gm_n60, gm_n63, gm_n602, gm_n576);
	nand (gm_n5974, gm_n72, in_20, in_19, gm_n5973, gm_n394);
	nand (gm_n5975, gm_n5974, gm_n5972, gm_n5971);
	nor (gm_n5976, gm_n5962, gm_n5854, gm_n5852, gm_n5975, gm_n5969);
	and (gm_n5977, gm_n806, gm_n146, in_18, gm_n5865);
	or (gm_n5978, gm_n90, gm_n78, in_9, gm_n2402, gm_n207);
	nor (gm_n5979, gm_n246, gm_n244, gm_n119, gm_n5978);
	nand (gm_n5980, gm_n64, in_16, gm_n59, gm_n1524, gm_n571);
	nor (gm_n5981, gm_n781, gm_n72, in_20, gm_n5980);
	nor (gm_n5982, gm_n5981, gm_n5979, gm_n5977);
	or (gm_n5983, gm_n95, gm_n90, in_10, gm_n362, gm_n99);
	nor (gm_n5984, gm_n244, gm_n212, in_18, gm_n5983);
	nand (gm_n5985, gm_n314, gm_n76, gm_n62, gm_n427, gm_n595);
	nor (gm_n5986, gm_n374, gm_n72, gm_n55, gm_n5985);
	nand (gm_n5987, in_14, gm_n78, gm_n62, gm_n3063, gm_n624);
	nor (gm_n5988, gm_n244, gm_n89, in_18, gm_n5987);
	nor (gm_n5989, gm_n5988, gm_n5986, gm_n5984);
	nand (gm_n5990, gm_n5976, gm_n5850, gm_n5848, gm_n5989, gm_n5982);
	nor (gm_n5991, gm_n667, in_13, gm_n62, gm_n462, gm_n257);
	nand (gm_n5992, gm_n104, gm_n72, gm_n55, gm_n5991, gm_n373);
	and (gm_n5993, gm_n90, gm_n76, gm_n59, gm_n1001, gm_n154);
	nand (gm_n5994, gm_n146, gm_n88, in_18, gm_n5993);
	nor (gm_n5995, gm_n358, in_13, in_9, gm_n432, gm_n344);
	nand (gm_n5996, gm_n327, gm_n72, in_17, gm_n5995, gm_n339);
	nand (gm_n5997, gm_n5996, gm_n5994, gm_n5992);
	and (gm_n5998, in_14, in_10, gm_n62, gm_n3063, gm_n1011);
	nand (gm_n5999, gm_n88, gm_n86, in_18, gm_n5998);
	nor (gm_n6000, gm_n344, gm_n76, in_9, gm_n481, gm_n480);
	nand (gm_n6001, gm_n255, gm_n72, gm_n55, gm_n6000, gm_n311);
	and (gm_n6002, gm_n233, gm_n75, gm_n60, gm_n2065, gm_n422);
	nand (gm_n6003, gm_n72, in_20, gm_n56, gm_n6002);
	nand (gm_n6004, gm_n6003, gm_n6001, gm_n5999);
	nor (gm_n6005, gm_n5990, gm_n5846, gm_n5844, gm_n6004, gm_n5997);
	or (gm_n6006, gm_n818, gm_n76, in_9, gm_n502, gm_n406);
	nor (gm_n6007, gm_n388, gm_n72, gm_n55, gm_n6006, gm_n256);
	or (gm_n6008, gm_n155, in_12, gm_n94, gm_n2769, gm_n276);
	nor (gm_n6009, in_21, in_20, in_16, gm_n6008, gm_n496);
	or (gm_n6010, gm_n358, gm_n76, gm_n62, gm_n796, gm_n667);
	nor (gm_n6011, gm_n184, gm_n72, gm_n55, gm_n6010, gm_n374);
	nor (gm_n6012, gm_n6011, gm_n6009, gm_n6007);
	or (gm_n6013, gm_n92, gm_n90, in_10, gm_n589, gm_n95);
	nor (gm_n6014, gm_n244, gm_n841, gm_n119, gm_n6013);
	nand (gm_n6015, gm_n79, in_16, in_12, gm_n936, gm_n571);
	nor (gm_n6016, gm_n219, in_21, in_20, gm_n6015);
	or (gm_n6017, gm_n431, gm_n76, gm_n62, gm_n443, gm_n345);
	nor (gm_n6018, gm_n256, gm_n72, in_17, gm_n6017, gm_n374);
	nor (gm_n6019, gm_n6018, gm_n6016, gm_n6014);
	nand (gm_n6020, gm_n6005, gm_n5843, gm_n5841, gm_n6019, gm_n6012);
	and (gm_n6021, gm_n125, in_13, gm_n62, gm_n579, gm_n126);
	nand (gm_n6022, gm_n174, in_21, in_17, gm_n6021, gm_n405);
	nor (gm_n6023, gm_n796, in_13, gm_n62, gm_n463, gm_n257);
	nand (gm_n6024, gm_n122, gm_n72, gm_n55, gm_n6023, gm_n206);
	nor (gm_n6025, gm_n431, gm_n76, in_9, gm_n621, gm_n502);
	nand (gm_n6026, gm_n104, in_21, gm_n55, gm_n6025, gm_n373);
	nand (gm_n6027, gm_n6026, gm_n6024, gm_n6022);
	nand (gm_n6028, gm_n327, in_21, in_17, gm_n1076, gm_n336);
	nor (gm_n6029, gm_n667, in_13, in_9, gm_n432, gm_n480);
	nand (gm_n6030, gm_n254, gm_n72, gm_n55, gm_n6029, gm_n595);
	nor (gm_n6031, gm_n168, gm_n60, in_11, gm_n842, gm_n283);
	nand (gm_n6032, gm_n72, in_20, in_19, gm_n6031, gm_n281);
	nand (gm_n6033, gm_n6032, gm_n6030, gm_n6028);
	nor (gm_n6034, gm_n6020, gm_n5840, gm_n5838, gm_n6033, gm_n6027);
	nor (gm_n6035, gm_n184, in_21, gm_n55, gm_n4424, gm_n620);
	nand (gm_n6036, gm_n733, gm_n73, in_12, gm_n1456, gm_n222);
	nor (gm_n6037, gm_n58, gm_n72, gm_n85, gm_n6036);
	nand (gm_n6038, gm_n1144, in_15, gm_n63, gm_n714, gm_n422);
	nor (gm_n6039, in_21, gm_n85, gm_n56, gm_n6038, gm_n269);
	nor (gm_n6040, gm_n6039, gm_n6037, gm_n6035);
	or (gm_n6041, gm_n461, in_13, in_9, gm_n502, gm_n866);
	nor (gm_n6042, gm_n313, in_21, gm_n55, gm_n6041, gm_n374);
	nand (gm_n6043, in_13, gm_n62, gm_n94, gm_n576, gm_n123);
	nor (gm_n6044, gm_n441, in_21, in_17, gm_n6043, gm_n375);
	nand (gm_n6045, gm_n110, in_13, in_9, gm_n341, gm_n123);
	nor (gm_n6046, gm_n105, gm_n72, in_17, gm_n6045, gm_n441);
	nor (gm_n6047, gm_n6046, gm_n6044, gm_n6042);
	nand (gm_n6048, gm_n6034, gm_n5836, gm_n5834, gm_n6047, gm_n6040);
	and (gm_n6049, gm_n90, in_10, gm_n62, gm_n825, gm_n1158);
	nand (gm_n6050, gm_n166, gm_n86, gm_n119, gm_n6049);
	nor (gm_n6051, gm_n461, gm_n76, in_9, gm_n1132, gm_n463);
	nand (gm_n6052, gm_n206, in_21, in_17, gm_n6051, gm_n405);
	nor (gm_n6053, gm_n431, in_13, gm_n62, gm_n743, gm_n596);
	nand (gm_n6054, gm_n104, in_21, in_17, gm_n6053, gm_n327);
	nand (gm_n6055, gm_n6054, gm_n6052, gm_n6050);
	nor (gm_n6056, gm_n431, gm_n76, gm_n62, gm_n1583, gm_n344);
	nand (gm_n6057, gm_n255, gm_n72, gm_n55, gm_n6056, gm_n373);
	nand (gm_n6058, gm_n199, gm_n131, gm_n119, gm_n4512, gm_n545);
	nand (gm_n6059, gm_n311, gm_n72, in_17, gm_n5703, gm_n595);
	nand (gm_n6060, gm_n6059, gm_n6058, gm_n6057);
	nor (gm_n6061, gm_n6048, gm_n5833, gm_n5831, gm_n6060, gm_n6055);
	nor (gm_n6062, gm_n121, in_21, in_17, gm_n839, gm_n620);
	or (gm_n6063, gm_n274, in_13, gm_n59, gm_n355);
	nor (gm_n6064, gm_n184, in_21, gm_n55, gm_n6063, gm_n620);
	or (gm_n6065, gm_n393, gm_n263, gm_n60, gm_n4917, gm_n643);
	nor (gm_n6066, in_21, gm_n85, in_19, gm_n6065);
	nor (gm_n6067, gm_n6066, gm_n6064, gm_n6062);
	nand (gm_n6068, gm_n392, gm_n79, in_15, gm_n998, gm_n281);
	nor (gm_n6069, gm_n72, in_20, in_19, gm_n6068);
	or (gm_n6070, gm_n605, gm_n147, in_14, gm_n842);
	nor (gm_n6071, gm_n1989, gm_n211, in_18, gm_n6070);
	or (gm_n6072, gm_n430, in_13, gm_n62, gm_n345, gm_n431);
	nor (gm_n6073, gm_n184, in_21, in_17, gm_n6072, gm_n479);
	nor (gm_n6074, gm_n6073, gm_n6071, gm_n6069);
	nand (gm_n6075, gm_n6061, gm_n5830, gm_n5828, gm_n6074, gm_n6067);
	nor (gm_n6076, gm_n90, in_10, gm_n62, gm_n3099, gm_n467);
	nand (gm_n6077, gm_n245, gm_n243, gm_n119, gm_n6076);
	nor (gm_n6078, gm_n293, gm_n274, gm_n60, gm_n2060, gm_n760);
	nand (gm_n6079, gm_n72, in_20, in_19, gm_n6078);
	or (gm_n6080, gm_n103, in_21, gm_n55, gm_n1540, gm_n105);
	nand (gm_n6081, gm_n6080, gm_n6079, gm_n6077);
	nor (gm_n6082, gm_n430, in_13, in_9, gm_n481, gm_n431);
	nand (gm_n6083, gm_n255, in_21, gm_n55, gm_n6082, gm_n327);
	nor (gm_n6084, gm_n461, gm_n76, in_9, gm_n743, gm_n430);
	nand (gm_n6085, gm_n311, gm_n72, in_17, gm_n6084, gm_n405);
	nor (gm_n6086, gm_n227, in_16, gm_n59, gm_n4967, gm_n263);
	nand (gm_n6087, gm_n138, in_21, in_20, gm_n6086);
	nand (gm_n6088, gm_n6087, gm_n6085, gm_n6083);
	nor (gm_n6089, gm_n6075, gm_n5826, gm_n5824, gm_n6088, gm_n6081);
	nand (gm_n6090, gm_n314, in_13, in_9, gm_n341, gm_n316);
	nor (gm_n6091, gm_n441, in_21, gm_n55, gm_n6090, gm_n313);
	or (gm_n6092, gm_n114, gm_n73, gm_n59, gm_n1519, gm_n213);
	nor (gm_n6093, gm_n219, in_21, in_20, gm_n6092);
	or (gm_n6094, gm_n90, gm_n78, gm_n62, gm_n3006, gm_n807);
	nor (gm_n6095, gm_n437, gm_n130, in_18, gm_n6094);
	nor (gm_n6096, gm_n6095, gm_n6093, gm_n6091);
	nand (gm_n6097, gm_n61, in_16, in_12, gm_n3454, gm_n79);
	nor (gm_n6098, gm_n219, in_21, in_20, gm_n6097);
	nand (gm_n6099, gm_n123, gm_n76, in_9, gm_n186, gm_n126);
	nor (gm_n6100, gm_n312, gm_n72, in_17, gm_n6099, gm_n375);
	nand (gm_n6101, gm_n110, in_13, in_9, gm_n579, gm_n186);
	nor (gm_n6102, gm_n620, in_21, in_17, gm_n6101, gm_n375);
	nor (gm_n6103, gm_n6102, gm_n6100, gm_n6098);
	nand (gm_n6104, gm_n6089, gm_n5822, gm_n5820, gm_n6103, gm_n6096);
	nor (gm_n6105, gm_n406, in_13, in_9, gm_n502, gm_n345);
	nand (gm_n6106, gm_n102, gm_n72, gm_n55, gm_n6105, gm_n339);
	nor (gm_n6107, gm_n461, in_13, gm_n62, gm_n597, gm_n443);
	nand (gm_n6108, gm_n254, in_21, in_17, gm_n6107, gm_n339);
	nor (gm_n6109, gm_n609, in_13, gm_n62, gm_n481, gm_n406);
	nand (gm_n6110, gm_n339, in_21, gm_n55, gm_n6109, gm_n373);
	nand (gm_n6111, gm_n6110, gm_n6108, gm_n6106);
	nor (gm_n6112, gm_n263, gm_n159, in_15, gm_n1519, gm_n447);
	nand (gm_n6113, gm_n72, gm_n85, in_19, gm_n6112);
	nand (gm_n6114, gm_n102, gm_n72, in_17, gm_n3341, gm_n339);
	nor (gm_n6115, gm_n461, in_13, gm_n62, gm_n730, gm_n256);
	nand (gm_n6116, gm_n102, in_21, gm_n55, gm_n6115);
	nand (gm_n6117, gm_n6116, gm_n6114, gm_n6113);
	nor (gm_n6118, gm_n6104, gm_n5818, gm_n5816, gm_n6117, gm_n6111);
	nand (gm_n6119, gm_n306, gm_n64, gm_n60, gm_n869, gm_n486);
	nor (gm_n6120, gm_n72, gm_n85, gm_n56, gm_n6119);
	nand (gm_n6121, gm_n192, in_15, in_11, gm_n3625, gm_n448);
	nor (gm_n6122, in_21, in_20, gm_n56, gm_n6121);
	nand (gm_n6123, gm_n532, in_14, in_10, gm_n829, gm_n335);
	nor (gm_n6124, gm_n244, gm_n212, gm_n119, gm_n6123);
	nor (gm_n6125, gm_n6124, gm_n6122, gm_n6120);
	and (gm_n6126, gm_n254, in_21, in_17, gm_n1497, gm_n1076);
	or (gm_n6127, gm_n290, gm_n155, in_15, gm_n2589, gm_n293);
	nor (gm_n6128, in_21, gm_n85, in_19, gm_n6127);
	nor (gm_n6129, gm_n841, gm_n87, in_18, gm_n3645);
	nor (gm_n6130, gm_n6129, gm_n6128, gm_n6126);
	nand (gm_n6131, gm_n6118, gm_n5814, gm_n5812, gm_n6130, gm_n6125);
	nor (gm_n6132, gm_n609, in_10, in_9, gm_n503, gm_n807);
	nand (gm_n6133, gm_n199, gm_n119, in_14, gm_n6132, gm_n323);
	nor (gm_n6134, gm_n147, gm_n95, in_10, gm_n389);
	nand (gm_n6135, gm_n254, gm_n72, in_17, gm_n6134, gm_n1076);
	nor (gm_n6136, gm_n248, in_14, gm_n78, gm_n438, gm_n369);
	nand (gm_n6137, gm_n323, gm_n129, gm_n119, gm_n6136);
	nand (gm_n6138, gm_n6137, gm_n6135, gm_n6133);
	nor (gm_n6139, gm_n514, in_13, in_9, gm_n463, gm_n796);
	nand (gm_n6140, gm_n254, in_21, in_17, gm_n6139, gm_n405);
	nor (gm_n6141, gm_n257, in_13, in_9, gm_n705, gm_n662);
	nand (gm_n6142, gm_n206, in_21, gm_n55, gm_n6141);
	nor (gm_n6143, gm_n193, gm_n60, gm_n63, gm_n770, gm_n271);
	nand (gm_n6144, gm_n72, gm_n85, in_19, gm_n6143, gm_n75);
	nand (gm_n6145, gm_n6144, gm_n6142, gm_n6140);
	nor (out_17, gm_n6138, gm_n6131, gm_n5811, gm_n6145);
	or (gm_n6147, gm_n92, in_14, gm_n78, gm_n589, gm_n148);
	nor (gm_n6148, gm_n531, gm_n89, gm_n119, gm_n6147);
	nor (gm_n6149, gm_n358, in_13, in_9, gm_n1583, gm_n344);
	nand (gm_n6150, gm_n102, in_21, in_17, gm_n6149, gm_n595);
	or (gm_n6151, gm_n406, gm_n76, in_9, gm_n462, gm_n344);
	nor (gm_n6152, gm_n441, in_21, gm_n55, gm_n6151, gm_n313);
	nand (gm_n6153, gm_n90, gm_n78, gm_n62, gm_n3587, gm_n600);
	nor (gm_n6154, gm_n244, gm_n167, gm_n119, gm_n6153);
	and (gm_n6155, gm_n713, gm_n90, in_10, gm_n722, gm_n490);
	nand (gm_n6156, gm_n131, gm_n129, in_18, gm_n6155);
	nor (gm_n6157, gm_n514, gm_n76, gm_n62, gm_n988, gm_n344);
	nand (gm_n6158, gm_n102, gm_n72, in_17, gm_n6157, gm_n1076);
	nand (gm_n6159, gm_n486, gm_n154, gm_n60, gm_n1531, gm_n869);
	nor (gm_n6160, gm_n72, gm_n85, gm_n56, gm_n6159);
	nand (gm_n6161, gm_n264, in_16, in_12, gm_n3886, gm_n949);
	nor (gm_n6162, gm_n139, gm_n72, in_20, gm_n6161);
	nand (gm_n6163, gm_n174, in_21, gm_n55, gm_n4530, gm_n523);
	nor (gm_n6164, gm_n359, gm_n76, in_9, gm_n443, gm_n480);
	nand (gm_n6165, gm_n174, gm_n72, in_17, gm_n6164, gm_n595);
	nand (gm_n6166, in_14, gm_n78, gm_n62, gm_n1198, gm_n624);
	nor (gm_n6167, gm_n437, gm_n244, in_18, gm_n6166);
	or (gm_n6168, gm_n155, in_16, in_12, gm_n1176, gm_n276);
	nor (gm_n6169, gm_n139, gm_n72, in_20, gm_n6168);
	nor (gm_n6170, gm_n95, gm_n90, gm_n78, gm_n149, gm_n133);
	nand (gm_n6171, gm_n243, gm_n131, gm_n119, gm_n6170);
	nand (gm_n6172, gm_n104, gm_n72, gm_n55, gm_n5716, gm_n254);
	or (gm_n6173, gm_n818, gm_n76, gm_n62, gm_n431, gm_n667);
	nor (gm_n6174, gm_n441, gm_n72, gm_n55, gm_n6173, gm_n328);
	or (gm_n6175, gm_n227, gm_n73, gm_n59, gm_n1223, gm_n297);
	nor (gm_n6176, gm_n219, in_21, in_20, gm_n6175);
	and (gm_n6177, gm_n90, gm_n78, gm_n62, gm_n1401, gm_n600);
	nand (gm_n6178, gm_n806, gm_n86, gm_n119, gm_n6177);
	nor (gm_n6179, gm_n114, gm_n73, in_12, gm_n1884, gm_n158);
	nand (gm_n6180, gm_n57, in_21, in_20, gm_n6179);
	nand (gm_n6181, gm_n405, in_13, in_9, gm_n615, gm_n314);
	nor (gm_n6182, gm_n103, in_21, gm_n55, gm_n6181);
	nand (gm_n6183, gm_n448, in_19, in_15, gm_n1068, gm_n545);
	nor (gm_n6184, gm_n6183, gm_n72, in_20);
	nor (gm_n6185, gm_n152, in_16, gm_n59, gm_n1689, gm_n155);
	nand (gm_n6186, gm_n179, in_21, gm_n85, gm_n6185);
	nor (gm_n6187, gm_n159, gm_n297, in_15, gm_n855, gm_n485);
	nand (gm_n6188, gm_n72, gm_n85, in_19, gm_n6187);
	or (gm_n6189, gm_n213, in_16, gm_n59, gm_n632, gm_n319);
	nor (gm_n6190, gm_n496, gm_n72, gm_n85, gm_n6189);
	or (gm_n6191, in_14, gm_n78, in_9, gm_n808, gm_n362);
	nor (gm_n6192, gm_n212, gm_n87, in_18, gm_n6191);
	nor (gm_n6193, gm_n572, gm_n67, gm_n90, gm_n2017, gm_n467);
	nand (gm_n6194, gm_n200, gm_n164, in_18, gm_n6193);
	nand (gm_n6195, gm_n125, gm_n76, in_9, gm_n402, gm_n316);
	or (gm_n6196, gm_n479, in_21, in_17, gm_n6195, gm_n662);
	or (gm_n6197, gm_n90, gm_n78, gm_n62, gm_n2198, gm_n807);
	nor (gm_n6198, gm_n1989, gm_n244, in_18, gm_n6197);
	or (gm_n6199, gm_n158, in_16, in_12, gm_n2589, gm_n319);
	nor (gm_n6200, gm_n219, in_21, gm_n85, gm_n6199);
	nor (gm_n6201, gm_n115, in_16, in_12, gm_n1542, gm_n319);
	nand (gm_n6202, gm_n138, gm_n72, gm_n85, gm_n6201);
	nor (gm_n6203, gm_n269, gm_n274, gm_n60, gm_n520, gm_n643);
	nand (gm_n6204, gm_n72, in_20, gm_n56, gm_n6203);
	nand (gm_n6205, gm_n281, gm_n233, gm_n60, gm_n2172, gm_n869);
	nor (gm_n6206, in_21, in_20, gm_n56, gm_n6205);
	nand (gm_n6207, gm_n187, gm_n76, gm_n62, gm_n1049, gm_n314);
	nor (gm_n6208, gm_n103, in_21, in_17, gm_n6207, gm_n184);
	nor (gm_n6209, gm_n114, gm_n73, gm_n59, gm_n2333, gm_n274);
	nand (gm_n6210, gm_n113, gm_n72, gm_n85, gm_n6209);
	nor (gm_n6211, gm_n190, in_16, gm_n59, gm_n2956, gm_n227);
	nand (gm_n6212, gm_n138, in_21, gm_n85, gm_n6211);
	nand (gm_n6213, in_13, gm_n59, gm_n63, gm_n601, gm_n1144);
	nor (gm_n6214, gm_n620, gm_n72, gm_n55, gm_n6213, gm_n662);
	or (gm_n6215, gm_n92, gm_n90, in_10, gm_n491, gm_n389);
	nor (gm_n6216, gm_n531, gm_n167, gm_n119, gm_n6215);
	nor (gm_n6217, gm_n220, gm_n73, gm_n59, gm_n4935, gm_n263);
	nand (gm_n6218, gm_n296, in_21, gm_n85, gm_n6217);
	or (gm_n6219, gm_n95, in_11, in_10, gm_n775);
	nor (gm_n6220, gm_n191, in_19, in_15, gm_n6219, gm_n193);
	nand (gm_n6221, gm_n6220, in_21, gm_n85);
	nor (gm_n6222, gm_n818, in_13, gm_n62, gm_n463, gm_n406);
	nand (gm_n6223, gm_n254, in_21, gm_n55, gm_n6222, gm_n255);
	nand (gm_n6224, gm_n179, in_21, in_20, gm_n2108);
	nor (gm_n6225, gm_n114, gm_n73, gm_n59, gm_n1284, gm_n213);
	nand (gm_n6226, gm_n179, gm_n72, in_20, gm_n6225);
	nand (gm_n6227, gm_n6223, gm_n6221, gm_n6218, gm_n6226, gm_n6224);
	nor (gm_n6228, gm_n90, gm_n78, in_9, gm_n1176, gm_n207);
	nand (gm_n6229, gm_n199, gm_n131, gm_n119, gm_n6228);
	nor (gm_n6230, gm_n263, in_16, in_12, gm_n2589, gm_n354);
	nand (gm_n6231, gm_n383, gm_n72, gm_n85, gm_n6230);
	nor (gm_n6232, gm_n263, gm_n73, gm_n59, gm_n1859, gm_n385);
	nand (gm_n6233, gm_n113, in_21, gm_n85, gm_n6232);
	nand (gm_n6234, gm_n6233, gm_n6231, gm_n6229);
	nor (gm_n6235, gm_n274, in_16, gm_n59, gm_n887, gm_n276);
	nand (gm_n6236, gm_n296, in_21, gm_n85, gm_n6235);
	nor (gm_n6237, gm_n393, gm_n213, gm_n60, gm_n1332, gm_n633);
	nand (gm_n6238, gm_n72, in_20, in_19, gm_n6237);
	nor (gm_n6239, gm_n114, gm_n73, gm_n59, gm_n705, gm_n213);
	nand (gm_n6240, gm_n495, in_21, gm_n85, gm_n6239);
	nand (gm_n6241, gm_n6240, gm_n6238, gm_n6236);
	nor (gm_n6242, gm_n6227, gm_n6216, gm_n6214, gm_n6241, gm_n6234);
	nand (gm_n6243, gm_n224, gm_n64, gm_n60, gm_n394, gm_n422);
	nor (gm_n6244, in_21, in_20, in_19, gm_n6243);
	or (gm_n6245, gm_n274, gm_n193, gm_n60, gm_n1173, gm_n393);
	nor (gm_n6246, gm_n72, in_20, gm_n56, gm_n6245);
	nand (gm_n6247, gm_n600, in_14, gm_n78, gm_n793, gm_n335);
	nor (gm_n6248, gm_n165, gm_n89, in_18, gm_n6247);
	nor (gm_n6249, gm_n6248, gm_n6246, gm_n6244);
	nand (gm_n6250, gm_n339, in_13, in_9, gm_n884, gm_n788);
	nor (gm_n6251, gm_n103, gm_n72, in_17, gm_n6250);
	nor (gm_n6252, gm_n217, gm_n211, gm_n119, gm_n246);
	nand (gm_n6253, gm_n64, gm_n73, gm_n59, gm_n2573, gm_n77);
	nor (gm_n6254, gm_n139, gm_n72, gm_n85, gm_n6253);
	nor (gm_n6255, gm_n6254, gm_n6252, gm_n6251);
	nand (gm_n6256, gm_n6242, gm_n6212, gm_n6210, gm_n6255, gm_n6249);
	and (gm_n6257, gm_n90, gm_n76, gm_n59, gm_n1947, gm_n222);
	nand (gm_n6258, gm_n348, gm_n131, in_18, gm_n6257);
	nor (gm_n6259, gm_n263, in_16, in_12, gm_n4967, gm_n276);
	nand (gm_n6260, gm_n57, in_21, gm_n85, gm_n6259);
	nand (gm_n6261, gm_n436, gm_n86, in_18, gm_n3046);
	nand (gm_n6262, gm_n6261, gm_n6260, gm_n6258);
	nor (gm_n6263, gm_n90, gm_n78, gm_n62, gm_n135, gm_n92);
	nand (gm_n6264, gm_n367, gm_n131, gm_n119, gm_n6263);
	nor (gm_n6265, gm_n297, in_16, gm_n59, gm_n474, gm_n354);
	nand (gm_n6266, gm_n138, in_21, in_20, gm_n6265);
	and (gm_n6267, gm_n90, gm_n78, in_9, gm_n1841, gm_n532);
	nand (gm_n6268, gm_n323, gm_n164, gm_n119, gm_n6267);
	nand (gm_n6269, gm_n6268, gm_n6266, gm_n6264);
	nor (gm_n6270, gm_n6256, gm_n6208, gm_n6206, gm_n6269, gm_n6262);
	or (gm_n6271, gm_n207, in_14, in_10, gm_n376, gm_n370);
	nor (gm_n6272, gm_n212, gm_n211, in_18, gm_n6271);
	nand (gm_n6273, gm_n76, gm_n62, gm_n94, gm_n576, gm_n314);
	nor (gm_n6274, gm_n312, gm_n72, gm_n55, gm_n6273, gm_n662);
	or (gm_n6275, gm_n158, in_16, gm_n59, gm_n3382, gm_n276);
	nor (gm_n6276, gm_n912, in_21, gm_n85, gm_n6275);
	nor (gm_n6277, gm_n6276, gm_n6274, gm_n6272);
	nand (gm_n6278, gm_n64, in_16, gm_n59, gm_n535, gm_n221);
	nor (gm_n6279, gm_n496, in_21, gm_n85, gm_n6278);
	nand (gm_n6280, gm_n78, gm_n62, in_8, gm_n2074, gm_n532);
	nor (gm_n6281, gm_n132, in_18, in_14, gm_n6280, gm_n824);
	nand (gm_n6282, gm_n64, in_16, in_12, gm_n2065, gm_n571);
	nor (gm_n6283, gm_n496, in_21, gm_n85, gm_n6282);
	nor (gm_n6284, gm_n6283, gm_n6281, gm_n6279);
	nand (gm_n6285, gm_n6270, gm_n6204, gm_n6202, gm_n6284, gm_n6277);
	nor (gm_n6286, gm_n263, gm_n73, in_12, gm_n2956, gm_n319);
	nand (gm_n6287, gm_n383, gm_n72, gm_n85, gm_n6286);
	nor (gm_n6288, gm_n115, in_12, gm_n94, gm_n939, gm_n152);
	nand (gm_n6289, in_21, gm_n85, in_16, gm_n6288, gm_n113);
	nor (gm_n6290, gm_n208, gm_n358, in_13, gm_n287, gm_n256);
	nand (gm_n6291, gm_n206, gm_n72, gm_n55, gm_n6290);
	nand (gm_n6292, gm_n6291, gm_n6289, gm_n6287);
	and (gm_n6293, gm_n126, in_13, in_9, gm_n341, gm_n579);
	nand (gm_n6294, gm_n104, gm_n72, gm_n55, gm_n6293, gm_n327);
	nor (gm_n6295, gm_n158, gm_n59, in_8, gm_n161, gm_n152);
	nand (gm_n6296, gm_n72, in_20, in_16, gm_n6295, gm_n495);
	nor (gm_n6297, gm_n90, in_10, gm_n62, gm_n520, gm_n362);
	nand (gm_n6298, gm_n146, gm_n131, in_18, gm_n6297);
	nand (gm_n6299, gm_n6298, gm_n6296, gm_n6294);
	nor (gm_n6300, gm_n6285, gm_n6200, gm_n6198, gm_n6299, gm_n6292);
	or (gm_n6301, gm_n274, gm_n74, gm_n60, gm_n1052, gm_n760);
	nor (gm_n6302, in_21, gm_n85, gm_n56, gm_n6301);
	nand (gm_n6303, gm_n77, in_16, in_12, gm_n950, gm_n222);
	nor (gm_n6304, gm_n384, in_21, gm_n85, gm_n6303);
	nand (gm_n6305, gm_n281, gm_n214, gm_n60, gm_n1569, gm_n422);
	nor (gm_n6306, gm_n72, gm_n85, in_19, gm_n6305);
	nor (gm_n6307, gm_n6306, gm_n6304, gm_n6302);
	or (gm_n6308, gm_n207, gm_n90, in_10, gm_n389, gm_n287);
	nor (gm_n6309, gm_n211, gm_n132, gm_n119, gm_n6308);
	nand (gm_n6310, in_14, in_10, in_9, gm_n1605, gm_n624);
	nor (gm_n6311, gm_n368, gm_n246, gm_n119, gm_n6310);
	and (gm_n6312, gm_n129, gm_n88, in_18, gm_n2799);
	nor (gm_n6313, gm_n6312, gm_n6311, gm_n6309);
	nand (gm_n6314, gm_n6300, gm_n6196, gm_n6194, gm_n6313, gm_n6307);
	nor (gm_n6315, gm_n461, in_13, gm_n62, gm_n988, gm_n463);
	nand (gm_n6316, gm_n523, gm_n72, gm_n55, gm_n6315, gm_n373);
	nor (gm_n6317, gm_n297, in_16, in_12, gm_n298, gm_n276);
	nand (gm_n6318, gm_n697, gm_n72, gm_n85, gm_n6317);
	nor (gm_n6319, gm_n358, gm_n76, gm_n62, gm_n621, gm_n344);
	nand (gm_n6320, gm_n120, in_21, in_17, gm_n6319, gm_n339);
	nand (gm_n6321, gm_n6320, gm_n6318, gm_n6316);
	nor (gm_n6322, gm_n247, in_14, gm_n78, gm_n467, gm_n350);
	nand (gm_n6323, gm_n323, gm_n86, in_18, gm_n6322);
	nor (gm_n6324, gm_n263, gm_n74, in_15, gm_n799, gm_n633);
	nand (gm_n6325, in_21, gm_n85, gm_n56, gm_n6324);
	nor (gm_n6326, gm_n406, in_13, gm_n62, gm_n1583, gm_n596);
	nand (gm_n6327, gm_n104, gm_n72, gm_n55, gm_n6326, gm_n206);
	nand (gm_n6328, gm_n6327, gm_n6325, gm_n6323);
	nor (gm_n6329, gm_n6314, gm_n6192, gm_n6190, gm_n6328, gm_n6321);
	nand (gm_n6330, gm_n214, gm_n73, in_12, gm_n3679, gm_n571);
	nor (gm_n6331, gm_n139, gm_n72, gm_n85, gm_n6330);
	nand (gm_n6332, gm_n334, in_14, gm_n78, gm_n722, gm_n1345);
	nor (gm_n6333, gm_n167, gm_n211, in_18, gm_n6332);
	or (gm_n6334, gm_n74, in_19, in_15, gm_n6219, gm_n643);
	nor (gm_n6335, gm_n6334, gm_n72, in_20);
	nor (gm_n6336, gm_n6335, gm_n6333, gm_n6331);
	or (gm_n6337, gm_n207, gm_n977, gm_n90, gm_n761);
	nor (gm_n6338, gm_n246, gm_n244, gm_n119, gm_n6337);
	or (gm_n6339, gm_n430, in_13, in_9, gm_n597, gm_n406);
	nor (gm_n6340, gm_n388, in_21, in_17, gm_n6339, gm_n256);
	nand (gm_n6341, gm_n142, in_16, gm_n59, gm_n571, gm_n214);
	nor (gm_n6342, gm_n58, gm_n72, gm_n85, gm_n6341);
	nor (gm_n6343, gm_n6342, gm_n6340, gm_n6338);
	nand (gm_n6344, gm_n6329, gm_n6188, gm_n6186, gm_n6343, gm_n6336);
	nor (gm_n6345, gm_n257, gm_n76, in_9, gm_n743, gm_n502);
	nand (gm_n6346, gm_n120, gm_n72, gm_n55, gm_n6345, gm_n1076);
	nor (gm_n6347, gm_n256, gm_n461, in_13, gm_n775, gm_n370);
	nand (gm_n6348, gm_n327, gm_n72, in_17, gm_n6347);
	nor (gm_n6349, gm_n196, gm_n158, gm_n60, gm_n633, gm_n485);
	nand (gm_n6350, in_21, gm_n85, gm_n56, gm_n6349);
	nand (gm_n6351, gm_n6350, gm_n6348, gm_n6346);
	nor (gm_n6352, gm_n133, in_14, gm_n78, gm_n438, gm_n376);
	nand (gm_n6353, gm_n367, gm_n245, gm_n119, gm_n6352);
	and (gm_n6354, gm_n532, in_14, gm_n78, gm_n793, gm_n1157);
	nand (gm_n6355, gm_n348, gm_n166, gm_n119, gm_n6354);
	nor (gm_n6356, gm_n95, in_14, in_10, gm_n369, gm_n286);
	nand (gm_n6357, gm_n436, gm_n367, in_18, gm_n6356);
	nand (gm_n6358, gm_n6357, gm_n6355, gm_n6353);
	nor (gm_n6359, gm_n6344, gm_n6184, gm_n6182, gm_n6358, gm_n6351);
	or (gm_n6360, in_14, gm_n78, in_9, gm_n2077, gm_n807);
	nor (gm_n6361, gm_n1989, gm_n824, in_18, gm_n6360);
	or (gm_n6362, gm_n514, in_13, gm_n62, gm_n1132, gm_n430);
	nor (gm_n6363, gm_n388, gm_n72, gm_n55, gm_n6362, gm_n328);
	or (gm_n6364, gm_n155, in_16, in_12, gm_n2357, gm_n319);
	nor (gm_n6365, gm_n912, gm_n72, gm_n85, gm_n6364);
	nor (gm_n6366, gm_n6365, gm_n6363, gm_n6361);
	and (gm_n6367, gm_n254, gm_n72, gm_n55, gm_n6082, gm_n339);
	or (gm_n6368, gm_n240, gm_n133, in_14, gm_n842);
	nor (gm_n6369, gm_n211, gm_n89, in_18, gm_n6368);
	nor (gm_n6370, gm_n184, gm_n72, in_17, gm_n5861, gm_n312);
	nor (gm_n6371, gm_n6370, gm_n6369, gm_n6367);
	nand (gm_n6372, gm_n6359, gm_n6180, gm_n6178, gm_n6371, gm_n6366);
	and (gm_n6373, gm_n64, in_16, in_12, gm_n2443, gm_n303);
	nand (gm_n6374, gm_n296, gm_n72, in_20, gm_n6373);
	and (gm_n6375, gm_n126, in_13, gm_n62, gm_n1049, gm_n185);
	nand (gm_n6376, gm_n102, gm_n72, in_17, gm_n6375, gm_n104);
	nor (gm_n6377, gm_n269, gm_n263, gm_n60, gm_n633, gm_n278);
	nand (gm_n6378, in_21, gm_n85, gm_n56, gm_n6377);
	nand (gm_n6379, gm_n6378, gm_n6376, gm_n6374);
	nor (gm_n6380, gm_n609, in_13, in_9, gm_n481, gm_n257);
	nand (gm_n6381, gm_n122, in_21, gm_n55, gm_n6380, gm_n327);
	nor (gm_n6382, gm_n430, in_13, in_9, gm_n462, gm_n442);
	nand (gm_n6383, gm_n104, gm_n72, in_17, gm_n6382, gm_n254);
	and (gm_n6384, gm_n187, in_13, in_9, gm_n402, gm_n341);
	nand (gm_n6385, gm_n122, in_21, in_17, gm_n6384, gm_n373);
	nand (gm_n6386, gm_n6385, gm_n6383, gm_n6381);
	nor (gm_n6387, gm_n6372, gm_n6176, gm_n6174, gm_n6386, gm_n6379);
	nand (gm_n6388, gm_n1076, gm_n76, gm_n62, gm_n2230, gm_n788);
	nor (gm_n6389, gm_n103, gm_n72, gm_n55, gm_n6388);
	or (gm_n6390, gm_n121, gm_n99, gm_n76, gm_n431, gm_n247);
	nor (gm_n6391, gm_n312, gm_n72, gm_n55, gm_n6390);
	or (gm_n6392, gm_n514, gm_n95, gm_n76, gm_n328, gm_n149);
	nor (gm_n6393, gm_n103, gm_n72, in_17, gm_n6392);
	nor (gm_n6394, gm_n6393, gm_n6391, gm_n6389);
	or (gm_n6395, gm_n213, gm_n168, gm_n60, gm_n2589, gm_n269);
	nor (gm_n6396, in_21, in_20, gm_n56, gm_n6395);
	nand (gm_n6397, gm_n90, in_10, in_9, gm_n1713, gm_n624);
	nor (gm_n6398, gm_n244, gm_n212, in_18, gm_n6397);
	or (gm_n6399, gm_n369, in_14, in_10, gm_n526, gm_n438);
	nor (gm_n6400, gm_n246, gm_n130, in_18, gm_n6399);
	nor (gm_n6401, gm_n6400, gm_n6398, gm_n6396);
	nand (gm_n6402, gm_n6387, gm_n6172, gm_n6171, gm_n6401, gm_n6394);
	nor (gm_n6403, gm_n461, gm_n76, in_9, gm_n359, gm_n430);
	nand (gm_n6404, gm_n122, gm_n72, in_17, gm_n6403, gm_n206);
	nor (gm_n6405, gm_n807, in_14, in_10, gm_n491, gm_n350);
	nand (gm_n6406, gm_n348, gm_n806, in_18, gm_n6405);
	nor (gm_n6407, gm_n406, in_13, in_9, gm_n1132, gm_n463);
	nand (gm_n6408, gm_n255, in_21, in_17, gm_n6407, gm_n373);
	nand (gm_n6409, gm_n6408, gm_n6406, gm_n6404);
	nor (gm_n6410, gm_n155, in_16, in_12, gm_n2029, gm_n354);
	nand (gm_n6411, gm_n495, in_21, in_20, gm_n6410);
	nor (gm_n6412, gm_n257, gm_n76, gm_n62, gm_n432, gm_n344);
	nand (gm_n6413, gm_n254, gm_n72, gm_n55, gm_n6412, gm_n339);
	nor (gm_n6414, gm_n430, gm_n76, gm_n62, gm_n1583, gm_n480);
	nand (gm_n6415, gm_n174, in_21, gm_n55, gm_n6414, gm_n1076);
	nand (gm_n6416, gm_n6415, gm_n6413, gm_n6411);
	nor (gm_n6417, gm_n6402, gm_n6169, gm_n6167, gm_n6416, gm_n6409);
	or (gm_n6418, gm_n514, in_13, in_9, gm_n743, gm_n463);
	nor (gm_n6419, gm_n313, in_21, gm_n55, gm_n6418, gm_n374);
	and (gm_n6420, gm_n102, gm_n72, gm_n55, gm_n6082, gm_n122);
	or (gm_n6421, gm_n358, gm_n76, gm_n62, gm_n1583, gm_n463);
	nor (gm_n6422, gm_n103, gm_n72, in_17, gm_n6421, gm_n328);
	nor (gm_n6423, gm_n6422, gm_n6420, gm_n6419);
	or (gm_n6424, gm_n807, in_14, gm_n78, gm_n526, gm_n370);
	nor (gm_n6425, gm_n246, gm_n824, in_18, gm_n6424);
	nand (gm_n6426, gm_n61, in_16, in_12, gm_n936, gm_n154);
	nor (gm_n6427, gm_n262, gm_n72, in_20, gm_n6426);
	nand (gm_n6428, gm_n110, in_13, in_9, gm_n402, gm_n341);
	nor (gm_n6429, gm_n121, gm_n72, gm_n55, gm_n6428, gm_n388);
	nor (gm_n6430, gm_n6429, gm_n6427, gm_n6425);
	nand (gm_n6431, gm_n6417, gm_n6165, gm_n6163, gm_n6430, gm_n6423);
	nand (gm_n6432, in_21, gm_n85, in_19, gm_n5472, gm_n379);
	nor (gm_n6433, in_14, in_10, in_9, gm_n2421, gm_n369);
	nand (gm_n6434, gm_n348, gm_n323, gm_n119, gm_n6433);
	nor (gm_n6435, gm_n228, gm_n977, in_14, gm_n362, gm_n238);
	nand (gm_n6436, gm_n243, gm_n166, gm_n119, gm_n6435);
	nand (gm_n6437, gm_n6436, gm_n6434, gm_n6432);
	nor (gm_n6438, gm_n259, gm_n90, in_10, gm_n491, gm_n362);
	nand (gm_n6439, gm_n166, gm_n146, in_18, gm_n6438);
	nor (gm_n6440, gm_n114, gm_n73, gm_n59, gm_n4967, gm_n263);
	nand (gm_n6441, gm_n113, gm_n72, gm_n85, gm_n6440);
	and (gm_n6442, in_14, in_10, gm_n62, gm_n1392, gm_n600);
	nand (gm_n6443, gm_n243, gm_n200, gm_n119, gm_n6442);
	nand (gm_n6444, gm_n6443, gm_n6441, gm_n6439);
	nor (gm_n6445, gm_n6431, gm_n6162, gm_n6160, gm_n6444, gm_n6437);
	or (gm_n6446, gm_n155, in_16, gm_n59, gm_n1923, gm_n385);
	nor (gm_n6447, gm_n139, gm_n72, gm_n85, gm_n6446);
	or (gm_n6448, gm_n609, in_13, in_9, gm_n359, gm_n431);
	nor (gm_n6449, gm_n479, gm_n72, gm_n55, gm_n6448, gm_n662);
	or (gm_n6450, gm_n461, in_13, in_9, gm_n988, gm_n443);
	nor (gm_n6451, gm_n313, gm_n72, gm_n55, gm_n6450, gm_n374);
	nor (gm_n6452, gm_n6451, gm_n6449, gm_n6447);
	or (gm_n6453, gm_n461, gm_n76, in_9, gm_n345, gm_n430);
	nor (gm_n6454, gm_n183, gm_n72, in_17, gm_n6453, gm_n313);
	nand (gm_n6455, gm_n392, gm_n233, in_15, gm_n1758, gm_n1101);
	nor (gm_n6456, gm_n72, in_20, gm_n56, gm_n6455);
	nand (gm_n6457, gm_n233, in_16, in_12, gm_n1135, gm_n303);
	nor (gm_n6458, gm_n219, gm_n72, in_20, gm_n6457);
	nor (gm_n6459, gm_n6458, gm_n6456, gm_n6454);
	nand (gm_n6460, gm_n6445, gm_n6158, gm_n6156, gm_n6459, gm_n6452);
	nand (gm_n6461, gm_n206, gm_n72, gm_n55, gm_n4476, gm_n339);
	nand (gm_n6462, gm_n367, gm_n88, gm_n119, gm_n1714);
	and (gm_n6463, in_13, gm_n62, gm_n94, gm_n601, gm_n123);
	nand (gm_n6464, gm_n254, in_21, in_17, gm_n6463, gm_n255);
	nand (gm_n6465, gm_n6464, gm_n6462, gm_n6461);
	nor (gm_n6466, gm_n190, in_16, gm_n59, gm_n385, gm_n135);
	nand (gm_n6467, gm_n179, gm_n72, in_20, gm_n6466);
	nand (gm_n6468, gm_n174, gm_n72, gm_n55, gm_n2914, gm_n523);
	nor (gm_n6469, gm_n485, gm_n158, gm_n60, gm_n2826, gm_n764);
	nand (gm_n6470, in_21, in_20, in_19, gm_n6469);
	nand (gm_n6471, gm_n6470, gm_n6468, gm_n6467);
	nor (gm_n6472, gm_n6460, gm_n6154, gm_n6152, gm_n6471, gm_n6465);
	nor (gm_n6473, in_14, in_10, gm_n62, gm_n1837, gm_n133);
	nand (gm_n6474, gm_n436, gm_n86, gm_n119, gm_n6473);
	nor (gm_n6475, gm_n190, gm_n73, in_12, gm_n1170, gm_n385);
	nand (gm_n6476, gm_n113, in_21, in_20, gm_n6475);
	nor (gm_n6477, gm_n213, gm_n73, in_12, gm_n1824, gm_n319);
	nand (gm_n6478, gm_n179, gm_n72, in_20, gm_n6477);
	nand (gm_n6479, gm_n6474, gm_n6472, gm_n6150, gm_n6478, gm_n6476);
	and (gm_n6480, gm_n77, gm_n73, in_12, gm_n626, gm_n233);
	nand (gm_n6481, gm_n697, in_21, in_20, gm_n6480);
	nor (gm_n6482, gm_n207, gm_n841, in_14, gm_n1382, gm_n980);
	nand (gm_n6483, gm_n6482, gm_n86, in_18);
	nor (gm_n6484, gm_n147, in_14, gm_n78, gm_n3786, gm_n287);
	nand (gm_n6485, gm_n243, gm_n131, in_18, gm_n6484);
	nand (gm_n6486, gm_n6485, gm_n6483, gm_n6481);
	or (gm_n6487, gm_n447, gm_n190, gm_n60, gm_n1751, gm_n760);
	nor (gm_n6488, gm_n72, gm_n85, in_19, gm_n6487);
	nor (out_18, gm_n6486, gm_n6479, gm_n6148, gm_n6488);
	or (gm_n6490, gm_n78, in_9, gm_n94, gm_n467, gm_n417);
	nor (gm_n6491, gm_n244, in_18, gm_n90, gm_n6490, gm_n437);
	nor (gm_n6492, gm_n90, gm_n78, in_9, gm_n1837, gm_n92);
	nand (gm_n6493, gm_n436, gm_n129, gm_n119, gm_n6492);
	or (gm_n6494, gm_n274, gm_n196, gm_n60, gm_n633, gm_n393);
	nor (gm_n6495, in_21, in_20, gm_n56, gm_n6494);
	or (gm_n6496, gm_n207, in_14, in_10, gm_n370, gm_n208);
	nor (gm_n6497, gm_n824, gm_n132, gm_n119, gm_n6496);
	and (gm_n6498, gm_n268, gm_n143, gm_n60, gm_n1186, gm_n545);
	nand (gm_n6499, in_21, in_20, gm_n56, gm_n6498);
	nor (gm_n6500, gm_n274, gm_n193, gm_n60, gm_n1052, gm_n485);
	nand (gm_n6501, gm_n72, in_20, gm_n56, gm_n6500);
	or (gm_n6502, gm_n95, in_14, in_10, gm_n369, gm_n208);
	nor (gm_n6503, gm_n244, gm_n89, gm_n119, gm_n6502);
	and (gm_n6504, gm_n383, in_21, in_20, gm_n5821);
	nor (gm_n6505, gm_n662, gm_n76, gm_n62, gm_n3721, gm_n406);
	nand (gm_n6506, gm_n254, gm_n72, in_17, gm_n6505);
	nor (gm_n6507, gm_n293, gm_n263, in_15, gm_n633, gm_n632);
	nand (gm_n6508, in_21, gm_n85, in_19, gm_n6507);
	or (gm_n6509, gm_n431, gm_n313, gm_n76, gm_n589, gm_n370);
	nor (gm_n6510, gm_n620, gm_n72, gm_n55, gm_n6509);
	or (gm_n6511, gm_n147, gm_n90, gm_n78, gm_n438, gm_n376);
	nor (gm_n6512, gm_n244, gm_n167, gm_n119, gm_n6511);
	and (gm_n6513, gm_n264, gm_n73, gm_n59, gm_n778, gm_n275);
	nand (gm_n6514, gm_n57, gm_n72, gm_n85, gm_n6513);
	nor (gm_n6515, gm_n90, in_10, gm_n62, gm_n2474, gm_n369);
	nand (gm_n6516, gm_n348, gm_n200, in_18, gm_n6515);
	and (gm_n6517, gm_n93, in_6, in_5, gm_n426);
	nand (gm_n6518, gm_n76, gm_n62, in_8, gm_n6517, gm_n314);
	nor (gm_n6519, gm_n183, gm_n72, in_17, gm_n6518, gm_n375);
	or (gm_n6520, gm_n152, gm_n73, in_12, gm_n3099, gm_n213);
	nor (gm_n6521, gm_n219, gm_n72, in_20, gm_n6520);
	and (gm_n6522, gm_n76, gm_n62, in_8, gm_n6517, gm_n579);
	nand (gm_n6523, gm_n120, in_21, gm_n55, gm_n6522, gm_n255);
	nor (gm_n6524, gm_n158, gm_n73, in_12, gm_n3006, gm_n385);
	nand (gm_n6525, gm_n138, gm_n72, in_20, gm_n6524);
	nor (gm_n6526, gm_n479, in_21, gm_n55, gm_n1231, gm_n256);
	nand (gm_n6527, gm_n106, in_13, gm_n62, gm_n341, gm_n126);
	nor (gm_n6528, gm_n312, in_21, gm_n55, gm_n6527, gm_n328);
	nor (gm_n6529, gm_n796, in_13, in_9, gm_n463, gm_n442);
	nand (gm_n6530, gm_n206, gm_n72, gm_n55, gm_n6529, gm_n405);
	nor (gm_n6531, in_14, gm_n78, in_9, gm_n1006, gm_n369);
	nand (gm_n6532, gm_n166, gm_n86, in_18, gm_n6531);
	or (gm_n6533, gm_n514, in_13, in_9, gm_n621, gm_n596);
	nor (gm_n6534, gm_n184, gm_n72, gm_n55, gm_n6533, gm_n479);
	or (gm_n6535, gm_n818, gm_n76, gm_n62, gm_n442, gm_n430);
	nor (gm_n6536, gm_n441, gm_n72, gm_n55, gm_n6535, gm_n184);
	and (gm_n6537, gm_n233, gm_n73, in_12, gm_n2276, gm_n303);
	nand (gm_n6538, gm_n296, in_21, gm_n85, gm_n6537);
	nor (gm_n6539, gm_n406, gm_n76, gm_n62, gm_n743, gm_n596);
	nand (gm_n6540, gm_n104, in_21, gm_n55, gm_n6539, gm_n174);
	or (gm_n6541, gm_n609, gm_n76, gm_n62, gm_n621, gm_n480);
	nor (gm_n6542, gm_n313, gm_n72, gm_n55, gm_n6541, gm_n374);
	or (gm_n6543, gm_n298, gm_n76, gm_n62, gm_n406, gm_n662);
	nor (gm_n6544, gm_n374, in_21, gm_n55, gm_n6543);
	nor (gm_n6545, gm_n430, in_13, in_9, gm_n432, gm_n257);
	nand (gm_n6546, gm_n523, gm_n72, in_17, gm_n6545, gm_n311);
	and (gm_n6547, gm_n61, gm_n73, in_12, gm_n1947, gm_n143);
	nand (gm_n6548, gm_n179, in_21, in_20, gm_n6547);
	nand (gm_n6549, gm_n90, gm_n78, gm_n62, gm_n884, gm_n1158);
	nor (gm_n6550, gm_n1989, gm_n165, gm_n119, gm_n6549);
	nand (gm_n6551, gm_n78, in_9, in_8, gm_n1263, gm_n713);
	nor (gm_n6552, gm_n167, in_18, in_14, gm_n6551, gm_n531);
	nor (gm_n6553, gm_n480, in_13, gm_n62, gm_n502, gm_n432);
	nand (gm_n6554, gm_n255, gm_n72, gm_n55, gm_n6553, gm_n327);
	nor (gm_n6555, gm_n213, gm_n159, in_15, gm_n399, gm_n393);
	nand (gm_n6556, in_21, in_20, in_19, gm_n6555);
	nor (gm_n6557, gm_n72, gm_n85, in_19, gm_n4422, gm_n393);
	nand (gm_n6558, gm_n78, in_9, gm_n94, gm_n1496, gm_n1011);
	nor (gm_n6559, gm_n165, gm_n119, in_14, gm_n6558, gm_n841);
	nor (gm_n6560, gm_n274, in_16, in_12, gm_n1150, gm_n319);
	nand (gm_n6561, gm_n495, gm_n72, in_20, gm_n6560);
	nor (gm_n6562, gm_n168, gm_n158, gm_n60, gm_n196, gm_n191);
	nand (gm_n6563, gm_n72, gm_n85, gm_n56, gm_n6562);
	nor (gm_n6564, in_14, gm_n78, in_9, gm_n1698, gm_n369);
	nand (gm_n6565, gm_n436, gm_n129, in_18, gm_n6564);
	nor (gm_n6566, in_14, in_10, in_9, gm_n3721, gm_n207);
	nand (gm_n6567, gm_n367, gm_n323, gm_n119, gm_n6566);
	nor (gm_n6568, gm_n375, gm_n76, in_9, gm_n511, gm_n480);
	nand (gm_n6569, gm_n206, gm_n72, in_17, gm_n6568);
	nand (gm_n6570, gm_n6565, gm_n6563, gm_n6561, gm_n6569, gm_n6567);
	nor (gm_n6571, gm_n158, in_16, gm_n59, gm_n354, gm_n180);
	nand (gm_n6572, gm_n495, gm_n72, gm_n85, gm_n6571);
	nor (gm_n6573, gm_n358, gm_n76, gm_n62, gm_n1132, gm_n344);
	nand (gm_n6574, gm_n120, in_21, in_17, gm_n6573, gm_n339);
	nor (gm_n6575, gm_n121, gm_n76, in_9, gm_n1664, gm_n406);
	nand (gm_n6576, gm_n206, in_21, gm_n55, gm_n6575);
	nand (gm_n6577, gm_n6576, gm_n6574, gm_n6572);
	nor (gm_n6578, gm_n90, in_10, gm_n62, gm_n3660, gm_n207);
	nand (gm_n6579, gm_n200, gm_n164, in_18, gm_n6578);
	nand (gm_n6580, gm_n327, gm_n72, in_17, gm_n1279, gm_n1076);
	nand (gm_n6581, gm_n200, gm_n146, gm_n119, gm_n3514);
	nand (gm_n6582, gm_n6581, gm_n6580, gm_n6579);
	nor (gm_n6583, gm_n6570, gm_n6559, gm_n6557, gm_n6582, gm_n6577);
	nor (gm_n6584, gm_n479, in_21, gm_n55, gm_n4584, gm_n662);
	nand (gm_n6585, gm_n733, gm_n73, in_12, gm_n1186, gm_n154);
	nor (gm_n6586, gm_n781, gm_n72, in_20, gm_n6585);
	or (gm_n6587, gm_n168, gm_n115, gm_n60, gm_n2008, gm_n485);
	nor (gm_n6588, in_21, gm_n85, gm_n56, gm_n6587);
	nor (gm_n6589, gm_n6588, gm_n6586, gm_n6584);
	or (gm_n6590, gm_n227, in_16, gm_n59, gm_n1689, gm_n263);
	nor (gm_n6591, gm_n139, gm_n72, gm_n85, gm_n6590);
	or (gm_n6592, gm_n240, gm_n60, gm_n63, gm_n770, gm_n760);
	nor (gm_n6593, in_21, in_20, in_19, gm_n6592, gm_n191);
	nand (gm_n6594, gm_n125, gm_n76, gm_n62, gm_n788, gm_n126);
	nor (gm_n6595, gm_n313, in_21, gm_n55, gm_n6594, gm_n620);
	nor (gm_n6596, gm_n6595, gm_n6593, gm_n6591);
	nand (gm_n6597, gm_n6583, gm_n6556, gm_n6554, gm_n6596, gm_n6589);
	and (gm_n6598, in_14, in_10, in_9, gm_n2416, gm_n624);
	nand (gm_n6599, gm_n245, gm_n164, gm_n119, gm_n6598);
	nor (gm_n6600, gm_n213, gm_n191, in_15, gm_n764, gm_n355);
	nand (gm_n6601, gm_n72, gm_n85, gm_n56, gm_n6600);
	or (gm_n6602, gm_n662, gm_n72, in_17, gm_n4654, gm_n374);
	nand (gm_n6603, gm_n6602, gm_n6601, gm_n6599);
	and (gm_n6604, gm_n448, gm_n214, gm_n60, gm_n1179, gm_n449);
	nand (gm_n6605, in_21, in_20, in_19, gm_n6604);
	nor (gm_n6606, gm_n461, gm_n76, in_9, gm_n988, gm_n430);
	nand (gm_n6607, gm_n102, gm_n72, gm_n55, gm_n6606, gm_n405);
	nand (gm_n6608, gm_n255, in_21, gm_n55, gm_n3762, gm_n311);
	nand (gm_n6609, gm_n6608, gm_n6607, gm_n6605);
	nor (gm_n6610, gm_n6597, gm_n6552, gm_n6550, gm_n6609, gm_n6603);
	or (gm_n6611, gm_n480, gm_n76, gm_n62, gm_n988, gm_n443);
	nor (gm_n6612, gm_n441, gm_n72, in_17, gm_n6611, gm_n328);
	nand (gm_n6613, gm_n233, gm_n73, gm_n59, gm_n1095, gm_n275);
	nor (gm_n6614, gm_n139, in_21, in_20, gm_n6613);
	or (gm_n6615, gm_n358, gm_n76, gm_n62, gm_n988, gm_n344);
	nor (gm_n6616, gm_n121, in_21, gm_n55, gm_n6615, gm_n441);
	nor (gm_n6617, gm_n6616, gm_n6614, gm_n6612);
	or (gm_n6618, gm_n133, gm_n90, in_10, gm_n589, gm_n438);
	nor (gm_n6619, gm_n212, gm_n211, gm_n119, gm_n6618);
	nand (gm_n6620, in_14, in_10, gm_n62, gm_n946, gm_n600);
	nor (gm_n6621, gm_n244, gm_n841, gm_n119, gm_n6620);
	or (gm_n6622, gm_n667, in_13, gm_n62, gm_n432, gm_n480);
	nor (gm_n6623, gm_n121, in_21, gm_n55, gm_n6622, gm_n479);
	nor (gm_n6624, gm_n6623, gm_n6621, gm_n6619);
	nand (gm_n6625, gm_n6610, gm_n6548, gm_n6546, gm_n6624, gm_n6617);
	nor (gm_n6626, gm_n240, in_15, gm_n63, gm_n770, gm_n643);
	nand (gm_n6627, gm_n72, gm_n85, in_19, gm_n6626, gm_n486);
	and (gm_n6628, in_14, in_10, in_9, gm_n2416, gm_n713);
	nand (gm_n6629, gm_n131, gm_n86, in_18, gm_n6628);
	nor (gm_n6630, gm_n190, in_16, in_12, gm_n2963, gm_n220);
	nand (gm_n6631, gm_n57, in_21, gm_n85, gm_n6630);
	nand (gm_n6632, gm_n6631, gm_n6629, gm_n6627);
	nor (gm_n6633, gm_n114, gm_n73, gm_n59, gm_n1514, gm_n263);
	nand (gm_n6634, gm_n383, gm_n72, gm_n85, gm_n6633);
	nand (gm_n6635, gm_n327, in_21, in_17, gm_n4407, gm_n595);
	nor (gm_n6636, gm_n121, gm_n76, gm_n62, gm_n808, gm_n442);
	nand (gm_n6637, gm_n373, in_21, in_17, gm_n6636);
	nand (gm_n6638, gm_n6637, gm_n6635, gm_n6634);
	nor (gm_n6639, gm_n6625, gm_n6544, gm_n6542, gm_n6638, gm_n6632);
	or (gm_n6640, gm_n213, in_16, gm_n59, gm_n1859, gm_n385);
	nor (gm_n6641, gm_n496, gm_n72, in_20, gm_n6640);
	nand (gm_n6642, gm_n176, in_15, in_11, gm_n449, gm_n1144);
	nor (gm_n6643, in_21, gm_n85, gm_n56, gm_n6642, gm_n1331);
	nor (gm_n6644, gm_n103, in_21, in_17, gm_n3443, gm_n313);
	nor (gm_n6645, gm_n6644, gm_n6643, gm_n6641);
	nand (gm_n6646, gm_n64, gm_n73, gm_n59, gm_n875, gm_n571);
	nor (gm_n6647, gm_n496, in_21, gm_n85, gm_n6646);
	and (gm_n6648, gm_n174, gm_n72, gm_n55, gm_n405, gm_n209);
	nand (gm_n6649, gm_n484, gm_n143, gm_n60, gm_n1758, gm_n268);
	nor (gm_n6650, gm_n72, in_20, in_19, gm_n6649);
	nor (gm_n6651, gm_n6650, gm_n6648, gm_n6647);
	nand (gm_n6652, gm_n6639, gm_n6540, gm_n6538, gm_n6651, gm_n6645);
	and (gm_n6653, gm_n79, in_16, gm_n59, gm_n2070, gm_n275);
	nand (gm_n6654, gm_n697, gm_n72, in_20, gm_n6653);
	nor (gm_n6655, gm_n191, gm_n159, in_15, gm_n799, gm_n263);
	nand (gm_n6656, in_21, gm_n85, in_19, gm_n6655);
	or (gm_n6657, gm_n103, in_21, in_17, gm_n3501, gm_n375);
	nand (gm_n6658, gm_n6657, gm_n6656, gm_n6654);
	nor (gm_n6659, gm_n90, in_10, in_9, gm_n399, gm_n207);
	nand (gm_n6660, gm_n348, gm_n200, gm_n119, gm_n6659);
	nor (gm_n6661, gm_n155, in_16, in_12, gm_n3929, gm_n319);
	nand (gm_n6662, gm_n138, in_21, in_20, gm_n6661);
	and (gm_n6663, gm_n77, in_16, in_12, gm_n1531, gm_n79);
	nand (gm_n6664, gm_n179, in_21, gm_n85, gm_n6663);
	nand (gm_n6665, gm_n6664, gm_n6662, gm_n6660);
	nor (gm_n6666, gm_n6652, gm_n6536, gm_n6534, gm_n6665, gm_n6658);
	nand (gm_n6667, gm_n79, gm_n73, in_12, gm_n5152, gm_n949);
	nor (gm_n6668, gm_n219, gm_n72, gm_n85, gm_n6667);
	nand (gm_n6669, gm_n61, in_16, in_12, gm_n1569, gm_n222);
	nor (gm_n6670, gm_n912, gm_n72, in_20, gm_n6669);
	nand (gm_n6671, gm_n90, gm_n78, in_9, gm_n2712, gm_n713);
	nor (gm_n6672, gm_n531, gm_n212, gm_n119, gm_n6671);
	nor (gm_n6673, gm_n6672, gm_n6670, gm_n6668);
	or (gm_n6674, gm_n818, in_13, in_9, gm_n442, gm_n430);
	nor (gm_n6675, gm_n374, gm_n72, gm_n55, gm_n6674, gm_n375);
	or (gm_n6676, gm_n514, in_13, gm_n62, gm_n621, gm_n443);
	nor (gm_n6677, gm_n256, in_21, in_17, gm_n6676, gm_n620);
	or (gm_n6678, gm_n358, gm_n76, in_9, gm_n502, gm_n796);
	nor (gm_n6679, gm_n103, in_21, in_17, gm_n6678, gm_n105);
	nor (gm_n6680, gm_n6679, gm_n6677, gm_n6675);
	nand (gm_n6681, gm_n6666, gm_n6532, gm_n6530, gm_n6680, gm_n6673);
	nor (gm_n6682, gm_n290, in_15, gm_n63, gm_n761, gm_n605);
	nand (gm_n6683, in_21, gm_n85, in_19, gm_n6682, gm_n75);
	nor (gm_n6684, gm_n257, gm_n76, in_9, gm_n2256, gm_n313);
	nand (gm_n6685, gm_n254, in_21, in_17, gm_n6684);
	nand (gm_n6686, gm_n245, gm_n146, gm_n119, gm_n1860);
	nand (gm_n6687, gm_n6686, gm_n6685, gm_n6683);
	nor (gm_n6688, in_14, in_10, gm_n62, gm_n4088, gm_n467);
	nand (gm_n6689, gm_n243, gm_n88, gm_n119, gm_n6688);
	nor (gm_n6690, gm_n667, gm_n76, in_9, gm_n481, gm_n406);
	nand (gm_n6691, gm_n102, in_21, in_17, gm_n6690, gm_n1076);
	and (gm_n6692, gm_n392, gm_n60, in_11, gm_n602, gm_n170);
	nand (gm_n6693, gm_n72, in_20, in_19, gm_n6692, gm_n75);
	nand (gm_n6694, gm_n6693, gm_n6691, gm_n6689);
	nor (gm_n6695, gm_n6681, gm_n6528, gm_n6526, gm_n6694, gm_n6687);
	or (gm_n6696, in_14, in_10, gm_n62, gm_n1661, gm_n807);
	nor (gm_n6697, gm_n824, gm_n167, in_18, gm_n6696);
	or (gm_n6698, gm_n141, gm_n194, in_14, gm_n807, gm_n240);
	nor (gm_n6699, gm_n531, gm_n89, in_18, gm_n6698);
	or (gm_n6700, gm_n667, in_13, gm_n62, gm_n1132, gm_n257);
	nor (gm_n6701, gm_n479, gm_n72, gm_n55, gm_n6700, gm_n313);
	nor (gm_n6702, gm_n6701, gm_n6699, gm_n6697);
	nor (gm_n6703, in_11, gm_n78, gm_n62, gm_n463, gm_n432);
	nand (gm_n6704, gm_n192, gm_n56, gm_n60, gm_n6703, gm_n486);
	nor (gm_n6705, gm_n6704, gm_n72, gm_n85);
	or (gm_n6706, gm_n207, gm_n90, in_10, gm_n350, gm_n247);
	nor (gm_n6707, gm_n368, gm_n1989, gm_n119, gm_n6706);
	or (gm_n6708, gm_n461, gm_n76, in_9, gm_n621, gm_n502);
	nor (gm_n6709, gm_n441, gm_n72, in_17, gm_n6708, gm_n662);
	nor (gm_n6710, gm_n6709, gm_n6707, gm_n6705);
	nand (gm_n6711, gm_n6695, gm_n6525, gm_n6523, gm_n6710, gm_n6702);
	nor (gm_n6712, gm_n158, in_16, gm_n59, gm_n320, gm_n220);
	nand (gm_n6713, gm_n697, gm_n72, in_20, gm_n6712);
	nor (gm_n6714, gm_n406, gm_n76, in_9, gm_n502, gm_n481);
	nand (gm_n6715, gm_n523, gm_n72, gm_n55, gm_n6714, gm_n327);
	and (gm_n6716, in_13, in_9, gm_n94, gm_n756, gm_n340);
	nand (gm_n6717, gm_n122, gm_n72, gm_n55, gm_n6716, gm_n174);
	nand (gm_n6718, gm_n6717, gm_n6715, gm_n6713);
	nand (gm_n6719, gm_n523, gm_n72, in_17, gm_n1155, gm_n311);
	nor (gm_n6720, gm_n212, gm_n909, in_14, gm_n369, gm_n240);
	nand (gm_n6721, gm_n6720, gm_n86, in_18);
	nor (gm_n6722, gm_n90, in_10, in_9, gm_n2402, gm_n362);
	nand (gm_n6723, gm_n436, gm_n146, in_18, gm_n6722);
	nand (gm_n6724, gm_n6723, gm_n6721, gm_n6719);
	nor (gm_n6725, gm_n6711, gm_n6521, gm_n6519, gm_n6724, gm_n6718);
	nor (gm_n6726, gm_n159, gm_n89, in_18, gm_n309, gm_n824);
	nand (gm_n6727, gm_n222, gm_n392, in_15, gm_n1161, gm_n394);
	nor (gm_n6728, in_21, in_20, in_19, gm_n6727);
	nand (gm_n6729, gm_n77, gm_n73, in_12, gm_n2860, gm_n154);
	nor (gm_n6730, gm_n58, gm_n72, gm_n85, gm_n6729);
	nor (gm_n6731, gm_n6730, gm_n6728, gm_n6726);
	or (gm_n6732, gm_n90, in_10, in_9, gm_n815, gm_n133);
	nor (gm_n6733, gm_n1989, gm_n211, gm_n119, gm_n6732);
	nor (gm_n6734, gm_n256, in_21, gm_n55, gm_n2094, gm_n374);
	and (gm_n6735, gm_n120, gm_n72, gm_n55, gm_n3109, gm_n523);
	nor (gm_n6736, gm_n6735, gm_n6734, gm_n6733);
	nand (gm_n6737, gm_n6725, gm_n6516, gm_n6514, gm_n6736, gm_n6731);
	nor (gm_n6738, gm_n149, gm_n90, gm_n78, gm_n362, gm_n349);
	nand (gm_n6739, gm_n348, gm_n806, gm_n119, gm_n6738);
	nor (gm_n6740, gm_n393, gm_n263, in_15, gm_n1016, gm_n764);
	nand (gm_n6741, in_21, gm_n85, gm_n56, gm_n6740);
	nor (gm_n6742, gm_n818, in_13, in_9, gm_n596, gm_n461);
	nand (gm_n6743, gm_n120, in_21, in_17, gm_n6742, gm_n523);
	nand (gm_n6744, gm_n6743, gm_n6741, gm_n6739);
	nor (gm_n6745, gm_n196, gm_n193, gm_n60, gm_n293, gm_n274);
	nand (gm_n6746, in_21, in_20, gm_n56, gm_n6745);
	nor (gm_n6747, gm_n324, gm_n155, in_15, gm_n633, gm_n485);
	nand (gm_n6748, in_21, in_20, gm_n56, gm_n6747);
	nor (gm_n6749, gm_n290, gm_n213, in_15, gm_n520, gm_n393);
	nand (gm_n6750, in_21, gm_n85, gm_n56, gm_n6749);
	nand (gm_n6751, gm_n6750, gm_n6748, gm_n6746);
	nor (gm_n6752, gm_n6737, gm_n6512, gm_n6510, gm_n6751, gm_n6744);
	or (gm_n6753, gm_n263, gm_n168, in_15, gm_n1223, gm_n485);
	nor (gm_n6754, gm_n72, in_20, in_19, gm_n6753);
	or (gm_n6755, gm_n393, gm_n158, in_15, gm_n1689, gm_n643);
	nor (gm_n6756, gm_n72, in_20, gm_n56, gm_n6755);
	and (gm_n6757, in_21, in_20, in_19, gm_n3688, gm_n281);
	nor (gm_n6758, gm_n6757, gm_n6756, gm_n6754);
	nand (gm_n6759, gm_n264, in_16, in_12, gm_n571, gm_n265);
	nor (gm_n6760, gm_n912, in_21, gm_n85, gm_n6759);
	and (gm_n6761, gm_n348, gm_n325, in_18, gm_n436);
	nand (gm_n6762, gm_n143, gm_n73, in_12, gm_n303, gm_n216);
	nor (gm_n6763, gm_n384, gm_n72, in_20, gm_n6762);
	nor (gm_n6764, gm_n6763, gm_n6761, gm_n6760);
	nand (gm_n6765, gm_n6752, gm_n6508, gm_n6506, gm_n6764, gm_n6758);
	nor (gm_n6766, gm_n447, gm_n158, in_15, gm_n1519, gm_n643);
	nand (gm_n6767, in_21, in_20, in_19, gm_n6766);
	nor (gm_n6768, in_14, in_10, gm_n62, gm_n832, gm_n362);
	nand (gm_n6769, gm_n367, gm_n200, gm_n119, gm_n6768);
	and (gm_n6770, gm_n484, gm_n60, in_11, gm_n1929, gm_n171);
	nand (gm_n6771, gm_n72, gm_n85, in_19, gm_n6770, gm_n281);
	nand (gm_n6772, gm_n6771, gm_n6769, gm_n6767);
	nor (gm_n6773, gm_n358, gm_n76, in_9, gm_n1583, gm_n443);
	nand (gm_n6774, gm_n102, in_21, in_17, gm_n6773, gm_n122);
	nand (gm_n6775, gm_n72, gm_n85, in_19, gm_n1752, gm_n394);
	nor (gm_n6776, gm_n480, in_13, gm_n62, gm_n502, gm_n462);
	nand (gm_n6777, gm_n104, gm_n72, gm_n55, gm_n6776, gm_n174);
	nand (gm_n6778, gm_n6777, gm_n6775, gm_n6774);
	nor (gm_n6779, gm_n6765, gm_n6504, gm_n6503, gm_n6778, gm_n6772);
	or (gm_n6780, gm_n283, in_15, in_11, gm_n981, gm_n290);
	nor (gm_n6781, in_21, in_20, gm_n56, gm_n6780, gm_n485);
	or (gm_n6782, gm_n190, gm_n73, gm_n59, gm_n135, gm_n227);
	nor (gm_n6783, gm_n781, gm_n72, in_20, gm_n6782);
	nand (gm_n6784, gm_n90, gm_n78, in_9, gm_n1531, gm_n91);
	nor (gm_n6785, gm_n212, gm_n165, in_18, gm_n6784);
	nor (gm_n6786, gm_n6785, gm_n6783, gm_n6781);
	nand (gm_n6787, gm_n264, in_16, gm_n59, gm_n586, gm_n275);
	nor (gm_n6788, gm_n912, gm_n72, gm_n85, gm_n6787);
	or (gm_n6789, gm_n514, in_13, gm_n62, gm_n462, gm_n596);
	nor (gm_n6790, gm_n121, gm_n72, gm_n55, gm_n6789, gm_n441);
	or (gm_n6791, gm_n147, gm_n90, gm_n78, gm_n491, gm_n248);
	nor (gm_n6792, gm_n1989, gm_n165, gm_n119, gm_n6791);
	nor (gm_n6793, gm_n6792, gm_n6790, gm_n6788);
	nand (gm_n6794, gm_n6779, gm_n6501, gm_n6499, gm_n6793, gm_n6786);
	nor (gm_n6795, gm_n461, in_13, gm_n62, gm_n743, gm_n430);
	nand (gm_n6796, gm_n122, in_21, in_17, gm_n6795, gm_n327);
	nand (gm_n6797, gm_n291, in_12, gm_n94, gm_n214, gm_n160);
	nor (gm_n6798, gm_n58, gm_n85, in_16, gm_n6797, gm_n354);
	nand (gm_n6799, gm_n6798, in_21);
	nor (gm_n6800, gm_n207, gm_n90, in_10, gm_n438, gm_n389);
	nand (gm_n6801, gm_n436, gm_n129, gm_n119, gm_n6800);
	nand (gm_n6802, gm_n6801, gm_n6799, gm_n6796);
	nor (gm_n6803, gm_n605, gm_n467, gm_n90, gm_n842);
	nand (gm_n6804, gm_n436, gm_n86, gm_n119, gm_n6803);
	nor (gm_n6805, gm_n239, gm_n60, gm_n63, gm_n2017, gm_n633);
	nand (gm_n6806, gm_n72, gm_n85, gm_n56, gm_n6805, gm_n448);
	nor (gm_n6807, gm_n115, in_16, in_12, gm_n1324, gm_n319);
	nand (gm_n6808, gm_n138, gm_n72, in_20, gm_n6807);
	nand (gm_n6809, gm_n6808, gm_n6806, gm_n6804);
	nor (gm_n6810, gm_n6794, gm_n6497, gm_n6495, gm_n6809, gm_n6802);
	nor (gm_n6811, gm_n406, in_13, in_9, gm_n743, gm_n502);
	nand (gm_n6812, gm_n122, gm_n72, gm_n55, gm_n6811, gm_n174);
	nand (gm_n6813, gm_n174, in_21, gm_n55, gm_n3588, gm_n523);
	nor (gm_n6814, gm_n461, gm_n76, gm_n62, gm_n502, gm_n359);
	nand (gm_n6815, gm_n174, in_21, in_17, gm_n6814, gm_n595);
	nand (gm_n6816, gm_n6812, gm_n6810, gm_n6493, gm_n6815, gm_n6813);
	and (gm_n6817, gm_n104, in_13, in_9, gm_n1359, gm_n314);
	nand (gm_n6818, gm_n373, in_21, in_17, gm_n6817);
	nand (gm_n6819, gm_n243, gm_n806, in_18, gm_n5323);
	and (gm_n6820, gm_n106, in_13, gm_n62, gm_n3679, gm_n339);
	nand (gm_n6821, gm_n311, in_21, in_17, gm_n6820);
	nand (gm_n6822, gm_n6821, gm_n6819, gm_n6818);
	or (gm_n6823, gm_n406, in_13, gm_n62, gm_n345, gm_n344);
	nor (gm_n6824, gm_n479, in_21, gm_n55, gm_n6823, gm_n375);
	nor (out_19, gm_n6822, gm_n6816, gm_n6491, gm_n6824);
	nand (gm_n6826, gm_n76, in_9, in_8, gm_n1496, gm_n579);
	nor (gm_n6827, gm_n183, gm_n72, gm_n55, gm_n6826, gm_n313);
	and (gm_n6828, gm_n255, in_13, in_9, gm_n615, gm_n340);
	nand (gm_n6829, gm_n102, gm_n72, in_17, gm_n6828);
	or (gm_n6830, gm_n114, gm_n73, gm_n59, gm_n2357, gm_n213);
	nor (gm_n6831, gm_n262, gm_n72, in_20, gm_n6830);
	or (gm_n6832, gm_n430, in_13, gm_n62, gm_n621, gm_n480);
	nor (gm_n6833, gm_n105, gm_n72, in_17, gm_n6832, gm_n388);
	and (gm_n6834, gm_n523, in_13, gm_n62, gm_n4926, gm_n788);
	nand (gm_n6835, gm_n254, in_21, in_17, gm_n6834);
	nor (gm_n6836, gm_n609, in_13, gm_n62, gm_n345, gm_n406);
	nand (gm_n6837, gm_n174, gm_n72, gm_n55, gm_n6836, gm_n1076);
	or (gm_n6838, gm_n190, gm_n59, in_8, gm_n508, gm_n152);
	nor (gm_n6839, in_21, gm_n85, gm_n73, gm_n6838, gm_n219);
	nand (gm_n6840, gm_n392, gm_n75, gm_n60, gm_n1841, gm_n222);
	nor (gm_n6841, in_21, in_20, gm_n56, gm_n6840);
	nor (gm_n6842, gm_n90, gm_n78, gm_n62, gm_n2474, gm_n369);
	nand (gm_n6843, gm_n806, gm_n129, gm_n119, gm_n6842);
	nor (gm_n6844, gm_n431, in_13, gm_n62, gm_n481, gm_n463);
	nand (gm_n6845, gm_n254, gm_n72, in_17, gm_n6844, gm_n595);
	nand (gm_n6846, gm_n123, gm_n76, in_9, gm_n3876, gm_n255);
	nor (gm_n6847, gm_n374, in_21, gm_n55, gm_n6846);
	or (gm_n6848, gm_n92, gm_n78, gm_n62, gm_n502, gm_n866);
	nor (gm_n6849, gm_n212, gm_n119, in_14, gm_n6848, gm_n368);
	nor (gm_n6850, gm_n247, in_14, in_10, gm_n467, gm_n350);
	nand (gm_n6851, gm_n166, gm_n164, in_18, gm_n6850);
	and (gm_n6852, gm_n77, in_16, gm_n59, gm_n936, gm_n79);
	nand (gm_n6853, gm_n113, gm_n72, gm_n85, gm_n6852);
	or (gm_n6854, gm_n147, gm_n90, gm_n78, gm_n775, gm_n349);
	nor (gm_n6855, gm_n368, gm_n212, gm_n119, gm_n6854);
	or (gm_n6856, gm_n287, in_14, in_10, gm_n526, gm_n362);
	nor (gm_n6857, gm_n841, gm_n211, in_18, gm_n6856);
	nor (gm_n6858, gm_n358, in_13, in_9, gm_n463, gm_n866);
	nand (gm_n6859, gm_n122, gm_n72, in_17, gm_n6858, gm_n206);
	nor (gm_n6860, gm_n90, gm_n78, in_9, gm_n835, gm_n369);
	nand (gm_n6861, gm_n146, gm_n131, gm_n119, gm_n6860);
	nand (gm_n6862, in_14, in_10, gm_n62, gm_n1001, gm_n91);
	nor (gm_n6863, gm_n824, gm_n89, gm_n119, gm_n6862);
	nand (gm_n6864, gm_n122, in_13, in_12, gm_n2885, gm_n264);
	nor (gm_n6865, gm_n479, in_21, in_17, gm_n6864);
	nor (gm_n6866, gm_n447, gm_n158, in_15, gm_n2931, gm_n633);
	nand (gm_n6867, gm_n72, gm_n85, in_19, gm_n6866);
	nor (gm_n6868, gm_n207, gm_n90, gm_n78, gm_n414, gm_n287);
	nand (gm_n6869, gm_n243, gm_n88, gm_n119, gm_n6868);
	nand (gm_n6870, gm_n579, gm_n1157, gm_n76, gm_n722, gm_n339);
	nor (gm_n6871, gm_n620, in_21, in_17, gm_n6870);
	or (gm_n6872, gm_n514, in_13, in_9, gm_n743, gm_n502);
	nor (gm_n6873, gm_n105, gm_n72, in_17, gm_n6872, gm_n441);
	nor (gm_n6874, gm_n514, in_13, in_9, gm_n2823, gm_n375);
	nand (gm_n6875, gm_n206, in_21, gm_n55, gm_n6874);
	and (gm_n6876, gm_n123, in_13, gm_n62, gm_n1049, gm_n187);
	nand (gm_n6877, gm_n405, in_21, in_17, gm_n6876, gm_n373);
	or (gm_n6878, gm_n259, gm_n90, in_10, gm_n362, gm_n349);
	nor (gm_n6879, gm_n1989, gm_n87, gm_n119, gm_n6878);
	nand (gm_n6880, gm_n79, in_16, in_12, gm_n803, gm_n949);
	nor (gm_n6881, gm_n496, gm_n72, in_20, gm_n6880);
	nor (gm_n6882, gm_n855, gm_n760, gm_n190);
	nand (gm_n6883, gm_n367, gm_n200, in_18, gm_n6882);
	nor (gm_n6884, gm_n406, in_13, in_9, gm_n597, gm_n443);
	nand (gm_n6885, gm_n102, gm_n72, gm_n55, gm_n6884, gm_n1076);
	or (gm_n6886, gm_n358, gm_n76, gm_n62, gm_n443, gm_n359);
	nor (gm_n6887, gm_n388, in_21, in_17, gm_n6886, gm_n256);
	or (gm_n6888, gm_n115, gm_n74, in_15, gm_n799, gm_n193);
	nor (gm_n6889, in_21, in_20, gm_n56, gm_n6888);
	nor (gm_n6890, gm_n114, in_12, in_8, gm_n913, gm_n213);
	nand (gm_n6891, gm_n72, gm_n85, in_16, gm_n6890, gm_n113);
	and (gm_n6892, gm_n949, gm_n79, gm_n59, gm_n1456);
	nand (gm_n6893, gm_n72, gm_n85, in_19, gm_n6892, gm_n379);
	nor (gm_n6894, gm_n313, in_21, in_17, gm_n6063, gm_n620);
	nand (gm_n6895, gm_n90, gm_n78, gm_n62, gm_n1401, gm_n532);
	nor (gm_n6896, gm_n1989, gm_n87, gm_n119, gm_n6895);
	nor (gm_n6897, gm_n297, gm_n73, in_12, gm_n4917, gm_n152);
	nand (gm_n6898, gm_n57, gm_n72, in_20, gm_n6897);
	nor (gm_n6899, gm_n256, in_13, gm_n62, gm_n480, gm_n329);
	nand (gm_n6900, gm_n206, in_21, gm_n55, gm_n6899);
	nor (gm_n6901, gm_n207, in_14, in_10, gm_n389, gm_n349);
	nand (gm_n6902, gm_n245, gm_n164, in_18, gm_n6901);
	nor (gm_n6903, gm_n115, gm_n73, in_12, gm_n657, gm_n354);
	nand (gm_n6904, gm_n697, gm_n72, gm_n85, gm_n6903);
	nor (gm_n6905, gm_n514, gm_n76, gm_n62, gm_n481, gm_n430);
	nand (gm_n6906, gm_n104, in_21, in_17, gm_n6905, gm_n120);
	nand (gm_n6907, gm_n6902, gm_n6900, gm_n6898, gm_n6906, gm_n6904);
	nor (gm_n6908, gm_n158, gm_n73, in_12, gm_n2029, gm_n385);
	nand (gm_n6909, gm_n495, in_21, in_20, gm_n6908);
	nor (gm_n6910, gm_n114, in_16, in_12, gm_n1719, gm_n213);
	nand (gm_n6911, gm_n697, in_21, gm_n85, gm_n6910);
	nor (gm_n6912, gm_n114, gm_n73, in_12, gm_n1125, gm_n190);
	nand (gm_n6913, gm_n113, gm_n72, in_20, gm_n6912);
	nand (gm_n6914, gm_n6913, gm_n6911, gm_n6909);
	and (gm_n6915, gm_n303, t_7, gm_n73);
	nand (gm_n6916, gm_n138, in_21, in_20, gm_n6915);
	nor (gm_n6917, gm_n90, in_13, in_12, gm_n1719, gm_n158);
	nand (gm_n6918, gm_n164, gm_n88, in_18, gm_n6917);
	nor (gm_n6919, gm_n76, in_9, in_8, gm_n842, gm_n431);
	nand (gm_n6920, gm_n311, in_21, gm_n55, gm_n6919, gm_n1076);
	nand (gm_n6921, gm_n6920, gm_n6918, gm_n6916);
	nor (gm_n6922, gm_n6907, gm_n6896, gm_n6894, gm_n6921, gm_n6914);
	or (gm_n6923, gm_n807, gm_n90, in_10, gm_n376, gm_n349);
	nor (gm_n6924, gm_n824, gm_n89, gm_n119, gm_n6923);
	nand (gm_n6925, gm_n2193, gm_n90, gm_n78, gm_n335, gm_n532);
	nor (gm_n6926, gm_n246, gm_n130, in_18, gm_n6925);
	nand (gm_n6927, gm_n222, gm_n379, gm_n60, gm_n751, gm_n449);
	nor (gm_n6928, gm_n72, in_20, in_19, gm_n6927);
	nor (gm_n6929, gm_n6928, gm_n6926, gm_n6924);
	or (gm_n6930, gm_n406, gm_n76, in_9, gm_n743, gm_n443);
	nor (gm_n6931, gm_n103, in_21, in_17, gm_n6930, gm_n662);
	nand (gm_n6932, gm_n721, gm_n90, gm_n78, gm_n793, gm_n1158);
	nor (gm_n6933, gm_n841, gm_n165, in_18, gm_n6932);
	or (gm_n6934, gm_n430, in_13, in_9, gm_n481, gm_n406);
	nor (gm_n6935, gm_n183, in_21, in_17, gm_n6934, gm_n256);
	nor (gm_n6936, gm_n6935, gm_n6933, gm_n6931);
	nand (gm_n6937, gm_n6922, gm_n6893, gm_n6891, gm_n6936, gm_n6929);
	nor (gm_n6938, gm_n297, gm_n73, gm_n59, gm_n552, gm_n319);
	nand (gm_n6939, gm_n495, in_21, in_20, gm_n6938);
	nor (gm_n6940, gm_n190, in_16, in_12, gm_n1542, gm_n354);
	nand (gm_n6941, gm_n697, in_21, in_20, gm_n6940);
	nor (gm_n6942, gm_n115, gm_n74, in_15, gm_n552, gm_n290);
	nand (gm_n6943, gm_n72, in_20, gm_n56, gm_n6942);
	nand (gm_n6944, gm_n6943, gm_n6941, gm_n6939);
	nor (gm_n6945, in_14, in_10, gm_n62, gm_n320, gm_n92);
	nand (gm_n6946, gm_n245, gm_n129, gm_n119, gm_n6945);
	nor (gm_n6947, gm_n359, in_13, in_9, gm_n502, gm_n442);
	nand (gm_n6948, gm_n254, gm_n72, in_17, gm_n6947, gm_n595);
	and (gm_n6949, in_14, gm_n78, gm_n62, gm_n626, gm_n532);
	nand (gm_n6950, gm_n806, gm_n199, gm_n119, gm_n6949);
	nand (gm_n6951, gm_n6950, gm_n6948, gm_n6946);
	nor (gm_n6952, gm_n6937, gm_n6889, gm_n6887, gm_n6951, gm_n6944);
	nor (gm_n6953, gm_n184, gm_n72, gm_n55, gm_n1199, gm_n312);
	nand (gm_n6954, gm_n264, in_16, gm_n59, gm_n1135, gm_n275);
	nor (gm_n6955, gm_n58, in_21, gm_n85, gm_n6954);
	nand (gm_n6956, gm_n126, in_13, gm_n62, gm_n1049, gm_n314);
	nor (gm_n6957, gm_n328, in_21, gm_n55, gm_n6956, gm_n374);
	nor (gm_n6958, gm_n6957, gm_n6955, gm_n6953);
	or (gm_n6959, gm_n514, gm_n76, gm_n62, gm_n988, gm_n430);
	nor (gm_n6960, gm_n313, gm_n72, in_17, gm_n6959, gm_n374);
	or (gm_n6961, gm_n159, gm_n56, in_15, gm_n5552, gm_n447);
	nor (gm_n6962, gm_n6961, gm_n72, in_20);
	or (gm_n6963, gm_n406, gm_n76, in_9, gm_n463, gm_n359);
	nor (gm_n6964, gm_n103, in_21, gm_n55, gm_n6963, gm_n121);
	nor (gm_n6965, gm_n6964, gm_n6962, gm_n6960);
	nand (gm_n6966, gm_n6952, gm_n6885, gm_n6883, gm_n6965, gm_n6958);
	nor (gm_n6967, gm_n227, gm_n73, in_12, gm_n511, gm_n213);
	nand (gm_n6968, gm_n113, gm_n72, in_20, gm_n6967);
	nor (gm_n6969, gm_n76, gm_n62, in_8, gm_n407, gm_n406);
	nand (gm_n6970, gm_n120, in_21, in_17, gm_n6969, gm_n405);
	and (gm_n6971, gm_n79, gm_n76, gm_n59, gm_n919);
	nand (gm_n6972, gm_n104, gm_n72, gm_n55, gm_n6971, gm_n327);
	nand (gm_n6973, gm_n6972, gm_n6970, gm_n6968);
	nor (gm_n6974, gm_n297, gm_n73, gm_n59, gm_n2077, gm_n276);
	nand (gm_n6975, gm_n57, gm_n72, in_20, gm_n6974);
	nor (gm_n6976, gm_n168, gm_n60, gm_n63, gm_n770, gm_n541);
	nand (gm_n6977, in_21, gm_n85, gm_n56, gm_n6976, gm_n448);
	and (gm_n6978, in_14, in_10, in_9, gm_n1001, gm_n532);
	nand (gm_n6979, gm_n245, gm_n146, gm_n119, gm_n6978);
	nand (gm_n6980, gm_n6979, gm_n6977, gm_n6975);
	nor (gm_n6981, gm_n6966, gm_n6881, gm_n6879, gm_n6980, gm_n6973);
	nand (gm_n6982, gm_n555, gm_n1011, gm_n176);
	nor (gm_n6983, gm_n824, gm_n119, gm_n90, gm_n6982, gm_n437);
	nor (gm_n6984, gm_n437, gm_n165, gm_n119, gm_n4995);
	or (gm_n6985, gm_n596, in_13, gm_n62, gm_n1583, gm_n480);
	nor (gm_n6986, gm_n183, gm_n72, gm_n55, gm_n6985, gm_n375);
	nor (gm_n6987, gm_n6986, gm_n6984, gm_n6983);
	or (gm_n6988, gm_n430, gm_n76, gm_n62, gm_n359, gm_n257);
	nor (gm_n6989, gm_n103, in_21, gm_n55, gm_n6988, gm_n662);
	nand (gm_n6990, gm_n2193, in_14, gm_n78, gm_n490, gm_n600);
	nor (gm_n6991, gm_n841, gm_n824, in_18, gm_n6990);
	nand (gm_n6992, gm_n214, gm_n73, gm_n59, gm_n612, gm_n949);
	nor (gm_n6993, gm_n139, gm_n72, gm_n85, gm_n6992);
	nor (gm_n6994, gm_n6993, gm_n6991, gm_n6989);
	nand (gm_n6995, gm_n6981, gm_n6877, gm_n6875, gm_n6994, gm_n6987);
	nor (gm_n6996, gm_n297, in_16, gm_n59, gm_n4917, gm_n319);
	nand (gm_n6997, gm_n179, gm_n72, in_20, gm_n6996);
	nand (gm_n6998, gm_n122, gm_n72, gm_n55, gm_n1932, gm_n174);
	and (gm_n6999, gm_n214, gm_n484, gm_n60, gm_n1179, gm_n268);
	nand (gm_n7000, gm_n72, gm_n85, in_19, gm_n6999);
	nand (gm_n7001, gm_n7000, gm_n6998, gm_n6997);
	or (gm_n7002, gm_n72, gm_n85, gm_n56, gm_n3988, gm_n447);
	nor (gm_n7003, in_14, gm_n59, in_8, gm_n2769, gm_n190);
	nand (gm_n7004, gm_n146, in_18, gm_n76, gm_n7003, gm_n436);
	nor (gm_n7005, gm_n358, gm_n76, gm_n62, gm_n432, gm_n344);
	nand (gm_n7006, gm_n102, in_21, gm_n55, gm_n7005, gm_n405);
	nand (gm_n7007, gm_n7006, gm_n7004, gm_n7002);
	nor (gm_n7008, gm_n6995, gm_n6873, gm_n6871, gm_n7007, gm_n7001);
	and (gm_n7009, gm_n72, gm_n85, in_19, gm_n5127, gm_n486);
	or (gm_n7010, gm_n115, in_16, in_12, gm_n1332, gm_n276);
	nor (gm_n7011, gm_n262, in_21, gm_n85, gm_n7010);
	or (gm_n7012, gm_n158, in_16, in_12, gm_n832, gm_n354);
	nor (gm_n7013, gm_n384, in_21, gm_n85, gm_n7012);
	nor (gm_n7014, gm_n7013, gm_n7011, gm_n7009);
	nand (gm_n7015, gm_n64, in_16, in_12, gm_n586, gm_n949);
	nor (gm_n7016, gm_n781, in_21, gm_n85, gm_n7015);
	or (gm_n7017, in_14, in_10, gm_n62, gm_n705, gm_n92);
	nor (gm_n7018, gm_n244, gm_n212, gm_n119, gm_n7017);
	or (gm_n7019, gm_n807, in_14, in_10, gm_n389, gm_n370);
	nor (gm_n7020, gm_n1989, gm_n824, in_18, gm_n7019);
	nor (gm_n7021, gm_n7020, gm_n7018, gm_n7016);
	nand (gm_n7022, gm_n7008, gm_n6869, gm_n6867, gm_n7021, gm_n7014);
	and (gm_n7023, gm_n90, gm_n78, in_9, gm_n1030, gm_n334);
	nand (gm_n7024, gm_n131, gm_n86, in_18, gm_n7023);
	and (gm_n7025, gm_n187, gm_n76, gm_n62, gm_n341, gm_n314);
	nand (gm_n7026, gm_n405, in_21, gm_n55, gm_n7025, gm_n373);
	nor (gm_n7027, gm_n297, gm_n73, in_12, gm_n2077, gm_n354);
	nand (gm_n7028, gm_n57, gm_n72, in_20, gm_n7027);
	nand (gm_n7029, gm_n7028, gm_n7026, gm_n7024);
	nor (gm_n7030, gm_n514, gm_n76, gm_n62, gm_n743, gm_n430);
	nand (gm_n7031, gm_n102, in_21, gm_n55, gm_n7030, gm_n122);
	nor (gm_n7032, gm_n514, gm_n76, in_9, gm_n597, gm_n596);
	nand (gm_n7033, gm_n104, in_21, gm_n55, gm_n7032, gm_n120);
	and (gm_n7034, in_14, gm_n78, in_9, gm_n2497, gm_n713);
	nand (gm_n7035, gm_n436, gm_n348, gm_n119, gm_n7034);
	nand (gm_n7036, gm_n7035, gm_n7033, gm_n7031);
	nor (gm_n7037, gm_n7022, gm_n6865, gm_n6863, gm_n7036, gm_n7029);
	or (gm_n7038, in_13, in_9, in_8, gm_n2769, gm_n442);
	nor (gm_n7039, gm_n620, gm_n72, gm_n55, gm_n7038, gm_n328);
	or (gm_n7040, gm_n90, gm_n78, gm_n62, gm_n654, gm_n133);
	nor (gm_n7041, gm_n246, gm_n87, in_18, gm_n7040);
	or (gm_n7042, gm_n259, in_14, in_10, gm_n370, gm_n362);
	nor (gm_n7043, gm_n246, gm_n87, gm_n119, gm_n7042);
	nor (gm_n7044, gm_n7043, gm_n7041, gm_n7039);
	or (gm_n7045, gm_n667, gm_n76, in_9, gm_n480, gm_n345);
	nor (gm_n7046, gm_n388, in_21, gm_n55, gm_n7045, gm_n662);
	nor (gm_n7047, in_21, in_20, gm_n56, gm_n2097, gm_n191);
	or (gm_n7048, gm_n263, in_12, in_8, gm_n2690, gm_n354);
	nor (gm_n7049, gm_n72, gm_n85, gm_n73, gm_n7048, gm_n262);
	nor (gm_n7050, gm_n7049, gm_n7047, gm_n7046);
	nand (gm_n7051, gm_n7037, gm_n6861, gm_n6859, gm_n7050, gm_n7044);
	nor (gm_n7052, gm_n246, gm_n274, in_18, gm_n2060, gm_n290);
	nand (gm_n7053, gm_n7052, gm_n348);
	nor (gm_n7054, gm_n293, gm_n190, in_15, gm_n932, gm_n633);
	nand (gm_n7055, gm_n72, gm_n85, in_19, gm_n7054);
	nor (gm_n7056, gm_n514, gm_n76, in_9, gm_n2198, gm_n313);
	nand (gm_n7057, gm_n174, gm_n72, in_17, gm_n7056);
	nand (gm_n7058, gm_n7057, gm_n7055, gm_n7053);
	and (gm_n7059, gm_n264, in_16, in_12, gm_n2646, gm_n275);
	nand (gm_n7060, gm_n383, gm_n72, gm_n85, gm_n7059);
	nand (gm_n7061, in_21, in_20, in_19, gm_n6626, gm_n281);
	nor (gm_n7062, gm_n191, in_19, gm_n60, gm_n5552, gm_n290);
	nand (gm_n7063, gm_n7062, gm_n72, gm_n85);
	nand (gm_n7064, gm_n7063, gm_n7061, gm_n7060);
	nor (gm_n7065, gm_n7051, gm_n6857, gm_n6855, gm_n7064, gm_n7058);
	nor (gm_n7066, gm_n165, in_18, gm_n55, gm_n1449);
	or (gm_n7067, gm_n514, gm_n76, gm_n62, gm_n730, gm_n184);
	nor (gm_n7068, gm_n620, in_21, gm_n55, gm_n7067);
	and (gm_n7069, gm_n72, in_20, gm_n56, gm_n4573, gm_n75);
	nor (gm_n7070, gm_n7069, gm_n7068, gm_n7066);
	or (gm_n7071, gm_n158, in_16, gm_n59, gm_n4437, gm_n276);
	nor (gm_n7072, gm_n496, in_21, gm_n85, gm_n7071);
	nand (gm_n7073, gm_n449, in_15, gm_n63, gm_n3818, gm_n1942);
	nor (gm_n7074, gm_n72, gm_n85, in_19, gm_n7073, gm_n269);
	nand (gm_n7075, gm_n449, gm_n264, in_15, gm_n2096, gm_n486);
	nor (gm_n7076, gm_n72, gm_n85, in_19, gm_n7075);
	nor (gm_n7077, gm_n7076, gm_n7074, gm_n7072);
	nand (gm_n7078, gm_n7065, gm_n6853, gm_n6851, gm_n7077, gm_n7070);
	and (gm_n7079, gm_n90, in_10, gm_n62, gm_n2443, gm_n1011);
	nand (gm_n7080, gm_n806, gm_n164, gm_n119, gm_n7079);
	nor (gm_n7081, gm_n461, in_13, in_9, gm_n743, gm_n344);
	nand (gm_n7082, gm_n104, gm_n72, gm_n55, gm_n7081, gm_n206);
	nor (gm_n7083, gm_n147, gm_n90, in_10, gm_n349, gm_n259);
	nand (gm_n7084, gm_n367, gm_n323, in_18, gm_n7083);
	nand (gm_n7085, gm_n7084, gm_n7082, gm_n7080);
	nand (gm_n7086, in_21, gm_n85, gm_n56, gm_n1525, gm_n75);
	nor (gm_n7087, gm_n406, gm_n76, in_9, gm_n988, gm_n502);
	nand (gm_n7088, gm_n311, gm_n72, in_17, gm_n7087, gm_n1076);
	and (gm_n7089, in_14, gm_n78, gm_n62, gm_n2608, gm_n532);
	nand (gm_n7090, gm_n245, gm_n129, gm_n119, gm_n7089);
	nand (gm_n7091, gm_n7090, gm_n7088, gm_n7086);
	nor (gm_n7092, gm_n7078, gm_n6849, gm_n6847, gm_n7091, gm_n7085);
	or (gm_n7093, gm_n358, in_13, in_9, gm_n988, gm_n430);
	nor (gm_n7094, gm_n256, in_21, in_17, gm_n7093, gm_n620);
	nand (gm_n7095, gm_n143, gm_n75, in_15, gm_n678, gm_n1398);
	nor (gm_n7096, in_21, gm_n85, in_19, gm_n7095);
	or (gm_n7097, gm_n431, in_13, in_9, gm_n597, gm_n596);
	nor (gm_n7098, gm_n183, gm_n72, gm_n55, gm_n7097, gm_n256);
	nor (gm_n7099, gm_n7098, gm_n7096, gm_n7094);
	nand (gm_n7100, gm_n143, in_16, in_12, gm_n991, gm_n275);
	nor (gm_n7101, gm_n262, in_21, gm_n85, gm_n7100);
	nand (gm_n7102, gm_n281, gm_n154, in_15, gm_n1531, gm_n422);
	nor (gm_n7103, in_21, in_20, in_19, gm_n7102);
	nand (gm_n7104, gm_n405, gm_n828, in_13, gm_n793, gm_n788);
	nor (gm_n7105, gm_n479, in_21, gm_n55, gm_n7104);
	nor (gm_n7106, gm_n7105, gm_n7103, gm_n7101);
	nand (gm_n7107, gm_n7092, gm_n6845, gm_n6843, gm_n7106, gm_n7099);
	nor (gm_n7108, gm_n99, gm_n90, in_10, gm_n148, gm_n147);
	nand (gm_n7109, gm_n348, gm_n323, gm_n119, gm_n7108);
	nand (gm_n7110, gm_n311, in_21, in_17, gm_n4924, gm_n339);
	nor (gm_n7111, in_14, in_10, gm_n62, gm_n821, gm_n207);
	nand (gm_n7112, gm_n806, gm_n146, gm_n119, gm_n7111);
	nand (gm_n7113, gm_n7112, gm_n7110, gm_n7109);
	and (gm_n7114, in_13, in_9, in_8, gm_n1929, gm_n123);
	nand (gm_n7115, gm_n120, gm_n72, in_17, gm_n7114, gm_n122);
	nor (gm_n7116, gm_n461, gm_n76, in_9, gm_n345, gm_n596);
	nand (gm_n7117, gm_n206, in_21, gm_n55, gm_n7116, gm_n595);
	nor (gm_n7118, gm_n358, gm_n76, gm_n62, gm_n443, gm_n345);
	nand (gm_n7119, gm_n405, gm_n72, gm_n55, gm_n7118, gm_n373);
	nand (gm_n7120, gm_n7119, gm_n7117, gm_n7115);
	nor (gm_n7121, gm_n7107, gm_n6841, gm_n6839, gm_n7120, gm_n7113);
	nor (gm_n7122, gm_n441, gm_n72, gm_n55, gm_n2321, gm_n375);
	and (gm_n7123, gm_n367, gm_n806, gm_n119, gm_n6917);
	nand (gm_n7124, in_14, gm_n78, gm_n62, gm_n1451, gm_n532);
	nor (gm_n7125, gm_n130, gm_n89, gm_n119, gm_n7124);
	nor (gm_n7126, gm_n7125, gm_n7123, gm_n7122);
	nand (gm_n7127, gm_n77, gm_n73, gm_n59, gm_n264, gm_n82);
	nor (gm_n7128, gm_n58, gm_n72, gm_n85, gm_n7127);
	nand (gm_n7129, gm_n484, gm_n64, in_15, gm_n486, gm_n306);
	nor (gm_n7130, in_21, gm_n85, in_19, gm_n7129);
	or (gm_n7131, gm_n158, gm_n60, gm_n94, gm_n633, gm_n508);
	nor (gm_n7132, gm_n72, in_20, in_19, gm_n7131, gm_n293);
	nor (gm_n7133, gm_n7132, gm_n7130, gm_n7128);
	nand (gm_n7134, gm_n7121, gm_n6837, gm_n6835, gm_n7133, gm_n7126);
	nor (gm_n7135, gm_n1331, gm_n158, gm_n60, gm_n2826, gm_n290);
	nand (gm_n7136, in_21, gm_n85, gm_n56, gm_n7135);
	nor (gm_n7137, gm_n115, in_16, gm_n59, gm_n887, gm_n152);
	nand (gm_n7138, gm_n296, in_21, in_20, gm_n7137);
	or (gm_n7139, gm_n121, gm_n72, gm_n55, gm_n3957, gm_n479);
	nand (gm_n7140, gm_n7139, gm_n7138, gm_n7136);
	nor (gm_n7141, gm_n358, in_13, gm_n62, gm_n1583, gm_n502);
	nand (gm_n7142, gm_n373, gm_n72, in_17, gm_n7141, gm_n1076);
	nand (gm_n7143, gm_n72, gm_n85, gm_n56, gm_n2372, gm_n1101);
	nor (gm_n7144, gm_n430, in_13, gm_n62, gm_n480, gm_n345);
	nand (gm_n7145, gm_n254, in_21, gm_n55, gm_n7144, gm_n595);
	nand (gm_n7146, gm_n7145, gm_n7143, gm_n7142);
	nor (gm_n7147, gm_n7134, gm_n6833, gm_n6831, gm_n7146, gm_n7140);
	nor (gm_n7148, gm_n257, gm_n76, gm_n62, gm_n743, gm_n344);
	nand (gm_n7149, gm_n174, in_21, in_17, gm_n7148, gm_n405);
	nor (gm_n7150, gm_n207, gm_n95, in_10, gm_n248);
	nand (gm_n7151, gm_n104, gm_n72, gm_n55, gm_n7150, gm_n254);
	and (gm_n7152, in_14, in_10, gm_n62, gm_n2416, gm_n334);
	nand (gm_n7153, gm_n199, gm_n166, in_18, gm_n7152);
	nand (gm_n7154, gm_n7149, gm_n7147, gm_n6829, gm_n7153, gm_n7151);
	or (gm_n7155, gm_n183, in_21, gm_n55, gm_n4435);
	nand (gm_n7156, gm_n245, gm_n164, in_18, gm_n6257);
	nor (gm_n7157, gm_n148, gm_n90, gm_n78, gm_n526, gm_n207);
	nand (gm_n7158, gm_n436, gm_n199, in_18, gm_n7157);
	nand (gm_n7159, gm_n7158, gm_n7156, gm_n7155);
	or (gm_n7160, gm_n207, in_14, in_10, gm_n491, gm_n259);
	nor (gm_n7161, gm_n368, gm_n132, gm_n119, gm_n7160);
	nor (out_20, gm_n7159, gm_n7154, gm_n6827, gm_n7161);
	or (gm_n7163, gm_n193, gm_n297, gm_n60, gm_n3382, gm_n447);
	nor (gm_n7164, in_21, in_20, in_19, gm_n7163);
	nor (gm_n7165, gm_n643, in_15, gm_n63, gm_n2017, gm_n770);
	nand (gm_n7166, in_21, gm_n85, in_19, gm_n7165, gm_n394);
	nor (gm_n7167, gm_n349, gm_n90, in_10, gm_n369, gm_n350);
	nand (gm_n7168, gm_n166, gm_n164, gm_n119, gm_n7167);
	or (gm_n7169, gm_n431, gm_n76, in_9, gm_n1583, gm_n344);
	nor (gm_n7170, gm_n184, gm_n72, in_17, gm_n7169, gm_n312);
	nand (gm_n7171, gm_n79, gm_n75, gm_n60, gm_n1179, gm_n392);
	nor (gm_n7172, gm_n72, gm_n85, gm_n56, gm_n7171);
	nor (gm_n7173, gm_n158, gm_n59, in_8, gm_n417, gm_n276);
	nand (gm_n7174, in_21, gm_n85, in_16, gm_n7173, gm_n57);
	nor (gm_n7175, gm_n259, gm_n90, in_10, gm_n349, gm_n807);
	nand (gm_n7176, gm_n436, gm_n164, in_18, gm_n7175);
	nand (gm_n7177, gm_n235, gm_n76, gm_n62, gm_n788, gm_n595);
	nor (gm_n7178, gm_n388, in_21, gm_n55, gm_n7177);
	or (gm_n7179, gm_n158, gm_n73, gm_n59, gm_n1260, gm_n220);
	nor (gm_n7180, gm_n384, in_21, gm_n85, gm_n7179);
	nor (gm_n7181, gm_n796, in_13, gm_n62, gm_n463, gm_n431);
	nand (gm_n7182, gm_n104, in_21, gm_n55, gm_n7181, gm_n254);
	nand (gm_n7183, gm_n122, in_21, in_17, gm_n6971, gm_n174);
	or (gm_n7184, gm_n514, gm_n76, in_9, gm_n359, gm_n609);
	nor (gm_n7185, gm_n388, gm_n72, in_17, gm_n7184, gm_n662);
	or (gm_n7186, gm_n190, in_16, gm_n59, gm_n4917, gm_n227);
	nor (gm_n7187, gm_n58, gm_n72, in_20, gm_n7186);
	nor (gm_n7188, gm_n287, in_14, gm_n78, gm_n389, gm_n369);
	nand (gm_n7189, gm_n166, gm_n86, gm_n119, gm_n7188);
	nand (gm_n7190, gm_n72, gm_n85, in_19, gm_n916);
	nand (gm_n7191, gm_n233, gm_n73, gm_n59, gm_n571, gm_n142);
	nor (gm_n7192, gm_n496, gm_n72, in_20, gm_n7191);
	and (gm_n7193, gm_n104, in_21, in_17, gm_n1313, gm_n174);
	nor (gm_n7194, gm_n430, gm_n76, gm_n62, gm_n1583, gm_n257);
	nand (gm_n7195, gm_n327, gm_n72, in_17, gm_n7194, gm_n339);
	nor (gm_n7196, gm_n227, in_16, in_12, gm_n278, gm_n297);
	nand (gm_n7197, gm_n113, gm_n72, gm_n85, gm_n7196);
	and (gm_n7198, gm_n436, gm_n129, in_18, gm_n1473);
	or (gm_n7199, gm_n90, in_10, gm_n62, gm_n207, gm_n203);
	nor (gm_n7200, gm_n244, gm_n167, gm_n119, gm_n7199);
	and (gm_n7201, in_14, gm_n78, gm_n62, gm_n946, gm_n334);
	nand (gm_n7202, gm_n348, gm_n200, in_18, gm_n7201);
	nor (gm_n7203, gm_n257, gm_n76, in_9, gm_n2474, gm_n328);
	nand (gm_n7204, gm_n373, in_21, gm_n55, gm_n7203);
	or (gm_n7205, gm_n293, gm_n158, in_15, gm_n3929, gm_n760);
	nor (gm_n7206, gm_n72, gm_n85, in_19, gm_n7205);
	nand (gm_n7207, gm_n106, in_13, in_9, gm_n126, gm_n125);
	nor (gm_n7208, gm_n441, gm_n72, gm_n55, gm_n7207, gm_n375);
	nor (gm_n7209, gm_n90, in_10, in_9, gm_n2244, gm_n92);
	nand (gm_n7210, gm_n131, gm_n129, in_18, gm_n7209);
	nand (gm_n7211, gm_n72, in_20, gm_n56, gm_n6892, gm_n394);
	or (gm_n7212, gm_n406, gm_n76, gm_n62, gm_n743, gm_n502);
	nor (gm_n7213, gm_n441, gm_n72, gm_n55, gm_n7212, gm_n256);
	or (gm_n7214, gm_n431, in_13, gm_n62, gm_n621, gm_n463);
	nor (gm_n7215, gm_n479, in_21, gm_n55, gm_n7214, gm_n256);
	nand (gm_n7216, gm_n436, gm_n164, gm_n119, gm_n6882);
	nor (gm_n7217, gm_n596, gm_n76, gm_n62, gm_n442, gm_n345);
	nand (gm_n7218, gm_n120, in_21, gm_n55, gm_n7217, gm_n523);
	or (gm_n7219, gm_n667, gm_n76, in_9, gm_n359, gm_n257);
	nor (gm_n7220, gm_n183, in_21, gm_n55, gm_n7219, gm_n662);
	or (gm_n7221, gm_n461, in_13, in_9, gm_n988, gm_n344);
	nor (gm_n7222, gm_n184, in_21, in_17, gm_n7221, gm_n312);
	nor (gm_n7223, gm_n193, gm_n297, gm_n60, gm_n562, gm_n293);
	nand (gm_n7224, in_21, in_20, gm_n56, gm_n7223);
	nor (gm_n7225, gm_n257, in_13, in_9, gm_n988, gm_n443);
	nand (gm_n7226, gm_n254, in_21, gm_n55, gm_n7225, gm_n595);
	nand (gm_n7227, gm_n222, in_16, in_12, gm_n2547, gm_n275);
	nor (gm_n7228, gm_n58, in_21, gm_n85, gm_n7227);
	nor (gm_n7229, gm_n159, gm_n60, gm_n63, gm_n2690, gm_n605);
	nand (gm_n7230, in_21, in_20, gm_n56, gm_n7229, gm_n1101);
	and (gm_n7231, in_14, in_10, gm_n62, gm_n1524, gm_n1011);
	nand (gm_n7232, gm_n245, gm_n199, in_18, gm_n7231);
	nor (gm_n7233, gm_n609, in_13, in_9, gm_n597, gm_n442);
	nand (gm_n7234, gm_n255, in_21, gm_n55, gm_n7233, gm_n373);
	nand (gm_n7235, gm_n7234, gm_n7232, gm_n7230);
	nand (gm_n7236, gm_n214, in_16, in_12, gm_n2547, gm_n275);
	nor (gm_n7237, gm_n496, gm_n72, in_20, gm_n7236);
	or (gm_n7238, gm_n807, in_10, in_9, gm_n503, gm_n463);
	nor (gm_n7239, gm_n211, gm_n119, gm_n90, gm_n7238, gm_n167);
	or (gm_n7240, gm_n190, in_16, in_12, gm_n1006, gm_n152);
	nor (gm_n7241, gm_n262, gm_n72, in_20, gm_n7240);
	nor (gm_n7242, gm_n7237, gm_n7235, gm_n7228, gm_n7241, gm_n7239);
	nor (gm_n7243, gm_n103, gm_n72, in_17, gm_n3300, gm_n121);
	or (gm_n7244, gm_n609, in_13, in_9, gm_n462, gm_n461);
	nor (gm_n7245, gm_n121, in_21, gm_n55, gm_n7244, gm_n479);
	or (gm_n7246, gm_n667, gm_n76, in_9, gm_n406, gm_n796);
	nor (gm_n7247, gm_n103, in_21, in_17, gm_n7246, gm_n105);
	nor (gm_n7248, gm_n7247, gm_n7245, gm_n7243);
	or (gm_n7249, gm_n596, gm_n76, in_9, gm_n621, gm_n442);
	nor (gm_n7250, gm_n620, in_21, gm_n55, gm_n7249, gm_n328);
	or (gm_n7251, gm_n662, gm_n76, in_9, gm_n1481, gm_n442);
	nor (gm_n7252, gm_n441, gm_n72, in_17, gm_n7251);
	nand (gm_n7253, gm_n187, in_13, in_9, gm_n1049, gm_n402);
	nor (gm_n7254, gm_n312, gm_n72, in_17, gm_n7253, gm_n662);
	nor (gm_n7255, gm_n7254, gm_n7252, gm_n7250);
	nand (gm_n7256, gm_n7242, gm_n7226, gm_n7224, gm_n7255, gm_n7248);
	and (gm_n7257, gm_n79, gm_n73, in_12, gm_n636, gm_n733);
	nand (gm_n7258, gm_n138, gm_n72, in_20, gm_n7257);
	nor (gm_n7259, gm_n297, gm_n74, gm_n60, gm_n4614, gm_n159);
	nand (gm_n7260, in_21, in_20, gm_n56, gm_n7259);
	and (gm_n7261, gm_n281, gm_n214, in_15, gm_n3886, gm_n869);
	nand (gm_n7262, in_21, gm_n85, in_19, gm_n7261);
	nand (gm_n7263, gm_n7262, gm_n7260, gm_n7258);
	nor (gm_n7264, gm_n227, gm_n73, in_12, gm_n1203, gm_n158);
	nand (gm_n7265, gm_n113, in_21, gm_n85, gm_n7264);
	and (gm_n7266, gm_n713, in_14, gm_n78, gm_n793, gm_n1345);
	nand (gm_n7267, gm_n436, gm_n243, gm_n119, gm_n7266);
	nor (gm_n7268, gm_n213, gm_n73, gm_n59, gm_n1671, gm_n220);
	nand (gm_n7269, gm_n57, gm_n72, in_20, gm_n7268);
	nand (gm_n7270, gm_n7269, gm_n7267, gm_n7265);
	nor (gm_n7271, gm_n7256, gm_n7222, gm_n7220, gm_n7270, gm_n7263);
	nand (gm_n7272, gm_n61, gm_n73, gm_n59, gm_n2283, gm_n264);
	nor (gm_n7273, gm_n262, in_21, in_20, gm_n7272);
	or (gm_n7274, gm_n293, gm_n213, gm_n60, gm_n1052, gm_n643);
	nor (gm_n7275, in_21, in_20, gm_n56, gm_n7274);
	nor (gm_n7276, gm_n441, in_21, in_17, gm_n6195, gm_n313);
	nor (gm_n7277, gm_n7276, gm_n7275, gm_n7273);
	or (gm_n7278, gm_n480, in_13, gm_n62, gm_n502, gm_n481);
	nor (gm_n7279, gm_n184, gm_n72, in_17, gm_n7278, gm_n374);
	or (gm_n7280, gm_n257, gm_n76, in_9, gm_n1132, gm_n463);
	nor (gm_n7281, gm_n103, in_21, in_17, gm_n7280, gm_n313);
	nand (gm_n7282, gm_n579, in_13, in_9, gm_n341, gm_n316);
	nor (gm_n7283, gm_n184, in_21, in_17, gm_n7282, gm_n620);
	nor (gm_n7284, gm_n7283, gm_n7281, gm_n7279);
	nand (gm_n7285, gm_n7271, gm_n7218, gm_n7216, gm_n7284, gm_n7277);
	nor (gm_n7286, gm_n667, gm_n76, gm_n62, gm_n462, gm_n480);
	nand (gm_n7287, gm_n254, gm_n72, in_17, gm_n7286, gm_n255);
	nand (gm_n7288, gm_n102, in_21, gm_n55, gm_n4246, gm_n595);
	nor (gm_n7289, gm_n148, in_14, gm_n78, gm_n350, gm_n207);
	nand (gm_n7290, gm_n164, gm_n131, in_18, gm_n7289);
	nand (gm_n7291, gm_n7290, gm_n7288, gm_n7287);
	and (gm_n7292, gm_n76, in_9, in_8, gm_n1496, gm_n402);
	nand (gm_n7293, gm_n327, in_21, gm_n55, gm_n7292, gm_n1076);
	nor (gm_n7294, gm_n190, in_16, in_12, gm_n765, gm_n319);
	nand (gm_n7295, gm_n697, gm_n72, gm_n85, gm_n7294);
	nand (gm_n7296, gm_n348, gm_n323, in_18, gm_n1676);
	nand (gm_n7297, gm_n7296, gm_n7295, gm_n7293);
	nor (gm_n7298, gm_n7285, gm_n7215, gm_n7213, gm_n7297, gm_n7291);
	or (gm_n7299, gm_n461, gm_n76, in_9, gm_n1583, gm_n463);
	nor (gm_n7300, gm_n103, gm_n72, gm_n55, gm_n7299, gm_n313);
	nand (gm_n7301, in_14, gm_n78, gm_n62, gm_n1012, gm_n1158);
	nor (gm_n7302, gm_n531, gm_n1989, gm_n119, gm_n7301);
	or (gm_n7303, gm_n430, gm_n76, in_9, gm_n988, gm_n406);
	nor (gm_n7304, gm_n312, gm_n72, in_17, gm_n7303, gm_n328);
	nor (gm_n7305, gm_n7304, gm_n7302, gm_n7300);
	nor (gm_n7306, gm_n103, in_21, gm_n55, gm_n3300, gm_n105);
	nand (gm_n7307, gm_n1101, gm_n56, in_15, gm_n6703, gm_n545);
	nor (gm_n7308, gm_n7307, in_21, gm_n85);
	nand (gm_n7309, gm_n600, in_14, gm_n78, gm_n333, gm_n995);
	nor (gm_n7310, gm_n368, gm_n89, gm_n119, gm_n7309);
	nor (gm_n7311, gm_n7310, gm_n7308, gm_n7306);
	nand (gm_n7312, gm_n7298, gm_n7211, gm_n7210, gm_n7311, gm_n7305);
	nor (gm_n7313, gm_n643, gm_n60, gm_n63, gm_n981, gm_n980);
	nand (gm_n7314, gm_n72, gm_n85, gm_n56, gm_n7313, gm_n394);
	and (gm_n7315, gm_n379, gm_n143, in_15, gm_n2276, gm_n192);
	nand (gm_n7316, in_21, gm_n85, gm_n56, gm_n7315);
	and (gm_n7317, gm_n125, gm_n76, in_9, gm_n316, gm_n579);
	nand (gm_n7318, gm_n174, gm_n72, in_17, gm_n7317, gm_n1076);
	nand (gm_n7319, gm_n7318, gm_n7316, gm_n7314);
	nor (gm_n7320, gm_n406, gm_n76, in_9, gm_n597, gm_n596);
	nand (gm_n7321, gm_n174, in_21, gm_n55, gm_n7320, gm_n255);
	nor (gm_n7322, gm_n92, in_10, gm_n62, gm_n462, gm_n344);
	nand (gm_n7323, gm_n166, gm_n119, gm_n90, gm_n7322, gm_n243);
	nor (gm_n7324, gm_n447, gm_n155, gm_n60, gm_n2333, gm_n643);
	nand (gm_n7325, gm_n72, in_20, gm_n56, gm_n7324);
	nand (gm_n7326, gm_n7325, gm_n7323, gm_n7321);
	nor (gm_n7327, gm_n7312, gm_n7208, gm_n7206, gm_n7326, gm_n7319);
	nor (gm_n7328, gm_n388, gm_n72, gm_n55, gm_n4491, gm_n328);
	or (gm_n7329, gm_n369, gm_n240, in_14, gm_n761);
	nor (gm_n7330, gm_n437, gm_n87, in_18, gm_n7329);
	nand (gm_n7331, gm_n123, gm_n76, in_9, gm_n316, gm_n186);
	nor (gm_n7332, gm_n183, in_21, gm_n55, gm_n7331, gm_n375);
	nor (gm_n7333, gm_n7332, gm_n7330, gm_n7328);
	or (gm_n7334, gm_n1331, gm_n158, gm_n60, gm_n2931, gm_n290);
	nor (gm_n7335, in_21, in_20, in_19, gm_n7334);
	nand (gm_n7336, gm_n126, gm_n76, gm_n62, gm_n402, gm_n341);
	nor (gm_n7337, gm_n103, in_21, gm_n55, gm_n7336, gm_n662);
	nand (gm_n7338, gm_n233, in_16, in_12, gm_n1179, gm_n571);
	nor (gm_n7339, gm_n384, gm_n72, in_20, gm_n7338);
	nor (gm_n7340, gm_n7339, gm_n7337, gm_n7335);
	nand (gm_n7341, gm_n7327, gm_n7204, gm_n7202, gm_n7340, gm_n7333);
	nor (gm_n7342, gm_n168, gm_n60, gm_n63, gm_n842, gm_n271);
	nand (gm_n7343, gm_n72, gm_n85, gm_n56, gm_n7342, gm_n448);
	and (gm_n7344, gm_n90, gm_n78, gm_n62, gm_n2605, gm_n1158);
	nand (gm_n7345, gm_n436, gm_n199, in_18, gm_n7344);
	nand (gm_n7346, gm_n255, gm_n72, in_17, gm_n804, gm_n327);
	nand (gm_n7347, gm_n7346, gm_n7345, gm_n7343);
	nor (gm_n7348, gm_n461, gm_n95, in_13, gm_n376, gm_n256);
	nand (gm_n7349, gm_n206, gm_n72, in_17, gm_n7348);
	and (gm_n7350, gm_n143, gm_n73, gm_n59, gm_n875, gm_n275);
	nand (gm_n7351, gm_n179, gm_n72, gm_n85, gm_n7350);
	nor (gm_n7352, gm_n155, gm_n73, gm_n59, gm_n1324, gm_n220);
	nand (gm_n7353, gm_n57, in_21, gm_n85, gm_n7352);
	nand (gm_n7354, gm_n7353, gm_n7351, gm_n7349);
	nor (gm_n7355, gm_n7341, gm_n7200, gm_n7198, gm_n7354, gm_n7347);
	or (gm_n7356, gm_n184, gm_n148, gm_n76, gm_n431, gm_n286);
	nor (gm_n7357, gm_n479, in_21, gm_n55, gm_n7356);
	nand (gm_n7358, gm_n125, in_13, gm_n62, gm_n185, gm_n126);
	nor (gm_n7359, gm_n441, in_21, gm_n55, gm_n7358, gm_n328);
	or (gm_n7360, gm_n227, gm_n73, gm_n59, gm_n1661, gm_n297);
	nor (gm_n7361, gm_n384, gm_n72, in_20, gm_n7360);
	nor (gm_n7362, gm_n7361, gm_n7359, gm_n7357);
	or (gm_n7363, gm_n461, gm_n99, gm_n76, gm_n438, gm_n256);
	nor (gm_n7364, gm_n620, in_21, gm_n55, gm_n7363);
	and (gm_n7365, gm_n254, in_21, in_17, gm_n693, gm_n595);
	or (gm_n7366, gm_n293, gm_n158, in_15, gm_n760, gm_n657);
	nor (gm_n7367, in_21, in_20, in_19, gm_n7366);
	nor (gm_n7368, gm_n7367, gm_n7365, gm_n7364);
	nand (gm_n7369, gm_n7355, gm_n7197, gm_n7195, gm_n7368, gm_n7362);
	nor (gm_n7370, gm_n259, gm_n90, gm_n78, gm_n491, gm_n369);
	nand (gm_n7371, gm_n367, gm_n166, gm_n119, gm_n7370);
	nand (gm_n7372, gm_n104, in_21, in_17, gm_n5463, gm_n327);
	nor (gm_n7373, gm_n431, in_13, gm_n62, gm_n503, gm_n596);
	nand (gm_n7374, gm_n523, in_21, in_17, gm_n7373, gm_n311);
	nand (gm_n7375, gm_n7374, gm_n7372, gm_n7371);
	nor (gm_n7376, gm_n158, gm_n73, gm_n59, gm_n4437, gm_n354);
	nand (gm_n7377, gm_n495, in_21, in_20, gm_n7376);
	nor (gm_n7378, gm_n480, in_13, in_9, gm_n743, gm_n502);
	nand (gm_n7379, gm_n104, in_21, gm_n55, gm_n7378, gm_n327);
	nor (gm_n7380, gm_n662, in_13, in_9, gm_n2823, gm_n442);
	nand (gm_n7381, gm_n102, in_21, in_17, gm_n7380);
	nand (gm_n7382, gm_n7381, gm_n7379, gm_n7377);
	nor (gm_n7383, gm_n7369, gm_n7193, gm_n7192, gm_n7382, gm_n7375);
	and (gm_n7384, gm_n120, in_21, in_17, gm_n5523, gm_n595);
	or (gm_n7385, gm_n313, in_13, in_9, gm_n3660, gm_n406);
	nor (gm_n7386, gm_n183, in_21, gm_n55, gm_n7385);
	nand (gm_n7387, in_14, in_10, gm_n62, gm_n2416, gm_n91);
	nor (gm_n7388, gm_n841, gm_n824, gm_n119, gm_n7387);
	nor (gm_n7389, gm_n7388, gm_n7386, gm_n7384);
	or (gm_n7390, gm_n358, gm_n76, gm_n62, gm_n1132, gm_n443);
	nor (gm_n7391, gm_n328, gm_n72, gm_n55, gm_n7390, gm_n374);
	or (gm_n7392, gm_n362, gm_n90, in_10, gm_n491, gm_n376);
	nor (gm_n7393, gm_n824, gm_n89, gm_n119, gm_n7392);
	or (gm_n7394, gm_n796, in_13, gm_n62, gm_n502, gm_n406);
	nor (gm_n7395, gm_n312, in_21, in_17, gm_n7394, gm_n313);
	nor (gm_n7396, gm_n7395, gm_n7393, gm_n7391);
	nand (gm_n7397, gm_n7383, gm_n7190, gm_n7189, gm_n7396, gm_n7389);
	nor (gm_n7398, gm_n609, gm_n76, gm_n62, gm_n481, gm_n480);
	nand (gm_n7399, gm_n104, gm_n72, gm_n55, gm_n7398, gm_n327);
	nor (gm_n7400, gm_n155, in_16, gm_n59, gm_n1906, gm_n276);
	nand (gm_n7401, gm_n57, gm_n72, in_20, gm_n7400);
	nor (gm_n7402, gm_n407, gm_n133, in_14, gm_n605);
	nand (gm_n7403, gm_n88, gm_n86, in_18, gm_n7402);
	nand (gm_n7404, gm_n7403, gm_n7401, gm_n7399);
	nor (gm_n7405, gm_n155, gm_n74, gm_n60, gm_n298, gm_n168);
	nand (gm_n7406, gm_n72, gm_n85, gm_n56, gm_n7405);
	and (gm_n7407, gm_n106, in_13, gm_n62, gm_n126, gm_n107);
	nand (gm_n7408, gm_n254, in_21, in_17, gm_n7407, gm_n405);
	or (gm_n7409, gm_n5886, gm_n368);
	nand (gm_n7410, gm_n7409, gm_n7408, gm_n7406);
	nor (gm_n7411, gm_n7397, gm_n7187, gm_n7185, gm_n7410, gm_n7404);
	or (gm_n7412, gm_n263, in_16, gm_n59, gm_n2357, gm_n276);
	nor (gm_n7413, gm_n496, in_21, gm_n85, gm_n7412);
	or (gm_n7414, gm_n406, in_13, in_9, gm_n502, gm_n432);
	nor (gm_n7415, gm_n121, gm_n72, gm_n55, gm_n7414, gm_n479);
	nor (gm_n7416, gm_n368, gm_n119, gm_n90, gm_n6982, gm_n437);
	nor (gm_n7417, gm_n7416, gm_n7415, gm_n7413);
	nand (gm_n7418, in_14, gm_n78, in_9, gm_n2916, gm_n334);
	nor (gm_n7419, gm_n244, gm_n167, in_18, gm_n7418);
	and (gm_n7420, gm_n595, gm_n72, in_17, gm_n6134, gm_n373);
	or (gm_n7421, gm_n406, gm_n76, in_9, gm_n503, gm_n344);
	nor (gm_n7422, gm_n103, in_21, gm_n55, gm_n7421, gm_n121);
	nor (gm_n7423, gm_n7422, gm_n7420, gm_n7419);
	nand (gm_n7424, gm_n7411, gm_n7183, gm_n7182, gm_n7423, gm_n7417);
	and (gm_n7425, gm_n91, gm_n88, gm_n90, gm_n1942, gm_n170);
	nand (gm_n7426, gm_n7425, gm_n86, gm_n119);
	nor (gm_n7427, gm_n480, in_13, in_9, gm_n502, gm_n481);
	nand (gm_n7428, gm_n122, gm_n72, in_17, gm_n7427, gm_n327);
	nor (gm_n7429, gm_n596, gm_n76, in_9, gm_n1583, gm_n442);
	nand (gm_n7430, gm_n174, in_21, gm_n55, gm_n7429, gm_n339);
	nand (gm_n7431, gm_n7430, gm_n7428, gm_n7426);
	nor (gm_n7432, gm_n297, gm_n73, in_12, gm_n1884, gm_n276);
	nand (gm_n7433, gm_n57, in_21, in_20, gm_n7432);
	nor (gm_n7434, gm_n114, in_16, gm_n59, gm_n695, gm_n190);
	nand (gm_n7435, gm_n697, in_21, gm_n85, gm_n7434);
	and (gm_n7436, gm_n264, in_16, in_12, gm_n2547, gm_n275);
	nand (gm_n7437, gm_n296, gm_n72, gm_n85, gm_n7436);
	nand (gm_n7438, gm_n7437, gm_n7435, gm_n7433);
	nor (gm_n7439, gm_n7424, gm_n7180, gm_n7178, gm_n7438, gm_n7431);
	or (gm_n7440, gm_n667, in_13, gm_n62, gm_n503, gm_n480);
	nor (gm_n7441, gm_n479, gm_n72, in_17, gm_n7440, gm_n256);
	nand (gm_n7442, gm_n484, gm_n75, in_15, gm_n615, gm_n264);
	nor (gm_n7443, gm_n72, gm_n85, gm_n56, gm_n7442);
	and (gm_n7444, gm_n72, in_20, in_19, gm_n1966, gm_n75);
	nor (gm_n7445, gm_n7444, gm_n7443, gm_n7441);
	or (gm_n7446, gm_n190, in_16, in_12, gm_n2730, gm_n152);
	nor (gm_n7447, gm_n781, in_21, in_20, gm_n7446);
	nand (gm_n7448, gm_n449, gm_n79, in_15, gm_n991);
	nor (gm_n7449, gm_n72, gm_n85, in_19, gm_n7448, gm_n191);
	nand (gm_n7450, gm_n423, gm_n233, in_15, gm_n545);
	nor (gm_n7451, gm_n72, gm_n85, in_19, gm_n7450, gm_n74);
	nor (gm_n7452, gm_n7451, gm_n7449, gm_n7447);
	nand (gm_n7453, gm_n7439, gm_n7176, gm_n7174, gm_n7452, gm_n7445);
	and (gm_n7454, gm_n264, gm_n73, in_12, gm_n612, gm_n571);
	nand (gm_n7455, gm_n495, gm_n72, in_20, gm_n7454);
	and (gm_n7456, gm_n91, gm_n90, gm_n78, gm_n793, gm_n2670);
	nand (gm_n7457, gm_n243, gm_n166, gm_n119, gm_n7456);
	and (gm_n7458, gm_n90, gm_n78, in_9, gm_n2646, gm_n624);
	nand (gm_n7459, gm_n323, gm_n164, in_18, gm_n7458);
	nand (gm_n7460, gm_n7459, gm_n7457, gm_n7455);
	nor (gm_n7461, gm_n158, in_16, in_12, gm_n320, gm_n385);
	nand (gm_n7462, gm_n113, in_21, gm_n85, gm_n7461);
	nor (gm_n7463, gm_n297, gm_n73, in_12, gm_n1906, gm_n385);
	nand (gm_n7464, gm_n138, gm_n72, gm_n85, gm_n7463);
	nor (gm_n7465, gm_n213, gm_n73, in_12, gm_n1923, gm_n385);
	nand (gm_n7466, gm_n179, in_21, gm_n85, gm_n7465);
	nand (gm_n7467, gm_n7466, gm_n7464, gm_n7462);
	nor (gm_n7468, gm_n7453, gm_n7172, gm_n7170, gm_n7467, gm_n7460);
	or (gm_n7469, gm_n213, gm_n73, gm_n59, gm_n1965, gm_n276);
	nor (gm_n7470, gm_n384, gm_n72, in_20, gm_n7469);
	or (gm_n7471, gm_n158, in_16, in_12, gm_n320, gm_n220);
	nor (gm_n7472, gm_n912, in_21, gm_n85, gm_n7471);
	or (gm_n7473, gm_n430, gm_n76, in_9, gm_n1132, gm_n431);
	nor (gm_n7474, gm_n479, gm_n72, gm_n55, gm_n7473, gm_n328);
	nor (gm_n7475, gm_n7474, gm_n7472, gm_n7470);
	nand (gm_n7476, gm_n233, in_16, gm_n59, gm_n1095, gm_n571);
	nor (gm_n7477, gm_n219, in_21, in_20, gm_n7476);
	or (gm_n7478, gm_n514, in_13, in_9, gm_n511, gm_n184);
	nor (gm_n7479, gm_n388, gm_n72, in_17, gm_n7478);
	nand (gm_n7480, gm_n185, in_13, gm_n62, gm_n471, gm_n339);
	nor (gm_n7481, gm_n620, in_21, gm_n55, gm_n7480);
	nor (gm_n7482, gm_n7481, gm_n7479, gm_n7477);
	nand (gm_n7483, gm_n7468, gm_n7168, gm_n7166, gm_n7482, gm_n7475);
	nor (gm_n7484, gm_n92, gm_n90, gm_n78, gm_n248, gm_n95);
	nand (gm_n7485, gm_n243, gm_n806, gm_n119, gm_n7484);
	and (gm_n7486, gm_n268, gm_n214, in_15, gm_n1531, gm_n545);
	nand (gm_n7487, in_21, gm_n85, gm_n56, gm_n7486);
	nor (gm_n7488, gm_n99, gm_n90, in_10, gm_n369, gm_n148);
	nand (gm_n7489, gm_n131, gm_n129, gm_n119, gm_n7488);
	nand (gm_n7490, gm_n7489, gm_n7487, gm_n7485);
	nor (gm_n7491, gm_n256, gm_n76, gm_n62, gm_n3315, gm_n480);
	nand (gm_n7492, gm_n120, in_21, in_17, gm_n7491);
	nor (gm_n7493, gm_n818, gm_n76, in_9, gm_n667, gm_n358);
	nand (gm_n7494, gm_n122, in_21, gm_n55, gm_n7493, gm_n373);
	nand (gm_n7495, gm_n102, in_21, gm_n55, gm_n4177, gm_n1076);
	nand (gm_n7496, gm_n7495, gm_n7494, gm_n7492);
	nor (out_21, gm_n7490, gm_n7483, gm_n7164, gm_n7496);
endmodule
