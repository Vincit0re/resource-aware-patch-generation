module top ( g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 , g98 , g99 , g100 , g101 , g102 , g103 , g104 , g105 , g106 , g107 , g108 , g109 , g110 , g111 , g112 , g113 , g114 , g115 , g116 , g117 , g118 , g119 , g120 , g121 , g122 , g123 , g124 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g136 , g137 , g138 , g139 , g140 , g141 , g142 , g143 , g144 , g145 , g146 , g147 , g148 , g149 , g150 , g151 , g152 , g153 , g154 , g155 , g156 , g157 , g158 , g159 , g160 , g161 , g162 , g163 , g164 , g165 , g166 , g167 , g168 , g169 , g170 , g171 , g172 , g173 , g174 , g175 , g176 , g177 , g178 , g179 , g180 , g181 , g182 , g183 , g184 , g185 , g186 , g187 , g188 , g189 , g190 , g191 , g192 , g193 , g194 , g195 , g196 , g197 , g198 , g199 , g200 , g201 , g202 , g203 , g204 , g205 , g206 , g207 , g208 , g209 , g210 , g211 , g212 , g213 , g214 , g215 , g216 , g217 , g218 , g219 , g220 );
input g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 , g98 , g99 , g100 , g101 , g102 , g103 , g104 , g105 , g106 , g107 , g108 , g109 , g110 , g111 , g112 , g113 , g114 , g115 , g116 , g117 , g118 , g119 , g120 , g121 , g122 , g123 , g124 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g136 , g137 , g138 , g139 , g140 , g141 , g142 , g143 , g144 , g145 , g146 , g147 , g148 , g149 , g150 , g151 , g152 , g153 , g154 , g155 , g156 ;
output g157 , g158 , g159 , g160 , g161 , g162 , g163 , g164 , g165 , g166 , g167 , g168 , g169 , g170 , g171 , g172 , g173 , g174 , g175 , g176 , g177 , g178 , g179 , g180 , g181 , g182 , g183 , g184 , g185 , g186 , g187 , g188 , g189 , g190 , g191 , g192 , g193 , g194 , g195 , g196 , g197 , g198 , g199 , g200 , g201 , g202 , g203 , g204 , g205 , g206 , g207 , g208 , g209 , g210 , g211 , g212 , g213 , g214 , g215 , g216 , g217 , g218 , g219 , g220 ;

wire g4669 , g4670 , g4671 , g4672 , g4673 , g4674 , g4675 , g4676 , g4677 , 
     g4678 , g4679 , g4680 , g4681 , g4682 , g4683 , g4684 , g4685 , g4686 , g4687 , 
     g4688 , g4689 , g4690 , g4691 , g4692 , g4693 , g4694 , g4695 , g4696 , g4697 , 
     g4698 , g4699 , g4700 , g4701 , g4702 , g4703 , g4704 , g4705 , g4706 , g4707 , 
     g4708 , g4709 , g4710 , g4711 , g4712 , g4713 , g4714 , g4715 , g4716 , g4717 , 
     g4718 , g4719 , g4720 , g4721 , g4722 , g4723 , g4724 , g4725 , g4726 , g4727 , 
     g4728 , g4729 , g4730 , g4731 , g4732 , g4733 , g4734 , g4735 , g4736 , g4737 , 
     g4738 , g4739 , g4740 , g4741 , g4742 , g4743 , g4744 , g4745 , g4746 , g4747 , 
     g4748 , g4749 , g4750 , g4751 , g4752 , g4753 , g4754 , g4755 , g4756 , g4757 , 
     g4758 , g4759 , g4760 , g4761 , g4762 , g4763 , g4764 , g4765 , g4766 , g4767 , 
     g4768 , g4769 , g4770 , g4771 , g4772 , g4773 , g4774 , g4775 , g4776 , g4777 , 
     g4778 , g4779 , g4780 , g4781 , g4782 , g4783 , g4784 , g4785 , g4786 , g4787 , 
     g4788 , g4789 , g4790 , g4791 , g4792 , g4793 , g4794 , g4795 , g4796 , g4797 , 
     g4798 , g4799 , g4800 , g4801 , g4802 , g4803 , g4804 , g4805 , g4806 , g4807 , 
     g4808 , g4809 , g4810 , g4811 , g4812 , g4813 , g4814 , g4815 , g4816 , g4817 , 
     g4818 , g4819 , g4820 , g4821 , g4822 , g4823 , g4824 , g4825 , g4826 , g4827 , 
     g4828 , g4829 , g4830 , g4831 , g4832 , g4833 , g4834 , g4835 , g4836 , g4837 , 
     g4838 , g4839 , g4840 , g4841 , g4842 , g4843 , g4844 , g4845 , g4846 , g4847 , 
     g4848 , g4849 , g4850 , g4851 , g4852 , g4853 , g4854 , g4855 , g4856 , g4857 , 
     g4858 , g4859 , g4860 , g4861 , g4862 , g4863 , g4864 , g4865 , g4866 , g4867 , 
     g4868 , g4869 , g4870 , g4871 , g4872 , g4873 , g4874 , g4875 , g4876 , g4877 , 
     g4878 , g4879 , g4880 , g4881 , g4882 , g4883 , g4884 , g4885 , g4886 , g4887 , 
     g4888 , g4889 , g442 , g443 , g444 , g445 , g446 , g447 , g448 , g449 , 
     g450 , g451 , g452 , g453 , g454 , g455 , g456 , g457 , g458 , g459 , 
     g460 , g461 , g462 , g463 , g464 , g465 , g466 , g467 , g468 , g469 , 
     g470 , g471 , g472 , g473 , g474 , g475 , g476 , g477 , g478 , g479 , 
     g480 , g481 , g482 , g483 , g484 , g485 , g486 , g487 , g488 , g489 , 
     g490 , g491 , g492 , g493 , g494 , g495 , g496 , g497 , g498 , g499 , 
     g500 , g501 , g502 , g503 , g504 , g505 , g506 , g507 , g508 , g509 , 
     g510 , g511 , g512 , g513 , g514 , g515 , g516 , g517 , g518 , g519 , 
     g520 , g521 , g522 , g523 , g524 , g525 , g526 , g527 , g528 , g529 , 
     g530 , g531 , g532 , g533 , g534 , g535 , g536 , g537 , g538 , g539 , 
     g540 , g541 , g542 , g543 , g544 , g545 , g546 , g547 , g548 , g549 , 
     g550 , g551 , g552 , g553 , g554 , g555 , g556 , g557 , g558 , g559 , 
     g560 , g561 , g562 , g563 , g564 , g565 , g566 , g567 , g568 , g569 , 
     g570 , g571 , g572 , g573 , g574 , g575 , g576 , g577 , g578 , g579 , 
     g580 , g581 , g582 , g583 , g584 , g585 , g586 , g587 , g588 , g589 , 
     g590 , g591 , g592 , g593 , g594 , g595 , g596 , g597 , g598 , g599 , 
     g600 , g601 , g602 , g603 , g604 , g605 , g606 , g607 , g608 , g609 , 
     g610 , g611 , g612 , g613 , g614 , g615 , g616 , g617 , g618 , g619 , 
     g620 , g621 , g622 , g623 , g624 , g625 , g626 , g627 , g628 , g629 , 
     g630 , g631 , g632 , g633 , g634 , g635 , g636 , g637 , g638 , g639 , 
     g640 , g641 , g642 , g643 , g644 , g645 , g646 , g647 , g648 , g649 , 
     g650 , g651 , g652 , g653 , g654 , g655 , g656 , g657 , g658 , g659 , 
     g660 , g661 , g662 , g663 , g664 , g665 , g666 , g667 , g668 , g669 , 
     g670 , g671 , g672 , g673 , g674 , g675 , g676 , g677 , g678 , g679 , 
     g680 , g681 , g682 , g683 , g684 , g685 , g686 , g687 , g688 , g689 , 
     g690 , g691 , g692 , g693 , g694 , g695 , g696 , g697 , g698 , g699 , 
     g700 , g701 , g702 , g703 , g704 , g705 , g706 , g707 , g708 , g709 , 
     g710 , g711 , g712 , g713 , g714 , g715 , g716 , g717 , g718 , g719 , 
     g720 , g721 , g722 , g723 , g724 , g725 , g726 , g727 , g728 , g729 , 
     g730 , g731 , g732 , g733 , g734 , g735 , g736 , g737 , g738 , g739 , 
     g740 , g741 , g742 , g743 , g744 , g745 , g746 , g747 , g748 , g749 , 
     g750 , g751 , g752 , g753 , g754 , g755 , g756 , g757 , g758 , g759 , 
     g760 , g761 , g762 , g763 , g764 , g765 , g766 , g767 , g768 , g769 , 
     g770 , g771 , g772 , g773 , g774 , g775 , g776 , g777 , g778 , g779 , 
     g780 , g781 , g782 , g783 , g784 , g785 , g786 , g787 , g788 , g789 , 
     g790 , g791 , g792 , g793 , g794 , g795 , g796 , g797 , g798 , g799 , 
     g800 , g801 , g802 , g803 , g804 , g805 , g806 , g807 , g808 , g809 , 
     g810 , g811 , g812 , g813 , g814 , g815 , g816 , g817 , g818 , g819 , 
     g820 , g821 , g822 , g823 , g824 , g825 , g826 , g827 , g828 , g829 , 
     g830 , g831 , g832 , g833 , g834 , g835 , g836 , g837 , g838 , g839 , 
     g840 , g841 , g842 , g843 , g844 , g845 , g846 , g847 , g848 , g849 , 
     g850 , g851 , g852 , g853 , g854 , g855 , g856 , g857 , g858 , g859 , 
     g860 , g861 , g862 , g863 , g864 , g865 , g866 , g867 , g868 , g869 , 
     g870 , g871 , g872 , g873 , g874 , g875 , g876 , g877 , g878 , g879 , 
     g880 , g881 , g882 , g883 , g884 , g885 , g886 , g887 , g888 , g889 , 
     g890 , g891 , g892 , g893 , g894 , g895 , g896 , g897 , g898 , g899 , 
     g900 , g901 , g902 , g903 , g904 , g905 , g906 , g907 , g908 , g909 , 
     g910 , g911 , g912 , g913 , g914 , g915 , g916 , g917 , g918 , g919 , 
     g920 , g921 , g922 , g923 , g924 , g925 , g926 , g927 , g928 , g929 , 
     g930 , g931 , g932 , g933 , g934 , g935 , g936 , g937 , g938 , g939 , 
     g940 , g941 , g942 , g943 , g944 , g945 , g946 , g947 , g948 , g949 , 
     g950 , g951 , g952 , g953 , g954 , g955 , g956 , g957 , g958 , g959 , 
     g960 , g961 , g962 , g963 , g964 , g965 , g966 , g967 , g968 , g969 , 
     g970 , g971 , g972 , g973 , g974 , g975 , g976 , g977 , g978 , g979 , 
     g980 , g981 , g982 , g983 , g984 , g985 , g986 , g987 , g988 , g989 , 
     g990 , g991 , g992 , g993 , g994 , g995 , g996 , g997 , g998 , g999 , 
     g1000 , g1001 , g1002 , g1003 , g1004 , g1005 , g1006 , g1007 , g1008 , g1009 , 
     g1010 , g1011 , g1012 , g1013 , g1014 , g1015 , g1016 , g1017 , g1018 , g1019 , 
     g1020 , g1021 , g1022 , g1023 , g1024 , g1025 , g1026 , g1027 , g1028 , g1029 , 
     g1030 , g1031 , g1032 , g1033 , g1034 , g1035 , g1036 , g1037 , g1038 , g1039 , 
     g1040 , g1041 , g1042 , g1043 , g1044 , g1045 , g1046 , g1047 , g1048 , g1049 , 
     g1050 , g1051 , g1052 , g1053 , g1054 , g1055 , g1056 , g1057 , g1058 , g1059 , 
     g1060 , g1061 , g1062 , g1063 , g1064 , g1065 , g1066 , g1067 , g1068 , g1069 , 
     g1070 , g1071 , g1072 , g1073 , g1074 , g1075 , g1076 , g1077 , g1078 , g1079 , 
     g1080 , g1081 , g1082 , g1083 , g1084 , g1085 , g1086 , g1087 , g1088 , g1089 , 
     g1090 , g1091 , g1092 , g1093 , g1094 , g1095 , g1096 , g1097 , g1098 , g1099 , 
     g1100 , g1101 , g1102 , g1103 , g1104 , g1105 , g1106 , g1107 , g1108 , g1109 , 
     g1110 , g1111 , g1112 , g1113 , g1114 , g1115 , g1116 , g1117 , g1118 , g1119 , 
     g1120 , g1121 , g1122 , g1123 , g1124 , g1125 , g1126 , g1127 , g1128 , g1129 , 
     g1130 , g1131 , g1132 , g1133 , g1134 , g1135 , g1136 , g1137 , g1138 , g1139 , 
     g1140 , g1141 , g1142 , g1143 , g1144 , g1145 , g1146 , g1147 , g1148 , g1149 , 
     g1150 , g1151 , g1152 , g1153 , g1154 , g1155 , g1156 , g1157 , g1158 , g1159 , 
     g1160 , g1161 , g1162 , g1163 , g1164 , g1165 , g1166 , g1167 , g1168 , g1169 , 
     g1170 , g1171 , g1172 , g1173 , g1174 , g1175 , g1176 , g1177 , g1178 , g1179 , 
     g1180 , g1181 , g1182 , g1183 , g1184 , g1185 , g1186 , g1187 , g1188 , g1189 , 
     g1190 , g1191 , g1192 , g1193 , g1194 , g1195 , g1196 , g1197 , g1198 , g1199 , 
     g1200 , g1201 , g1202 , g1203 , g1204 , g1205 , g1206 , g1207 , g1208 , g1209 , 
     g1210 , g1211 , g1212 , g1213 , g1214 , g1215 , g1216 , g1217 , g1218 , g1219 , 
     g1220 , g1221 , g1222 , g1223 , g1224 , g1225 , g1226 , g1227 , g1228 , g1229 , 
     g1230 , g1231 , g1232 , g1233 , g1234 , g1235 , g1236 , g1237 , g1238 , g1239 , 
     g1240 , g1241 , g1242 , g1243 , g1244 , g1245 , g1246 , g1247 , g1248 , g1249 , 
     g1250 , g1251 , g1252 , g1253 , g1254 , g1255 , g1256 , g1257 , g1258 , g1259 , 
     g1260 , g1261 , g1262 , g1263 , g1264 , g1265 , g1266 , g1267 , g1268 , g1269 , 
     g1270 , g1271 , g1272 , g1273 , g1274 , g1275 , g1276 , g1277 , g1278 , g1279 , 
     g1280 , g1281 , g1282 , g1283 , g1284 , g1285 , g1286 , g1287 , g1288 , g1289 , 
     g1290 , g1291 , g1292 , g1293 , g1294 , g1295 , g1296 , g1297 , g1298 , g1299 , 
     g1300 , g1301 , g1302 , g1303 , g1304 , g1305 , g1306 , g1307 , g1308 , g1309 , 
     g1310 , g1311 , g1312 , g1313 , g1314 , g1315 , g1316 , g1317 , g1318 , g1319 , 
     g1320 , g1321 , g1322 , g1323 , g1324 , g1325 , g1326 , g1327 , g1328 , g1329 , 
     g1330 , g1331 , g1332 , g1333 , g1334 , g1335 , g1336 , g1337 , g1338 , g1339 , 
     g1340 , g1341 , g1342 , g1343 , g1344 , g1345 , g1346 , g1347 , g1348 , g1349 , 
     g1350 , g1351 , g1352 , g1353 , g1354 , g1355 , g1356 , g1357 , g1358 , g1359 , 
     g1360 , g1361 , g1362 , g1363 , g1364 , g1365 , g1366 , g1367 , g1368 , g1369 , 
     g1370 , g1371 , g1372 , g1373 , g1374 , g1375 , g1376 , g1377 ;
buf ( g4669 , g0 );
buf ( g4670 , g1 );
buf ( g4671 , g2 );
buf ( g4672 , g3 );
buf ( g4673 , g4 );
buf ( g4674 , g5 );
buf ( g4675 , g6 );
buf ( g4676 , g7 );
buf ( g4677 , g8 );
buf ( g4678 , g9 );
buf ( g4679 , g10 );
buf ( g4680 , g11 );
buf ( g4681 , g12 );
buf ( g4682 , g13 );
buf ( g4683 , g14 );
buf ( g4684 , g15 );
buf ( g4685 , g16 );
buf ( g4686 , g17 );
buf ( g4687 , g18 );
buf ( g4688 , g19 );
buf ( g4689 , g20 );
buf ( g4690 , g21 );
buf ( g4691 , g22 );
buf ( g4692 , g23 );
buf ( g4693 , g24 );
buf ( g4694 , g25 );
buf ( g4695 , g26 );
buf ( g4696 , g27 );
buf ( g4697 , g28 );
buf ( g4698 , g29 );
buf ( g4699 , g30 );
buf ( g4700 , g31 );
buf ( g4701 , g32 );
buf ( g4702 , g33 );
buf ( g4703 , g34 );
buf ( g4704 , g35 );
buf ( g4705 , g36 );
buf ( g4706 , g37 );
buf ( g4707 , g38 );
buf ( g4708 , g39 );
buf ( g4709 , g40 );
buf ( g4710 , g41 );
buf ( g4711 , g42 );
buf ( g4712 , g43 );
buf ( g4713 , g44 );
buf ( g4714 , g45 );
buf ( g4715 , g46 );
buf ( g4716 , g47 );
buf ( g4717 , g48 );
buf ( g4718 , g49 );
buf ( g4719 , g50 );
buf ( g4720 , g51 );
buf ( g4721 , g52 );
buf ( g4722 , g53 );
buf ( g4723 , g54 );
buf ( g4724 , g55 );
buf ( g4725 , g56 );
buf ( g4726 , g57 );
buf ( g4727 , g58 );
buf ( g4728 , g59 );
buf ( g4729 , g60 );
buf ( g4730 , g61 );
buf ( g4731 , g62 );
buf ( g4732 , g63 );
buf ( g4733 , g64 );
buf ( g4734 , g65 );
buf ( g4735 , g66 );
buf ( g4736 , g67 );
buf ( g4737 , g68 );
buf ( g4738 , g69 );
buf ( g4739 , g70 );
buf ( g4740 , g71 );
buf ( g4741 , g72 );
buf ( g4742 , g73 );
buf ( g4743 , g74 );
buf ( g4744 , g75 );
buf ( g4745 , g76 );
buf ( g4746 , g77 );
buf ( g4747 , g78 );
buf ( g4748 , g79 );
buf ( g4749 , g80 );
buf ( g4750 , g81 );
buf ( g4751 , g82 );
buf ( g4752 , g83 );
buf ( g4753 , g84 );
buf ( g4754 , g85 );
buf ( g4755 , g86 );
buf ( g4756 , g87 );
buf ( g4757 , g88 );
buf ( g4758 , g89 );
buf ( g4759 , g90 );
buf ( g4760 , g91 );
buf ( g4761 , g92 );
buf ( g4762 , g93 );
buf ( g4763 , g94 );
buf ( g4764 , g95 );
buf ( g4765 , g96 );
buf ( g4766 , g97 );
buf ( g4767 , g98 );
buf ( g4768 , g99 );
buf ( g4769 , g100 );
buf ( g4770 , g101 );
buf ( g4771 , g102 );
buf ( g4772 , g103 );
buf ( g4773 , g104 );
buf ( g4774 , g105 );
buf ( g4775 , g106 );
buf ( g4776 , g107 );
buf ( g4777 , g108 );
buf ( g4778 , g109 );
buf ( g4779 , g110 );
buf ( g4780 , g111 );
buf ( g4781 , g112 );
buf ( g4782 , g113 );
buf ( g4783 , g114 );
buf ( g4784 , g115 );
buf ( g4785 , g116 );
buf ( g4786 , g117 );
buf ( g4787 , g118 );
buf ( g4788 , g119 );
buf ( g4789 , g120 );
buf ( g4790 , g121 );
buf ( g4791 , g122 );
buf ( g4792 , g123 );
buf ( g4793 , g124 );
buf ( g4794 , g125 );
buf ( g4795 , g126 );
buf ( g4796 , g127 );
buf ( g4797 , g128 );
buf ( g4798 , g129 );
buf ( g4799 , g130 );
buf ( g4800 , g131 );
buf ( g4801 , g132 );
buf ( g4802 , g133 );
buf ( g4803 , g134 );
buf ( g4804 , g135 );
buf ( g4805 , g136 );
buf ( g4806 , g137 );
buf ( g4807 , g138 );
buf ( g4808 , g139 );
buf ( g4809 , g140 );
buf ( g4810 , g141 );
buf ( g4811 , g142 );
buf ( g4812 , g143 );
buf ( g4813 , g144 );
buf ( g4814 , g145 );
buf ( g4815 , g146 );
buf ( g4816 , g147 );
buf ( g4817 , g148 );
buf ( g4818 , g149 );
buf ( g4819 , g150 );
buf ( g4820 , g151 );
buf ( g4821 , g152 );
buf ( g4822 , g153 );
buf ( g4823 , g154 );
buf ( g4824 , g155 );
buf ( g4825 , g156 );
buf ( g157 , g4826 );
buf ( g158 , g4827 );
buf ( g159 , g4828 );
buf ( g160 , g4829 );
buf ( g161 , g4830 );
buf ( g162 , g4831 );
buf ( g163 , g4832 );
buf ( g164 , g4833 );
buf ( g165 , g4834 );
buf ( g166 , g4835 );
buf ( g167 , g4836 );
buf ( g168 , g4837 );
buf ( g169 , g4838 );
buf ( g170 , g4839 );
buf ( g171 , g4840 );
buf ( g172 , g4841 );
buf ( g173 , g4842 );
buf ( g174 , g4843 );
buf ( g175 , g4844 );
buf ( g176 , g4845 );
buf ( g177 , g4846 );
buf ( g178 , g4847 );
buf ( g179 , g4848 );
buf ( g180 , g4849 );
buf ( g181 , g4850 );
buf ( g182 , g4851 );
buf ( g183 , g4852 );
buf ( g184 , g4853 );
buf ( g185 , g4854 );
buf ( g186 , g4855 );
buf ( g187 , g4856 );
buf ( g188 , g4857 );
buf ( g189 , g4858 );
buf ( g190 , g4859 );
buf ( g191 , g4860 );
buf ( g192 , g4861 );
buf ( g193 , g4862 );
buf ( g194 , g4863 );
buf ( g195 , g4864 );
buf ( g196 , g4865 );
buf ( g197 , g4866 );
buf ( g198 , g4867 );
buf ( g199 , g4868 );
buf ( g200 , g4869 );
buf ( g201 , g4870 );
buf ( g202 , g4871 );
buf ( g203 , g4872 );
buf ( g204 , g4873 );
buf ( g205 , g4874 );
buf ( g206 , g4875 );
buf ( g207 , g4876 );
buf ( g208 , g4877 );
buf ( g209 , g4878 );
buf ( g210 , g4879 );
buf ( g211 , g4880 );
buf ( g212 , g4881 );
buf ( g213 , g4882 );
buf ( g214 , g4883 );
buf ( g215 , g4884 );
buf ( g216 , g4885 );
buf ( g217 , g4886 );
buf ( g218 , g4887 );
buf ( g219 , g4888 );
buf ( g220 , g4889 );
buf ( g4826 , g4783 );
buf ( g4827 , g4783 );
buf ( g4828 , g4783 );
buf ( g4829 , g4792 );
buf ( g4830 , g4792 );
buf ( g4831 , g4805 );
buf ( g4832 , g4805 );
buf ( g4833 , g4805 );
buf ( g4834 , g1004 );
buf ( g4835 , g1001 );
buf ( g4836 , g995 );
buf ( g4837 , g998 );
buf ( g4838 , g1002 );
buf ( g4839 , g1000 );
buf ( g4840 , g997 );
buf ( g4841 , g994 );
buf ( g4842 , g992 );
buf ( g4843 , g993 );
buf ( g4844 , g4783 );
buf ( g4845 , g1344 );
buf ( g4846 , g1357 );
buf ( g4847 , g1350 );
buf ( g4848 , g1358 );
buf ( g4849 , g990 );
buf ( g4850 , g991 );
buf ( g4851 , g958 );
buf ( g4852 , g1126 );
buf ( g4853 , g784 );
buf ( g4854 , g1146 );
buf ( g4855 , g807 );
buf ( g4856 , g653 );
buf ( g4857 , g589 );
buf ( g4858 , g983 );
buf ( g4859 , g1352 );
buf ( g4860 , g989 );
buf ( g4861 , g975 );
buf ( g4862 , g590 );
buf ( g4863 , g1199 );
buf ( g4864 , g1245 );
buf ( g4865 , g732 );
buf ( g4866 , g1135 );
buf ( g4867 , g457 );
buf ( g4868 , g1356 );
buf ( g4869 , g1356 );
buf ( g4870 , g1348 );
buf ( g4871 , g1348 );
buf ( g4872 , g1343 );
buf ( g4873 , g1017 );
buf ( g4874 , g1017 );
buf ( g4875 , g1325 );
buf ( g4876 , g1240 );
buf ( g4877 , g923 );
buf ( g4878 , g971 );
buf ( g4879 , g821 );
buf ( g4880 , g820 );
buf ( g4881 , g902 );
buf ( g4882 , g1197 );
buf ( g4883 , g1338 );
buf ( g4884 , g1338 );
buf ( g4885 , g1339 );
buf ( g4886 , g1377 );
buf ( g4887 , 1'b0 );
buf ( g4888 , g1244 );
buf ( g4889 , g1243 );
not ( g445 , g4680 );
nand ( g446 , g4788 , g4785 );
not ( g447 , g4722 );
nor ( g448 , g446 , g447 );
not ( g449 , g448 );
not ( g450 , g4788 );
nand ( g451 , g450 , g4785 , g4701 );
not ( g452 , g4712 );
nor ( g453 , g452 , g4785 );
nand ( g454 , g453 , g4788 );
nor ( g455 , g4788 , g4785 );
nand ( g456 , g455 , g4733 );
nand ( g457 , g449 , g451 , g454 , g456 );
not ( g458 , g457 );
or ( g459 , g445 , g458 );
not ( g460 , g4680 );
nand ( g461 , g460 , g4686 );
nand ( g462 , g459 , g461 );
nor ( g463 , g462 , g4802 );
not ( g464 , g463 );
not ( g465 , g4769 );
not ( g466 , g4814 );
nor ( g467 , g466 , g4813 );
nand ( g468 , g465 , g467 );
not ( g469 , g468 );
not ( g470 , g4779 );
nor ( g471 , g4813 , g4814 );
nand ( g472 , g470 , g471 );
not ( g473 , g472 );
or ( g474 , g469 , g473 );
nand ( g475 , g474 , g4691 );
not ( g476 , g4759 );
nand ( g477 , g476 , g4813 , g4814 );
not ( g478 , g4814 );
not ( g479 , g4749 );
nand ( g480 , g478 , g479 , g4813 );
or ( g481 , g4691 , g4693 );
nand ( g482 , g477 , g480 , g481 );
not ( g483 , g4691 );
nand ( g484 , g483 , g481 );
nand ( g485 , g482 , g484 );
nand ( g486 , g475 , g485 , g4807 );
not ( g487 , g4765 );
not ( g488 , g4814 );
nor ( g489 , g488 , g4813 );
nand ( g490 , g487 , g489 );
not ( g491 , g4745 );
not ( g492 , g4813 );
nor ( g493 , g492 , g4814 );
nand ( g494 , g491 , g493 );
not ( g495 , g4813 );
not ( g496 , g4814 );
nor ( g497 , g495 , g496 );
not ( g498 , g4755 );
nand ( g499 , g497 , g498 );
not ( g500 , g4775 );
nor ( g501 , g4813 , g4814 );
nand ( g502 , g500 , g501 );
nand ( g503 , g490 , g494 , g499 , g502 );
and ( g504 , g503 , g4691 );
or ( g505 , g4690 , g4691 );
nand ( g506 , g505 , g4677 );
nor ( g507 , g504 , g506 );
and ( g508 , g464 , g486 , g507 );
not ( g509 , g4801 );
not ( g510 , g4680 );
not ( g511 , g4734 );
nor ( g512 , g511 , g4785 , g4788 );
nand ( g513 , g4788 , g4785 );
not ( g514 , g4723 );
nor ( g515 , g513 , g514 );
nor ( g516 , g512 , g515 );
not ( g517 , g516 );
not ( g518 , g4788 );
nand ( g519 , g518 , g4702 );
and ( g520 , g4785 , g519 );
not ( g521 , g4785 );
nand ( g522 , g4713 , g4788 );
and ( g523 , g521 , g522 );
nor ( g524 , g520 , g523 );
nor ( g525 , g517 , g524 );
not ( g526 , g525 );
or ( g527 , g510 , g526 );
or ( g528 , g4674 , g4680 );
nand ( g529 , g527 , g528 );
and ( g530 , g509 , g529 );
and ( g531 , g462 , g4802 );
nor ( g532 , g530 , g531 );
not ( g533 , g4680 );
not ( g534 , g4739 );
nor ( g535 , g534 , g4785 );
not ( g536 , g4788 );
nand ( g537 , g535 , g536 );
not ( g538 , g4788 );
nand ( g539 , g4785 , g538 , g4707 );
not ( g540 , g4785 );
nand ( g541 , g540 , g4788 , g4717 );
nand ( g542 , g4788 , g4728 , g4785 );
nand ( g543 , g537 , g539 , g541 , g542 );
not ( g544 , g543 );
or ( g545 , g533 , g544 );
nand ( g546 , g460 , g4682 );
nand ( g547 , g545 , g546 );
and ( g548 , g547 , g4796 );
not ( g549 , g547 );
not ( g550 , g4796 );
and ( g551 , g549 , g550 );
nor ( g552 , g548 , g551 );
not ( g553 , g4691 );
not ( g554 , g4813 );
not ( g555 , g4763 );
nand ( g556 , g554 , g555 , g4814 );
not ( g557 , g4753 );
nand ( g558 , g557 , g4813 , g4814 );
nor ( g559 , g4814 , g4743 );
nand ( g560 , g559 , g4813 );
not ( g561 , g4814 );
not ( g562 , g4773 );
nand ( g563 , g561 , g495 , g562 );
nand ( g564 , g556 , g558 , g560 , g563 );
not ( g565 , g564 );
or ( g566 , g553 , g565 );
or ( g567 , g4687 , g4691 );
nand ( g568 , g566 , g567 );
not ( g569 , g4803 );
and ( g570 , g568 , g569 );
not ( g571 , g568 );
and ( g572 , g571 , g4803 );
nor ( g573 , g570 , g572 );
nand ( g574 , g508 , g532 , g552 , g573 );
not ( g575 , g4680 );
not ( g576 , g4785 );
nor ( g577 , g576 , g4788 );
not ( g578 , g4706 );
nand ( g579 , g577 , g578 );
not ( g580 , g4788 );
nor ( g581 , g580 , g4785 );
not ( g582 , g4716 );
nand ( g583 , g581 , g582 );
not ( g584 , g4738 );
nor ( g585 , g4785 , g4788 );
nand ( g586 , g584 , g585 );
not ( g587 , g4727 );
nand ( g588 , g587 , g4788 , g4785 );
nand ( g589 , g579 , g583 , g586 , g588 );
not ( g590 , g589 );
not ( g591 , g590 );
or ( g592 , g575 , g591 );
nand ( g593 , g460 , g4673 );
nand ( g594 , g592 , g593 );
not ( g595 , g594 );
not ( g596 , g4797 );
and ( g597 , g595 , g596 );
and ( g598 , g594 , g4797 );
nor ( g599 , g597 , g598 );
not ( g600 , g4691 );
not ( g601 , g4814 );
and ( g602 , g4813 , g4757 );
not ( g603 , g4813 );
and ( g604 , g603 , g4767 );
nor ( g605 , g602 , g604 );
nor ( g606 , g601 , g605 );
nor ( g607 , g4814 , g4813 );
nand ( g608 , g607 , g4777 );
not ( g609 , g4814 );
nand ( g610 , g609 , g4747 , g4813 );
nand ( g611 , g608 , g610 );
nor ( g612 , g606 , g611 );
not ( g613 , g612 );
or ( g614 , g600 , g613 );
or ( g615 , g4691 , g4694 );
nand ( g616 , g614 , g615 );
not ( g617 , g616 );
not ( g618 , g4809 );
not ( g619 , g618 );
and ( g620 , g617 , g619 );
not ( g621 , g529 );
and ( g622 , g621 , g4801 );
nor ( g623 , g620 , g622 );
not ( g624 , g4680 );
not ( g625 , g4785 );
not ( g626 , g4731 );
not ( g627 , g4788 );
nand ( g628 , g625 , g626 , g627 );
not ( g629 , g4699 );
not ( g630 , g4788 );
nand ( g631 , g629 , g630 , g4785 );
not ( g632 , g4785 );
not ( g633 , g4710 );
nand ( g634 , g632 , g633 , g4788 );
not ( g635 , g4720 );
nand ( g636 , g635 , g4788 , g4785 );
nand ( g637 , g628 , g631 , g634 , g636 );
not ( g638 , g637 );
or ( g639 , g624 , g638 );
or ( g640 , g4680 , g4681 );
nand ( g641 , g639 , g640 );
xnor ( g642 , g641 , g4793 );
not ( g643 , g4680 );
not ( g644 , g4715 );
nand ( g645 , g581 , g644 );
not ( g646 , g4705 );
nand ( g647 , g577 , g646 );
not ( g648 , g4737 );
nor ( g649 , g4785 , g4788 );
nand ( g650 , g648 , g649 );
not ( g651 , g4726 );
nand ( g652 , g651 , g4785 , g4788 );
nand ( g653 , g645 , g647 , g650 , g652 );
not ( g654 , g653 );
or ( g655 , g643 , g654 );
or ( g656 , g4680 , g4683 );
nand ( g657 , g655 , g656 );
not ( g658 , g4798 );
and ( g659 , g657 , g658 );
not ( g660 , g657 );
and ( g661 , g660 , g4798 );
nor ( g662 , g659 , g661 );
nand ( g663 , g599 , g623 , g642 , g662 );
nor ( g664 , g574 , g663 );
not ( g665 , g4680 );
nor ( g666 , g4788 , g4740 );
not ( g667 , g4785 );
nand ( g668 , g666 , g667 );
not ( g669 , g4708 );
not ( g670 , g4788 );
nand ( g671 , g669 , g670 , g4785 );
not ( g672 , g4729 );
nand ( g673 , g672 , g4788 , g4785 );
not ( g674 , g4718 );
nand ( g675 , g667 , g674 , g4788 );
nand ( g676 , g668 , g671 , g673 , g675 );
not ( g677 , g676 );
not ( g678 , g677 );
not ( g679 , g678 );
or ( g680 , g665 , g679 );
or ( g681 , g4672 , g4680 );
nand ( g682 , g680 , g681 );
not ( g683 , g682 );
and ( g684 , g683 , g4794 );
not ( g685 , g4804 );
not ( g686 , g685 );
not ( g687 , g4691 );
not ( g688 , g4761 );
nand ( g689 , g688 , g4813 , g4814 );
not ( g690 , g4771 );
nand ( g691 , g690 , g489 );
not ( g692 , g4781 );
nand ( g693 , g692 , g501 );
not ( g694 , g4751 );
nand ( g695 , g694 , g466 , g4813 );
nand ( g696 , g689 , g691 , g693 , g695 );
not ( g697 , g696 );
or ( g698 , g687 , g697 );
or ( g699 , g4691 , g4692 );
nand ( g700 , g698 , g699 );
not ( g701 , g700 );
or ( g702 , g686 , g701 );
not ( g703 , g4691 );
not ( g704 , g4770 );
not ( g705 , g4814 );
nor ( g706 , g705 , g4813 );
nand ( g707 , g704 , g706 );
nor ( g708 , g4814 , g4750 );
nand ( g709 , g708 , g4813 );
not ( g710 , g4760 );
nand ( g711 , g710 , g4813 , g4814 );
not ( g712 , g4780 );
nor ( g713 , g4814 , g4813 );
nand ( g714 , g712 , g713 );
nand ( g715 , g707 , g709 , g711 , g714 );
not ( g716 , g715 );
or ( g717 , g703 , g716 );
or ( g718 , g4691 , g4688 );
nand ( g719 , g717 , g718 );
not ( g720 , g4806 );
or ( g721 , g719 , g720 );
nand ( g722 , g702 , g721 );
nor ( g723 , g684 , g722 );
not ( g724 , g4680 );
nand ( g725 , g4703 , g4785 );
nor ( g726 , g725 , g4788 );
not ( g727 , g726 );
not ( g728 , g4785 );
nand ( g729 , g728 , g4735 );
nand ( g730 , g728 , g4788 );
nand ( g731 , g4788 , g4724 );
nand ( g732 , g727 , g729 , g730 , g731 );
not ( g733 , g732 );
or ( g734 , g724 , g733 );
nand ( g735 , g460 , g4685 );
nand ( g736 , g734 , g735 );
and ( g737 , g736 , g4800 );
not ( g738 , g736 );
not ( g739 , g4800 );
and ( g740 , g738 , g739 );
nor ( g741 , g737 , g740 );
not ( g742 , g700 );
nand ( g743 , g742 , g4804 );
and ( g744 , g741 , g743 );
and ( g745 , g720 , g719 );
and ( g746 , g616 , g618 );
nor ( g747 , g745 , g746 );
nand ( g748 , g723 , g744 , g747 );
nand ( g749 , g475 , g485 );
not ( g750 , g4807 );
and ( g751 , g749 , g750 );
and ( g752 , g4813 , g4758 );
not ( g753 , g4813 );
and ( g754 , g753 , g4768 );
nor ( g755 , g752 , g754 );
nand ( g756 , g755 , g4814 );
not ( g757 , g756 );
and ( g758 , g4813 , g4748 );
not ( g759 , g4813 );
and ( g760 , g759 , g4778 );
nor ( g761 , g758 , g760 );
nand ( g762 , g761 , g466 );
not ( g763 , g762 );
or ( g764 , g757 , g763 );
nand ( g765 , g764 , g4691 );
or ( g766 , g4691 , g4689 );
nand ( g767 , g765 , g766 );
not ( g768 , g4808 );
xnor ( g769 , g767 , g768 );
nor ( g770 , g751 , g769 );
not ( g771 , g4794 );
nand ( g772 , g682 , g771 );
nand ( g773 , g4814 , g4813 );
nor ( g774 , g773 , g4756 );
not ( g775 , g774 );
nor ( g776 , g4814 , g4746 );
nand ( g777 , g776 , g4813 );
not ( g778 , g4813 );
not ( g779 , g4766 );
nand ( g780 , g778 , g779 , g4814 );
nor ( g781 , g4814 , g4813 );
not ( g782 , g4776 );
nand ( g783 , g781 , g782 );
nand ( g784 , g775 , g777 , g780 , g783 );
and ( g785 , g784 , g4691 );
nor ( g786 , g4691 , g4695 );
nor ( g787 , g785 , g786 );
and ( g788 , g787 , g4810 );
not ( g789 , g787 );
not ( g790 , g4810 );
and ( g791 , g789 , g790 );
nor ( g792 , g788 , g791 );
not ( g793 , g4680 );
nand ( g794 , g4788 , g4785 );
not ( g795 , g794 );
not ( g796 , g4725 );
and ( g797 , g795 , g796 );
nor ( g798 , g4788 , g4736 );
and ( g799 , g798 , g728 );
nor ( g800 , g797 , g799 );
not ( g801 , g4714 );
not ( g802 , g4785 );
nand ( g803 , g801 , g802 , g4788 );
not ( g804 , g4788 );
not ( g805 , g4704 );
nand ( g806 , g804 , g805 , g4785 );
nand ( g807 , g800 , g803 , g806 );
not ( g808 , g807 );
or ( g809 , g793 , g808 );
or ( g810 , g4680 , g4684 );
nand ( g811 , g809 , g810 );
not ( g812 , g811 );
not ( g813 , g4799 );
not ( g814 , g813 );
and ( g815 , g812 , g814 );
and ( g816 , g811 , g813 );
nor ( g817 , g815 , g816 );
nand ( g818 , g770 , g772 , g792 , g817 );
nor ( g819 , g748 , g818 );
nand ( g820 , g664 , g819 );
not ( g821 , g820 );
not ( g822 , g611 );
not ( g823 , g4813 );
nand ( g824 , g823 , g4767 , g4814 );
nand ( g825 , g4813 , g4757 , g4814 );
nand ( g826 , g824 , g825 , g4698 );
not ( g827 , g826 );
not ( g828 , g4748 );
nand ( g829 , g828 , g4813 );
not ( g830 , g4813 );
not ( g831 , g4778 );
nand ( g832 , g830 , g831 );
nor ( g833 , g4795 , g4814 );
nand ( g834 , g829 , g832 , g833 );
nor ( g835 , g4813 , g4768 );
not ( g836 , g835 );
not ( g837 , g4758 );
nand ( g838 , g837 , g4813 );
not ( g839 , g4795 );
nand ( g840 , g836 , g838 , g839 , g4814 );
nand ( g841 , g822 , g827 , g834 , g840 );
not ( g842 , g841 );
not ( g843 , g842 );
not ( g844 , g715 );
nand ( g845 , g844 , g4806 );
nand ( g846 , g4802 , g457 );
nand ( g847 , g560 , g563 );
not ( g848 , g847 );
not ( g849 , g556 );
not ( g850 , g849 );
nand ( g851 , g848 , g850 , g558 , g4803 );
nand ( g852 , g845 , g846 , g851 );
not ( g853 , g852 );
or ( g854 , g843 , g853 );
not ( g855 , g841 );
nand ( g856 , g689 , g693 );
not ( g857 , g856 );
and ( g858 , g691 , g695 );
nand ( g859 , g857 , g858 );
nor ( g860 , g859 , g685 );
nand ( g861 , g855 , g860 );
nand ( g862 , g854 , g861 );
not ( g863 , g862 );
not ( g864 , g4790 );
not ( g865 , g864 );
nand ( g866 , g678 , g4786 );
not ( g867 , g866 );
or ( g868 , g865 , g867 );
buf ( g869 , g637 );
not ( g870 , g869 );
nand ( g871 , g870 , g4790 );
nand ( g872 , g868 , g871 );
not ( g873 , g4709 );
nand ( g874 , g873 , g4785 , g538 );
not ( g875 , g4741 );
nor ( g876 , g4785 , g4788 );
nand ( g877 , g875 , g876 );
not ( g878 , g4788 );
not ( g879 , g878 );
nor ( g880 , g4785 , g4719 );
nand ( g881 , g879 , g880 );
not ( g882 , g4730 );
nand ( g883 , g882 , g4785 , g4788 );
nand ( g884 , g874 , g877 , g881 , g883 );
not ( g885 , g884 );
not ( g886 , g4785 );
nand ( g887 , g886 , g633 , g4788 );
nor ( g888 , g4785 , g4731 );
nand ( g889 , g878 , g888 );
nand ( g890 , g635 , g4785 , g4788 );
nand ( g891 , g887 , g631 , g889 , g890 );
not ( g892 , g891 );
or ( g893 , g885 , g892 );
not ( g894 , g884 );
not ( g895 , g891 );
nand ( g896 , g894 , g895 );
nand ( g897 , g893 , g896 );
not ( g898 , g897 );
and ( g899 , g872 , g898 );
not ( g900 , g872 );
and ( g901 , g900 , g897 );
nor ( g902 , g899 , g901 );
and ( g903 , g4810 , g4809 );
not ( g904 , g4810 );
and ( g905 , g904 , g618 );
or ( g906 , g903 , g905 );
xnor ( g907 , g4807 , g4808 );
xor ( g908 , g906 , g907 );
not ( g909 , g908 );
or ( g910 , g720 , g4825 );
not ( g911 , g4825 );
or ( g912 , g911 , g4806 );
nand ( g913 , g910 , g912 );
not ( g914 , g913 );
xnor ( g915 , g4811 , g4812 );
not ( g916 , g915 );
or ( g917 , g914 , g916 );
or ( g918 , g915 , g913 );
nand ( g919 , g917 , g918 );
not ( g920 , g919 );
or ( g921 , g909 , g920 );
or ( g922 , g919 , g908 );
nand ( g923 , g921 , g922 );
not ( g924 , g923 );
xor ( g925 , g4796 , g4801 );
xor ( g926 , g4804 , g4802 );
and ( g927 , g925 , g926 );
not ( g928 , g925 );
not ( g929 , g926 );
and ( g930 , g928 , g929 );
nor ( g931 , g927 , g930 );
not ( g932 , g4800 );
not ( g933 , g813 );
or ( g934 , g932 , g933 );
nand ( g935 , g739 , g4799 );
nand ( g936 , g934 , g935 );
not ( g937 , g936 );
and ( g938 , g931 , g937 );
not ( g939 , g931 );
and ( g940 , g939 , g936 );
nor ( g941 , g938 , g940 );
and ( g942 , g4803 , g4824 );
not ( g943 , g4803 );
not ( g944 , g4824 );
and ( g945 , g943 , g944 );
or ( g946 , g942 , g945 );
xor ( g947 , g4797 , g4798 );
xor ( g948 , g946 , g947 );
and ( g949 , g941 , g948 );
not ( g950 , g941 );
not ( g951 , g948 );
and ( g952 , g950 , g951 );
nor ( g953 , g949 , g952 );
nand ( g954 , g4700 , g4732 , g4744 , g4774 );
and ( g955 , g954 , g4815 );
nand ( g956 , g4711 , g4721 , g4754 , g4764 );
and ( g957 , g956 , g4787 );
nor ( g958 , g955 , g957 );
nand ( g959 , g924 , g953 , g958 );
not ( g960 , g750 );
not ( g961 , g543 );
not ( g962 , g961 );
or ( g963 , g960 , g962 );
nand ( g964 , g963 , g4806 );
nor ( g965 , g611 , g826 );
nand ( g966 , g834 , g840 );
nand ( g967 , g965 , g966 );
not ( g968 , g967 );
or ( g969 , g961 , g678 );
nand ( g970 , g964 , g968 , g969 );
not ( g971 , g953 );
nand ( g972 , g707 , g709 , g711 , g714 );
xor ( g973 , g972 , g696 );
not ( g974 , g973 );
buf ( g975 , g543 );
nor ( g976 , g975 , g4697 );
not ( g977 , g550 );
not ( g978 , g961 );
or ( g979 , g977 , g978 );
nand ( g980 , g979 , g4794 );
not ( g981 , g637 );
nand ( g982 , g981 , g677 );
nand ( g983 , g869 , g4790 );
buf ( g984 , g884 );
not ( g985 , g984 );
and ( g986 , g4669 , g4671 );
nand ( g987 , g4784 , g4789 );
nor ( g988 , g986 , g987 );
nand ( g989 , g988 , g958 );
nor ( g990 , g954 , g956 );
not ( g991 , g990 );
nand ( g992 , g4808 , g4809 , g4807 , g4810 );
nand ( g993 , g4789 , g4670 , g4679 );
not ( g994 , g4754 );
not ( g995 , g4732 );
not ( g996 , g4820 );
not ( g997 , g4711 );
not ( g998 , g4744 );
not ( g999 , g4819 );
not ( g1000 , g4764 );
not ( g1001 , g4774 );
not ( g1002 , g4721 );
not ( g1003 , g4697 );
not ( g1004 , g4700 );
not ( g1005 , g4676 );
nand ( g1006 , g670 , g669 , g4785 );
not ( g1007 , g4729 );
nand ( g1008 , g1007 , g4788 , g4785 );
not ( g1009 , g4785 );
nand ( g1010 , g1009 , g674 , g4788 );
nand ( g1011 , g668 , g1006 , g1008 , g1010 );
not ( g1012 , g1011 );
nor ( g1013 , g1012 , g4786 );
and ( g1014 , g4791 , g1013 );
not ( g1015 , g4791 );
and ( g1016 , g1015 , g869 );
nor ( g1017 , g1014 , g1016 );
not ( g1018 , g794 );
not ( g1019 , g4725 );
and ( g1020 , g1018 , g1019 );
and ( g1021 , g798 , g728 );
nor ( g1022 , g1020 , g1021 );
not ( g1023 , g1022 );
not ( g1024 , g4788 );
nand ( g1025 , g1024 , g805 , g4785 );
nand ( g1026 , g576 , g801 , g4788 );
nand ( g1027 , g1025 , g1026 );
not ( g1028 , g1027 );
not ( g1029 , g1028 );
or ( g1030 , g1023 , g1029 );
not ( g1031 , g448 );
nand ( g1032 , g1031 , g456 , g451 , g454 );
nand ( g1033 , g1030 , g1032 );
not ( g1034 , g455 );
not ( g1035 , g4733 );
or ( g1036 , g1034 , g1035 );
nand ( g1037 , g4788 , g4785 , g4722 );
nand ( g1038 , g1036 , g1037 );
not ( g1039 , g1038 );
nor ( g1040 , g452 , g4785 );
and ( g1041 , g1040 , g4788 );
nand ( g1042 , g4785 , g4701 );
nor ( g1043 , g1042 , g4788 );
nor ( g1044 , g1041 , g1043 );
nand ( g1045 , g1039 , g1028 , g1044 , g1022 );
nand ( g1046 , g1033 , g1045 );
not ( g1047 , g732 );
nand ( g1048 , g4713 , g4788 );
nor ( g1049 , g1048 , g4785 );
not ( g1050 , g1049 );
nand ( g1051 , g4702 , g4785 , g536 );
nand ( g1052 , g1050 , g516 , g1051 );
not ( g1053 , g1052 );
or ( g1054 , g1047 , g1053 );
not ( g1055 , g4724 );
nand ( g1056 , g1055 , g4785 );
and ( g1057 , g1056 , g4788 );
nor ( g1058 , g1057 , g1049 );
nand ( g1059 , g4785 , g4788 );
not ( g1060 , g1059 );
not ( g1061 , g514 );
and ( g1062 , g1060 , g1061 );
not ( g1063 , g4734 );
nor ( g1064 , g1063 , g4785 , g4788 );
nor ( g1065 , g1062 , g1064 );
nand ( g1066 , g4703 , g4785 );
not ( g1067 , g1066 );
not ( g1068 , g4788 );
and ( g1069 , g1067 , g1068 );
and ( g1070 , g728 , g4735 );
nor ( g1071 , g1069 , g1070 );
nand ( g1072 , g1058 , g1065 , g1071 , g1051 );
nand ( g1073 , g1054 , g1072 );
xor ( g1074 , g1046 , g1073 );
buf ( g1075 , g1074 );
not ( g1076 , g1011 );
not ( g1077 , g891 );
or ( g1078 , g1076 , g1077 );
nand ( g1079 , g1078 , g982 );
and ( g1080 , g1079 , g984 );
not ( g1081 , g1079 );
and ( g1082 , g1081 , g985 );
nor ( g1083 , g1080 , g1082 );
and ( g1084 , g1083 , g976 );
not ( g1085 , g1083 );
and ( g1086 , g975 , g1003 );
and ( g1087 , g1085 , g1086 );
nor ( g1088 , g1084 , g1087 );
not ( g1089 , g975 );
xnor ( g1090 , g1089 , g1083 );
nand ( g1091 , g480 , g477 , g472 , g468 );
not ( g1092 , g4756 );
nand ( g1093 , g1092 , g4814 , g4813 );
nand ( g1094 , g780 , g777 , g783 , g1093 );
not ( g1095 , g1094 );
and ( g1096 , g1091 , g1095 );
not ( g1097 , g1091 );
and ( g1098 , g1097 , g1094 );
nor ( g1099 , g1096 , g1098 );
not ( g1100 , g1099 );
and ( g1101 , g4821 , g4820 );
not ( g1102 , g4821 );
and ( g1103 , g1102 , g996 );
nor ( g1104 , g1101 , g1103 );
and ( g1105 , g4794 , g4817 );
not ( g1106 , g4794 );
not ( g1107 , g4817 );
and ( g1108 , g1106 , g1107 );
nor ( g1109 , g1105 , g1108 );
and ( g1110 , g1104 , g1109 );
not ( g1111 , g1104 );
not ( g1112 , g1109 );
and ( g1113 , g1111 , g1112 );
nor ( g1114 , g1110 , g1113 );
and ( g1115 , g4793 , g4818 );
not ( g1116 , g4793 );
not ( g1117 , g4818 );
and ( g1118 , g1116 , g1117 );
nor ( g1119 , g1115 , g1118 );
not ( g1120 , g4747 );
not ( g1121 , g4813 );
nor ( g1122 , g1121 , g4814 );
not ( g1123 , g1122 );
or ( g1124 , g1120 , g1123 );
nand ( g1125 , g1124 , g608 );
nor ( g1126 , g1125 , g606 );
or ( g1127 , g564 , g1126 );
nand ( g1128 , g1126 , g564 );
nand ( g1129 , g1127 , g1128 );
and ( g1130 , g1129 , g1100 );
not ( g1131 , g1129 );
and ( g1132 , g1131 , g1099 );
nor ( g1133 , g1130 , g1132 );
nand ( g1134 , g4800 , g732 );
not ( g1135 , g525 );
nand ( g1136 , g1135 , g4801 );
and ( g1137 , g1134 , g1136 );
nor ( g1138 , g1137 , g1005 );
not ( g1139 , g4814 );
and ( g1140 , g4813 , g4758 );
not ( g1141 , g4813 );
and ( g1142 , g1141 , g4768 );
nor ( g1143 , g1140 , g1142 );
not ( g1144 , g1143 );
or ( g1145 , g1139 , g1144 );
nand ( g1146 , g1145 , g762 );
not ( g1147 , g4814 );
not ( g1148 , g4752 );
and ( g1149 , g4813 , g1148 );
not ( g1150 , g4813 );
not ( g1151 , g4782 );
and ( g1152 , g1150 , g1151 );
nor ( g1153 , g1149 , g1152 );
and ( g1154 , g1147 , g1153 );
not ( g1155 , g1147 );
not ( g1156 , g4762 );
and ( g1157 , g4813 , g1156 );
not ( g1158 , g4813 );
not ( g1159 , g4772 );
and ( g1160 , g1158 , g1159 );
nor ( g1161 , g1157 , g1160 );
and ( g1162 , g1155 , g1161 );
nor ( g1163 , g1154 , g1162 );
and ( g1164 , g1146 , g1163 );
not ( g1165 , g1146 );
and ( g1166 , g4813 , g4752 );
not ( g1167 , g4813 );
and ( g1168 , g1167 , g4782 );
or ( g1169 , g1166 , g1168 );
and ( g1170 , g1147 , g1169 );
not ( g1171 , g1147 );
and ( g1172 , g4813 , g4762 );
not ( g1173 , g4813 );
and ( g1174 , g1173 , g4772 );
or ( g1175 , g1172 , g1174 );
and ( g1176 , g1171 , g1175 );
or ( g1177 , g1170 , g1176 );
and ( g1178 , g1165 , g1177 );
nor ( g1179 , g1164 , g1178 );
and ( g1180 , g1179 , g503 );
not ( g1181 , g1179 );
not ( g1182 , g503 );
and ( g1183 , g1181 , g1182 );
nor ( g1184 , g1180 , g1183 );
not ( g1185 , g973 );
nand ( g1186 , g1184 , g1185 );
not ( g1187 , g1186 );
not ( g1188 , g1184 );
not ( g1189 , g974 );
nand ( g1190 , g1188 , g1189 );
not ( g1191 , g1190 );
or ( g1192 , g1187 , g1191 );
nor ( g1193 , g1133 , g4697 );
nand ( g1194 , g1192 , g1193 );
not ( g1195 , g4697 );
nand ( g1196 , g1190 , g1133 , g1186 , g1195 );
nand ( g1197 , g1194 , g1196 );
not ( g1198 , g1074 );
not ( g1199 , g653 );
not ( g1200 , g1199 );
not ( g1201 , g590 );
or ( g1202 , g1200 , g1201 );
nand ( g1203 , g653 , g589 );
nand ( g1204 , g1202 , g1203 );
nor ( g1205 , g1204 , g4697 );
nand ( g1206 , g1198 , g1205 );
nand ( g1207 , g1074 , g1204 , g1003 );
nand ( g1208 , g1088 , g1206 , g1207 );
not ( g1209 , g1204 );
not ( g1210 , g1074 );
or ( g1211 , g1209 , g1210 );
or ( g1212 , g1074 , g1204 );
nand ( g1213 , g1211 , g1212 );
not ( g1214 , g1213 );
not ( g1215 , g1090 );
or ( g1216 , g1214 , g1215 );
nand ( g1217 , g1216 , g1208 );
xnor ( g1218 , g4823 , g4822 );
not ( g1219 , g1218 );
and ( g1220 , g4816 , g999 );
not ( g1221 , g4816 );
and ( g1222 , g1221 , g4819 );
or ( g1223 , g1220 , g1222 );
not ( g1224 , g1223 );
or ( g1225 , g1219 , g1224 );
not ( g1226 , g1223 );
not ( g1227 , g1218 );
nand ( g1228 , g1226 , g1227 );
nand ( g1229 , g1225 , g1228 );
not ( g1230 , g1229 );
and ( g1231 , g1114 , g1119 );
not ( g1232 , g1114 );
not ( g1233 , g1119 );
and ( g1234 , g1232 , g1233 );
nor ( g1235 , g1231 , g1234 );
nor ( g1236 , g1230 , g1235 );
not ( g1237 , g1235 );
or ( g1238 , g1237 , g1229 );
nand ( g1239 , g1238 , g4678 );
nor ( g1240 , g1236 , g1239 );
or ( g1241 , g959 , g1240 );
nor ( g1242 , g1197 , g1241 );
nand ( g1243 , g1217 , g1242 );
not ( g1244 , g1243 );
not ( g1245 , g807 );
not ( g1246 , g1245 );
not ( g1247 , g4809 );
nand ( g1248 , g965 , g966 );
not ( g1249 , g1248 );
not ( g1250 , g1249 );
or ( g1251 , g1247 , g1250 );
or ( g1252 , g658 , g1249 );
nand ( g1253 , g1251 , g1252 );
nand ( g1254 , g1253 , g1199 );
nor ( g1255 , g678 , g771 );
and ( g1256 , g859 , g685 );
buf ( g1257 , g715 );
and ( g1258 , g1257 , g720 );
nor ( g1259 , g1256 , g1258 );
xor ( g1260 , g961 , g866 );
xnor ( g1261 , g1260 , g897 );
not ( g1262 , g1261 );
and ( g1263 , g1198 , g4791 );
nand ( g1264 , g1262 , g1263 );
not ( g1265 , g968 );
nand ( g1266 , g1265 , g980 , g969 );
nand ( g1267 , g1266 , g970 );
buf ( g1268 , g1248 );
or ( g1269 , g4801 , g1135 );
not ( g1270 , g732 );
nand ( g1271 , g1270 , g1136 , g739 );
nand ( g1272 , g1269 , g1271 );
nand ( g1273 , g1268 , g1138 );
nand ( g1274 , g813 , g1248 );
not ( g1275 , g1249 );
not ( g1276 , g790 );
or ( g1277 , g1275 , g1276 );
nand ( g1278 , g1277 , g1274 );
or ( g1279 , g1278 , g1246 );
nand ( g1280 , g1279 , g1254 );
nand ( g1281 , g863 , g1273 );
not ( g1282 , g4807 );
not ( g1283 , g968 );
or ( g1284 , g1282 , g1283 );
nand ( g1285 , g967 , g4796 );
nand ( g1286 , g1284 , g1285 );
not ( g1287 , g1011 );
nand ( g1288 , g1286 , g1287 );
and ( g1289 , g1267 , g1288 );
nor ( g1290 , g1249 , g1255 , g4793 );
not ( g1291 , g1290 );
not ( g1292 , g870 );
not ( g1293 , g1292 );
or ( g1294 , g1291 , g1293 );
and ( g1295 , g1287 , g4806 );
nor ( g1296 , g1295 , g4804 );
nand ( g1297 , g1292 , g1296 , g1249 );
nand ( g1298 , g1294 , g1297 );
nor ( g1299 , g1289 , g1298 );
not ( g1300 , g1286 );
buf ( g1301 , g975 );
not ( g1302 , g1301 );
or ( g1303 , g1300 , g1302 );
not ( g1304 , g4797 );
not ( g1305 , g1304 );
not ( g1306 , g1268 );
or ( g1307 , g1305 , g1306 );
not ( g1308 , g4808 );
nand ( g1309 , g1308 , g1249 );
nand ( g1310 , g1307 , g1309 );
buf ( g1311 , g589 );
or ( g1312 , g1310 , g1311 );
nand ( g1313 , g1303 , g1312 );
or ( g1314 , g1299 , g1313 );
not ( g1315 , g1253 );
nand ( g1316 , g4676 , g653 );
not ( g1317 , g1316 );
and ( g1318 , g1315 , g1317 );
and ( g1319 , g1310 , g1311 );
nor ( g1320 , g1318 , g1319 );
nand ( g1321 , g1314 , g1320 );
or ( g1322 , g4811 , g1182 );
and ( g1323 , g1182 , g4811 );
nor ( g1324 , g1323 , g4812 );
nand ( g1325 , g1322 , g1324 );
not ( g1326 , g457 );
nor ( g1327 , g4803 , g4802 );
nand ( g1328 , g1326 , g1327 );
not ( g1329 , g558 );
nor ( g1330 , g1329 , g847 , g849 );
and ( g1331 , g1328 , g1330 );
not ( g1332 , g4802 );
nand ( g1333 , g1332 , g1326 );
and ( g1334 , g1333 , g4803 );
nor ( g1335 , g1331 , g1334 );
nand ( g1336 , g1261 , g1075 , g4791 );
or ( g1337 , g984 , g4791 );
nand ( g1338 , g1336 , g1264 , g1337 );
not ( g1339 , g1217 );
not ( g1340 , g4786 );
not ( g1341 , g864 );
or ( g1342 , g1340 , g1341 );
nand ( g1343 , g1342 , g1011 );
and ( g1344 , g4742 , g4783 );
and ( g1345 , g4791 , g653 );
not ( g1346 , g4791 );
and ( g1347 , g1346 , g1089 );
nor ( g1348 , g1345 , g1347 );
nand ( g1349 , g1278 , g1273 , g807 );
nand ( g1350 , g4787 , g4675 , g4789 );
not ( g1351 , g987 );
nand ( g1352 , g4696 , g1351 , g958 );
and ( g1353 , g4791 , g589 );
not ( g1354 , g4791 );
and ( g1355 , g1354 , g1011 );
nor ( g1356 , g1353 , g1355 );
nand ( g1357 , g4675 , g4789 );
nand ( g1358 , g4815 , g4675 , g4789 );
and ( g1359 , g1280 , g4676 );
nor ( g1360 , g1359 , g1281 );
not ( g1361 , g1360 );
not ( g1362 , g1321 );
or ( g1363 , g1361 , g1362 );
not ( g1364 , g1268 );
not ( g1365 , g1272 );
or ( g1366 , g1364 , g1365 );
nand ( g1367 , g1366 , g1349 );
nor ( g1368 , g862 , g1005 );
and ( g1369 , g1367 , g1368 );
not ( g1370 , g861 );
not ( g1371 , g1335 );
or ( g1372 , g1370 , g1371 );
nand ( g1373 , g1372 , g1259 );
and ( g1374 , g842 , g845 );
and ( g1375 , g1373 , g1374 );
nor ( g1376 , g1369 , g1375 );
nand ( g1377 , g1363 , g1376 );
endmodule

