module top ( g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 , g98 , g99 , g100 , g101 , g102 , g103 , g104 , g105 , g106 , g107 , g108 , g109 , g110 , g111 , g112 , g113 , g114 , g115 , g116 , g117 , g118 , g119 , g120 , g121 , g122 , g123 , g124 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g136 , g137 , g138 , g139 , g140 , g141 , g142 , g143 , g144 , g145 , g146 , g147 , g148 , g149 , g150 , g151 , g152 , g153 , g154 , g155 , g156 , g157 , g158 , g159 , g160 , g161 , g162 , g163 , g164 , g165 , g166 , g167 , g168 , g169 , g170 , g171 , g172 , g173 , g174 , g175 , g176 , g177 , g178 , g179 , g180 , g181 , g182 , g183 , g184 , g185 , g186 , g187 , g188 , g189 , g190 , g191 , g192 , g193 , g194 , g195 , g196 , g197 , g198 , g199 , g200 , g201 , g202 , g203 , g204 , g205 , g206 , g207 , g208 , g209 , g210 , g211 );
input g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 , g98 , g99 , g100 , g101 , g102 , g103 , g104 , g105 , g106 , g107 , g108 , g109 , g110 , g111 , g112 , g113 , g114 , g115 , g116 , g117 , g118 , g119 , g120 , g121 , g122 , g123 , g124 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g136 , g137 , g138 , g139 , g140 , g141 , g142 , g143 , g144 , g145 , g146 , g147 , g148 , g149 , g150 , g151 , g152 , g153 , g154 , g155 , g156 , g157 , g158 , g159 , g160 , g161 , g162 , g163 , g164 , g165 , g166 , g167 , g168 , g169 , g170 , g171 , g172 , g173 , g174 , g175 , g176 , g177 , g178 , g179 , g180 , g181 , g182 , g183 , g184 , g185 , g186 , g187 , g188 , g189 , g190 , g191 , g192 , g193 , g194 , g195 , g196 , g197 ;
output g198 , g199 , g200 , g201 , g202 , g203 , g204 , g205 , g206 , g207 , g208 , g209 , g210 , g211 ;

wire n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , 
     n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , 
     n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , 
     n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , 
     n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , 
     n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , 
     n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , 
     n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , 
     n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , 
     n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , 
     n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , 
     n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , 
     n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , 
     n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , 
     n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , 
     n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , 
     n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , 
     n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , 
     n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , 
     n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , 
     n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , 
     n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , 
     n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , 
     n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , 
     n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , 
     n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , 
     n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , 
     n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , 
     n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , 
     n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , 
     n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , 
     n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , 
     n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , 
     n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , 
     n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , 
     n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , 
     n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , 
     n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , 
     n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , 
     n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , 
     n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , 
     n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , 
     n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , 
     n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , 
     n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , 
     n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , 
     n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , 
     n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , 
     n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , 
     n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , 
     n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , 
     n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , 
     n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , 
     n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , 
     n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , 
     n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , 
     n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , 
     n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , 
     n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , 
     n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , 
     n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , 
     n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , 
     n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , 
     n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , 
     n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , 
     n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , 
     n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , 
     n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , 
     n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , 
     n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , 
     n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , 
     n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , 
     n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , 
     n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , 
     n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , 
     n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , 
     n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , 
     n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , 
     n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , 
     n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , 
     n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , 
     n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , 
     n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , 
     n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , 
     n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , 
     n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , 
     n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , 
     n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , 
     n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , 
     n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , 
     n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , 
     n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , 
     n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , 
     n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , 
     n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , 
     n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , 
     n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , 
     n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , 
     n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , 
     n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , 
     n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , 
     n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , 
     n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , 
     n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , 
     n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , 
     n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , 
     n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , 
     n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , 
     n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , 
     n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , 
     n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , 
     n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , 
     n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , 
     n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , 
     n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , 
     n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , 
     n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , 
     n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , 
     n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , 
     n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , 
     n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , 
     n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , 
     n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , 
     n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , 
     n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , 
     n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , 
     n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , 
     n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , 
     n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , 
     n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , 
     n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , 
     n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , 
     n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , 
     n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , 
     n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , 
     n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , 
     n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , 
     n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , 
     n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , 
     n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , 
     n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , 
     n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , 
     n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , 
     n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , 
     n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , 
     n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , 
     n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , 
     n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , 
     n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , 
     n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , 
     n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , 
     n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , 
     n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , 
     n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , 
     n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , 
     n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , 
     n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , 
     n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , 
     n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , 
     n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , 
     n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , 
     n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , 
     n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , 
     n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , 
     n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , 
     n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , 
     n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , 
     n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , 
     n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , 
     n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , 
     n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , 
     n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , 
     n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , 
     n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , 
     n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , 
     n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , 
     n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , 
     n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , 
     n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , 
     n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , 
     n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , 
     n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , 
     n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , 
     n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , 
     n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , 
     n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , 
     n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , 
     n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , 
     n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , 
     n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , 
     n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , 
     n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , 
     n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , 
     n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , 
     n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , 
     n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , 
     n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , 
     n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , 
     n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , 
     n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , 
     n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , 
     n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , 
     n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , 
     n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , 
     n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , 
     n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , 
     n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , 
     n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , 
     n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , 
     n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , 
     n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , 
     n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , 
     n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , 
     n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , 
     n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , 
     n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , 
     n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , 
     n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , 
     n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , 
     n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , 
     n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , 
     n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , 
     n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , 
     n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , 
     n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , 
     n2250 ;
buf ( n1 , g0 );
buf ( n2 , g1 );
buf ( n3 , g2 );
buf ( n4 , g3 );
buf ( n5 , g4 );
buf ( n6 , g5 );
buf ( n7 , g6 );
buf ( n8 , g7 );
buf ( n9 , g8 );
buf ( n10 , g9 );
buf ( n11 , g10 );
buf ( n12 , g11 );
buf ( n13 , g12 );
buf ( n14 , g13 );
buf ( n15 , g14 );
buf ( n16 , g15 );
buf ( n17 , g16 );
buf ( n18 , g17 );
buf ( n19 , g18 );
buf ( n20 , g19 );
buf ( n21 , g20 );
buf ( n22 , g21 );
buf ( n23 , g22 );
buf ( n24 , g23 );
buf ( n25 , g24 );
buf ( n26 , g25 );
buf ( n27 , g26 );
buf ( n28 , g27 );
buf ( n29 , g28 );
buf ( n30 , g29 );
buf ( n31 , g30 );
buf ( n32 , g31 );
buf ( n33 , g32 );
buf ( n34 , g33 );
buf ( n35 , g34 );
buf ( n36 , g35 );
buf ( n37 , g36 );
buf ( n38 , g37 );
buf ( n39 , g38 );
buf ( n40 , g39 );
buf ( n41 , g40 );
buf ( n42 , g41 );
buf ( n43 , g42 );
buf ( n44 , g43 );
buf ( n45 , g44 );
buf ( n46 , g45 );
buf ( n47 , g46 );
buf ( n48 , g47 );
buf ( n49 , g48 );
buf ( n50 , g49 );
buf ( n51 , g50 );
buf ( n52 , g51 );
buf ( n53 , g52 );
buf ( n54 , g53 );
buf ( n55 , g54 );
buf ( n56 , g55 );
buf ( n57 , g56 );
buf ( n58 , g57 );
buf ( n59 , g58 );
buf ( n60 , g59 );
buf ( n61 , g60 );
buf ( n62 , g61 );
buf ( n63 , g62 );
buf ( n64 , g63 );
buf ( n65 , g64 );
buf ( n66 , g65 );
buf ( n67 , g66 );
buf ( n68 , g67 );
buf ( n69 , g68 );
buf ( n70 , g69 );
buf ( n71 , g70 );
buf ( n72 , g71 );
buf ( n73 , g72 );
buf ( n74 , g73 );
buf ( n75 , g74 );
buf ( n76 , g75 );
buf ( n77 , g76 );
buf ( n78 , g77 );
buf ( n79 , g78 );
buf ( n80 , g79 );
buf ( n81 , g80 );
buf ( n82 , g81 );
buf ( n83 , g82 );
buf ( n84 , g83 );
buf ( n85 , g84 );
buf ( n86 , g85 );
buf ( n87 , g86 );
buf ( n88 , g87 );
buf ( n89 , g88 );
buf ( n90 , g89 );
buf ( n91 , g90 );
buf ( n92 , g91 );
buf ( n93 , g92 );
buf ( n94 , g93 );
buf ( n95 , g94 );
buf ( n96 , g95 );
buf ( n97 , g96 );
buf ( n98 , g97 );
buf ( n99 , g98 );
buf ( n100 , g99 );
buf ( n101 , g100 );
buf ( n102 , g101 );
buf ( n103 , g102 );
buf ( n104 , g103 );
buf ( n105 , g104 );
buf ( n106 , g105 );
buf ( n107 , g106 );
buf ( n108 , g107 );
buf ( n109 , g108 );
buf ( n110 , g109 );
buf ( n111 , g110 );
buf ( n112 , g111 );
buf ( n113 , g112 );
buf ( n114 , g113 );
buf ( n115 , g114 );
buf ( n116 , g115 );
buf ( n117 , g116 );
buf ( n118 , g117 );
buf ( n119 , g118 );
buf ( n120 , g119 );
buf ( n121 , g120 );
buf ( n122 , g121 );
buf ( n123 , g122 );
buf ( n124 , g123 );
buf ( n125 , g124 );
buf ( n126 , g125 );
buf ( n127 , g126 );
buf ( n128 , g127 );
buf ( n129 , g128 );
buf ( n130 , g129 );
buf ( n131 , g130 );
buf ( n132 , g131 );
buf ( n133 , g132 );
buf ( n134 , g133 );
buf ( n135 , g134 );
buf ( n136 , g135 );
buf ( n137 , g136 );
buf ( n138 , g137 );
buf ( n139 , g138 );
buf ( n140 , g139 );
buf ( n141 , g140 );
buf ( n142 , g141 );
buf ( n143 , g142 );
buf ( n144 , g143 );
buf ( n145 , g144 );
buf ( n146 , g145 );
buf ( n147 , g146 );
buf ( n148 , g147 );
buf ( n149 , g148 );
buf ( n150 , g149 );
buf ( n151 , g150 );
buf ( n152 , g151 );
buf ( n153 , g152 );
buf ( n154 , g153 );
buf ( n155 , g154 );
buf ( n156 , g155 );
buf ( n157 , g156 );
buf ( n158 , g157 );
buf ( n159 , g158 );
buf ( n160 , g159 );
buf ( n161 , g160 );
buf ( n162 , g161 );
buf ( n163 , g162 );
buf ( n164 , g163 );
buf ( n165 , g164 );
buf ( n166 , g165 );
buf ( n167 , g166 );
buf ( n168 , g167 );
buf ( n169 , g168 );
buf ( n170 , g169 );
buf ( n171 , g170 );
buf ( n172 , g171 );
buf ( n173 , g172 );
buf ( n174 , g173 );
buf ( n175 , g174 );
buf ( n176 , g175 );
buf ( n177 , g176 );
buf ( n178 , g177 );
buf ( n179 , g178 );
buf ( n180 , g179 );
buf ( n181 , g180 );
buf ( n182 , g181 );
buf ( n183 , g182 );
buf ( n184 , g183 );
buf ( n185 , g184 );
buf ( n186 , g185 );
buf ( n187 , g186 );
buf ( n188 , g187 );
buf ( n189 , g188 );
buf ( n190 , g189 );
buf ( n191 , g190 );
buf ( n192 , g191 );
buf ( n193 , g192 );
buf ( n194 , g193 );
buf ( n195 , g194 );
buf ( n196 , g195 );
buf ( n197 , g196 );
buf ( n198 , g197 );
buf ( g198 , n199 );
buf ( g199 , n200 );
buf ( g200 , n201 );
buf ( g201 , n202 );
buf ( g202 , n203 );
buf ( g203 , n204 );
buf ( g204 , n205 );
buf ( g205 , n206 );
buf ( g206 , n207 );
buf ( g207 , n208 );
buf ( g208 , n209 );
buf ( g209 , n210 );
buf ( g210 , n211 );
buf ( g211 , n212 );
buf ( n199 , n2250 );
buf ( n200 , n2248 );
buf ( n201 , n2247 );
buf ( n202 , n1582 );
buf ( n203 , n635 );
buf ( n204 , n2245 );
buf ( n205 , n2244 );
buf ( n206 , n2245 );
buf ( n207 , n2245 );
buf ( n208 , n1208 );
buf ( n209 , n67 );
buf ( n210 , n70 );
buf ( n211 , n73 );
buf ( n212 , n78 );
not ( n215 , n119 );
not ( n216 , n120 );
and ( n217 , n215 , n216 );
and ( n218 , n1 , n217 );
not ( n219 , n218 );
and ( n220 , n3 , n219 );
not ( n221 , n3 );
and ( n222 , n1 , n221 );
and ( n223 , n119 , n120 );
not ( n224 , n223 );
and ( n225 , n222 , n224 );
not ( n226 , n225 );
not ( n227 , n40 );
and ( n228 , n6 , n227 );
not ( n229 , n228 );
not ( n230 , n6 );
and ( n231 , n230 , n142 );
not ( n232 , n231 );
and ( n233 , n229 , n232 );
not ( n234 , n6 );
and ( n235 , n234 , n42 );
not ( n236 , n235 );
and ( n237 , n6 , n181 );
not ( n238 , n237 );
and ( n239 , n236 , n238 );
and ( n240 , n233 , n239 );
not ( n241 , n240 );
not ( n242 , n43 );
and ( n243 , n6 , n242 );
not ( n244 , n243 );
not ( n245 , n6 );
and ( n246 , n245 , n141 );
not ( n247 , n246 );
and ( n248 , n244 , n247 );
not ( n249 , n248 );
not ( n250 , n6 );
and ( n251 , n250 , n45 );
not ( n252 , n251 );
and ( n253 , n6 , n180 );
not ( n254 , n253 );
and ( n255 , n252 , n254 );
not ( n256 , n255 );
and ( n257 , n249 , n256 );
not ( n258 , n257 );
not ( n259 , n233 );
not ( n260 , n239 );
and ( n261 , n259 , n260 );
not ( n262 , n261 );
and ( n263 , n258 , n262 );
and ( n264 , n248 , n255 );
not ( n265 , n264 );
not ( n266 , n46 );
and ( n267 , n6 , n266 );
not ( n268 , n267 );
not ( n269 , n6 );
and ( n270 , n269 , n140 );
not ( n271 , n270 );
and ( n272 , n268 , n271 );
not ( n273 , n272 );
not ( n274 , n6 );
and ( n275 , n274 , n48 );
not ( n276 , n275 );
and ( n277 , n6 , n179 );
not ( n278 , n277 );
and ( n279 , n276 , n278 );
not ( n280 , n279 );
and ( n281 , n273 , n280 );
not ( n282 , n281 );
not ( n283 , n51 );
and ( n284 , n6 , n283 );
not ( n285 , n284 );
not ( n286 , n6 );
and ( n287 , n286 , n139 );
not ( n288 , n287 );
and ( n289 , n285 , n288 );
not ( n290 , n6 );
and ( n291 , n290 , n50 );
not ( n292 , n291 );
and ( n293 , n6 , n178 );
not ( n294 , n293 );
and ( n295 , n292 , n294 );
and ( n296 , n289 , n295 );
not ( n297 , n296 );
and ( n298 , n272 , n279 );
not ( n299 , n298 );
and ( n300 , n297 , n299 );
not ( n301 , n289 );
not ( n302 , n295 );
and ( n303 , n301 , n302 );
not ( n304 , n303 );
not ( n305 , n52 );
and ( n306 , n6 , n305 );
not ( n307 , n306 );
not ( n308 , n6 );
and ( n309 , n308 , n149 );
not ( n310 , n309 );
and ( n311 , n307 , n310 );
not ( n312 , n6 );
and ( n313 , n312 , n54 );
not ( n314 , n313 );
and ( n315 , n6 , n187 );
not ( n316 , n315 );
and ( n317 , n314 , n316 );
and ( n318 , n311 , n317 );
not ( n319 , n318 );
not ( n320 , n311 );
not ( n321 , n317 );
and ( n322 , n320 , n321 );
not ( n323 , n322 );
not ( n324 , n55 );
and ( n325 , n6 , n324 );
not ( n326 , n325 );
not ( n327 , n6 );
and ( n328 , n327 , n148 );
not ( n329 , n328 );
and ( n330 , n326 , n329 );
not ( n331 , n330 );
not ( n332 , n6 );
and ( n333 , n332 , n57 );
not ( n334 , n333 );
and ( n335 , n6 , n186 );
not ( n336 , n335 );
and ( n337 , n334 , n336 );
not ( n338 , n337 );
and ( n339 , n331 , n338 );
not ( n340 , n339 );
and ( n341 , n323 , n340 );
not ( n342 , n58 );
and ( n343 , n6 , n342 );
not ( n344 , n343 );
not ( n345 , n6 );
and ( n346 , n345 , n147 );
not ( n347 , n346 );
and ( n348 , n344 , n347 );
not ( n349 , n6 );
and ( n350 , n349 , n60 );
not ( n351 , n350 );
and ( n352 , n6 , n185 );
not ( n353 , n352 );
and ( n354 , n351 , n353 );
and ( n355 , n348 , n354 );
not ( n356 , n355 );
and ( n357 , n330 , n337 );
not ( n358 , n357 );
and ( n359 , n356 , n358 );
not ( n360 , n348 );
not ( n361 , n354 );
and ( n362 , n360 , n361 );
not ( n363 , n362 );
not ( n364 , n61 );
and ( n365 , n6 , n364 );
not ( n366 , n365 );
not ( n367 , n6 );
and ( n368 , n367 , n146 );
not ( n369 , n368 );
and ( n370 , n366 , n369 );
not ( n371 , n370 );
not ( n372 , n6 );
and ( n373 , n372 , n63 );
not ( n374 , n373 );
and ( n375 , n6 , n184 );
not ( n376 , n375 );
and ( n377 , n374 , n376 );
not ( n378 , n377 );
and ( n379 , n371 , n378 );
not ( n380 , n379 );
and ( n381 , n363 , n380 );
not ( n382 , n64 );
and ( n383 , n6 , n382 );
not ( n384 , n383 );
not ( n385 , n6 );
and ( n386 , n385 , n145 );
not ( n387 , n386 );
and ( n388 , n384 , n387 );
not ( n389 , n388 );
not ( n390 , n6 );
and ( n391 , n390 , n66 );
not ( n392 , n391 );
and ( n393 , n6 , n183 );
not ( n394 , n393 );
and ( n395 , n392 , n394 );
not ( n396 , n395 );
and ( n397 , n389 , n396 );
and ( n398 , n370 , n377 );
not ( n399 , n398 );
and ( n400 , n397 , n399 );
not ( n401 , n400 );
and ( n402 , n381 , n401 );
not ( n403 , n402 );
and ( n404 , n359 , n403 );
not ( n405 , n404 );
and ( n406 , n341 , n405 );
not ( n407 , n406 );
and ( n408 , n319 , n407 );
not ( n409 , n408 );
and ( n410 , n304 , n409 );
not ( n411 , n410 );
and ( n412 , n300 , n411 );
not ( n413 , n412 );
and ( n414 , n282 , n413 );
not ( n415 , n414 );
and ( n416 , n265 , n415 );
not ( n417 , n416 );
and ( n418 , n263 , n417 );
not ( n419 , n418 );
and ( n420 , n241 , n419 );
not ( n421 , n156 );
not ( n422 , n6 );
not ( n423 , n93 );
and ( n424 , n422 , n423 );
and ( n425 , n421 , n424 );
not ( n426 , n425 );
and ( n427 , n198 , n426 );
not ( n428 , n427 );
not ( n429 , n88 );
and ( n430 , n6 , n429 );
not ( n431 , n430 );
not ( n432 , n6 );
and ( n433 , n432 , n157 );
not ( n434 , n433 );
and ( n435 , n431 , n434 );
not ( n436 , n435 );
not ( n437 , n6 );
and ( n438 , n437 , n90 );
not ( n439 , n438 );
and ( n440 , n6 , n194 );
not ( n441 , n440 );
and ( n442 , n439 , n441 );
not ( n443 , n442 );
and ( n444 , n436 , n443 );
not ( n445 , n444 );
not ( n446 , n6 );
and ( n447 , n446 , n156 );
and ( n448 , n93 , n447 );
not ( n449 , n448 );
and ( n450 , n445 , n449 );
and ( n451 , n428 , n450 );
not ( n452 , n451 );
not ( n453 , n85 );
and ( n454 , n6 , n453 );
not ( n455 , n454 );
not ( n456 , n6 );
and ( n457 , n456 , n158 );
not ( n458 , n457 );
and ( n459 , n455 , n458 );
not ( n460 , n6 );
and ( n461 , n460 , n87 );
not ( n462 , n461 );
and ( n463 , n6 , n195 );
not ( n464 , n463 );
and ( n465 , n462 , n464 );
and ( n466 , n459 , n465 );
not ( n467 , n466 );
and ( n468 , n435 , n442 );
not ( n469 , n468 );
and ( n470 , n467 , n469 );
and ( n471 , n452 , n470 );
not ( n472 , n471 );
not ( n473 , n459 );
not ( n474 , n465 );
and ( n475 , n473 , n474 );
not ( n476 , n475 );
not ( n477 , n82 );
and ( n478 , n6 , n477 );
not ( n479 , n478 );
not ( n480 , n6 );
and ( n481 , n480 , n159 );
not ( n482 , n481 );
and ( n483 , n479 , n482 );
not ( n484 , n483 );
not ( n485 , n6 );
and ( n486 , n485 , n84 );
not ( n487 , n486 );
and ( n488 , n6 , n196 );
not ( n489 , n488 );
and ( n490 , n487 , n489 );
not ( n491 , n490 );
and ( n492 , n484 , n491 );
not ( n493 , n492 );
and ( n494 , n476 , n493 );
and ( n495 , n472 , n494 );
not ( n496 , n495 );
and ( n497 , n483 , n490 );
not ( n498 , n497 );
not ( n499 , n79 );
and ( n500 , n6 , n499 );
not ( n501 , n500 );
not ( n502 , n6 );
and ( n503 , n502 , n160 );
not ( n504 , n503 );
and ( n505 , n501 , n504 );
not ( n506 , n6 );
and ( n507 , n506 , n81 );
not ( n508 , n507 );
and ( n509 , n6 , n197 );
not ( n510 , n509 );
and ( n511 , n508 , n510 );
and ( n512 , n505 , n511 );
not ( n513 , n512 );
and ( n514 , n498 , n513 );
and ( n515 , n496 , n514 );
not ( n516 , n515 );
not ( n517 , n78 );
and ( n518 , n6 , n517 );
not ( n519 , n518 );
not ( n520 , n6 );
and ( n521 , n520 , n150 );
not ( n522 , n521 );
and ( n523 , n519 , n522 );
not ( n524 , n523 );
not ( n525 , n6 );
and ( n526 , n525 , n77 );
not ( n527 , n526 );
and ( n528 , n6 , n188 );
not ( n529 , n528 );
and ( n530 , n527 , n529 );
not ( n531 , n530 );
and ( n532 , n524 , n531 );
not ( n533 , n532 );
not ( n534 , n505 );
not ( n535 , n511 );
and ( n536 , n534 , n535 );
not ( n537 , n536 );
and ( n538 , n533 , n537 );
and ( n539 , n516 , n538 );
not ( n540 , n539 );
and ( n541 , n523 , n530 );
not ( n542 , n541 );
not ( n543 , n73 );
and ( n544 , n6 , n543 );
not ( n545 , n544 );
not ( n546 , n6 );
and ( n547 , n546 , n151 );
not ( n548 , n547 );
and ( n549 , n545 , n548 );
not ( n550 , n549 );
not ( n551 , n6 );
and ( n552 , n551 , n75 );
not ( n553 , n552 );
and ( n554 , n6 , n189 );
not ( n555 , n554 );
and ( n556 , n553 , n555 );
not ( n557 , n556 );
and ( n558 , n550 , n557 );
not ( n559 , n558 );
and ( n560 , n542 , n559 );
not ( n561 , n70 );
and ( n562 , n6 , n561 );
not ( n563 , n562 );
not ( n564 , n6 );
and ( n565 , n564 , n152 );
not ( n566 , n565 );
and ( n567 , n563 , n566 );
not ( n568 , n6 );
and ( n569 , n568 , n72 );
not ( n570 , n569 );
and ( n571 , n6 , n190 );
not ( n572 , n571 );
and ( n573 , n570 , n572 );
and ( n574 , n567 , n573 );
not ( n575 , n574 );
and ( n576 , n549 , n556 );
not ( n577 , n576 );
and ( n578 , n575 , n577 );
and ( n579 , n560 , n578 );
and ( n580 , n540 , n579 );
not ( n581 , n580 );
not ( n582 , n574 );
and ( n583 , n558 , n582 );
not ( n584 , n583 );
not ( n585 , n567 );
not ( n586 , n573 );
and ( n587 , n585 , n586 );
not ( n588 , n587 );
not ( n589 , n67 );
and ( n590 , n6 , n589 );
not ( n591 , n590 );
not ( n592 , n6 );
and ( n593 , n592 , n153 );
not ( n594 , n593 );
and ( n595 , n591 , n594 );
not ( n596 , n595 );
not ( n597 , n6 );
and ( n598 , n597 , n69 );
not ( n599 , n598 );
and ( n600 , n6 , n191 );
not ( n601 , n600 );
and ( n602 , n599 , n601 );
not ( n603 , n602 );
and ( n604 , n596 , n603 );
not ( n605 , n604 );
and ( n606 , n588 , n605 );
and ( n607 , n584 , n606 );
and ( n608 , n581 , n607 );
not ( n609 , n608 );
and ( n610 , n300 , n341 );
and ( n611 , n359 , n381 );
and ( n612 , n610 , n611 );
and ( n613 , n388 , n395 );
not ( n614 , n613 );
not ( n615 , n398 );
and ( n616 , n595 , n602 );
not ( n617 , n616 );
and ( n618 , n615 , n617 );
and ( n619 , n614 , n618 );
not ( n620 , n281 );
not ( n621 , n303 );
and ( n622 , n620 , n621 );
not ( n623 , n318 );
not ( n624 , n397 );
and ( n625 , n623 , n624 );
and ( n626 , n622 , n625 );
not ( n627 , n240 );
not ( n628 , n264 );
and ( n629 , n627 , n628 );
and ( n630 , n263 , n629 );
and ( n631 , n626 , n630 );
and ( n632 , n619 , n631 );
and ( n633 , n612 , n632 );
and ( n634 , n609 , n633 );
or ( n635 , n420 , n634 );
not ( n636 , n6 );
and ( n637 , n636 , n136 );
not ( n638 , n637 );
not ( n639 , n31 );
and ( n640 , n6 , n639 );
not ( n641 , n640 );
and ( n642 , n638 , n641 );
not ( n643 , n642 );
not ( n644 , n6 );
and ( n645 , n644 , n32 );
not ( n646 , n645 );
and ( n647 , n6 , n175 );
not ( n648 , n647 );
and ( n649 , n646 , n648 );
not ( n650 , n649 );
and ( n651 , n643 , n650 );
not ( n652 , n651 );
not ( n653 , n6 );
and ( n654 , n653 , n135 );
not ( n655 , n654 );
not ( n656 , n34 );
and ( n657 , n6 , n656 );
not ( n658 , n657 );
and ( n659 , n655 , n658 );
not ( n660 , n6 );
and ( n661 , n660 , n35 );
not ( n662 , n661 );
and ( n663 , n6 , n174 );
not ( n664 , n663 );
and ( n665 , n662 , n664 );
and ( n666 , n659 , n665 );
not ( n667 , n666 );
and ( n668 , n642 , n649 );
not ( n669 , n668 );
and ( n670 , n667 , n669 );
not ( n671 , n6 );
and ( n672 , n671 , n134 );
not ( n673 , n672 );
not ( n674 , n37 );
and ( n675 , n6 , n674 );
not ( n676 , n675 );
and ( n677 , n673 , n676 );
not ( n678 , n677 );
not ( n679 , n6 );
and ( n680 , n679 , n38 );
not ( n681 , n680 );
and ( n682 , n6 , n173 );
not ( n683 , n682 );
and ( n684 , n681 , n683 );
not ( n685 , n684 );
and ( n686 , n678 , n685 );
not ( n687 , n686 );
not ( n688 , n659 );
not ( n689 , n665 );
and ( n690 , n688 , n689 );
not ( n691 , n690 );
and ( n692 , n687 , n691 );
not ( n693 , n692 );
and ( n694 , n670 , n693 );
not ( n695 , n694 );
and ( n696 , n652 , n695 );
not ( n697 , n6 );
and ( n698 , n697 , n130 );
not ( n699 , n698 );
not ( n700 , n20 );
and ( n701 , n6 , n700 );
not ( n702 , n701 );
and ( n703 , n699 , n702 );
not ( n704 , n703 );
and ( n705 , n8 , n9 );
not ( n706 , n705 );
not ( n707 , n170 );
and ( n708 , n6 , n707 );
not ( n709 , n708 );
and ( n710 , n706 , n709 );
and ( n711 , n704 , n710 );
not ( n712 , n711 );
not ( n713 , n6 );
and ( n714 , n713 , n129 );
not ( n715 , n714 );
not ( n716 , n22 );
and ( n717 , n6 , n716 );
not ( n718 , n717 );
and ( n719 , n715 , n718 );
not ( n720 , n719 );
not ( n721 , n705 );
not ( n722 , n169 );
and ( n723 , n6 , n722 );
not ( n724 , n723 );
and ( n725 , n721 , n724 );
and ( n726 , n720 , n725 );
not ( n727 , n726 );
and ( n728 , n712 , n727 );
not ( n729 , n6 );
and ( n730 , n729 , n138 );
not ( n731 , n730 );
not ( n732 , n26 );
and ( n733 , n6 , n732 );
not ( n734 , n733 );
and ( n735 , n731 , n734 );
not ( n736 , n705 );
not ( n737 , n177 );
and ( n738 , n6 , n737 );
not ( n739 , n738 );
and ( n740 , n736 , n739 );
not ( n741 , n740 );
and ( n742 , n735 , n741 );
not ( n743 , n742 );
not ( n744 , n6 );
and ( n745 , n744 , n128 );
not ( n746 , n745 );
not ( n747 , n25 );
and ( n748 , n6 , n747 );
not ( n749 , n748 );
and ( n750 , n746 , n749 );
not ( n751 , n705 );
not ( n752 , n168 );
and ( n753 , n6 , n752 );
not ( n754 , n753 );
and ( n755 , n751 , n754 );
not ( n756 , n755 );
and ( n757 , n750 , n756 );
not ( n758 , n757 );
and ( n759 , n743 , n758 );
and ( n760 , n728 , n759 );
not ( n761 , n735 );
and ( n762 , n761 , n740 );
not ( n763 , n762 );
not ( n764 , n6 );
and ( n765 , n764 , n137 );
not ( n766 , n765 );
not ( n767 , n28 );
and ( n768 , n6 , n767 );
not ( n769 , n768 );
and ( n770 , n766 , n769 );
not ( n771 , n770 );
not ( n772 , n6 );
and ( n773 , n772 , n29 );
not ( n774 , n773 );
and ( n775 , n6 , n176 );
not ( n776 , n775 );
and ( n777 , n774 , n776 );
not ( n778 , n777 );
and ( n779 , n771 , n778 );
not ( n780 , n779 );
and ( n781 , n763 , n780 );
and ( n782 , n781 , n670 );
and ( n783 , n760 , n782 );
and ( n784 , n677 , n684 );
not ( n785 , n784 );
not ( n786 , n750 );
and ( n787 , n786 , n755 );
not ( n788 , n787 );
and ( n789 , n770 , n777 );
not ( n790 , n789 );
and ( n791 , n788 , n790 );
and ( n792 , n785 , n791 );
not ( n793 , n710 );
and ( n794 , n703 , n793 );
not ( n795 , n794 );
not ( n796 , n6 );
and ( n797 , n796 , n131 );
not ( n798 , n797 );
not ( n799 , n18 );
and ( n800 , n6 , n799 );
not ( n801 , n800 );
and ( n802 , n798 , n801 );
not ( n803 , n705 );
not ( n804 , n171 );
and ( n805 , n6 , n804 );
not ( n806 , n805 );
and ( n807 , n803 , n806 );
not ( n808 , n807 );
and ( n809 , n802 , n808 );
not ( n810 , n809 );
and ( n811 , n795 , n810 );
not ( n812 , n802 );
and ( n813 , n812 , n807 );
not ( n814 , n813 );
not ( n815 , n725 );
and ( n816 , n719 , n815 );
not ( n817 , n816 );
and ( n818 , n814 , n817 );
and ( n819 , n811 , n818 );
and ( n820 , n792 , n819 );
and ( n821 , n783 , n820 );
and ( n822 , n696 , n821 );
and ( n823 , n635 , n822 );
not ( n824 , n823 );
not ( n825 , n813 );
not ( n826 , n816 );
not ( n827 , n787 );
not ( n828 , n696 );
not ( n829 , n789 );
and ( n830 , n828 , n829 );
not ( n831 , n830 );
and ( n832 , n781 , n831 );
not ( n833 , n832 );
and ( n834 , n759 , n833 );
not ( n835 , n834 );
and ( n836 , n827 , n835 );
not ( n837 , n836 );
and ( n838 , n826 , n837 );
not ( n839 , n838 );
and ( n840 , n728 , n839 );
not ( n841 , n840 );
and ( n842 , n811 , n841 );
not ( n843 , n842 );
and ( n844 , n825 , n843 );
and ( n845 , n824 , n844 );
not ( n846 , n845 );
not ( n847 , n705 );
not ( n848 , n6 );
and ( n849 , n848 , n123 );
not ( n850 , n849 );
not ( n851 , n16 );
and ( n852 , n6 , n851 );
not ( n853 , n852 );
and ( n854 , n850 , n853 );
not ( n855 , n6 );
and ( n856 , n855 , n124 );
not ( n857 , n856 );
not ( n858 , n14 );
and ( n859 , n6 , n858 );
not ( n860 , n859 );
and ( n861 , n857 , n860 );
not ( n862 , n861 );
not ( n863 , n164 );
and ( n864 , n6 , n863 );
not ( n865 , n864 );
and ( n866 , n862 , n865 );
not ( n867 , n866 );
and ( n868 , n854 , n867 );
not ( n869 , n868 );
and ( n870 , n847 , n869 );
not ( n871 , n870 );
not ( n872 , n6 );
and ( n873 , n872 , n126 );
not ( n874 , n873 );
not ( n875 , n10 );
and ( n876 , n6 , n875 );
not ( n877 , n876 );
and ( n878 , n874 , n877 );
not ( n879 , n878 );
not ( n880 , n705 );
not ( n881 , n166 );
and ( n882 , n6 , n881 );
not ( n883 , n882 );
and ( n884 , n880 , n883 );
and ( n885 , n879 , n884 );
not ( n886 , n885 );
not ( n887 , n6 );
and ( n888 , n887 , n125 );
not ( n889 , n888 );
not ( n890 , n12 );
and ( n891 , n6 , n890 );
not ( n892 , n891 );
and ( n893 , n889 , n892 );
not ( n894 , n893 );
not ( n895 , n705 );
not ( n896 , n165 );
and ( n897 , n6 , n896 );
not ( n898 , n897 );
and ( n899 , n895 , n898 );
and ( n900 , n894 , n899 );
not ( n901 , n900 );
and ( n902 , n886 , n901 );
not ( n903 , n6 );
and ( n904 , n903 , n127 );
not ( n905 , n904 );
not ( n906 , n5 );
and ( n907 , n906 , n6 );
not ( n908 , n907 );
and ( n909 , n905 , n908 );
not ( n910 , n909 );
not ( n911 , n705 );
not ( n912 , n167 );
and ( n913 , n6 , n912 );
not ( n914 , n913 );
and ( n915 , n911 , n914 );
and ( n916 , n910 , n915 );
not ( n917 , n916 );
and ( n918 , n705 , n854 );
not ( n919 , n918 );
and ( n920 , n917 , n919 );
and ( n921 , n902 , n920 );
not ( n922 , n899 );
and ( n923 , n893 , n922 );
not ( n924 , n923 );
not ( n925 , n705 );
not ( n926 , n864 );
and ( n927 , n925 , n926 );
not ( n928 , n927 );
and ( n929 , n861 , n928 );
not ( n930 , n929 );
and ( n931 , n924 , n930 );
not ( n932 , n884 );
and ( n933 , n878 , n932 );
not ( n934 , n933 );
not ( n935 , n915 );
and ( n936 , n909 , n935 );
not ( n937 , n936 );
and ( n938 , n934 , n937 );
and ( n939 , n931 , n938 );
and ( n940 , n921 , n939 );
and ( n941 , n871 , n940 );
and ( n942 , n846 , n941 );
not ( n943 , n942 );
not ( n944 , n916 );
and ( n945 , n931 , n870 );
not ( n946 , n945 );
and ( n947 , n902 , n946 );
not ( n948 , n947 );
and ( n949 , n938 , n948 );
not ( n950 , n949 );
and ( n951 , n944 , n950 );
and ( n952 , n943 , n951 );
not ( n953 , n952 );
and ( n954 , n226 , n953 );
not ( n955 , n255 );
and ( n956 , n317 , n955 );
not ( n957 , n956 );
not ( n958 , n317 );
and ( n959 , n958 , n255 );
not ( n960 , n959 );
and ( n961 , n957 , n960 );
and ( n962 , n395 , n961 );
not ( n963 , n962 );
not ( n964 , n395 );
not ( n965 , n961 );
and ( n966 , n964 , n965 );
not ( n967 , n966 );
and ( n968 , n963 , n967 );
not ( n969 , n968 );
and ( n970 , n295 , n969 );
not ( n971 , n970 );
not ( n972 , n295 );
and ( n973 , n972 , n968 );
not ( n974 , n973 );
and ( n975 , n971 , n974 );
and ( n976 , n279 , n975 );
not ( n977 , n976 );
not ( n978 , n279 );
not ( n979 , n975 );
and ( n980 , n978 , n979 );
not ( n981 , n980 );
and ( n982 , n977 , n981 );
not ( n983 , n982 );
and ( n984 , n354 , n983 );
not ( n985 , n984 );
not ( n986 , n354 );
and ( n987 , n986 , n982 );
not ( n988 , n987 );
and ( n989 , n985 , n988 );
not ( n990 , n6 );
and ( n991 , n990 , n116 );
not ( n992 , n991 );
and ( n993 , n6 , n182 );
not ( n994 , n993 );
and ( n995 , n992 , n994 );
not ( n996 , n377 );
and ( n997 , n337 , n996 );
not ( n998 , n997 );
not ( n999 , n337 );
and ( n1000 , n999 , n377 );
not ( n1001 , n1000 );
and ( n1002 , n998 , n1001 );
and ( n1003 , n995 , n1002 );
not ( n1004 , n1003 );
not ( n1005 , n995 );
not ( n1006 , n1002 );
and ( n1007 , n1005 , n1006 );
not ( n1008 , n1007 );
and ( n1009 , n1004 , n1008 );
not ( n1010 , n1009 );
and ( n1011 , n239 , n1010 );
not ( n1012 , n1011 );
not ( n1013 , n239 );
and ( n1014 , n1013 , n1009 );
not ( n1015 , n1014 );
and ( n1016 , n1012 , n1015 );
and ( n1017 , n989 , n1016 );
not ( n1018 , n1017 );
not ( n1019 , n989 );
not ( n1020 , n1016 );
and ( n1021 , n1019 , n1020 );
not ( n1022 , n1021 );
and ( n1023 , n1018 , n1022 );
and ( n1024 , n710 , n805 );
not ( n1025 , n1024 );
and ( n1026 , n708 , n807 );
not ( n1027 , n1026 );
and ( n1028 , n1025 , n1027 );
not ( n1029 , n1028 );
and ( n1030 , n777 , n1029 );
not ( n1031 , n1030 );
not ( n1032 , n777 );
and ( n1033 , n1032 , n1028 );
not ( n1034 , n1033 );
and ( n1035 , n1031 , n1034 );
not ( n1036 , n6 );
and ( n1037 , n1036 , n113 );
not ( n1038 , n1037 );
and ( n1039 , n6 , n172 );
not ( n1040 , n1039 );
and ( n1041 , n1038 , n1040 );
not ( n1042 , n1041 );
and ( n1043 , n649 , n1042 );
not ( n1044 , n1043 );
not ( n1045 , n649 );
and ( n1046 , n1045 , n1041 );
not ( n1047 , n1046 );
and ( n1048 , n1044 , n1047 );
and ( n1049 , n755 , n723 );
not ( n1050 , n1049 );
and ( n1051 , n753 , n725 );
not ( n1052 , n1051 );
and ( n1053 , n1050 , n1052 );
not ( n1054 , n1053 );
and ( n1055 , n740 , n1054 );
not ( n1056 , n1055 );
not ( n1057 , n740 );
and ( n1058 , n1057 , n1053 );
not ( n1059 , n1058 );
and ( n1060 , n1056 , n1059 );
and ( n1061 , n1060 , n665 );
not ( n1062 , n1061 );
not ( n1063 , n1060 );
not ( n1064 , n665 );
and ( n1065 , n1063 , n1064 );
not ( n1066 , n1065 );
and ( n1067 , n1062 , n1066 );
not ( n1068 , n1067 );
and ( n1069 , n1048 , n1068 );
not ( n1070 , n1069 );
not ( n1071 , n1048 );
and ( n1072 , n1071 , n1067 );
not ( n1073 , n1072 );
and ( n1074 , n1070 , n1073 );
and ( n1075 , n684 , n1074 );
not ( n1076 , n1075 );
not ( n1077 , n684 );
not ( n1078 , n1074 );
and ( n1079 , n1077 , n1078 );
not ( n1080 , n1079 );
and ( n1081 , n1076 , n1080 );
not ( n1082 , n1081 );
and ( n1083 , n1035 , n1082 );
not ( n1084 , n1083 );
not ( n1085 , n1035 );
and ( n1086 , n1085 , n1081 );
not ( n1087 , n1086 );
not ( n1088 , n442 );
and ( n1089 , n556 , n1088 );
not ( n1090 , n1089 );
not ( n1091 , n556 );
and ( n1092 , n1091 , n442 );
not ( n1093 , n1092 );
and ( n1094 , n1090 , n1093 );
not ( n1095 , n490 );
and ( n1096 , n602 , n1095 );
not ( n1097 , n1096 );
not ( n1098 , n602 );
and ( n1099 , n1098 , n490 );
not ( n1100 , n1099 );
and ( n1101 , n1097 , n1100 );
not ( n1102 , n6 );
and ( n1103 , n1102 , n118 );
not ( n1104 , n1103 );
and ( n1105 , n6 , n192 );
not ( n1106 , n1105 );
and ( n1107 , n1104 , n1106 );
not ( n1108 , n1107 );
and ( n1109 , n573 , n1108 );
not ( n1110 , n1109 );
not ( n1111 , n573 );
and ( n1112 , n1111 , n1107 );
not ( n1113 , n1112 );
and ( n1114 , n1110 , n1113 );
and ( n1115 , n1101 , n1114 );
not ( n1116 , n1115 );
not ( n1117 , n1101 );
not ( n1118 , n1114 );
and ( n1119 , n1117 , n1118 );
not ( n1120 , n1119 );
and ( n1121 , n1116 , n1120 );
not ( n1122 , n424 );
not ( n1123 , n193 );
and ( n1124 , n6 , n1123 );
not ( n1125 , n1124 );
and ( n1126 , n1122 , n1125 );
not ( n1127 , n511 );
and ( n1128 , n1126 , n1127 );
not ( n1129 , n1128 );
not ( n1130 , n1126 );
and ( n1131 , n1130 , n511 );
not ( n1132 , n1131 );
and ( n1133 , n1129 , n1132 );
not ( n1134 , n1133 );
and ( n1135 , n1121 , n1134 );
not ( n1136 , n1135 );
not ( n1137 , n1121 );
and ( n1138 , n1137 , n1133 );
not ( n1139 , n1138 );
and ( n1140 , n1136 , n1139 );
and ( n1141 , n1094 , n1140 );
not ( n1142 , n1141 );
not ( n1143 , n1094 );
not ( n1144 , n1140 );
and ( n1145 , n1143 , n1144 );
not ( n1146 , n1145 );
and ( n1147 , n1142 , n1146 );
not ( n1148 , n530 );
and ( n1149 , n465 , n1148 );
not ( n1150 , n1149 );
not ( n1151 , n465 );
and ( n1152 , n1151 , n530 );
not ( n1153 , n1152 );
and ( n1154 , n1150 , n1153 );
not ( n1155 , n1154 );
and ( n1156 , n1147 , n1155 );
not ( n1157 , n1156 );
and ( n1158 , n884 , n913 );
not ( n1159 , n1158 );
and ( n1160 , n882 , n915 );
not ( n1161 , n1160 );
and ( n1162 , n1159 , n1161 );
not ( n1163 , n1162 );
and ( n1164 , n927 , n897 );
not ( n1165 , n1164 );
and ( n1166 , n864 , n899 );
not ( n1167 , n1166 );
and ( n1168 , n1165 , n1167 );
not ( n1169 , n1168 );
not ( n1170 , n163 );
not ( n1171 , n161 );
not ( n1172 , n162 );
and ( n1173 , n1171 , n1172 );
not ( n1174 , n1173 );
and ( n1175 , n161 , n162 );
not ( n1176 , n1175 );
and ( n1177 , n1174 , n1176 );
and ( n1178 , n1170 , n1177 );
not ( n1179 , n1178 );
not ( n1180 , n705 );
and ( n1181 , n6 , n1180 );
not ( n1182 , n1177 );
and ( n1183 , n163 , n1182 );
not ( n1184 , n1183 );
and ( n1185 , n1181 , n1184 );
and ( n1186 , n1179 , n1185 );
and ( n1187 , n1169 , n1186 );
not ( n1188 , n1187 );
not ( n1189 , n1186 );
and ( n1190 , n1168 , n1189 );
not ( n1191 , n1190 );
and ( n1192 , n1188 , n1191 );
and ( n1193 , n1163 , n1192 );
not ( n1194 , n1193 );
not ( n1195 , n1192 );
and ( n1196 , n1162 , n1195 );
not ( n1197 , n1196 );
and ( n1198 , n1194 , n1197 );
not ( n1199 , n1198 );
not ( n1200 , n1147 );
and ( n1201 , n1200 , n1154 );
not ( n1202 , n1201 );
and ( n1203 , n1199 , n1202 );
and ( n1204 , n1157 , n1203 );
and ( n1205 , n1087 , n1204 );
and ( n1206 , n1084 , n1205 );
not ( n1207 , n1206 );
or ( n1208 , n1023 , n1207 );
not ( n1209 , n1208 );
not ( n1210 , n1037 );
and ( n1211 , n6 , n114 );
not ( n1212 , n1211 );
and ( n1213 , n1210 , n1212 );
not ( n1214 , n705 );
not ( n1215 , n27 );
and ( n1216 , n6 , n1215 );
and ( n1217 , n1214 , n1216 );
not ( n1218 , n705 );
not ( n1219 , n21 );
and ( n1220 , n6 , n1219 );
not ( n1221 , n1220 );
and ( n1222 , n1218 , n1221 );
not ( n1223 , n19 );
and ( n1224 , n6 , n1223 );
not ( n1225 , n1224 );
and ( n1226 , n1222 , n1225 );
not ( n1227 , n1226 );
not ( n1228 , n21 );
not ( n1229 , n705 );
and ( n1230 , n1229 , n1224 );
and ( n1231 , n1228 , n1230 );
not ( n1232 , n1231 );
and ( n1233 , n1227 , n1232 );
not ( n1234 , n1233 );
and ( n1235 , n1217 , n1234 );
not ( n1236 , n1235 );
not ( n1237 , n1217 );
and ( n1238 , n1237 , n1233 );
not ( n1239 , n1238 );
and ( n1240 , n1236 , n1239 );
and ( n1241 , n1213 , n1240 );
not ( n1242 , n1241 );
not ( n1243 , n1213 );
not ( n1244 , n1240 );
and ( n1245 , n1243 , n1244 );
not ( n1246 , n1245 );
and ( n1247 , n1242 , n1246 );
not ( n1248 , n680 );
and ( n1249 , n6 , n39 );
not ( n1250 , n1249 );
and ( n1251 , n1248 , n1250 );
not ( n1252 , n661 );
and ( n1253 , n6 , n36 );
not ( n1254 , n1253 );
and ( n1255 , n1252 , n1254 );
not ( n1256 , n645 );
and ( n1257 , n6 , n33 );
not ( n1258 , n1257 );
and ( n1259 , n1256 , n1258 );
not ( n1260 , n773 );
and ( n1261 , n6 , n30 );
not ( n1262 , n1261 );
and ( n1263 , n1260 , n1262 );
not ( n1264 , n23 );
and ( n1265 , n6 , n1264 );
not ( n1266 , n705 );
not ( n1267 , n24 );
and ( n1268 , n6 , n1267 );
not ( n1269 , n1268 );
and ( n1270 , n1266 , n1269 );
and ( n1271 , n1265 , n1270 );
not ( n1272 , n1271 );
not ( n1273 , n705 );
not ( n1274 , n1265 );
and ( n1275 , n1273 , n1274 );
and ( n1276 , n1275 , n1268 );
not ( n1277 , n1276 );
and ( n1278 , n1272 , n1277 );
not ( n1279 , n1278 );
and ( n1280 , n1263 , n1279 );
not ( n1281 , n1280 );
not ( n1282 , n1263 );
and ( n1283 , n1282 , n1278 );
not ( n1284 , n1283 );
and ( n1285 , n1281 , n1284 );
and ( n1286 , n1259 , n1285 );
not ( n1287 , n1286 );
not ( n1288 , n1259 );
not ( n1289 , n1285 );
and ( n1290 , n1288 , n1289 );
not ( n1291 , n1290 );
and ( n1292 , n1287 , n1291 );
not ( n1293 , n1292 );
and ( n1294 , n1255 , n1293 );
not ( n1295 , n1294 );
not ( n1296 , n1255 );
and ( n1297 , n1296 , n1292 );
not ( n1298 , n1297 );
and ( n1299 , n1295 , n1298 );
and ( n1300 , n1251 , n1299 );
not ( n1301 , n1300 );
not ( n1302 , n1251 );
not ( n1303 , n1299 );
and ( n1304 , n1302 , n1303 );
not ( n1305 , n1304 );
and ( n1306 , n1301 , n1305 );
and ( n1307 , n1247 , n1306 );
not ( n1308 , n1307 );
not ( n1309 , n1247 );
not ( n1310 , n1306 );
and ( n1311 , n1309 , n1310 );
not ( n1312 , n1311 );
and ( n1313 , n111 , n112 );
not ( n1314 , n1313 );
not ( n1315 , n111 );
not ( n1316 , n112 );
and ( n1317 , n1315 , n1316 );
not ( n1318 , n1317 );
and ( n1319 , n1314 , n1318 );
and ( n1320 , n1181 , n1319 );
not ( n1321 , n11 );
and ( n1322 , n6 , n1321 );
not ( n1323 , n15 );
and ( n1324 , n6 , n1323 );
not ( n1325 , n1324 );
and ( n1326 , n1322 , n1325 );
not ( n1327 , n1326 );
not ( n1328 , n1322 );
and ( n1329 , n1328 , n1324 );
not ( n1330 , n1329 );
and ( n1331 , n1327 , n1330 );
not ( n1332 , n13 );
and ( n1333 , n6 , n1332 );
not ( n1334 , n17 );
and ( n1335 , n6 , n1334 );
not ( n1336 , n1335 );
not ( n1337 , n7 );
and ( n1338 , n6 , n1337 );
not ( n1339 , n1338 );
and ( n1340 , n1336 , n1339 );
not ( n1341 , n1340 );
and ( n1342 , n1335 , n1338 );
not ( n1343 , n1342 );
and ( n1344 , n1341 , n1343 );
not ( n1345 , n1344 );
and ( n1346 , n1333 , n1345 );
not ( n1347 , n1346 );
not ( n1348 , n1333 );
and ( n1349 , n1348 , n1344 );
not ( n1350 , n1349 );
and ( n1351 , n1347 , n1350 );
and ( n1352 , n1331 , n1351 );
not ( n1353 , n1352 );
not ( n1354 , n1331 );
not ( n1355 , n1351 );
and ( n1356 , n1354 , n1355 );
not ( n1357 , n1356 );
and ( n1358 , n1353 , n1357 );
not ( n1359 , n1358 );
and ( n1360 , n1320 , n1359 );
not ( n1361 , n1360 );
not ( n1362 , n705 );
not ( n1363 , n1320 );
and ( n1364 , n1362 , n1363 );
and ( n1365 , n1358 , n1364 );
not ( n1366 , n1365 );
and ( n1367 , n1361 , n1366 );
and ( n1368 , n1312 , n1367 );
and ( n1369 , n1308 , n1368 );
not ( n1370 , n1369 );
and ( n1371 , n6 , n89 );
not ( n1372 , n1371 );
not ( n1373 , n438 );
and ( n1374 , n1372 , n1373 );
and ( n1375 , n6 , n76 );
not ( n1376 , n1375 );
not ( n1377 , n526 );
and ( n1378 , n1376 , n1377 );
and ( n1379 , n6 , n83 );
not ( n1380 , n1379 );
not ( n1381 , n486 );
and ( n1382 , n1380 , n1381 );
not ( n1383 , n1103 );
and ( n1384 , n6 , n117 );
not ( n1385 , n1384 );
and ( n1386 , n1383 , n1385 );
not ( n1387 , n1386 );
and ( n1388 , n1382 , n1387 );
not ( n1389 , n1388 );
not ( n1390 , n1382 );
and ( n1391 , n1390 , n1386 );
not ( n1392 , n1391 );
and ( n1393 , n1389 , n1392 );
not ( n1394 , n1393 );
and ( n1395 , n1378 , n1394 );
not ( n1396 , n1395 );
not ( n1397 , n1378 );
and ( n1398 , n1397 , n1393 );
not ( n1399 , n1398 );
and ( n1400 , n1396 , n1399 );
and ( n1401 , n1374 , n1400 );
not ( n1402 , n1401 );
not ( n1403 , n1374 );
not ( n1404 , n1400 );
and ( n1405 , n1403 , n1404 );
not ( n1406 , n1405 );
and ( n1407 , n1402 , n1406 );
not ( n1408 , n1407 );
and ( n1409 , n6 , n68 );
not ( n1410 , n1409 );
not ( n1411 , n598 );
and ( n1412 , n1410 , n1411 );
not ( n1413 , n1412 );
and ( n1414 , n6 , n74 );
not ( n1415 , n1414 );
not ( n1416 , n552 );
and ( n1417 , n1415 , n1416 );
and ( n1418 , n6 , n71 );
not ( n1419 , n1418 );
not ( n1420 , n569 );
and ( n1421 , n1419 , n1420 );
and ( n1422 , n6 , n80 );
not ( n1423 , n1422 );
not ( n1424 , n507 );
and ( n1425 , n1423 , n1424 );
and ( n1426 , n6 , n86 );
not ( n1427 , n1426 );
not ( n1428 , n461 );
and ( n1429 , n1427 , n1428 );
not ( n1430 , n424 );
not ( n1431 , n92 );
and ( n1432 , n6 , n1431 );
not ( n1433 , n1432 );
and ( n1434 , n1430 , n1433 );
not ( n1435 , n1434 );
and ( n1436 , n1429 , n1435 );
not ( n1437 , n1436 );
not ( n1438 , n1429 );
and ( n1439 , n1438 , n1434 );
not ( n1440 , n1439 );
and ( n1441 , n1437 , n1440 );
not ( n1442 , n1441 );
and ( n1443 , n1425 , n1442 );
not ( n1444 , n1443 );
not ( n1445 , n1425 );
and ( n1446 , n1445 , n1441 );
not ( n1447 , n1446 );
and ( n1448 , n1444 , n1447 );
and ( n1449 , n1421 , n1448 );
not ( n1450 , n1449 );
not ( n1451 , n1421 );
not ( n1452 , n1448 );
and ( n1453 , n1451 , n1452 );
not ( n1454 , n1453 );
and ( n1455 , n1450 , n1454 );
not ( n1456 , n1455 );
and ( n1457 , n1417 , n1456 );
not ( n1458 , n1457 );
not ( n1459 , n1417 );
and ( n1460 , n1459 , n1455 );
not ( n1461 , n1460 );
and ( n1462 , n1458 , n1461 );
not ( n1463 , n1462 );
and ( n1464 , n1413 , n1463 );
not ( n1465 , n1464 );
and ( n1466 , n1412 , n1462 );
not ( n1467 , n1466 );
and ( n1468 , n1465 , n1467 );
and ( n1469 , n1408 , n1468 );
not ( n1470 , n1469 );
not ( n1471 , n1468 );
and ( n1472 , n1407 , n1471 );
not ( n1473 , n1472 );
and ( n1474 , n1470 , n1473 );
not ( n1475 , n1474 );
and ( n1476 , n6 , n49 );
not ( n1477 , n1476 );
not ( n1478 , n291 );
and ( n1479 , n1477 , n1478 );
and ( n1480 , n6 , n47 );
not ( n1481 , n1480 );
not ( n1482 , n275 );
and ( n1483 , n1481 , n1482 );
and ( n1484 , n6 , n56 );
not ( n1485 , n1484 );
not ( n1486 , n333 );
and ( n1487 , n1485 , n1486 );
and ( n1488 , n6 , n53 );
not ( n1489 , n1488 );
not ( n1490 , n313 );
and ( n1491 , n1489 , n1490 );
and ( n1492 , n6 , n62 );
not ( n1493 , n1492 );
not ( n1494 , n373 );
and ( n1495 , n1493 , n1494 );
and ( n1496 , n6 , n65 );
not ( n1497 , n1496 );
not ( n1498 , n391 );
and ( n1499 , n1497 , n1498 );
not ( n1500 , n1499 );
and ( n1501 , n1495 , n1500 );
not ( n1502 , n1501 );
not ( n1503 , n1495 );
and ( n1504 , n1503 , n1499 );
not ( n1505 , n1504 );
and ( n1506 , n1502 , n1505 );
and ( n1507 , n1491 , n1506 );
not ( n1508 , n1507 );
not ( n1509 , n1491 );
not ( n1510 , n1506 );
and ( n1511 , n1509 , n1510 );
not ( n1512 , n1511 );
and ( n1513 , n1508 , n1512 );
not ( n1514 , n1513 );
and ( n1515 , n1487 , n1514 );
not ( n1516 , n1515 );
not ( n1517 , n1487 );
and ( n1518 , n1517 , n1513 );
not ( n1519 , n1518 );
and ( n1520 , n1516 , n1519 );
and ( n1521 , n1483 , n1520 );
not ( n1522 , n1521 );
not ( n1523 , n1483 );
not ( n1524 , n1520 );
and ( n1525 , n1523 , n1524 );
not ( n1526 , n1525 );
and ( n1527 , n1522 , n1526 );
not ( n1528 , n1527 );
and ( n1529 , n1479 , n1528 );
not ( n1530 , n1529 );
not ( n1531 , n1479 );
and ( n1532 , n1531 , n1527 );
not ( n1533 , n1532 );
and ( n1534 , n1530 , n1533 );
and ( n1535 , n6 , n44 );
not ( n1536 , n1535 );
not ( n1537 , n251 );
and ( n1538 , n1536 , n1537 );
not ( n1539 , n991 );
and ( n1540 , n6 , n115 );
not ( n1541 , n1540 );
and ( n1542 , n1539 , n1541 );
and ( n1543 , n6 , n59 );
not ( n1544 , n1543 );
not ( n1545 , n350 );
and ( n1546 , n1544 , n1545 );
and ( n1547 , n6 , n41 );
not ( n1548 , n1547 );
not ( n1549 , n235 );
and ( n1550 , n1548 , n1549 );
not ( n1551 , n1550 );
and ( n1552 , n1546 , n1551 );
not ( n1553 , n1552 );
not ( n1554 , n1546 );
and ( n1555 , n1554 , n1550 );
not ( n1556 , n1555 );
and ( n1557 , n1553 , n1556 );
and ( n1558 , n1542 , n1557 );
not ( n1559 , n1558 );
not ( n1560 , n1542 );
not ( n1561 , n1557 );
and ( n1562 , n1560 , n1561 );
not ( n1563 , n1562 );
and ( n1564 , n1559 , n1563 );
not ( n1565 , n1564 );
and ( n1566 , n1538 , n1565 );
not ( n1567 , n1566 );
not ( n1568 , n1538 );
and ( n1569 , n1568 , n1564 );
not ( n1570 , n1569 );
and ( n1571 , n1567 , n1570 );
and ( n1572 , n1534 , n1571 );
not ( n1573 , n1572 );
not ( n1574 , n1534 );
not ( n1575 , n1571 );
and ( n1576 , n1574 , n1575 );
not ( n1577 , n1576 );
and ( n1578 , n1573 , n1577 );
not ( n1579 , n1578 );
and ( n1580 , n1475 , n1579 );
not ( n1581 , n1580 );
or ( n1582 , n1370 , n1581 );
not ( n1583 , n1582 );
and ( n1584 , n99 , n100 );
and ( n1585 , n101 , n102 );
and ( n1586 , n1584 , n1585 );
and ( n1587 , n95 , n96 );
and ( n1588 , n97 , n98 );
and ( n1589 , n1587 , n1588 );
and ( n1590 , n1586 , n1589 );
and ( n1591 , n107 , n108 );
and ( n1592 , n109 , n110 );
and ( n1593 , n1591 , n1592 );
and ( n1594 , n103 , n104 );
and ( n1595 , n105 , n106 );
and ( n1596 , n1594 , n1595 );
and ( n1597 , n1593 , n1596 );
and ( n1598 , n1590 , n1597 );
and ( n1599 , n1583 , n1598 );
and ( n1600 , n1209 , n1599 );
not ( n1601 , n133 );
and ( n1602 , n6 , n1601 );
not ( n1603 , n1602 );
not ( n1604 , n6 );
and ( n1605 , n1604 , n132 );
not ( n1606 , n1605 );
and ( n1607 , n1603 , n1606 );
not ( n1608 , n659 );
and ( n1609 , n719 , n1608 );
not ( n1610 , n1609 );
not ( n1611 , n719 );
and ( n1612 , n1611 , n659 );
not ( n1613 , n1612 );
and ( n1614 , n1610 , n1613 );
and ( n1615 , n1607 , n1614 );
not ( n1616 , n1615 );
not ( n1617 , n1607 );
not ( n1618 , n1614 );
and ( n1619 , n1617 , n1618 );
not ( n1620 , n1619 );
and ( n1621 , n1616 , n1620 );
not ( n1622 , n750 );
and ( n1623 , n642 , n1622 );
not ( n1624 , n1623 );
not ( n1625 , n642 );
and ( n1626 , n1625 , n750 );
not ( n1627 , n1626 );
and ( n1628 , n1624 , n1627 );
and ( n1629 , n703 , n1628 );
not ( n1630 , n1629 );
not ( n1631 , n703 );
not ( n1632 , n1628 );
and ( n1633 , n1631 , n1632 );
not ( n1634 , n1633 );
and ( n1635 , n1630 , n1634 );
not ( n1636 , n1635 );
and ( n1637 , n770 , n1636 );
not ( n1638 , n1637 );
not ( n1639 , n770 );
and ( n1640 , n1639 , n1635 );
not ( n1641 , n1640 );
and ( n1642 , n1638 , n1641 );
and ( n1643 , n677 , n1642 );
not ( n1644 , n1643 );
not ( n1645 , n677 );
not ( n1646 , n1642 );
and ( n1647 , n1645 , n1646 );
not ( n1648 , n1647 );
and ( n1649 , n1644 , n1648 );
not ( n1650 , n1649 );
and ( n1651 , n735 , n1650 );
not ( n1652 , n1651 );
not ( n1653 , n735 );
and ( n1654 , n1653 , n1649 );
not ( n1655 , n1654 );
and ( n1656 , n1652 , n1655 );
and ( n1657 , n802 , n1656 );
not ( n1658 , n1657 );
not ( n1659 , n802 );
not ( n1660 , n1656 );
and ( n1661 , n1659 , n1660 );
not ( n1662 , n1661 );
and ( n1663 , n1658 , n1662 );
and ( n1664 , n1621 , n1663 );
not ( n1665 , n1664 );
not ( n1666 , n447 );
not ( n1667 , n91 );
and ( n1668 , n6 , n1667 );
not ( n1669 , n1668 );
and ( n1670 , n1666 , n1669 );
not ( n1671 , n459 );
and ( n1672 , n1670 , n1671 );
not ( n1673 , n1672 );
not ( n1674 , n1670 );
and ( n1675 , n1674 , n459 );
not ( n1676 , n1675 );
and ( n1677 , n1673 , n1676 );
not ( n1678 , n1677 );
and ( n1679 , n595 , n1678 );
not ( n1680 , n1679 );
not ( n1681 , n595 );
and ( n1682 , n1681 , n1677 );
not ( n1683 , n1682 );
and ( n1684 , n1680 , n1683 );
and ( n1685 , n435 , n1684 );
not ( n1686 , n1685 );
not ( n1687 , n435 );
not ( n1688 , n1684 );
and ( n1689 , n1687 , n1688 );
not ( n1690 , n1689 );
and ( n1691 , n1686 , n1690 );
not ( n1692 , n1691 );
and ( n1693 , n505 , n1692 );
not ( n1694 , n1693 );
not ( n1695 , n505 );
and ( n1696 , n1695 , n1691 );
not ( n1697 , n1696 );
and ( n1698 , n1694 , n1697 );
and ( n1699 , n523 , n1698 );
not ( n1700 , n1699 );
not ( n1701 , n523 );
not ( n1702 , n1698 );
and ( n1703 , n1701 , n1702 );
not ( n1704 , n1703 );
and ( n1705 , n1700 , n1704 );
not ( n1706 , n154 );
and ( n1707 , n6 , n1706 );
not ( n1708 , n1707 );
not ( n1709 , n6 );
and ( n1710 , n1709 , n155 );
not ( n1711 , n1710 );
and ( n1712 , n1708 , n1711 );
not ( n1713 , n1712 );
and ( n1714 , n483 , n1713 );
not ( n1715 , n1714 );
not ( n1716 , n483 );
and ( n1717 , n1716 , n1712 );
not ( n1718 , n1717 );
and ( n1719 , n1715 , n1718 );
not ( n1720 , n1719 );
and ( n1721 , n549 , n1720 );
not ( n1722 , n1721 );
not ( n1723 , n549 );
and ( n1724 , n1723 , n1719 );
not ( n1725 , n1724 );
and ( n1726 , n1722 , n1725 );
not ( n1727 , n1726 );
and ( n1728 , n567 , n1727 );
not ( n1729 , n1728 );
not ( n1730 , n567 );
and ( n1731 , n1730 , n1726 );
not ( n1732 , n1731 );
and ( n1733 , n1729 , n1732 );
not ( n1734 , n1733 );
and ( n1735 , n1705 , n1734 );
not ( n1736 , n1735 );
not ( n1737 , n1705 );
and ( n1738 , n1737 , n1733 );
not ( n1739 , n1738 );
and ( n1740 , n1736 , n1739 );
not ( n1741 , n1740 );
not ( n1742 , n6 );
not ( n1743 , n121 );
and ( n1744 , n1742 , n1743 );
not ( n1745 , n1744 );
and ( n1746 , n6 , n122 );
not ( n1747 , n1746 );
and ( n1748 , n1745 , n1747 );
not ( n1749 , n878 );
and ( n1750 , n1748 , n1749 );
not ( n1751 , n1750 );
not ( n1752 , n1748 );
and ( n1753 , n1752 , n878 );
not ( n1754 , n1753 );
and ( n1755 , n1751 , n1754 );
not ( n1756 , n893 );
and ( n1757 , n909 , n1756 );
not ( n1758 , n1757 );
not ( n1759 , n909 );
and ( n1760 , n1759 , n893 );
not ( n1761 , n1760 );
and ( n1762 , n1758 , n1761 );
and ( n1763 , n1755 , n1762 );
not ( n1764 , n1763 );
not ( n1765 , n1755 );
not ( n1766 , n1762 );
and ( n1767 , n1765 , n1766 );
not ( n1768 , n1767 );
and ( n1769 , n1764 , n1768 );
not ( n1770 , n2 );
not ( n1771 , n4 );
and ( n1772 , n1770 , n1771 );
not ( n1773 , n1772 );
and ( n1774 , n2 , n4 );
not ( n1775 , n1774 );
and ( n1776 , n1773 , n1775 );
not ( n1777 , n1776 );
and ( n1778 , n6 , n1777 );
not ( n1779 , n1778 );
not ( n1780 , n6 );
not ( n1781 , n217 );
not ( n1782 , n223 );
and ( n1783 , n1781 , n1782 );
not ( n1784 , n1783 );
and ( n1785 , n1780 , n1784 );
not ( n1786 , n1785 );
and ( n1787 , n1779 , n1786 );
not ( n1788 , n1787 );
and ( n1789 , n1769 , n1788 );
not ( n1790 , n1789 );
not ( n1791 , n1769 );
and ( n1792 , n1791 , n1787 );
not ( n1793 , n1792 );
and ( n1794 , n1790 , n1793 );
not ( n1795 , n1794 );
and ( n1796 , n861 , n1795 );
not ( n1797 , n1796 );
not ( n1798 , n861 );
and ( n1799 , n1798 , n1794 );
not ( n1800 , n1799 );
and ( n1801 , n1797 , n1800 );
and ( n1802 , n854 , n1801 );
not ( n1803 , n1802 );
not ( n1804 , n854 );
not ( n1805 , n1801 );
and ( n1806 , n1804 , n1805 );
not ( n1807 , n1806 );
and ( n1808 , n1803 , n1807 );
not ( n1809 , n1808 );
not ( n1810 , n272 );
and ( n1811 , n388 , n1810 );
not ( n1812 , n1811 );
not ( n1813 , n388 );
and ( n1814 , n1813 , n272 );
not ( n1815 , n1814 );
and ( n1816 , n1812 , n1815 );
not ( n1817 , n6 );
not ( n1818 , n144 );
and ( n1819 , n1817 , n1818 );
not ( n1820 , n1819 );
and ( n1821 , n6 , n143 );
not ( n1822 , n1821 );
and ( n1823 , n1820 , n1822 );
not ( n1824 , n330 );
and ( n1825 , n1823 , n1824 );
not ( n1826 , n1825 );
not ( n1827 , n1823 );
and ( n1828 , n1827 , n330 );
not ( n1829 , n1828 );
and ( n1830 , n1826 , n1829 );
and ( n1831 , n370 , n1830 );
not ( n1832 , n1831 );
not ( n1833 , n370 );
not ( n1834 , n1830 );
and ( n1835 , n1833 , n1834 );
not ( n1836 , n1835 );
and ( n1837 , n1832 , n1836 );
not ( n1838 , n1837 );
not ( n1839 , n311 );
and ( n1840 , n289 , n1839 );
not ( n1841 , n1840 );
not ( n1842 , n289 );
and ( n1843 , n1842 , n311 );
not ( n1844 , n1843 );
and ( n1845 , n1841 , n1844 );
and ( n1846 , n233 , n1845 );
not ( n1847 , n1846 );
not ( n1848 , n233 );
not ( n1849 , n1845 );
and ( n1850 , n1848 , n1849 );
not ( n1851 , n1850 );
and ( n1852 , n1847 , n1851 );
not ( n1853 , n248 );
and ( n1854 , n348 , n1853 );
not ( n1855 , n1854 );
not ( n1856 , n348 );
and ( n1857 , n1856 , n248 );
not ( n1858 , n1857 );
and ( n1859 , n1855 , n1858 );
not ( n1860 , n1859 );
and ( n1861 , n1852 , n1860 );
not ( n1862 , n1861 );
not ( n1863 , n1852 );
and ( n1864 , n1863 , n1859 );
not ( n1865 , n1864 );
and ( n1866 , n1862 , n1865 );
not ( n1867 , n1866 );
and ( n1868 , n1838 , n1867 );
not ( n1869 , n1868 );
and ( n1870 , n1837 , n1866 );
not ( n1871 , n1870 );
and ( n1872 , n1869 , n1871 );
not ( n1873 , n1872 );
and ( n1874 , n1816 , n1873 );
not ( n1875 , n1874 );
not ( n1876 , n1816 );
and ( n1877 , n1876 , n1872 );
not ( n1878 , n1877 );
and ( n1879 , n1875 , n1878 );
not ( n1880 , n1879 );
and ( n1881 , n1809 , n1880 );
and ( n1882 , n1741 , n1881 );
and ( n1883 , n1665 , n1882 );
not ( n1884 , n1621 );
not ( n1885 , n1663 );
and ( n1886 , n1884 , n1885 );
not ( n1887 , n94 );
not ( n1888 , n93 );
not ( n1889 , n6 );
and ( n1890 , n1889 , n91 );
and ( n1891 , n1888 , n1890 );
not ( n1892 , n1891 );
not ( n1893 , n6 );
not ( n1894 , n91 );
and ( n1895 , n1893 , n1894 );
and ( n1896 , n93 , n1895 );
not ( n1897 , n1896 );
and ( n1898 , n1892 , n1897 );
and ( n1899 , n1887 , n1898 );
not ( n1900 , n1898 );
and ( n1901 , n94 , n1900 );
and ( n1902 , n1 , n1774 );
not ( n1903 , n1902 );
and ( n1904 , n3 , n1903 );
not ( n1905 , n1904 );
not ( n1906 , n1772 );
and ( n1907 , n222 , n1906 );
not ( n1908 , n1907 );
not ( n1909 , n705 );
not ( n1910 , n1338 );
and ( n1911 , n1909 , n1910 );
not ( n1912 , n1911 );
and ( n1913 , n5 , n1912 );
not ( n1914 , n1913 );
and ( n1915 , n1908 , n1914 );
not ( n1916 , n10 );
not ( n1917 , n705 );
not ( n1918 , n1322 );
and ( n1919 , n1917 , n1918 );
and ( n1920 , n1916 , n1919 );
not ( n1921 , n1920 );
not ( n1922 , n5 );
and ( n1923 , n1922 , n1911 );
not ( n1924 , n1923 );
and ( n1925 , n1921 , n1924 );
not ( n1926 , n1919 );
and ( n1927 , n10 , n1926 );
not ( n1928 , n1927 );
not ( n1929 , n705 );
not ( n1930 , n1333 );
and ( n1931 , n1929 , n1930 );
not ( n1932 , n1931 );
and ( n1933 , n12 , n1932 );
not ( n1934 , n1933 );
and ( n1935 , n1928 , n1934 );
not ( n1936 , n14 );
not ( n1937 , n705 );
not ( n1938 , n1324 );
and ( n1939 , n1937 , n1938 );
and ( n1940 , n1936 , n1939 );
not ( n1941 , n1940 );
not ( n1942 , n12 );
and ( n1943 , n1942 , n1931 );
not ( n1944 , n1943 );
and ( n1945 , n1941 , n1944 );
not ( n1946 , n16 );
not ( n1947 , n705 );
not ( n1948 , n1335 );
and ( n1949 , n1947 , n1948 );
and ( n1950 , n1946 , n1949 );
not ( n1951 , n1939 );
and ( n1952 , n14 , n1951 );
not ( n1953 , n1952 );
and ( n1954 , n1950 , n1953 );
not ( n1955 , n1954 );
and ( n1956 , n1945 , n1955 );
not ( n1957 , n1956 );
and ( n1958 , n1935 , n1957 );
not ( n1959 , n1958 );
and ( n1960 , n1925 , n1959 );
not ( n1961 , n1960 );
and ( n1962 , n1915 , n1961 );
not ( n1963 , n1962 );
and ( n1964 , n1905 , n1963 );
and ( n1965 , n85 , n1429 );
not ( n1966 , n1965 );
not ( n1967 , n88 );
not ( n1968 , n1374 );
and ( n1969 , n1967 , n1968 );
not ( n1970 , n1969 );
and ( n1971 , n88 , n1374 );
not ( n1972 , n1971 );
not ( n1973 , n1891 );
and ( n1974 , n94 , n1973 );
not ( n1975 , n1974 );
not ( n1976 , n1896 );
and ( n1977 , n1975 , n1976 );
not ( n1978 , n1977 );
and ( n1979 , n1972 , n1978 );
not ( n1980 , n1979 );
and ( n1981 , n1970 , n1980 );
not ( n1982 , n1981 );
and ( n1983 , n1966 , n1982 );
not ( n1984 , n1983 );
not ( n1985 , n85 );
not ( n1986 , n1429 );
and ( n1987 , n1985 , n1986 );
not ( n1988 , n1987 );
not ( n1989 , n82 );
not ( n1990 , n1382 );
and ( n1991 , n1989 , n1990 );
not ( n1992 , n1991 );
and ( n1993 , n1988 , n1992 );
and ( n1994 , n1984 , n1993 );
not ( n1995 , n1994 );
and ( n1996 , n82 , n1382 );
not ( n1997 , n1996 );
and ( n1998 , n79 , n1425 );
not ( n1999 , n1998 );
and ( n2000 , n1997 , n1999 );
and ( n2001 , n1995 , n2000 );
not ( n2002 , n2001 );
not ( n2003 , n79 );
not ( n2004 , n1425 );
and ( n2005 , n2003 , n2004 );
not ( n2006 , n2005 );
not ( n2007 , n78 );
not ( n2008 , n1378 );
and ( n2009 , n2007 , n2008 );
not ( n2010 , n2009 );
and ( n2011 , n2006 , n2010 );
and ( n2012 , n2002 , n2011 );
not ( n2013 , n2012 );
and ( n2014 , n73 , n1417 );
not ( n2015 , n2014 );
and ( n2016 , n78 , n1378 );
not ( n2017 , n2016 );
and ( n2018 , n70 , n1421 );
not ( n2019 , n2018 );
and ( n2020 , n2017 , n2019 );
and ( n2021 , n2015 , n2020 );
and ( n2022 , n2013 , n2021 );
not ( n2023 , n2022 );
not ( n2024 , n2018 );
not ( n2025 , n73 );
not ( n2026 , n1417 );
and ( n2027 , n2025 , n2026 );
and ( n2028 , n2024 , n2027 );
not ( n2029 , n2028 );
not ( n2030 , n70 );
not ( n2031 , n1421 );
and ( n2032 , n2030 , n2031 );
not ( n2033 , n2032 );
not ( n2034 , n67 );
not ( n2035 , n1412 );
and ( n2036 , n2034 , n2035 );
not ( n2037 , n2036 );
and ( n2038 , n2033 , n2037 );
and ( n2039 , n2029 , n2038 );
and ( n2040 , n2023 , n2039 );
not ( n2041 , n2040 );
and ( n2042 , n61 , n1495 );
not ( n2043 , n2042 );
not ( n2044 , n64 );
not ( n2045 , n1499 );
and ( n2046 , n2044 , n2045 );
and ( n2047 , n2043 , n2046 );
not ( n2048 , n2047 );
not ( n2049 , n61 );
not ( n2050 , n1495 );
and ( n2051 , n2049 , n2050 );
not ( n2052 , n2051 );
not ( n2053 , n58 );
not ( n2054 , n1546 );
and ( n2055 , n2053 , n2054 );
not ( n2056 , n2055 );
and ( n2057 , n2052 , n2056 );
and ( n2058 , n2048 , n2057 );
and ( n2059 , n52 , n1491 );
not ( n2060 , n2059 );
not ( n2061 , n2042 );
and ( n2062 , n2060 , n2061 );
and ( n2063 , n67 , n1412 );
not ( n2064 , n2063 );
and ( n2065 , n64 , n1499 );
not ( n2066 , n2065 );
and ( n2067 , n2064 , n2066 );
and ( n2068 , n2062 , n2067 );
not ( n2069 , n55 );
not ( n2070 , n1487 );
and ( n2071 , n2069 , n2070 );
not ( n2072 , n2071 );
not ( n2073 , n52 );
not ( n2074 , n1491 );
and ( n2075 , n2073 , n2074 );
not ( n2076 , n2075 );
and ( n2077 , n2072 , n2076 );
and ( n2078 , n58 , n1546 );
not ( n2079 , n2078 );
and ( n2080 , n55 , n1487 );
not ( n2081 , n2080 );
and ( n2082 , n2079 , n2081 );
and ( n2083 , n2077 , n2082 );
and ( n2084 , n2068 , n2083 );
and ( n2085 , n2058 , n2084 );
and ( n2086 , n2041 , n2085 );
not ( n2087 , n2086 );
not ( n2088 , n51 );
not ( n2089 , n1479 );
and ( n2090 , n2088 , n2089 );
not ( n2091 , n2090 );
not ( n2092 , n2059 );
not ( n2093 , n2058 );
and ( n2094 , n2082 , n2093 );
not ( n2095 , n2094 );
and ( n2096 , n2077 , n2095 );
not ( n2097 , n2096 );
and ( n2098 , n2092 , n2097 );
not ( n2099 , n2098 );
and ( n2100 , n2091 , n2099 );
and ( n2101 , n2087 , n2100 );
not ( n2102 , n2101 );
and ( n2103 , n40 , n1550 );
not ( n2104 , n2103 );
and ( n2105 , n43 , n1538 );
not ( n2106 , n2105 );
and ( n2107 , n2104 , n2106 );
and ( n2108 , n46 , n1483 );
not ( n2109 , n2108 );
and ( n2110 , n51 , n1479 );
not ( n2111 , n2110 );
and ( n2112 , n2109 , n2111 );
and ( n2113 , n2107 , n2112 );
and ( n2114 , n2102 , n2113 );
not ( n2115 , n2114 );
not ( n2116 , n40 );
not ( n2117 , n1550 );
and ( n2118 , n2116 , n2117 );
not ( n2119 , n2118 );
not ( n2120 , n43 );
not ( n2121 , n1538 );
and ( n2122 , n2120 , n2121 );
not ( n2123 , n2122 );
not ( n2124 , n46 );
not ( n2125 , n1483 );
and ( n2126 , n2124 , n2125 );
not ( n2127 , n2126 );
and ( n2128 , n2123 , n2127 );
not ( n2129 , n2128 );
and ( n2130 , n2107 , n2129 );
not ( n2131 , n2130 );
and ( n2132 , n2119 , n2131 );
and ( n2133 , n2115 , n2132 );
not ( n2134 , n2133 );
not ( n2135 , n34 );
not ( n2136 , n1255 );
and ( n2137 , n2135 , n2136 );
not ( n2138 , n2137 );
not ( n2139 , n37 );
not ( n2140 , n1251 );
and ( n2141 , n2139 , n2140 );
not ( n2142 , n2141 );
and ( n2143 , n2138 , n2142 );
not ( n2144 , n1270 );
and ( n2145 , n25 , n2144 );
not ( n2146 , n2145 );
not ( n2147 , n1275 );
and ( n2148 , n22 , n2147 );
not ( n2149 , n2148 );
and ( n2150 , n2146 , n2149 );
and ( n2151 , n2143 , n2150 );
not ( n2152 , n26 );
and ( n2153 , n2152 , n1217 );
not ( n2154 , n2153 );
not ( n2155 , n25 );
and ( n2156 , n2155 , n1270 );
not ( n2157 , n2156 );
and ( n2158 , n2154 , n2157 );
and ( n2159 , n31 , n1259 );
not ( n2160 , n2159 );
and ( n2161 , n34 , n1255 );
not ( n2162 , n2161 );
and ( n2163 , n2160 , n2162 );
and ( n2164 , n2158 , n2163 );
and ( n2165 , n2151 , n2164 );
not ( n2166 , n1263 );
and ( n2167 , n28 , n2166 );
not ( n2168 , n2167 );
not ( n2169 , n28 );
and ( n2170 , n2169 , n1263 );
not ( n2171 , n2170 );
not ( n2172 , n1217 );
and ( n2173 , n26 , n2172 );
not ( n2174 , n2173 );
and ( n2175 , n2171 , n2174 );
and ( n2176 , n2168 , n2175 );
and ( n2177 , n37 , n1251 );
not ( n2178 , n2177 );
not ( n2179 , n18 );
and ( n2180 , n2179 , n1230 );
not ( n2181 , n2180 );
not ( n2182 , n31 );
not ( n2183 , n1259 );
and ( n2184 , n2182 , n2183 );
not ( n2185 , n2184 );
and ( n2186 , n2181 , n2185 );
and ( n2187 , n2178 , n2186 );
not ( n2188 , n1222 );
and ( n2189 , n20 , n2188 );
not ( n2190 , n2189 );
not ( n2191 , n1230 );
and ( n2192 , n18 , n2191 );
not ( n2193 , n2192 );
and ( n2194 , n2190 , n2193 );
not ( n2195 , n20 );
and ( n2196 , n2195 , n1222 );
not ( n2197 , n2196 );
not ( n2198 , n22 );
and ( n2199 , n2198 , n1275 );
not ( n2200 , n2199 );
and ( n2201 , n2197 , n2200 );
and ( n2202 , n2194 , n2201 );
and ( n2203 , n2187 , n2202 );
and ( n2204 , n2176 , n2203 );
and ( n2205 , n2165 , n2204 );
and ( n2206 , n2134 , n2205 );
not ( n2207 , n2206 );
not ( n2208 , n2180 );
not ( n2209 , n2143 );
and ( n2210 , n2209 , n2163 );
not ( n2211 , n2210 );
not ( n2212 , n2184 );
and ( n2213 , n28 , n2212 );
and ( n2214 , n2211 , n2213 );
not ( n2215 , n2214 );
and ( n2216 , n2176 , n2215 );
not ( n2217 , n2216 );
and ( n2218 , n2158 , n2217 );
not ( n2219 , n2218 );
and ( n2220 , n2150 , n2219 );
not ( n2221 , n2220 );
and ( n2222 , n2201 , n2221 );
not ( n2223 , n2222 );
and ( n2224 , n2194 , n2223 );
not ( n2225 , n2224 );
and ( n2226 , n2208 , n2225 );
and ( n2227 , n2207 , n2226 );
not ( n2228 , n2227 );
not ( n2229 , n1950 );
not ( n2230 , n1952 );
and ( n2231 , n2229 , n2230 );
not ( n2232 , n1949 );
and ( n2233 , n16 , n2232 );
not ( n2234 , n2233 );
not ( n2235 , n1904 );
and ( n2236 , n2234 , n2235 );
and ( n2237 , n2231 , n2236 );
and ( n2238 , n1935 , n1915 );
and ( n2239 , n1925 , n1945 );
and ( n2240 , n2238 , n2239 );
and ( n2241 , n2237 , n2240 );
and ( n2242 , n2228 , n2241 );
not ( n2243 , n1883 );
or ( n2244 , n1886 , n2243 );
or ( n2245 , n954 , n220 );
not ( n2246 , n1600 );
or ( n2247 , n2244 , n2246 );
or ( n2248 , n1901 , n1899 );
not ( n2249 , n1964 );
or ( n2250 , n2242 , n2249 );
endmodule

