module top (out_0, out_1, out_2, out_3, out_4, out_5, out_6, out_7, out_8, out_9, out_10, new_out1, new_out2, new_out3, new_out4, new_out5, in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27, in_28, in_29, in_30, in_31);
	input in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27, in_28, in_29, in_30, in_31;
	output out_0, out_1, out_2, out_3, out_4, out_5, out_6, out_7, out_8, out_9, out_10, out_11, new_out1, new_out2, new_out3, new_out4, new_out5;
	wire gm_n100, gm_n1000, gm_n1001, gm_n1002, gm_n1003, gm_n1004, gm_n1005, gm_n1006, gm_n1007, gm_n1008, gm_n1009, gm_n101, gm_n1010, gm_n1011, gm_n1012, gm_n1013, gm_n1014, gm_n1015, gm_n1016, gm_n1017, gm_n1018, gm_n1019, gm_n102, gm_n1020, gm_n1021, gm_n1022, gm_n1023, gm_n1024, gm_n1025, gm_n1026, gm_n1027, gm_n1028, gm_n1029, gm_n103, gm_n1030, gm_n1031, gm_n1032, gm_n1033, gm_n1034, gm_n1035, gm_n1036, gm_n1037, gm_n1038, gm_n1039, gm_n104, gm_n1040, gm_n1041, gm_n1042, gm_n1043, gm_n1044, gm_n1045, gm_n1046, gm_n1047, gm_n1048, gm_n1049, gm_n105, gm_n1050, gm_n1051, gm_n1052, gm_n1053, gm_n1054, gm_n1055, gm_n1056, gm_n1057, gm_n1058, gm_n1059, gm_n106, gm_n1060, gm_n1061, gm_n1062, gm_n1063, gm_n1064, gm_n1065, gm_n1066, gm_n1067, gm_n1068, gm_n1069, gm_n107, gm_n1070, gm_n1071, gm_n1072, gm_n1073, gm_n1074, gm_n1075, gm_n1076, gm_n1077, gm_n1078, gm_n1079, gm_n108, gm_n1080, gm_n1081, gm_n1082, gm_n1083, gm_n1084, gm_n1085, gm_n1086, gm_n1087, gm_n1088, gm_n1089, gm_n109, gm_n1090, gm_n1091, gm_n1092, gm_n1093, gm_n1094, gm_n1095, gm_n1096, gm_n1097, gm_n1098, gm_n1099, gm_n110, gm_n1100, gm_n1101, gm_n1102, gm_n1103, gm_n1104, gm_n1105, gm_n1106, gm_n1107, gm_n1108, gm_n1109, gm_n111, gm_n1110, gm_n1111, gm_n1112, gm_n1113, gm_n1114, gm_n1115, gm_n1116, gm_n1117, gm_n1118, gm_n1119, gm_n112, gm_n1120, gm_n1121, gm_n1122, gm_n1123, gm_n1124, gm_n1125, gm_n1126, gm_n1127, gm_n1128, gm_n1129, gm_n113, gm_n1130, gm_n1131, gm_n1132, gm_n1133, gm_n1134, gm_n1135, gm_n1136, gm_n1137, gm_n1138, gm_n1139, gm_n114, gm_n1140, gm_n1141, gm_n1142, gm_n1143, gm_n1144, gm_n1145, gm_n1146, gm_n1147, gm_n1148, gm_n1149, gm_n115, gm_n1150, gm_n1151, gm_n1152, gm_n1153, gm_n1154, gm_n1155, gm_n1156, gm_n1157, gm_n1158, gm_n1159, gm_n116, gm_n1160, gm_n1161, gm_n1162, gm_n1163, gm_n1164, gm_n1165, gm_n1166, gm_n1167, gm_n1168, gm_n1169, gm_n117, gm_n1170, gm_n1171, gm_n1172, gm_n1173, gm_n1174, gm_n1175, gm_n1176, gm_n1177, gm_n1178, gm_n1179, gm_n118, gm_n1180, gm_n1181, gm_n1182, gm_n1183, gm_n1184, gm_n1185, gm_n1186, gm_n1187, gm_n1188, gm_n1189, gm_n119, gm_n1190, gm_n1191, gm_n1192, gm_n1193, gm_n1194, gm_n1195, gm_n1196, gm_n1197, gm_n1198, gm_n1199, gm_n120, gm_n1200, gm_n1201, gm_n1202, gm_n1203, gm_n1204, gm_n1205, gm_n1206, gm_n1207, gm_n1208, gm_n1209, gm_n121, gm_n1211, gm_n1212, gm_n1213, gm_n1214, gm_n1215, gm_n1216, gm_n1217, gm_n1218, gm_n1219, gm_n122, gm_n1220, gm_n1221, gm_n1222, gm_n1223, gm_n1224, gm_n1225, gm_n1226, gm_n1227, gm_n1228, gm_n1229, gm_n123, gm_n1230, gm_n1231, gm_n1232, gm_n1233, gm_n1234, gm_n1235, gm_n1236, gm_n1237, gm_n1238, gm_n1239, gm_n124, gm_n1240, gm_n1241, gm_n1242, gm_n1243, gm_n1244, gm_n1245, gm_n1246, gm_n1247, gm_n1248, gm_n1249, gm_n125, gm_n1250, gm_n1251, gm_n1252, gm_n1253, gm_n1254, gm_n1255, gm_n1256, gm_n1257, gm_n1258, gm_n1259, gm_n126, gm_n1260, gm_n1261, gm_n1262, gm_n1263, gm_n1264, gm_n1265, gm_n1266, gm_n1267, gm_n1268, gm_n1269, gm_n127, gm_n1270, gm_n1271, gm_n1272, gm_n1273, gm_n1274, gm_n1275, gm_n1276, gm_n1277, gm_n1278, gm_n1279, gm_n128, gm_n1280, gm_n1281, gm_n1282, gm_n1283, gm_n1284, gm_n1285, gm_n1286, gm_n1287, gm_n1288, gm_n1289, gm_n129, gm_n1290, gm_n1291, gm_n1292, gm_n1293, gm_n1294, gm_n1295, gm_n1296, gm_n1297, gm_n1298, gm_n1299, gm_n130, gm_n1300, gm_n1301, gm_n1302, gm_n1303, gm_n1304, gm_n1305, gm_n1306, gm_n1307, gm_n1308, gm_n1309, gm_n131, gm_n1310, gm_n1311, gm_n1312, gm_n1313, gm_n1314, gm_n1315, gm_n1316, gm_n1317, gm_n1318, gm_n1319, gm_n132, gm_n1320, gm_n1321, gm_n1322, gm_n1323, gm_n1324, gm_n1325, gm_n1326, gm_n1327, gm_n1328, gm_n1329, gm_n133, gm_n1330, gm_n1331, gm_n1332, gm_n1333, gm_n1334, gm_n1335, gm_n1336, gm_n1337, gm_n1338, gm_n1339, gm_n134, gm_n1340, gm_n1341, gm_n1342, gm_n1343, gm_n1344, gm_n1345, gm_n1346, gm_n1347, gm_n1348, gm_n1349, gm_n135, gm_n1350, gm_n1351, gm_n1352, gm_n1353, gm_n1354, gm_n1355, gm_n1356, gm_n1357, gm_n1358, gm_n1359, gm_n136, gm_n1360, gm_n1361, gm_n1362, gm_n1363, gm_n1364, gm_n1365, gm_n1366, gm_n1367, gm_n1368, gm_n1369, gm_n137, gm_n1370, gm_n1371, gm_n1372, gm_n1373, gm_n1374, gm_n1375, gm_n1376, gm_n1377, gm_n1378, gm_n1379, gm_n138, gm_n1380, gm_n1381, gm_n1382, gm_n1383, gm_n1384, gm_n1385, gm_n1386, gm_n1387, gm_n1388, gm_n1389, gm_n139, gm_n1390, gm_n1391, gm_n1392, gm_n1393, gm_n1394, gm_n1395, gm_n1396, gm_n1397, gm_n1398, gm_n1399, gm_n140, gm_n1400, gm_n1401, gm_n1402, gm_n1403, gm_n1404, gm_n1405, gm_n1406, gm_n1407, gm_n1408, gm_n1409, gm_n141, gm_n1410, gm_n1411, gm_n1412, gm_n1413, gm_n1414, gm_n1416, gm_n1417, gm_n1418, gm_n1419, gm_n142, gm_n1420, gm_n1421, gm_n1422, gm_n1423, gm_n1424, gm_n1425, gm_n1426, gm_n1427, gm_n1428, gm_n1429, gm_n143, gm_n1430, gm_n1431, gm_n1432, gm_n1433, gm_n1434, gm_n1435, gm_n1436, gm_n1437, gm_n1438, gm_n1439, gm_n144, gm_n1440, gm_n1441, gm_n1442, gm_n1443, gm_n1444, gm_n1445, gm_n1446, gm_n1447, gm_n1448, gm_n1449, gm_n145, gm_n1450, gm_n1451, gm_n1452, gm_n1453, gm_n1454, gm_n1455, gm_n1456, gm_n1457, gm_n1458, gm_n1459, gm_n146, gm_n1460, gm_n1461, gm_n1462, gm_n1463, gm_n1464, gm_n1465, gm_n1466, gm_n1467, gm_n1468, gm_n1469, gm_n147, gm_n1470, gm_n1471, gm_n1472, gm_n1473, gm_n1474, gm_n1475, gm_n1476, gm_n1477, gm_n1478, gm_n1479, gm_n148, gm_n1480, gm_n1481, gm_n1482, gm_n1483, gm_n1484, gm_n1485, gm_n1486, gm_n1487, gm_n1488, gm_n1489, gm_n149, gm_n1490, gm_n1491, gm_n1492, gm_n1493, gm_n1494, gm_n1495, gm_n1496, gm_n1497, gm_n1498, gm_n1499, gm_n150, gm_n1500, gm_n1501, gm_n1502, gm_n1503, gm_n1504, gm_n1505, gm_n1506, gm_n1507, gm_n1508, gm_n1509, gm_n151, gm_n1510, gm_n1511, gm_n1512, gm_n1513, gm_n1514, gm_n1515, gm_n1516, gm_n1517, gm_n1518, gm_n1519, gm_n152, gm_n1520, gm_n1521, gm_n1522, gm_n1523, gm_n1524, gm_n1525, gm_n1526, gm_n1527, gm_n1528, gm_n1529, gm_n153, gm_n1530, gm_n1531, gm_n1532, gm_n1533, gm_n1534, gm_n1535, gm_n1536, gm_n1537, gm_n1538, gm_n1539, gm_n154, gm_n1540, gm_n1541, gm_n1542, gm_n1543, gm_n1544, gm_n1545, gm_n1546, gm_n1547, gm_n1548, gm_n1549, gm_n155, gm_n1550, gm_n1551, gm_n1552, gm_n1553, gm_n1554, gm_n1555, gm_n1556, gm_n1557, gm_n1558, gm_n1559, gm_n156, gm_n1560, gm_n1561, gm_n1562, gm_n1563, gm_n1564, gm_n1565, gm_n1566, gm_n1567, gm_n1568, gm_n1569, gm_n157, gm_n1570, gm_n1571, gm_n1572, gm_n1573, gm_n1574, gm_n1575, gm_n1576, gm_n1577, gm_n1578, gm_n1579, gm_n158, gm_n1580, gm_n1581, gm_n1582, gm_n1583, gm_n1584, gm_n1585, gm_n1586, gm_n1587, gm_n1588, gm_n1589, gm_n159, gm_n1590, gm_n1591, gm_n1592, gm_n1593, gm_n1594, gm_n1595, gm_n1596, gm_n1597, gm_n1598, gm_n1599, gm_n160, gm_n1600, gm_n1601, gm_n1602, gm_n1603, gm_n1604, gm_n1605, gm_n1606, gm_n1607, gm_n1609, gm_n161, gm_n1610, gm_n1611, gm_n1612, gm_n1613, gm_n1614, gm_n1615, gm_n1616, gm_n1617, gm_n1618, gm_n1619, gm_n162, gm_n1620, gm_n1621, gm_n1622, gm_n1623, gm_n1624, gm_n1625, gm_n1626, gm_n1627, gm_n1628, gm_n1629, gm_n163, gm_n1630, gm_n1631, gm_n1632, gm_n1633, gm_n1634, gm_n1635, gm_n1636, gm_n1637, gm_n1638, gm_n1639, gm_n164, gm_n1640, gm_n1641, gm_n1642, gm_n1643, gm_n1644, gm_n1645, gm_n1646, gm_n1647, gm_n1648, gm_n1649, gm_n165, gm_n1650, gm_n1651, gm_n1652, gm_n1653, gm_n1654, gm_n1655, gm_n1656, gm_n1657, gm_n1658, gm_n1659, gm_n166, gm_n1660, gm_n1661, gm_n1662, gm_n1663, gm_n1664, gm_n1665, gm_n1666, gm_n1667, gm_n1668, gm_n1669, gm_n167, gm_n1670, gm_n1671, gm_n1672, gm_n1673, gm_n1674, gm_n1675, gm_n1676, gm_n1677, gm_n1678, gm_n1679, gm_n168, gm_n1680, gm_n1681, gm_n1682, gm_n1683, gm_n1684, gm_n1685, gm_n1686, gm_n1687, gm_n1688, gm_n1689, gm_n169, gm_n1690, gm_n1691, gm_n1692, gm_n1693, gm_n1694, gm_n1695, gm_n1696, gm_n1697, gm_n1698, gm_n1699, gm_n170, gm_n1700, gm_n1701, gm_n1702, gm_n1703, gm_n1704, gm_n1705, gm_n1706, gm_n1707, gm_n1708, gm_n1709, gm_n171, gm_n1710, gm_n1711, gm_n1712, gm_n1713, gm_n1714, gm_n1715, gm_n1716, gm_n1717, gm_n1718, gm_n1719, gm_n172, gm_n1720, gm_n1721, gm_n1722, gm_n1723, gm_n1724, gm_n1725, gm_n1726, gm_n1727, gm_n1728, gm_n1729, gm_n173, gm_n1730, gm_n1731, gm_n1732, gm_n1733, gm_n1734, gm_n1735, gm_n1736, gm_n1737, gm_n1738, gm_n1739, gm_n174, gm_n1740, gm_n1741, gm_n1742, gm_n1743, gm_n1744, gm_n1745, gm_n1746, gm_n1747, gm_n1748, gm_n1749, gm_n175, gm_n1750, gm_n1751, gm_n1752, gm_n1753, gm_n1754, gm_n1755, gm_n1756, gm_n1757, gm_n1758, gm_n1759, gm_n176, gm_n1760, gm_n1761, gm_n1762, gm_n1763, gm_n1764, gm_n1765, gm_n1766, gm_n1767, gm_n1768, gm_n1769, gm_n177, gm_n1770, gm_n1771, gm_n1772, gm_n1773, gm_n1774, gm_n1775, gm_n1776, gm_n1777, gm_n1778, gm_n1779, gm_n178, gm_n1780, gm_n1781, gm_n1782, gm_n1783, gm_n1784, gm_n1785, gm_n1786, gm_n1787, gm_n1788, gm_n1789, gm_n179, gm_n1790, gm_n1791, gm_n1792, gm_n1793, gm_n1794, gm_n1795, gm_n1796, gm_n1797, gm_n1798, gm_n1799, gm_n180, gm_n1800, gm_n1801, gm_n1802, gm_n1803, gm_n1804, gm_n1805, gm_n1806, gm_n1807, gm_n1808, gm_n1809, gm_n181, gm_n1810, gm_n1811, gm_n1812, gm_n1813, gm_n1814, gm_n1816, gm_n1817, gm_n1818, gm_n1819, gm_n182, gm_n1820, gm_n1821, gm_n1822, gm_n1823, gm_n1824, gm_n1825, gm_n1826, gm_n1827, gm_n1828, gm_n1829, gm_n183, gm_n1830, gm_n1831, gm_n1832, gm_n1833, gm_n1834, gm_n1835, gm_n1836, gm_n1837, gm_n1838, gm_n1839, gm_n184, gm_n1840, gm_n1841, gm_n1842, gm_n1843, gm_n1844, gm_n1845, gm_n1846, gm_n1847, gm_n1848, gm_n1849, gm_n185, gm_n1850, gm_n1851, gm_n1852, gm_n1853, gm_n1854, gm_n1855, gm_n1856, gm_n1857, gm_n1858, gm_n1859, gm_n186, gm_n1860, gm_n1861, gm_n1862, gm_n1863, gm_n1864, gm_n1865, gm_n1866, gm_n1867, gm_n1868, gm_n1869, gm_n187, gm_n1870, gm_n1871, gm_n1872, gm_n1873, gm_n1874, gm_n1875, gm_n1876, gm_n1877, gm_n1878, gm_n1879, gm_n188, gm_n1880, gm_n1881, gm_n1882, gm_n1883, gm_n1884, gm_n1885, gm_n1886, gm_n1887, gm_n1888, gm_n1889, gm_n189, gm_n1890, gm_n1891, gm_n1892, gm_n1893, gm_n1894, gm_n1895, gm_n1896, gm_n1897, gm_n1898, gm_n1899, gm_n190, gm_n1900, gm_n1901, gm_n1902, gm_n1903, gm_n1904, gm_n1905, gm_n1906, gm_n1907, gm_n1908, gm_n1909, gm_n191, gm_n1910, gm_n1911, gm_n1912, gm_n1913, gm_n1914, gm_n1915, gm_n1916, gm_n1917, gm_n1918, gm_n1919, gm_n192, gm_n1920, gm_n1921, gm_n1922, gm_n1923, gm_n1924, gm_n1925, gm_n1926, gm_n1927, gm_n1928, gm_n1929, gm_n193, gm_n1930, gm_n1931, gm_n1932, gm_n1933, gm_n1934, gm_n1935, gm_n1936, gm_n1937, gm_n1938, gm_n1939, gm_n194, gm_n1940, gm_n1941, gm_n1942, gm_n1943, gm_n1944, gm_n1945, gm_n1946, gm_n1947, gm_n1948, gm_n1949, gm_n195, gm_n1950, gm_n1951, gm_n1952, gm_n1953, gm_n1954, gm_n1955, gm_n1956, gm_n1957, gm_n1958, gm_n1959, gm_n196, gm_n1960, gm_n1961, gm_n1962, gm_n1963, gm_n1964, gm_n1965, gm_n1966, gm_n1967, gm_n1968, gm_n1969, gm_n197, gm_n1970, gm_n1971, gm_n1972, gm_n1973, gm_n1974, gm_n1975, gm_n1976, gm_n1977, gm_n1978, gm_n1979, gm_n198, gm_n1980, gm_n1981, gm_n1982, gm_n1983, gm_n1984, gm_n1985, gm_n1986, gm_n1987, gm_n1988, gm_n1989, gm_n199, gm_n1990, gm_n1991, gm_n1992, gm_n1993, gm_n1994, gm_n1995, gm_n1996, gm_n1997, gm_n1998, gm_n1999, gm_n200, gm_n2000, gm_n2001, gm_n2002, gm_n2003, gm_n2004, gm_n2005, gm_n2006, gm_n2007, gm_n2008, gm_n201, gm_n2010, gm_n2011, gm_n2012, gm_n2013, gm_n2014, gm_n2015, gm_n2016, gm_n2017, gm_n2018, gm_n2019, gm_n202, gm_n2020, gm_n2021, gm_n2022, gm_n2023, gm_n2024, gm_n2025, gm_n2026, gm_n2027, gm_n2028, gm_n2029, gm_n203, gm_n2030, gm_n2031, gm_n2032, gm_n2033, gm_n2034, gm_n2035, gm_n2036, gm_n2037, gm_n2038, gm_n2039, gm_n204, gm_n2040, gm_n2041, gm_n2042, gm_n2043, gm_n2044, gm_n2045, gm_n2046, gm_n2047, gm_n2048, gm_n2049, gm_n205, gm_n2050, gm_n2051, gm_n2052, gm_n2053, gm_n2054, gm_n2055, gm_n2056, gm_n2057, gm_n2058, gm_n2059, gm_n206, gm_n2060, gm_n2061, gm_n2062, gm_n2063, gm_n2064, gm_n2065, gm_n2066, gm_n2067, gm_n2068, gm_n2069, gm_n207, gm_n2070, gm_n2071, gm_n2072, gm_n2073, gm_n2074, gm_n2075, gm_n2076, gm_n2077, gm_n2078, gm_n2079, gm_n208, gm_n2080, gm_n2081, gm_n2082, gm_n2083, gm_n2084, gm_n2085, gm_n2086, gm_n2087, gm_n2088, gm_n2089, gm_n209, gm_n2090, gm_n2091, gm_n2092, gm_n2093, gm_n2094, gm_n2095, gm_n2096, gm_n2097, gm_n2098, gm_n2099, gm_n210, gm_n2100, gm_n2101, gm_n2102, gm_n2103, gm_n2104, gm_n2105, gm_n2106, gm_n2107, gm_n2108, gm_n2109, gm_n211, gm_n2110, gm_n2111, gm_n2112, gm_n2113, gm_n2114, gm_n2115, gm_n2116, gm_n2117, gm_n2118, gm_n2119, gm_n212, gm_n2120, gm_n2121, gm_n2122, gm_n2123, gm_n2124, gm_n2125, gm_n2126, gm_n2127, gm_n2128, gm_n2129, gm_n213, gm_n2130, gm_n2131, gm_n2132, gm_n2133, gm_n2134, gm_n2135, gm_n2136, gm_n2137, gm_n2138, gm_n2139, gm_n214, gm_n2140, gm_n2141, gm_n2142, gm_n2143, gm_n2144, gm_n2145, gm_n2146, gm_n2147, gm_n2148, gm_n2149, gm_n215, gm_n2150, gm_n2151, gm_n2152, gm_n2153, gm_n2154, gm_n2155, gm_n2156, gm_n2157, gm_n2158, gm_n2159, gm_n216, gm_n2160, gm_n2161, gm_n2162, gm_n2163, gm_n2164, gm_n2165, gm_n2166, gm_n2167, gm_n2168, gm_n2169, gm_n217, gm_n2170, gm_n2171, gm_n2172, gm_n2173, gm_n2174, gm_n2175, gm_n2176, gm_n2177, gm_n2178, gm_n2179, gm_n218, gm_n2180, gm_n2181, gm_n2182, gm_n2183, gm_n2184, gm_n2185, gm_n2186, gm_n2187, gm_n2188, gm_n2189, gm_n219, gm_n2190, gm_n2191, gm_n2192, gm_n2193, gm_n2194, gm_n2195, gm_n2196, gm_n2197, gm_n2198, gm_n2199, gm_n220, gm_n2200, gm_n2201, gm_n2202, gm_n2203, gm_n2205, gm_n2206, gm_n2207, gm_n2208, gm_n2209, gm_n221, gm_n2210, gm_n2211, gm_n2212, gm_n2213, gm_n2214, gm_n2215, gm_n2216, gm_n2217, gm_n2218, gm_n2219, gm_n222, gm_n2220, gm_n2221, gm_n2222, gm_n2223, gm_n2224, gm_n2225, gm_n2226, gm_n2227, gm_n2228, gm_n2229, gm_n223, gm_n2230, gm_n2231, gm_n2232, gm_n2233, gm_n2234, gm_n2235, gm_n2236, gm_n2237, gm_n2238, gm_n2239, gm_n224, gm_n2240, gm_n2241, gm_n2242, gm_n2243, gm_n2244, gm_n2245, gm_n2246, gm_n2247, gm_n2248, gm_n2249, gm_n225, gm_n2250, gm_n2251, gm_n2252, gm_n2253, gm_n2254, gm_n2255, gm_n2256, gm_n2257, gm_n2258, gm_n2259, gm_n226, gm_n2260, gm_n2261, gm_n2262, gm_n2263, gm_n2264, gm_n2265, gm_n2266, gm_n2267, gm_n2268, gm_n2269, gm_n227, gm_n2270, gm_n2271, gm_n2272, gm_n2273, gm_n2274, gm_n2275, gm_n2276, gm_n2277, gm_n2278, gm_n2279, gm_n228, gm_n2280, gm_n2281, gm_n2282, gm_n2283, gm_n2284, gm_n2285, gm_n2286, gm_n2287, gm_n2288, gm_n2289, gm_n229, gm_n2290, gm_n2291, gm_n2292, gm_n2293, gm_n2294, gm_n2295, gm_n2296, gm_n2297, gm_n2298, gm_n2299, gm_n230, gm_n2300, gm_n2301, gm_n2302, gm_n2303, gm_n2304, gm_n2305, gm_n2306, gm_n2307, gm_n2308, gm_n2309, gm_n231, gm_n2310, gm_n2311, gm_n2312, gm_n2313, gm_n2314, gm_n2315, gm_n2316, gm_n2317, gm_n2318, gm_n2319, gm_n232, gm_n2320, gm_n2321, gm_n2322, gm_n2323, gm_n2324, gm_n2325, gm_n2326, gm_n2327, gm_n2328, gm_n2329, gm_n233, gm_n2330, gm_n2331, gm_n2332, gm_n2333, gm_n2334, gm_n2335, gm_n2336, gm_n2337, gm_n2338, gm_n2339, gm_n234, gm_n2340, gm_n2341, gm_n2342, gm_n2343, gm_n2344, gm_n2345, gm_n2346, gm_n2347, gm_n2348, gm_n2349, gm_n235, gm_n2350, gm_n2351, gm_n2352, gm_n2353, gm_n2354, gm_n2355, gm_n2356, gm_n2357, gm_n2358, gm_n2359, gm_n236, gm_n2360, gm_n2361, gm_n2362, gm_n2363, gm_n2364, gm_n2365, gm_n2366, gm_n2367, gm_n2368, gm_n2369, gm_n237, gm_n2370, gm_n2371, gm_n2372, gm_n2373, gm_n2374, gm_n2375, gm_n2376, gm_n2377, gm_n2378, gm_n2379, gm_n238, gm_n2380, gm_n2381, gm_n2382, gm_n2383, gm_n2384, gm_n2385, gm_n2386, gm_n2387, gm_n2388, gm_n239, gm_n2390, gm_n2391, gm_n2392, gm_n2393, gm_n2394, gm_n2395, gm_n2396, gm_n2397, gm_n2398, gm_n2399, gm_n240, gm_n2400, gm_n2401, gm_n2402, gm_n2403, gm_n2404, gm_n2405, gm_n2406, gm_n2407, gm_n2408, gm_n2409, gm_n241, gm_n2410, gm_n2411, gm_n2412, gm_n2413, gm_n2414, gm_n2415, gm_n2416, gm_n2417, gm_n2418, gm_n2419, gm_n242, gm_n2420, gm_n2421, gm_n2422, gm_n2423, gm_n2424, gm_n2425, gm_n2426, gm_n2427, gm_n2428, gm_n2429, gm_n243, gm_n2430, gm_n2431, gm_n2432, gm_n2433, gm_n2434, gm_n2435, gm_n2436, gm_n2437, gm_n2438, gm_n2439, gm_n244, gm_n2440, gm_n2441, gm_n2442, gm_n2443, gm_n2444, gm_n2445, gm_n2446, gm_n2447, gm_n2448, gm_n2449, gm_n245, gm_n2450, gm_n2451, gm_n2452, gm_n2453, gm_n2454, gm_n2455, gm_n2456, gm_n2457, gm_n2458, gm_n2459, gm_n246, gm_n2460, gm_n2461, gm_n2462, gm_n2463, gm_n2464, gm_n2465, gm_n2466, gm_n2467, gm_n2468, gm_n2469, gm_n247, gm_n2470, gm_n2471, gm_n2472, gm_n2473, gm_n2474, gm_n2475, gm_n2476, gm_n2477, gm_n2478, gm_n2479, gm_n248, gm_n2480, gm_n2481, gm_n2482, gm_n2483, gm_n2484, gm_n2485, gm_n2486, gm_n2487, gm_n2488, gm_n2489, gm_n249, gm_n2490, gm_n2491, gm_n2492, gm_n2493, gm_n2494, gm_n2495, gm_n2496, gm_n2497, gm_n2498, gm_n2499, gm_n250, gm_n2500, gm_n2501, gm_n2502, gm_n2503, gm_n2504, gm_n2505, gm_n2506, gm_n2507, gm_n2508, gm_n2509, gm_n251, gm_n2510, gm_n2511, gm_n2512, gm_n2513, gm_n2514, gm_n2515, gm_n2516, gm_n2517, gm_n2518, gm_n2519, gm_n252, gm_n2520, gm_n2521, gm_n2522, gm_n2523, gm_n2524, gm_n2525, gm_n2526, gm_n2527, gm_n2528, gm_n2529, gm_n253, gm_n2530, gm_n2531, gm_n2532, gm_n2533, gm_n2534, gm_n2535, gm_n2536, gm_n2537, gm_n2538, gm_n2539, gm_n254, gm_n2540, gm_n2541, gm_n2542, gm_n2543, gm_n2544, gm_n2545, gm_n2546, gm_n2547, gm_n2548, gm_n2549, gm_n255, gm_n2550, gm_n2551, gm_n2552, gm_n2553, gm_n2554, gm_n2555, gm_n2556, gm_n2557, gm_n2558, gm_n2559, gm_n256, gm_n2560, gm_n2561, gm_n2562, gm_n2563, gm_n2564, gm_n2565, gm_n2566, gm_n2567, gm_n2568, gm_n2569, gm_n257, gm_n2570, gm_n2571, gm_n2572, gm_n2573, gm_n2574, gm_n2575, gm_n2577, gm_n2578, gm_n2579, gm_n258, gm_n2580, gm_n2581, gm_n2582, gm_n2583, gm_n2584, gm_n2585, gm_n2586, gm_n2587, gm_n2588, gm_n2589, gm_n259, gm_n2590, gm_n2591, gm_n2592, gm_n2593, gm_n2594, gm_n2595, gm_n2596, gm_n2597, gm_n2598, gm_n2599, gm_n260, gm_n2600, gm_n2601, gm_n2602, gm_n2603, gm_n2604, gm_n2605, gm_n2606, gm_n2607, gm_n2608, gm_n2609, gm_n261, gm_n2610, gm_n2611, gm_n2612, gm_n2613, gm_n2614, gm_n2615, gm_n2616, gm_n2617, gm_n2618, gm_n2619, gm_n262, gm_n2620, gm_n2621, gm_n2622, gm_n2623, gm_n2624, gm_n2625, gm_n2626, gm_n2627, gm_n2628, gm_n2629, gm_n263, gm_n2630, gm_n2631, gm_n2632, gm_n2633, gm_n2634, gm_n2635, gm_n2636, gm_n2637, gm_n2638, gm_n2639, gm_n264, gm_n2640, gm_n2641, gm_n2642, gm_n2643, gm_n2644, gm_n2645, gm_n2646, gm_n2647, gm_n2648, gm_n2649, gm_n265, gm_n2650, gm_n2651, gm_n2652, gm_n2653, gm_n2654, gm_n2655, gm_n2656, gm_n2657, gm_n2658, gm_n2659, gm_n266, gm_n2660, gm_n2661, gm_n2662, gm_n2663, gm_n2664, gm_n2665, gm_n2666, gm_n2667, gm_n2668, gm_n2669, gm_n267, gm_n2670, gm_n2671, gm_n2672, gm_n2673, gm_n2674, gm_n2675, gm_n2676, gm_n2677, gm_n2678, gm_n2679, gm_n268, gm_n2680, gm_n2681, gm_n2682, gm_n2683, gm_n2684, gm_n2685, gm_n2686, gm_n2687, gm_n2688, gm_n2689, gm_n269, gm_n2690, gm_n2691, gm_n2692, gm_n2693, gm_n2694, gm_n2695, gm_n2696, gm_n2697, gm_n2698, gm_n2699, gm_n270, gm_n2700, gm_n2701, gm_n2702, gm_n2703, gm_n2704, gm_n2705, gm_n2706, gm_n2707, gm_n2708, gm_n2709, gm_n271, gm_n2710, gm_n2711, gm_n2712, gm_n2713, gm_n2714, gm_n2715, gm_n2716, gm_n2717, gm_n2718, gm_n2719, gm_n272, gm_n2720, gm_n2721, gm_n2722, gm_n2723, gm_n2724, gm_n2725, gm_n2726, gm_n2727, gm_n2728, gm_n2729, gm_n273, gm_n2730, gm_n2731, gm_n2732, gm_n2733, gm_n2734, gm_n2735, gm_n2736, gm_n2737, gm_n2738, gm_n2739, gm_n274, gm_n2740, gm_n2741, gm_n2742, gm_n2743, gm_n2744, gm_n2745, gm_n2746, gm_n2747, gm_n2748, gm_n2749, gm_n275, gm_n2750, gm_n2751, gm_n2752, gm_n2753, gm_n2754, gm_n2755, gm_n2756, gm_n2757, gm_n2758, gm_n2759, gm_n276, gm_n2760, gm_n2761, gm_n2762, gm_n2764, gm_n2765, gm_n2766, gm_n2767, gm_n2768, gm_n2769, gm_n277, gm_n2770, gm_n2771, gm_n2772, gm_n2773, gm_n2774, gm_n2775, gm_n2776, gm_n2777, gm_n2778, gm_n2779, gm_n278, gm_n2780, gm_n2781, gm_n2782, gm_n2783, gm_n2784, gm_n2785, gm_n2786, gm_n2787, gm_n2788, gm_n2789, gm_n279, gm_n2790, gm_n2791, gm_n2792, gm_n2793, gm_n2794, gm_n2795, gm_n2796, gm_n2797, gm_n2798, gm_n2799, gm_n280, gm_n2800, gm_n2801, gm_n2802, gm_n2803, gm_n2804, gm_n2805, gm_n2806, gm_n2807, gm_n2808, gm_n2809, gm_n281, gm_n2810, gm_n2811, gm_n2812, gm_n2813, gm_n2814, gm_n2815, gm_n2816, gm_n2817, gm_n2818, gm_n2819, gm_n282, gm_n2820, gm_n2821, gm_n2822, gm_n2823, gm_n2824, gm_n2825, gm_n2826, gm_n2827, gm_n2828, gm_n2829, gm_n283, gm_n2830, gm_n2831, gm_n2832, gm_n2833, gm_n2834, gm_n2835, gm_n2836, gm_n2837, gm_n2838, gm_n2839, gm_n284, gm_n2840, gm_n2841, gm_n2842, gm_n2843, gm_n2844, gm_n2845, gm_n2846, gm_n2847, gm_n2848, gm_n2849, gm_n285, gm_n2850, gm_n2851, gm_n2852, gm_n2853, gm_n2854, gm_n2855, gm_n2856, gm_n2857, gm_n2858, gm_n2859, gm_n286, gm_n2860, gm_n2861, gm_n2862, gm_n2863, gm_n2864, gm_n2865, gm_n2866, gm_n2867, gm_n2868, gm_n2869, gm_n287, gm_n2870, gm_n2871, gm_n2872, gm_n2873, gm_n2874, gm_n2875, gm_n2876, gm_n2877, gm_n2878, gm_n2879, gm_n288, gm_n2880, gm_n2881, gm_n2882, gm_n2883, gm_n2884, gm_n2885, gm_n2886, gm_n2887, gm_n2888, gm_n2889, gm_n289, gm_n2890, gm_n2891, gm_n2892, gm_n2893, gm_n2894, gm_n2895, gm_n2896, gm_n2897, gm_n2898, gm_n2899, gm_n290, gm_n2900, gm_n2901, gm_n2902, gm_n2903, gm_n2904, gm_n2905, gm_n2906, gm_n2907, gm_n2908, gm_n2909, gm_n291, gm_n2910, gm_n2911, gm_n2912, gm_n2913, gm_n2914, gm_n2915, gm_n2916, gm_n2917, gm_n2918, gm_n2919, gm_n292, gm_n2920, gm_n2921, gm_n2922, gm_n2923, gm_n2924, gm_n2925, gm_n2926, gm_n2927, gm_n2928, gm_n2929, gm_n293, gm_n2930, gm_n2931, gm_n2932, gm_n2933, gm_n2934, gm_n2935, gm_n2936, gm_n2937, gm_n2938, gm_n2939, gm_n294, gm_n2940, gm_n2941, gm_n2942, gm_n2943, gm_n2944, gm_n2945, gm_n2946, gm_n2947, gm_n2948, gm_n2949, gm_n295, gm_n2950, gm_n2951, gm_n2952, gm_n2953, gm_n2954, gm_n2955, gm_n2956, gm_n2957, gm_n2958, gm_n2959, gm_n296, gm_n2960, gm_n2961, gm_n2962, gm_n2963, gm_n2964, gm_n2965, gm_n2966, gm_n2967, gm_n2968, gm_n2969, gm_n297, gm_n2970, gm_n2971, gm_n2972, gm_n2973, gm_n2974, gm_n2975, gm_n2976, gm_n2977, gm_n2978, gm_n2979, gm_n298, gm_n2980, gm_n2981, gm_n2982, gm_n2983, gm_n2984, gm_n2985, gm_n2986, gm_n2987, gm_n2988, gm_n2989, gm_n299, gm_n2990, gm_n2991, gm_n2992, gm_n2993, gm_n2994, gm_n2995, gm_n2996, gm_n2997, gm_n2998, gm_n2999, gm_n300, gm_n3000, gm_n3001, gm_n3002, gm_n3003, gm_n3004, gm_n3005, gm_n3006, gm_n3007, gm_n3008, gm_n3009, gm_n301, gm_n3010, gm_n3011, gm_n3012, gm_n3013, gm_n3014, gm_n3015, gm_n3016, gm_n3017, gm_n3018, gm_n3019, gm_n302, gm_n3020, gm_n3021, gm_n3022, gm_n3023, gm_n3024, gm_n3025, gm_n3026, gm_n3027, gm_n3028, gm_n3029, gm_n303, gm_n3030, gm_n3031, gm_n3032, gm_n3033, gm_n3034, gm_n3035, gm_n3036, gm_n3037, gm_n3038, gm_n3039, gm_n304, gm_n3040, gm_n3041, gm_n3042, gm_n3043, gm_n3044, gm_n3045, gm_n3046, gm_n3047, gm_n3048, gm_n3049, gm_n305, gm_n3050, gm_n3051, gm_n3052, gm_n3053, gm_n3054, gm_n3055, gm_n3056, gm_n3057, gm_n3058, gm_n3059, gm_n306, gm_n3060, gm_n3061, gm_n3062, gm_n3063, gm_n3064, gm_n3065, gm_n3066, gm_n3067, gm_n3068, gm_n3069, gm_n307, gm_n3070, gm_n3071, gm_n3072, gm_n3073, gm_n3074, gm_n3075, gm_n3076, gm_n3077, gm_n3078, gm_n3079, gm_n308, gm_n3080, gm_n3081, gm_n3082, gm_n3083, gm_n3084, gm_n3085, gm_n3086, gm_n3087, gm_n3088, gm_n3089, gm_n309, gm_n3090, gm_n3091, gm_n3092, gm_n3093, gm_n3094, gm_n3095, gm_n3096, gm_n3097, gm_n3098, gm_n3099, gm_n310, gm_n3100, gm_n3101, gm_n3102, gm_n3103, gm_n3104, gm_n3105, gm_n3106, gm_n3107, gm_n3108, gm_n3109, gm_n311, gm_n3110, gm_n3111, gm_n3112, gm_n3113, gm_n3114, gm_n3115, gm_n3116, gm_n3117, gm_n3118, gm_n3119, gm_n312, gm_n3120, gm_n3121, gm_n3123, gm_n3124, gm_n3125, gm_n3126, gm_n3127, gm_n3128, gm_n3129, gm_n313, gm_n3130, gm_n3131, gm_n3132, gm_n3133, gm_n3134, gm_n3135, gm_n3136, gm_n3137, gm_n3138, gm_n3139, gm_n314, gm_n3140, gm_n3141, gm_n3142, gm_n3143, gm_n3144, gm_n3145, gm_n3146, gm_n3147, gm_n3148, gm_n3149, gm_n315, gm_n3150, gm_n3151, gm_n3152, gm_n3153, gm_n3154, gm_n3155, gm_n3156, gm_n3157, gm_n3158, gm_n3159, gm_n316, gm_n3160, gm_n3161, gm_n3162, gm_n3163, gm_n3164, gm_n3165, gm_n3166, gm_n3167, gm_n3168, gm_n3169, gm_n317, gm_n3170, gm_n3171, gm_n3172, gm_n3173, gm_n3174, gm_n3175, gm_n3176, gm_n3177, gm_n3178, gm_n3179, gm_n318, gm_n3180, gm_n3181, gm_n3182, gm_n3183, gm_n3184, gm_n3185, gm_n3186, gm_n3187, gm_n3188, gm_n3189, gm_n319, gm_n3190, gm_n3191, gm_n3192, gm_n3193, gm_n3194, gm_n3195, gm_n3196, gm_n3197, gm_n3198, gm_n3199, gm_n320, gm_n3200, gm_n3201, gm_n3202, gm_n3203, gm_n3204, gm_n3205, gm_n3206, gm_n3207, gm_n3208, gm_n3209, gm_n321, gm_n3210, gm_n3211, gm_n3212, gm_n3213, gm_n3214, gm_n3215, gm_n3216, gm_n3217, gm_n3218, gm_n3219, gm_n322, gm_n3220, gm_n3221, gm_n3222, gm_n3223, gm_n3224, gm_n3225, gm_n3226, gm_n3227, gm_n3228, gm_n3229, gm_n323, gm_n3230, gm_n3231, gm_n3232, gm_n3233, gm_n3234, gm_n3235, gm_n3236, gm_n3237, gm_n3238, gm_n3239, gm_n324, gm_n3240, gm_n3241, gm_n3242, gm_n3243, gm_n3244, gm_n3245, gm_n3246, gm_n3247, gm_n3248, gm_n3249, gm_n325, gm_n3250, gm_n3251, gm_n3252, gm_n3253, gm_n3254, gm_n3255, gm_n3256, gm_n3257, gm_n3258, gm_n3259, gm_n326, gm_n3260, gm_n3261, gm_n3262, gm_n3263, gm_n3264, gm_n3265, gm_n3266, gm_n3267, gm_n3268, gm_n3269, gm_n327, gm_n3270, gm_n3271, gm_n3272, gm_n3273, gm_n3274, gm_n3275, gm_n3276, gm_n3277, gm_n3278, gm_n3279, gm_n328, gm_n3280, gm_n3281, gm_n3282, gm_n3283, gm_n3284, gm_n3285, gm_n3286, gm_n3287, gm_n3288, gm_n3289, gm_n329, gm_n3290, gm_n3291, gm_n3292, gm_n3293, gm_n3294, gm_n3295, gm_n3296, gm_n3297, gm_n3298, gm_n3299, gm_n330, gm_n3300, gm_n3301, gm_n3302, gm_n3303, gm_n3304, gm_n3305, gm_n3306, gm_n3307, gm_n3308, gm_n3309, gm_n331, gm_n3310, gm_n3311, gm_n3312, gm_n3313, gm_n3314, gm_n3315, gm_n3316, gm_n3317, gm_n3318, gm_n3319, gm_n332, gm_n3320, gm_n3321, gm_n3322, gm_n3323, gm_n3324, gm_n3325, gm_n3326, gm_n3327, gm_n3328, gm_n3329, gm_n333, gm_n3330, gm_n3331, gm_n3332, gm_n3333, gm_n3334, gm_n3335, gm_n3336, gm_n3337, gm_n3338, gm_n3339, gm_n334, gm_n3340, gm_n3341, gm_n3342, gm_n3343, gm_n3344, gm_n3345, gm_n3346, gm_n3347, gm_n3348, gm_n3349, gm_n335, gm_n3350, gm_n3351, gm_n3352, gm_n3353, gm_n3354, gm_n3355, gm_n3356, gm_n3357, gm_n3358, gm_n3359, gm_n336, gm_n3360, gm_n3361, gm_n3362, gm_n3363, gm_n3364, gm_n3365, gm_n3366, gm_n3367, gm_n3368, gm_n3369, gm_n337, gm_n3370, gm_n3371, gm_n3372, gm_n3373, gm_n3374, gm_n3375, gm_n3376, gm_n3377, gm_n3378, gm_n3379, gm_n338, gm_n3380, gm_n3381, gm_n3382, gm_n3383, gm_n3384, gm_n3385, gm_n3386, gm_n3387, gm_n3388, gm_n3389, gm_n339, gm_n3390, gm_n3391, gm_n3392, gm_n3393, gm_n3394, gm_n3395, gm_n3396, gm_n3397, gm_n3398, gm_n3399, gm_n340, gm_n3400, gm_n3401, gm_n3402, gm_n3403, gm_n3404, gm_n3405, gm_n3406, gm_n3407, gm_n3408, gm_n3409, gm_n341, gm_n3410, gm_n3411, gm_n3412, gm_n3413, gm_n3414, gm_n3415, gm_n3416, gm_n3417, gm_n3418, gm_n3419, gm_n342, gm_n3420, gm_n3421, gm_n3422, gm_n3423, gm_n3424, gm_n3425, gm_n3426, gm_n3427, gm_n3428, gm_n3429, gm_n343, gm_n3430, gm_n3431, gm_n3432, gm_n3433, gm_n3434, gm_n3435, gm_n3436, gm_n3437, gm_n3438, gm_n3439, gm_n344, gm_n3440, gm_n3441, gm_n3442, gm_n3443, gm_n3444, gm_n3445, gm_n3446, gm_n3447, gm_n3448, gm_n3449, gm_n345, gm_n3450, gm_n3451, gm_n3452, gm_n3453, gm_n3454, gm_n3455, gm_n3456, gm_n3457, gm_n3458, gm_n3459, gm_n346, gm_n3460, gm_n3461, gm_n3462, gm_n3463, gm_n3464, gm_n3465, gm_n3466, gm_n3467, gm_n3468, gm_n3469, gm_n347, gm_n3470, gm_n3471, gm_n3472, gm_n3473, gm_n3474, gm_n3475, gm_n3476, gm_n3477, gm_n3478, gm_n348, gm_n3480, gm_n3481, gm_n3482, gm_n3483, gm_n3484, gm_n3485, gm_n3486, gm_n3487, gm_n3488, gm_n3489, gm_n349, gm_n3490, gm_n3491, gm_n3492, gm_n3493, gm_n3494, gm_n3495, gm_n3496, gm_n3497, gm_n3498, gm_n3499, gm_n350, gm_n3500, gm_n3501, gm_n3502, gm_n3503, gm_n3504, gm_n3505, gm_n3506, gm_n3507, gm_n3508, gm_n3509, gm_n351, gm_n3510, gm_n3511, gm_n3512, gm_n3513, gm_n3514, gm_n3515, gm_n3516, gm_n3517, gm_n3518, gm_n3519, gm_n352, gm_n3520, gm_n3521, gm_n3522, gm_n3523, gm_n3524, gm_n3525, gm_n3526, gm_n3527, gm_n3528, gm_n3529, gm_n353, gm_n3530, gm_n3531, gm_n3532, gm_n3533, gm_n3534, gm_n3535, gm_n3536, gm_n3537, gm_n3538, gm_n3539, gm_n354, gm_n3540, gm_n3541, gm_n3542, gm_n3543, gm_n3544, gm_n3545, gm_n3546, gm_n3547, gm_n3548, gm_n3549, gm_n355, gm_n3550, gm_n3551, gm_n3552, gm_n3553, gm_n3554, gm_n3555, gm_n3556, gm_n3557, gm_n3558, gm_n3559, gm_n356, gm_n3560, gm_n3561, gm_n3562, gm_n3563, gm_n3564, gm_n3565, gm_n3566, gm_n3567, gm_n3568, gm_n3569, gm_n357, gm_n3570, gm_n3571, gm_n3572, gm_n3573, gm_n3574, gm_n3575, gm_n3576, gm_n3577, gm_n3578, gm_n3579, gm_n358, gm_n3580, gm_n3581, gm_n3582, gm_n3583, gm_n3584, gm_n3585, gm_n3586, gm_n3587, gm_n3588, gm_n3589, gm_n359, gm_n3590, gm_n3591, gm_n3592, gm_n3593, gm_n3594, gm_n3595, gm_n3596, gm_n3597, gm_n3598, gm_n3599, gm_n360, gm_n3600, gm_n3601, gm_n3602, gm_n3603, gm_n3604, gm_n3605, gm_n3606, gm_n3607, gm_n3608, gm_n3609, gm_n361, gm_n3610, gm_n3611, gm_n3612, gm_n3613, gm_n3614, gm_n3615, gm_n3616, gm_n3617, gm_n3618, gm_n3619, gm_n362, gm_n3620, gm_n3621, gm_n3622, gm_n3623, gm_n3624, gm_n3625, gm_n3626, gm_n3627, gm_n3628, gm_n3629, gm_n363, gm_n3630, gm_n3631, gm_n3632, gm_n3633, gm_n3634, gm_n3635, gm_n3636, gm_n3637, gm_n3638, gm_n3639, gm_n364, gm_n3640, gm_n3641, gm_n3642, gm_n3643, gm_n3644, gm_n3645, gm_n3646, gm_n3647, gm_n3648, gm_n3649, gm_n365, gm_n3650, gm_n3651, gm_n3652, gm_n3653, gm_n3654, gm_n3655, gm_n3656, gm_n3657, gm_n3658, gm_n3659, gm_n366, gm_n3660, gm_n3661, gm_n3662, gm_n3663, gm_n3664, gm_n3665, gm_n3666, gm_n3667, gm_n3668, gm_n3669, gm_n367, gm_n3670, gm_n3671, gm_n3672, gm_n3673, gm_n3674, gm_n3675, gm_n3676, gm_n3677, gm_n3678, gm_n3679, gm_n368, gm_n3680, gm_n3681, gm_n3682, gm_n3683, gm_n3684, gm_n3685, gm_n3686, gm_n3687, gm_n3688, gm_n3689, gm_n369, gm_n3690, gm_n3691, gm_n3692, gm_n3693, gm_n3694, gm_n3695, gm_n3696, gm_n3697, gm_n3698, gm_n3699, gm_n370, gm_n3700, gm_n3701, gm_n3702, gm_n3703, gm_n3704, gm_n3705, gm_n3706, gm_n3707, gm_n3708, gm_n3709, gm_n371, gm_n3710, gm_n3711, gm_n3712, gm_n3713, gm_n3714, gm_n3715, gm_n3716, gm_n3717, gm_n3718, gm_n3719, gm_n372, gm_n3720, gm_n3721, gm_n3722, gm_n3723, gm_n3724, gm_n3725, gm_n3726, gm_n3727, gm_n3728, gm_n3729, gm_n373, gm_n3730, gm_n3731, gm_n3732, gm_n3733, gm_n3734, gm_n3735, gm_n3736, gm_n3737, gm_n3738, gm_n3739, gm_n374, gm_n3740, gm_n3741, gm_n3742, gm_n3743, gm_n3744, gm_n3745, gm_n3746, gm_n3747, gm_n3748, gm_n3749, gm_n375, gm_n3750, gm_n3751, gm_n3752, gm_n3753, gm_n3754, gm_n3755, gm_n3756, gm_n3757, gm_n3758, gm_n3759, gm_n376, gm_n3760, gm_n3761, gm_n3762, gm_n3763, gm_n3764, gm_n3765, gm_n3766, gm_n3767, gm_n3768, gm_n3769, gm_n377, gm_n3770, gm_n3771, gm_n3772, gm_n3773, gm_n3774, gm_n3775, gm_n3776, gm_n3777, gm_n3778, gm_n3779, gm_n378, gm_n3780, gm_n3781, gm_n3782, gm_n3783, gm_n3784, gm_n3785, gm_n3786, gm_n3787, gm_n3788, gm_n3789, gm_n379, gm_n3790, gm_n3791, gm_n3792, gm_n3793, gm_n3794, gm_n3795, gm_n3796, gm_n3797, gm_n3798, gm_n3799, gm_n380, gm_n3800, gm_n3801, gm_n3802, gm_n3803, gm_n3804, gm_n3805, gm_n3806, gm_n3807, gm_n3808, gm_n3809, gm_n381, gm_n3810, gm_n3811, gm_n3812, gm_n3813, gm_n3814, gm_n3815, gm_n3816, gm_n3817, gm_n3818, gm_n3819, gm_n382, gm_n3820, gm_n3821, gm_n3822, gm_n3823, gm_n3824, gm_n3825, gm_n3826, gm_n3827, gm_n3828, gm_n3829, gm_n383, gm_n3830, gm_n3831, gm_n3832, gm_n3833, gm_n3834, gm_n3835, gm_n3836, gm_n3837, gm_n3838, gm_n3839, gm_n384, gm_n3840, gm_n3841, gm_n3842, gm_n3843, gm_n3844, gm_n3846, gm_n3847, gm_n3848, gm_n3849, gm_n385, gm_n3850, gm_n3851, gm_n3852, gm_n3853, gm_n3854, gm_n3855, gm_n3856, gm_n3857, gm_n3858, gm_n3859, gm_n386, gm_n3860, gm_n3861, gm_n3862, gm_n3863, gm_n3864, gm_n3865, gm_n3866, gm_n3867, gm_n3868, gm_n3869, gm_n387, gm_n3870, gm_n3871, gm_n3872, gm_n3873, gm_n3874, gm_n3875, gm_n3876, gm_n3877, gm_n3878, gm_n3879, gm_n388, gm_n3880, gm_n3881, gm_n3882, gm_n3883, gm_n3884, gm_n3885, gm_n3886, gm_n3887, gm_n3888, gm_n3889, gm_n389, gm_n3890, gm_n3891, gm_n3892, gm_n3893, gm_n3894, gm_n3895, gm_n3896, gm_n3897, gm_n3898, gm_n3899, gm_n390, gm_n3900, gm_n3901, gm_n3902, gm_n3903, gm_n3904, gm_n3905, gm_n3906, gm_n3907, gm_n3908, gm_n3909, gm_n391, gm_n3910, gm_n3911, gm_n3912, gm_n3913, gm_n3914, gm_n3915, gm_n3916, gm_n3917, gm_n3918, gm_n3919, gm_n392, gm_n3920, gm_n3921, gm_n3922, gm_n3923, gm_n3924, gm_n3925, gm_n3926, gm_n3927, gm_n3928, gm_n3929, gm_n393, gm_n3930, gm_n3931, gm_n3932, gm_n3933, gm_n3934, gm_n3935, gm_n3936, gm_n3937, gm_n3938, gm_n3939, gm_n394, gm_n3940, gm_n3941, gm_n3942, gm_n3943, gm_n3944, gm_n3945, gm_n3946, gm_n3947, gm_n3948, gm_n3949, gm_n395, gm_n3950, gm_n3951, gm_n3952, gm_n3953, gm_n3954, gm_n3955, gm_n3956, gm_n3957, gm_n3958, gm_n3959, gm_n396, gm_n3960, gm_n3961, gm_n3962, gm_n3963, gm_n3964, gm_n3965, gm_n3966, gm_n3967, gm_n3968, gm_n3969, gm_n397, gm_n3970, gm_n3971, gm_n3972, gm_n3973, gm_n3974, gm_n3975, gm_n3976, gm_n3977, gm_n3978, gm_n3979, gm_n398, gm_n3980, gm_n3981, gm_n3982, gm_n3983, gm_n3984, gm_n3985, gm_n3986, gm_n3987, gm_n3988, gm_n3989, gm_n399, gm_n3990, gm_n3991, gm_n3992, gm_n3993, gm_n3994, gm_n3995, gm_n3996, gm_n3997, gm_n3998, gm_n3999, gm_n400, gm_n4000, gm_n4001, gm_n4002, gm_n4003, gm_n4004, gm_n4005, gm_n4006, gm_n4007, gm_n4008, gm_n4009, gm_n401, gm_n4010, gm_n4011, gm_n4012, gm_n4013, gm_n4014, gm_n4015, gm_n4016, gm_n4017, gm_n4018, gm_n4019, gm_n402, gm_n4020, gm_n4021, gm_n4022, gm_n4023, gm_n4024, gm_n4025, gm_n4026, gm_n4027, gm_n4028, gm_n4029, gm_n403, gm_n4030, gm_n4031, gm_n4032, gm_n4033, gm_n4034, gm_n4035, gm_n4036, gm_n4037, gm_n4038, gm_n4039, gm_n404, gm_n4040, gm_n4041, gm_n4042, gm_n4043, gm_n4044, gm_n4045, gm_n4046, gm_n4047, gm_n4048, gm_n4049, gm_n405, gm_n4050, gm_n4051, gm_n4052, gm_n4053, gm_n4054, gm_n4055, gm_n4056, gm_n4057, gm_n4058, gm_n4059, gm_n406, gm_n4060, gm_n4061, gm_n4062, gm_n4063, gm_n4064, gm_n4065, gm_n4066, gm_n4067, gm_n4068, gm_n4069, gm_n407, gm_n4070, gm_n4071, gm_n4072, gm_n4073, gm_n4074, gm_n4075, gm_n4076, gm_n4077, gm_n4078, gm_n4079, gm_n408, gm_n4080, gm_n4081, gm_n4082, gm_n4083, gm_n4084, gm_n4085, gm_n4086, gm_n4087, gm_n4088, gm_n4089, gm_n409, gm_n4090, gm_n4091, gm_n4092, gm_n4093, gm_n4094, gm_n4095, gm_n4096, gm_n4097, gm_n4098, gm_n4099, gm_n410, gm_n4100, gm_n4101, gm_n4102, gm_n4103, gm_n4104, gm_n4105, gm_n4106, gm_n4107, gm_n4108, gm_n4109, gm_n411, gm_n4110, gm_n4111, gm_n4112, gm_n4113, gm_n4114, gm_n4115, gm_n4116, gm_n4117, gm_n4118, gm_n4119, gm_n412, gm_n4120, gm_n4121, gm_n4122, gm_n4123, gm_n4124, gm_n4125, gm_n4126, gm_n4127, gm_n4128, gm_n4129, gm_n413, gm_n4130, gm_n4131, gm_n4132, gm_n4133, gm_n4134, gm_n4135, gm_n4136, gm_n4137, gm_n4138, gm_n4139, gm_n414, gm_n4140, gm_n4141, gm_n4142, gm_n4143, gm_n4144, gm_n4145, gm_n4146, gm_n4147, gm_n4148, gm_n4149, gm_n415, gm_n4150, gm_n4151, gm_n4152, gm_n4153, gm_n4154, gm_n4155, gm_n4156, gm_n4157, gm_n4158, gm_n4159, gm_n416, gm_n4160, gm_n4161, gm_n4162, gm_n4163, gm_n4164, gm_n4165, gm_n4166, gm_n4167, gm_n4168, gm_n4169, gm_n417, gm_n4170, gm_n4171, gm_n4172, gm_n4173, gm_n4174, gm_n4175, gm_n4176, gm_n4177, gm_n4178, gm_n4179, gm_n418, gm_n4180, gm_n4181, gm_n4182, gm_n4183, gm_n4184, gm_n4185, gm_n4186, gm_n4187, gm_n4188, gm_n4189, gm_n419, gm_n4190, gm_n4191, gm_n4192, gm_n4193, gm_n4194, gm_n4196, gm_n420, gm_n421, gm_n422, gm_n423, gm_n424, gm_n425, gm_n426, gm_n427, gm_n428, gm_n429, gm_n430, gm_n431, gm_n432, gm_n433, gm_n434, gm_n435, gm_n436, gm_n437, gm_n438, gm_n439, gm_n440, gm_n441, gm_n442, gm_n443, gm_n444, gm_n445, gm_n446, gm_n447, gm_n448, gm_n449, gm_n450, gm_n451, gm_n452, gm_n453, gm_n454, gm_n455, gm_n456, gm_n457, gm_n458, gm_n459, gm_n460, gm_n461, gm_n462, gm_n463, gm_n464, gm_n465, gm_n466, gm_n467, gm_n468, gm_n469, gm_n470, gm_n471, gm_n472, gm_n473, gm_n474, gm_n475, gm_n476, gm_n477, gm_n478, gm_n479, gm_n480, gm_n481, gm_n482, gm_n483, gm_n484, gm_n485, gm_n486, gm_n487, gm_n488, gm_n489, gm_n490, gm_n491, gm_n492, gm_n493, gm_n494, gm_n495, gm_n496, gm_n497, gm_n498, gm_n499, gm_n50, gm_n500, gm_n501, gm_n502, gm_n504, gm_n505, gm_n506, gm_n507, gm_n508, gm_n509, gm_n51, gm_n510, gm_n511, gm_n512, gm_n513, gm_n514, gm_n515, gm_n516, gm_n517, gm_n518, gm_n519, gm_n52, gm_n520, gm_n521, gm_n522, gm_n523, gm_n524, gm_n525, gm_n526, gm_n527, gm_n528, gm_n529, gm_n53, gm_n530, gm_n531, gm_n532, gm_n533, gm_n534, gm_n535, gm_n536, gm_n537, gm_n538, gm_n539, gm_n54, gm_n540, gm_n541, gm_n542, gm_n543, gm_n544, gm_n545, gm_n546, gm_n547, gm_n548, gm_n549, gm_n55, gm_n550, gm_n551, gm_n552, gm_n553, gm_n554, gm_n555, gm_n556, gm_n557, gm_n558, gm_n559, gm_n56, gm_n560, gm_n561, gm_n562, gm_n563, gm_n564, gm_n565, gm_n566, gm_n567, gm_n568, gm_n569, gm_n57, gm_n570, gm_n571, gm_n572, gm_n573, gm_n574, gm_n575, gm_n576, gm_n577, gm_n578, gm_n579, gm_n58, gm_n580, gm_n581, gm_n582, gm_n583, gm_n584, gm_n585, gm_n586, gm_n587, gm_n588, gm_n589, gm_n59, gm_n590, gm_n591, gm_n592, gm_n593, gm_n594, gm_n595, gm_n596, gm_n597, gm_n598, gm_n599, gm_n60, gm_n600, gm_n601, gm_n602, gm_n603, gm_n604, gm_n605, gm_n606, gm_n607, gm_n608, gm_n609, gm_n61, gm_n610, gm_n611, gm_n612, gm_n613, gm_n614, gm_n615, gm_n616, gm_n617, gm_n618, gm_n619, gm_n62, gm_n620, gm_n621, gm_n622, gm_n623, gm_n624, gm_n625, gm_n626, gm_n627, gm_n628, gm_n629, gm_n63, gm_n630, gm_n631, gm_n632, gm_n633, gm_n634, gm_n635, gm_n636, gm_n637, gm_n638, gm_n639, gm_n64, gm_n640, gm_n641, gm_n642, gm_n643, gm_n644, gm_n645, gm_n646, gm_n647, gm_n648, gm_n649, gm_n65, gm_n650, gm_n651, gm_n652, gm_n653, gm_n654, gm_n655, gm_n656, gm_n657, gm_n658, gm_n659, gm_n66, gm_n660, gm_n661, gm_n662, gm_n663, gm_n664, gm_n665, gm_n666, gm_n667, gm_n668, gm_n669, gm_n67, gm_n670, gm_n671, gm_n672, gm_n673, gm_n674, gm_n675, gm_n676, gm_n677, gm_n678, gm_n679, gm_n68, gm_n680, gm_n681, gm_n682, gm_n683, gm_n684, gm_n685, gm_n686, gm_n687, gm_n688, gm_n689, gm_n69, gm_n690, gm_n691, gm_n692, gm_n693, gm_n694, gm_n695, gm_n696, gm_n697, gm_n698, gm_n699, gm_n70, gm_n700, gm_n701, gm_n702, gm_n703, gm_n704, gm_n705, gm_n706, gm_n707, gm_n708, gm_n709, gm_n71, gm_n710, gm_n711, gm_n712, gm_n713, gm_n714, gm_n715, gm_n716, gm_n717, gm_n718, gm_n719, gm_n72, gm_n720, gm_n721, gm_n722, gm_n723, gm_n724, gm_n725, gm_n726, gm_n727, gm_n728, gm_n729, gm_n73, gm_n730, gm_n731, gm_n732, gm_n733, gm_n734, gm_n735, gm_n736, gm_n737, gm_n738, gm_n739, gm_n74, gm_n740, gm_n741, gm_n742, gm_n743, gm_n744, gm_n745, gm_n746, gm_n747, gm_n748, gm_n749, gm_n75, gm_n750, gm_n751, gm_n752, gm_n753, gm_n754, gm_n755, gm_n756, gm_n757, gm_n758, gm_n759, gm_n76, gm_n760, gm_n761, gm_n762, gm_n763, gm_n764, gm_n765, gm_n766, gm_n767, gm_n768, gm_n769, gm_n77, gm_n770, gm_n771, gm_n772, gm_n773, gm_n774, gm_n775, gm_n776, gm_n777, gm_n778, gm_n78, gm_n780, gm_n781, gm_n782, gm_n783, gm_n784, gm_n785, gm_n786, gm_n787, gm_n788, gm_n789, gm_n79, gm_n790, gm_n791, gm_n792, gm_n793, gm_n794, gm_n795, gm_n796, gm_n797, gm_n798, gm_n799, gm_n80, gm_n800, gm_n801, gm_n802, gm_n803, gm_n804, gm_n805, gm_n806, gm_n807, gm_n808, gm_n809, gm_n81, gm_n810, gm_n811, gm_n812, gm_n813, gm_n814, gm_n815, gm_n816, gm_n817, gm_n818, gm_n819, gm_n82, gm_n820, gm_n821, gm_n822, gm_n823, gm_n824, gm_n825, gm_n826, gm_n827, gm_n828, gm_n829, gm_n83, gm_n830, gm_n831, gm_n832, gm_n833, gm_n834, gm_n835, gm_n836, gm_n837, gm_n838, gm_n839, gm_n84, gm_n840, gm_n841, gm_n842, gm_n843, gm_n844, gm_n845, gm_n846, gm_n847, gm_n848, gm_n849, gm_n85, gm_n850, gm_n851, gm_n852, gm_n853, gm_n854, gm_n855, gm_n856, gm_n857, gm_n858, gm_n859, gm_n86, gm_n860, gm_n861, gm_n862, gm_n863, gm_n864, gm_n865, gm_n866, gm_n867, gm_n868, gm_n869, gm_n87, gm_n870, gm_n871, gm_n872, gm_n873, gm_n874, gm_n875, gm_n876, gm_n877, gm_n878, gm_n879, gm_n88, gm_n880, gm_n881, gm_n882, gm_n883, gm_n884, gm_n885, gm_n886, gm_n887, gm_n888, gm_n889, gm_n89, gm_n890, gm_n891, gm_n892, gm_n893, gm_n894, gm_n895, gm_n896, gm_n897, gm_n898, gm_n899, gm_n90, gm_n900, gm_n901, gm_n902, gm_n903, gm_n904, gm_n905, gm_n906, gm_n907, gm_n908, gm_n909, gm_n91, gm_n910, gm_n911, gm_n912, gm_n913, gm_n914, gm_n915, gm_n916, gm_n917, gm_n918, gm_n919, gm_n92, gm_n920, gm_n921, gm_n922, gm_n923, gm_n924, gm_n925, gm_n926, gm_n927, gm_n928, gm_n929, gm_n93, gm_n930, gm_n931, gm_n932, gm_n933, gm_n934, gm_n935, gm_n936, gm_n937, gm_n938, gm_n939, gm_n94, gm_n940, gm_n941, gm_n942, gm_n943, gm_n944, gm_n945, gm_n946, gm_n947, gm_n948, gm_n949, gm_n95, gm_n950, gm_n951, gm_n952, gm_n953, gm_n954, gm_n955, gm_n956, gm_n957, gm_n958, gm_n959, gm_n96, gm_n960, gm_n961, gm_n962, gm_n963, gm_n964, gm_n965, gm_n966, gm_n967, gm_n968, gm_n969, gm_n97, gm_n970, gm_n971, gm_n972, gm_n973, gm_n974, gm_n975, gm_n976, gm_n977, gm_n978, gm_n979, gm_n98, gm_n980, gm_n981, gm_n982, gm_n983, gm_n984, gm_n985, gm_n986, gm_n987, gm_n988, gm_n989, gm_n99, gm_n990, gm_n991, gm_n992, gm_n993, gm_n994, gm_n995, gm_n997, gm_n998, gm_n999;
	not (gm_n50, in_31);
	nand (gm_n51, in_30, in_29, in_28);
	not (gm_n52, in_24);
	not (gm_n53, in_25);
	nand (gm_n54, in_26, gm_n53, gm_n52);
	not (gm_n55, gm_n54);
	not (gm_n56, in_13);
	nand (gm_n57, in_14, gm_n56, in_12);
	not (gm_n58, in_11);
	not (gm_n59, in_1);
	not (gm_n60, in_3);
	nor (gm_n61, in_2, gm_n59, in_0, in_4, gm_n60);
	not (gm_n62, in_5);
	nor (gm_n63, in_7, in_6, gm_n62);
	not (gm_n64, in_8);
	not (gm_n65, in_9);
	nor (gm_n66, in_10, gm_n65, gm_n64);
	nand (gm_n67, gm_n63, gm_n61, gm_n58, gm_n66);
	not (gm_n68, in_16);
	nor (gm_n69, in_18, in_17, gm_n68);
	not (gm_n70, gm_n69);
	nor (gm_n71, gm_n57, in_19, in_15, gm_n70, gm_n67);
	not (gm_n72, in_20);
	nor (gm_n73, in_22, in_21, gm_n72);
	nand (gm_n74, gm_n55, in_27, in_23, gm_n73, gm_n71);
	nor (gm_n75, gm_n74, gm_n51, gm_n50);
	not (gm_n76, in_29);
	nor (gm_n77, gm_n50, in_30, gm_n76);
	not (gm_n78, in_28);
	nor (gm_n79, in_27, in_26, in_25);
	not (gm_n80, gm_n79);
	not (gm_n81, in_21);
	not (gm_n82, in_22);
	nor (gm_n83, in_23, gm_n82, gm_n81);
	not (gm_n84, gm_n83);
	nor (gm_n85, in_19, in_18, in_17);
	and (gm_n86, in_15, in_14, in_13);
	not (gm_n87, in_10);
	nand (gm_n88, gm_n58, gm_n87, in_9);
	nand (gm_n89, in_7, in_6, gm_n62);
	not (gm_n90, in_0);
	nand (gm_n91, in_2, gm_n59, gm_n90, in_4, in_3);
	nor (gm_n92, gm_n88, in_12, in_8, gm_n91, gm_n89);
	nand (gm_n93, gm_n85, gm_n72, gm_n68, gm_n92, gm_n86);
	nor (gm_n94, gm_n80, gm_n78, gm_n52, gm_n93, gm_n84);
	nand (gm_n95, gm_n94, gm_n77);
	not (gm_n96, in_30);
	nor (gm_n97, gm_n50, gm_n96, in_29);
	not (gm_n98, in_26);
	nor (gm_n99, in_27, gm_n98, in_25);
	and (gm_n100, in_23, in_22, in_21);
	not (gm_n101, gm_n100);
	not (gm_n102, in_19);
	nand (gm_n103, gm_n102, in_18, in_17);
	not (gm_n104, in_14);
	not (gm_n105, in_15);
	nand (gm_n106, gm_n105, gm_n104, in_13);
	nand (gm_n107, in_11, in_10, gm_n65);
	nor (gm_n108, in_2, in_1, in_0, in_4, gm_n60);
	not (gm_n109, in_7);
	nor (gm_n110, gm_n109, in_6, gm_n62);
	nand (gm_n111, gm_n110, gm_n108);
	or (gm_n112, gm_n106, in_12, in_8, gm_n111, gm_n107);
	nor (gm_n113, gm_n101, in_20, gm_n68, gm_n112, gm_n103);
	nand (gm_n114, gm_n97, gm_n78, in_24, gm_n113, gm_n99);
	not (gm_n115, gm_n51);
	not (gm_n116, in_17);
	nand (gm_n117, in_18, gm_n116, gm_n68);
	nor (gm_n118, gm_n104, in_13, in_12);
	nand (gm_n119, in_10, in_9, gm_n64);
	not (gm_n120, gm_n119);
	not (gm_n121, in_6);
	nor (gm_n122, in_7, gm_n121, in_5);
	not (gm_n123, in_4);
	nor (gm_n124, in_2, gm_n59, gm_n90, gm_n123, gm_n60);
	nand (gm_n125, gm_n120, gm_n118, in_11, gm_n124, gm_n122);
	nor (gm_n126, in_22, gm_n81, in_20);
	not (gm_n127, gm_n126);
	nor (gm_n128, gm_n117, in_19, gm_n105, gm_n127, gm_n125);
	nor (gm_n129, in_26, gm_n53, gm_n52);
	nand (gm_n130, gm_n115, in_27, in_23, gm_n129, gm_n128);
	nor (gm_n131, gm_n130, gm_n50);
	or (gm_n132, in_31, in_30, in_29);
	not (gm_n133, in_27);
	nor (gm_n134, gm_n133, in_26, in_25);
	not (gm_n135, gm_n134);
	not (gm_n136, in_18);
	nor (gm_n137, gm_n102, gm_n136, in_17);
	nor (gm_n138, in_15, in_14, in_13);
	not (gm_n139, gm_n138);
	and (gm_n140, in_7, in_6, in_5);
	and (gm_n141, in_2, in_1, in_0);
	nand (gm_n142, gm_n140, gm_n123, gm_n60, gm_n141);
	nor (gm_n143, gm_n88, in_12, in_8, gm_n142, gm_n139);
	nand (gm_n144, gm_n100, in_20, in_16, gm_n143, gm_n137);
	nor (gm_n145, gm_n132, in_28, in_24, gm_n144, gm_n135);
	nor (gm_n146, gm_n105, gm_n104, in_13);
	and (gm_n147, in_11, in_10, in_9);
	nor (gm_n148, in_7, in_6, gm_n62, gm_n91, in_8);
	and (gm_n149, gm_n146, in_16, in_12, gm_n148, gm_n147);
	nand (gm_n150, gm_n149, in_17);
	nand (gm_n151, in_20, in_19, gm_n136);
	nand (gm_n152, in_24, in_23, gm_n82);
	nor (gm_n153, gm_n150, gm_n53, gm_n81, gm_n152, gm_n151);
	nor (gm_n154, in_28, in_27, gm_n98);
	nand (gm_n155, gm_n50, gm_n96, gm_n76, gm_n154, gm_n153);
	nand (gm_n156, in_19, gm_n136, gm_n116);
	not (gm_n157, in_12);
	nand (gm_n158, in_15, gm_n104, gm_n56);
	or (gm_n159, in_11, in_10, in_9);
	nand (gm_n160, in_2, in_1, gm_n90, in_4, in_3);
	or (gm_n161, gm_n160, gm_n89, in_8);
	or (gm_n162, gm_n158, in_16, gm_n157, gm_n161, gm_n159);
	nor (gm_n163, gm_n84, in_24, gm_n72, gm_n162, gm_n156);
	nand (gm_n164, gm_n99, gm_n77, in_28, gm_n163);
	nor (gm_n165, in_22, gm_n81, gm_n72);
	nor (gm_n166, gm_n136, in_17, gm_n68);
	not (gm_n167, gm_n147);
	nand (gm_n168, in_15, gm_n104, in_13);
	nand (gm_n169, in_2, in_1, gm_n90, gm_n123, gm_n60);
	or (gm_n170, in_7, in_6, gm_n62, gm_n169, in_8);
	nor (gm_n171, gm_n168, gm_n167, in_12, gm_n170);
	nand (gm_n172, gm_n165, in_23, in_19, gm_n171, gm_n166);
	nor (gm_n173, gm_n98, gm_n53, in_24);
	not (gm_n174, gm_n173);
	nor (gm_n175, gm_n51, in_31, gm_n133, gm_n174, gm_n172);
	not (gm_n176, gm_n97);
	nor (gm_n177, in_27, gm_n98, gm_n53);
	not (gm_n178, gm_n137);
	nand (gm_n179, gm_n105, in_14, in_13);
	nor (gm_n180, gm_n58, gm_n87, in_9);
	nand (gm_n181, gm_n61, in_12, in_8, gm_n110, gm_n180);
	nor (gm_n182, gm_n178, in_20, gm_n68, gm_n181, gm_n179);
	nor (gm_n183, in_23, in_22, gm_n81);
	nand (gm_n184, gm_n177, gm_n78, gm_n52, gm_n183, gm_n182);
	nor (gm_n185, gm_n184, gm_n176);
	nor (gm_n186, in_31, in_30, gm_n76);
	not (gm_n187, gm_n85);
	nor (gm_n188, in_11, in_10, gm_n65);
	nor (gm_n189, in_15, in_14, gm_n56);
	and (gm_n190, gm_n122, gm_n61, gm_n64);
	nand (gm_n191, gm_n188, in_16, gm_n157, gm_n190, gm_n189);
	nor (gm_n192, gm_n84, in_24, gm_n72, gm_n191, gm_n187);
	nand (gm_n193, gm_n186, gm_n79, gm_n78, gm_n192);
	not (gm_n194, gm_n132);
	not (gm_n195, in_23);
	nor (gm_n196, gm_n195, gm_n82, in_21);
	not (gm_n197, gm_n196);
	nor (gm_n198, in_15, gm_n104, in_13);
	not (gm_n199, in_2);
	nor (gm_n200, gm_n199, in_1, gm_n90, gm_n123, in_3);
	and (gm_n201, gm_n140, in_12, in_8, gm_n200, gm_n147);
	nand (gm_n202, gm_n137, gm_n72, gm_n68, gm_n201, gm_n198);
	nor (gm_n203, gm_n135, in_28, gm_n52, gm_n202, gm_n197);
	nand (gm_n204, gm_n203, gm_n194);
	nor (gm_n205, in_31, gm_n96, in_29);
	not (gm_n206, gm_n205);
	and (gm_n207, in_27, in_26, in_25);
	not (gm_n208, gm_n207);
	nor (gm_n209, gm_n195, in_22, gm_n81);
	nor (gm_n210, gm_n109, gm_n121, in_5);
	nor (gm_n211, gm_n199, in_1, in_0, in_4, gm_n60);
	and (gm_n212, gm_n211, gm_n210, gm_n64);
	and (gm_n213, gm_n180, in_16, in_12, gm_n212, gm_n138);
	nand (gm_n214, gm_n85, in_24, gm_n72, gm_n213, gm_n209);
	nor (gm_n215, gm_n208, gm_n206, gm_n78, gm_n214);
	not (gm_n216, gm_n99);
	nor (gm_n217, gm_n50, in_30, in_29);
	not (gm_n218, gm_n217);
	not (gm_n219, gm_n156);
	nor (gm_n220, gm_n195, in_22, in_21);
	nand (gm_n221, gm_n105, in_14, gm_n56);
	nand (gm_n222, gm_n58, in_10, in_9);
	nand (gm_n223, in_7, in_6, in_5);
	nand (gm_n224, in_2, gm_n59, gm_n90, in_4, gm_n60);
	or (gm_n225, gm_n224, gm_n223, gm_n64);
	nor (gm_n226, gm_n221, gm_n68, gm_n157, gm_n225, gm_n222);
	nand (gm_n227, gm_n219, in_24, in_20, gm_n226, gm_n220);
	nor (gm_n228, gm_n218, gm_n216, gm_n78, gm_n227);
	not (gm_n229, gm_n77);
	nor (gm_n230, in_19, gm_n136, in_17);
	nor (gm_n231, gm_n105, in_14, in_13);
	nor (gm_n232, in_11, gm_n87, in_9);
	and (gm_n233, in_8, gm_n123, gm_n60, gm_n141, gm_n122);
	and (gm_n234, gm_n231, in_16, in_12, gm_n233, gm_n232);
	nand (gm_n235, gm_n209, in_24, gm_n72, gm_n234, gm_n230);
	nor (gm_n236, gm_n80, gm_n229, in_28, gm_n235);
	not (gm_n237, gm_n103);
	nor (gm_n238, in_2, gm_n59, gm_n90, in_4, in_3);
	and (gm_n239, gm_n140, gm_n157, gm_n64, gm_n238, gm_n232);
	and (gm_n240, gm_n237, gm_n72, in_16, gm_n239, gm_n138);
	nand (gm_n241, gm_n100, in_28, gm_n52, gm_n240, gm_n207);
	nor (gm_n242, gm_n241, gm_n176);
	not (gm_n243, gm_n177);
	not (gm_n244, gm_n86);
	nand (gm_n245, gm_n58, in_10, gm_n65);
	nand (gm_n246, in_7, gm_n121, in_5);
	or (gm_n247, gm_n160, gm_n246, gm_n64);
	nor (gm_n248, gm_n244, gm_n68, in_12, gm_n247, gm_n245);
	nand (gm_n249, gm_n237, in_24, gm_n72, gm_n248, gm_n196);
	nor (gm_n250, gm_n243, gm_n176, gm_n78, gm_n249);
	nor (gm_n251, gm_n236, gm_n228, gm_n215, gm_n250, gm_n242);
	nor (gm_n252, in_23, gm_n82, in_21);
	nand (gm_n253, in_11, gm_n87, in_9);
	nand (gm_n254, gm_n199, in_1, gm_n90, gm_n123, gm_n60);
	or (gm_n255, gm_n254, gm_n223, in_8);
	nor (gm_n256, gm_n244, gm_n68, gm_n157, gm_n255, gm_n253);
	nand (gm_n257, gm_n85, in_24, in_20, gm_n256, gm_n252);
	nor (gm_n258, gm_n135, gm_n229, gm_n78, gm_n257);
	nor (gm_n259, in_27, in_26, gm_n53);
	not (gm_n260, gm_n259);
	nor (gm_n261, in_23, in_22, in_21);
	nor (gm_n262, gm_n109, in_6, in_5);
	nor (gm_n263, in_2, gm_n59, in_0, gm_n123, in_3);
	nand (gm_n264, gm_n263, gm_n262, gm_n64);
	nor (gm_n265, gm_n168, gm_n68, in_12, gm_n264, gm_n245);
	nand (gm_n266, gm_n230, gm_n52, gm_n72, gm_n265, gm_n261);
	nor (gm_n267, gm_n260, gm_n229, gm_n78, gm_n266);
	not (gm_n268, gm_n186);
	nor (gm_n269, gm_n102, in_18, gm_n116);
	not (gm_n270, gm_n159);
	nand (gm_n271, in_2, in_1, gm_n90, in_4, gm_n60);
	nor (gm_n272, in_7, in_6, gm_n62, gm_n271, in_8);
	and (gm_n273, gm_n189, in_16, gm_n157, gm_n272, gm_n270);
	nand (gm_n274, gm_n100, in_24, gm_n72, gm_n273, gm_n269);
	nor (gm_n275, gm_n268, gm_n243, gm_n78, gm_n274);
	nor (gm_n276, gm_n275, gm_n267, gm_n258);
	nor (gm_n277, in_7, in_6, gm_n62, gm_n254, gm_n64);
	and (gm_n278, gm_n231, in_16, gm_n157, gm_n277, gm_n232);
	nand (gm_n279, gm_n137, in_24, in_20, gm_n278, gm_n220);
	nor (gm_n280, gm_n208, gm_n176, in_28, gm_n279);
	nor (gm_n281, in_2, in_1, in_0, gm_n123, gm_n60);
	nand (gm_n282, gm_n281, gm_n140);
	nor (gm_n283, gm_n168, in_12, gm_n64, gm_n282, gm_n253);
	nand (gm_n284, gm_n196, gm_n72, in_16, gm_n283, gm_n230);
	nor (gm_n285, gm_n135, in_28, gm_n52, gm_n284, gm_n206);
	nand (gm_n286, in_11, gm_n87, gm_n65);
	nand (gm_n287, in_8, in_4, gm_n60, gm_n141, gm_n210);
	nor (gm_n288, gm_n179, gm_n68, in_12, gm_n287, gm_n286);
	nand (gm_n289, gm_n209, gm_n52, gm_n72, gm_n288, gm_n269);
	nor (gm_n290, gm_n260, gm_n206, in_28, gm_n289);
	nor (gm_n291, gm_n290, gm_n285, gm_n280);
	nand (gm_n292, gm_n251, gm_n204, gm_n193, gm_n291, gm_n276);
	and (gm_n293, in_22, in_21, in_20);
	not (gm_n294, gm_n293);
	nand (gm_n295, gm_n199, gm_n59, in_0, gm_n123, gm_n60);
	nor (gm_n296, gm_n295, gm_n246);
	nor (gm_n297, gm_n87, in_9, in_8);
	nand (gm_n298, gm_n118, gm_n105, gm_n58, gm_n297, gm_n296);
	nor (gm_n299, in_18, gm_n116, in_16);
	not (gm_n300, gm_n299);
	nor (gm_n301, gm_n294, in_23, gm_n102, gm_n300, gm_n298);
	nor (gm_n302, in_26, in_25, in_24);
	or (gm_n303, in_30, in_29, in_28);
	not (gm_n304, gm_n303);
	nand (gm_n305, gm_n301, in_31, in_27, gm_n304, gm_n302);
	nor (gm_n306, gm_n96, in_29, in_28);
	nor (gm_n307, gm_n98, in_25, gm_n52);
	nor (gm_n308, in_7, in_6, in_5);
	nor (gm_n309, gm_n199, in_1, gm_n90, gm_n123, gm_n60);
	and (gm_n310, gm_n309, gm_n308);
	and (gm_n311, in_14, in_13, in_12);
	nand (gm_n312, gm_n120, gm_n105, gm_n58, gm_n311, gm_n310);
	nor (gm_n313, gm_n82, gm_n81, in_20);
	not (gm_n314, gm_n313);
	nor (gm_n315, gm_n117, gm_n195, gm_n102, gm_n314, gm_n312);
	nand (gm_n316, gm_n306, gm_n50, in_27, gm_n315, gm_n307);
	nor (gm_n317, in_2, in_1, in_0, in_3);
	nand (gm_n318, gm_n121, in_5, in_4, gm_n317, gm_n109);
	nand (gm_n319, gm_n87, gm_n65, in_8);
	or (gm_n320, gm_n56, in_12, in_11, gm_n319, gm_n318);
	nor (gm_n321, in_16, gm_n105, gm_n104);
	not (gm_n322, gm_n321);
	nand (gm_n323, in_20, in_19, in_18);
	or (gm_n324, gm_n320, gm_n81, gm_n116, gm_n323, gm_n322);
	and (gm_n325, in_24, in_23, in_22);
	not (gm_n326, gm_n325);
	nor (gm_n327, in_28, in_27, in_26);
	not (gm_n328, gm_n327);
	nor (gm_n329, gm_n324, in_29, in_25, gm_n328, gm_n326);
	nand (gm_n330, gm_n329, gm_n50, in_30);
	nand (gm_n331, gm_n330, gm_n316, gm_n305);
	not (gm_n332, gm_n166);
	nor (gm_n333, gm_n104, in_13, gm_n157);
	and (gm_n334, gm_n121, gm_n62, in_4, gm_n317, in_7);
	nand (gm_n335, gm_n333, in_15, in_11, gm_n334, gm_n120);
	nor (gm_n336, gm_n82, in_21, gm_n72);
	not (gm_n337, gm_n336);
	nor (gm_n338, gm_n332, gm_n195, in_19, gm_n337, gm_n335);
	nor (gm_n339, gm_n96, gm_n76, in_28);
	nand (gm_n340, gm_n307, in_31, in_27, gm_n339, gm_n338);
	nor (gm_n341, gm_n58, in_10, in_9);
	and (gm_n342, gm_n211, gm_n63, gm_n64);
	nand (gm_n343, gm_n138, gm_n68, gm_n157, gm_n342, gm_n341);
	nor (gm_n344, gm_n103, gm_n52, in_20, gm_n343, gm_n197);
	nand (gm_n345, gm_n259, gm_n77, gm_n78, gm_n344);
	nor (gm_n346, gm_n58, in_10, gm_n65);
	nand (gm_n347, gm_n109, in_6, in_5);
	nor (gm_n348, gm_n347, gm_n295, in_8);
	nand (gm_n349, gm_n146, in_16, gm_n157, gm_n348, gm_n346);
	nor (gm_n350, gm_n103, gm_n52, gm_n72, gm_n349, gm_n197);
	nand (gm_n351, gm_n134, gm_n194, gm_n78, gm_n350);
	nand (gm_n352, gm_n351, gm_n345, gm_n340);
	nor (gm_n353, gm_n292, gm_n185, gm_n175, gm_n352, gm_n331);
	nor (gm_n354, in_11, gm_n87, gm_n65);
	nand (gm_n355, gm_n199, gm_n59, gm_n90, in_4, in_3);
	nor (gm_n356, gm_n355, gm_n246, gm_n64);
	and (gm_n357, gm_n138, gm_n68, in_12, gm_n356, gm_n354);
	nand (gm_n358, gm_n230, in_24, in_20, gm_n357, gm_n261);
	nor (gm_n359, gm_n243, gm_n229, gm_n78, gm_n358);
	not (gm_n360, gm_n306);
	nor (gm_n361, in_22, in_21, in_20);
	nor (gm_n362, in_18, in_17, in_16);
	not (gm_n363, gm_n362);
	nor (gm_n364, in_2, in_1, in_0, in_4, in_3);
	nand (gm_n365, gm_n87, in_9, gm_n64, gm_n364, gm_n308);
	nand (gm_n366, gm_n104, in_13, in_12);
	nor (gm_n367, gm_n363, gm_n105, in_11, gm_n366, gm_n365);
	nand (gm_n368, gm_n55, in_23, gm_n102, gm_n367, gm_n361);
	nor (gm_n369, gm_n360, gm_n50, gm_n133, gm_n368);
	nor (gm_n370, gm_n133, gm_n98, in_25);
	not (gm_n371, gm_n370);
	nand (gm_n372, gm_n124, gm_n63, gm_n64);
	nor (gm_n373, gm_n168, in_16, gm_n157, gm_n372, gm_n222);
	nand (gm_n374, gm_n237, in_24, gm_n72, gm_n373, gm_n252);
	nor (gm_n375, gm_n371, gm_n229, in_28, gm_n374);
	nor (gm_n376, gm_n375, gm_n369, gm_n359);
	nor (gm_n377, gm_n271, gm_n246, in_8);
	and (gm_n378, gm_n198, in_16, in_12, gm_n377, gm_n346);
	nand (gm_n379, gm_n83, in_24, gm_n72, gm_n378, gm_n137);
	nor (gm_n380, gm_n218, gm_n243, gm_n78, gm_n379);
	nand (gm_n381, gm_n364, gm_n140, gm_n64);
	nor (gm_n382, gm_n244, in_16, in_12, gm_n381, gm_n88);
	nand (gm_n383, gm_n137, in_24, in_20, gm_n382, gm_n196);
	nor (gm_n384, gm_n260, gm_n132, gm_n78, gm_n383);
	or (gm_n385, in_7, in_6, in_5);
	or (gm_n386, gm_n385, gm_n271);
	nor (gm_n387, gm_n179, gm_n157, in_8, gm_n386, gm_n253);
	nand (gm_n388, gm_n85, gm_n72, in_16, gm_n387, gm_n100);
	nor (gm_n389, gm_n206, gm_n78, gm_n52, gm_n388, gm_n208);
	nor (gm_n390, gm_n389, gm_n384, gm_n380);
	nand (gm_n391, gm_n353, gm_n164, gm_n155, gm_n390, gm_n376);
	nor (gm_n392, gm_n96, in_29, gm_n78);
	nor (gm_n393, in_26, in_25, gm_n52);
	and (gm_n394, in_18, in_17, in_16);
	not (gm_n395, gm_n394);
	nand (gm_n396, in_10, gm_n65, in_8);
	nor (gm_n397, in_2, in_1, gm_n90, in_4, in_3);
	nand (gm_n398, gm_n397, gm_n210);
	nand (gm_n399, gm_n104, gm_n56, in_12);
	or (gm_n400, gm_n396, gm_n105, gm_n58, gm_n399, gm_n398);
	nor (gm_n401, gm_n294, gm_n195, gm_n102, gm_n400, gm_n395);
	nand (gm_n402, gm_n392, in_31, gm_n133, gm_n401, gm_n393);
	nor (gm_n403, in_2, gm_n59, gm_n90, gm_n123, in_3);
	and (gm_n404, gm_n270, gm_n157, in_8, gm_n403, gm_n308);
	nor (gm_n405, in_16, gm_n105, in_14);
	nor (gm_n406, in_20, in_19, gm_n136);
	and (gm_n407, gm_n404, in_17, gm_n56, gm_n406, gm_n405);
	nor (gm_n408, in_24, in_23, in_22);
	nor (gm_n409, gm_n78, in_27, gm_n98);
	and (gm_n410, gm_n407, gm_n53, in_21, gm_n409, gm_n408);
	nand (gm_n411, gm_n50, gm_n96, in_29, gm_n410);
	not (gm_n412, gm_n252);
	not (gm_n413, gm_n269);
	and (gm_n414, gm_n210, gm_n61, gm_n64);
	nand (gm_n415, gm_n86, in_16, in_12, gm_n414, gm_n354);
	nor (gm_n416, gm_n412, gm_n52, gm_n72, gm_n415, gm_n413);
	nand (gm_n417, gm_n370, gm_n194, gm_n78, gm_n416);
	nand (gm_n418, gm_n417, gm_n411, gm_n402);
	and (gm_n419, gm_n308, gm_n200, gm_n64);
	nand (gm_n420, gm_n86, in_16, in_12, gm_n419, gm_n270);
	nor (gm_n421, gm_n156, gm_n52, gm_n72, gm_n420, gm_n197);
	nand (gm_n422, gm_n99, gm_n77, in_28, gm_n421);
	not (gm_n423, gm_n165);
	and (gm_n424, gm_n262, gm_n200);
	nor (gm_n425, in_10, in_9, in_8);
	nand (gm_n426, in_14, in_13, gm_n157);
	not (gm_n427, gm_n426);
	nand (gm_n428, gm_n424, in_15, gm_n58, gm_n427, gm_n425);
	nor (gm_n429, gm_n423, gm_n195, gm_n102, gm_n428, gm_n363);
	nand (gm_n430, gm_n307, in_31, gm_n133, gm_n429, gm_n392);
	not (gm_n431, gm_n361);
	nand (gm_n432, gm_n87, in_9, gm_n64);
	nand (gm_n433, in_6, gm_n62, in_4, gm_n317, in_7);
	or (gm_n434, gm_n57, in_15, gm_n58, gm_n433, gm_n432);
	nor (gm_n435, gm_n431, gm_n195, gm_n102, gm_n434, gm_n395);
	nand (gm_n436, gm_n96, in_29, in_28);
	not (gm_n437, gm_n436);
	nand (gm_n438, gm_n393, in_31, in_27, gm_n437, gm_n435);
	nand (gm_n439, gm_n438, gm_n430, gm_n422);
	nor (gm_n440, gm_n391, gm_n145, gm_n131, gm_n439, gm_n418);
	nand (gm_n441, gm_n180, gm_n157, in_8, gm_n200, gm_n110);
	nor (gm_n442, gm_n187, in_20, in_16, gm_n441, gm_n221);
	nand (gm_n443, gm_n100, in_28, in_24, gm_n442, gm_n370);
	nor (gm_n444, gm_n443, gm_n206);
	nand (gm_n445, gm_n122, gm_n108, gm_n64);
	nor (gm_n446, gm_n179, in_16, gm_n157, gm_n445, gm_n222);
	nand (gm_n447, gm_n100, gm_n52, gm_n72, gm_n446, gm_n237);
	nor (gm_n448, gm_n208, gm_n268, gm_n78, gm_n447);
	nor (gm_n449, gm_n87, in_9, gm_n64);
	nor (gm_n450, in_2, gm_n59, gm_n90, in_4, gm_n60);
	nand (gm_n451, gm_n110, gm_n333, in_11, gm_n450, gm_n449);
	nor (gm_n452, gm_n136, gm_n116, in_16);
	not (gm_n453, gm_n452);
	nor (gm_n454, gm_n423, gm_n102, in_15, gm_n453, gm_n451);
	and (gm_n455, in_26, in_25, in_24);
	nand (gm_n456, gm_n306, in_27, in_23, gm_n455, gm_n454);
	nor (gm_n457, gm_n456, in_31);
	nor (gm_n458, gm_n457, gm_n448, gm_n444);
	not (gm_n459, gm_n230);
	nand (gm_n460, gm_n346, in_12, in_8, gm_n403, gm_n308);
	nor (gm_n461, gm_n158, gm_n72, in_16, gm_n460, gm_n459);
	nor (gm_n462, gm_n133, in_26, gm_n53);
	nand (gm_n463, gm_n220, in_28, in_24, gm_n462, gm_n461);
	nor (gm_n464, gm_n463, gm_n218);
	nand (gm_n465, in_2, in_1, in_0, in_4, in_3);
	nor (gm_n466, gm_n465, gm_n223, in_8);
	and (gm_n467, gm_n138, gm_n68, in_12, gm_n466, gm_n270);
	nand (gm_n468, gm_n237, gm_n52, in_20, gm_n467, gm_n261);
	nor (gm_n469, gm_n371, gm_n218, gm_n78, gm_n468);
	or (gm_n470, gm_n385, gm_n254, in_8);
	nor (gm_n471, gm_n139, gm_n68, gm_n157, gm_n470, gm_n167);
	nor (gm_n472, in_19, in_18, gm_n116);
	nand (gm_n473, gm_n100, gm_n52, gm_n72, gm_n472, gm_n471);
	nor (gm_n474, in_31, gm_n96, gm_n76);
	not (gm_n475, gm_n474);
	nor (gm_n476, gm_n473, gm_n135, in_28, gm_n475);
	nor (gm_n477, gm_n476, gm_n469, gm_n464);
	nand (gm_n478, gm_n440, gm_n114, gm_n95, gm_n477, gm_n458);
	nand (gm_n479, gm_n62, gm_n123, gm_n60, gm_n141, gm_n121);
	nor (gm_n480, in_9, gm_n64, in_7, gm_n479, gm_n87);
	and (gm_n481, in_13, in_12, in_11);
	nor (gm_n482, gm_n116, gm_n68, in_15);
	nand (gm_n483, gm_n480, gm_n136, in_14, gm_n482, gm_n481);
	nor (gm_n484, in_21, in_20, in_19);
	not (gm_n485, gm_n484);
	nand (gm_n486, gm_n53, in_24, gm_n195);
	nor (gm_n487, gm_n483, in_26, in_22, gm_n486, gm_n485);
	nor (gm_n488, gm_n76, in_28, in_27);
	nand (gm_n489, gm_n487, in_31, gm_n96, gm_n488);
	nand (gm_n490, gm_n231, gm_n68, gm_n157, gm_n419, gm_n341);
	nor (gm_n491, gm_n197, gm_n52, gm_n72, gm_n490, gm_n413);
	and (gm_n492, in_31, in_30, in_29);
	nand (gm_n493, gm_n491, gm_n207, gm_n78, gm_n492);
	or (gm_n494, gm_n158, in_16, in_12, gm_n287, gm_n253);
	nor (gm_n495, gm_n197, gm_n52, in_20, gm_n494, gm_n413);
	nand (gm_n496, gm_n207, gm_n97, in_28, gm_n495);
	nand (gm_n497, gm_n496, gm_n493, gm_n489);
	nor (gm_n498, in_2, in_1, gm_n90, gm_n123, in_3);
	nand (gm_n499, gm_n498, gm_n140);
	nor (gm_n500, gm_n106, gm_n157, in_8, gm_n499, gm_n253);
	nand (gm_n501, gm_n85, in_20, in_16, gm_n500, gm_n220);
	nor (gm_n502, gm_n206, in_28, in_24, gm_n501, gm_n371);
	nor (out_0, gm_n497, gm_n478, gm_n75, gm_n502);
	nand (gm_n504, in_15, in_14, gm_n56);
	nor (gm_n505, gm_n504, in_16, in_12, gm_n445, gm_n159);
	nand (gm_n506, gm_n83, in_24, gm_n72, gm_n505, gm_n219);
	nor (gm_n507, gm_n218, gm_n208, gm_n78, gm_n506);
	nor (gm_n508, in_30, gm_n76, in_28);
	nor (gm_n509, gm_n82, in_21, in_20);
	not (gm_n510, gm_n509);
	nor (gm_n511, in_7, gm_n121, gm_n62);
	and (gm_n512, gm_n511, gm_n211, gm_n64);
	nand (gm_n513, gm_n299, gm_n341, in_15, gm_n512, gm_n427);
	nor (gm_n514, gm_n54, gm_n195, in_19, gm_n513, gm_n510);
	nand (gm_n515, gm_n508, in_31, in_27, gm_n514);
	not (gm_n516, gm_n220);
	and (gm_n517, in_19, in_18, in_17);
	nor (gm_n518, gm_n89, in_12, in_8, gm_n286, gm_n224);
	nand (gm_n519, gm_n138, in_20, in_16, gm_n518, gm_n517);
	nor (gm_n520, gm_n208, gm_n78, in_24, gm_n519, gm_n516);
	nand (gm_n521, gm_n520, gm_n77);
	nand (gm_n522, gm_n200, gm_n63, gm_n64);
	nor (gm_n523, gm_n158, gm_n68, in_12, gm_n522, gm_n286);
	nand (gm_n524, gm_n137, in_24, gm_n72, gm_n523, gm_n196);
	nor (gm_n525, gm_n208, gm_n229, gm_n78, gm_n524);
	nor (gm_n526, gm_n72, in_19, gm_n136);
	not (gm_n527, gm_n526);
	and (gm_n528, in_16, in_15, in_14);
	not (gm_n529, gm_n528);
	nand (gm_n530, in_5, gm_n123, gm_n60, gm_n141, gm_n121);
	nand (gm_n531, gm_n157, in_11, in_10);
	or (gm_n532, in_9, gm_n64, gm_n109, gm_n531, gm_n530);
	nor (gm_n533, gm_n527, gm_n116, in_13, gm_n532, gm_n529);
	nor (gm_n534, gm_n52, in_23, gm_n82);
	nand (gm_n535, gm_n78, in_27, gm_n98);
	not (gm_n536, gm_n535);
	nand (gm_n537, gm_n533, gm_n53, in_21, gm_n536, gm_n534);
	nor (gm_n538, gm_n50, in_30, gm_n76, gm_n537);
	and (gm_n539, in_2, in_1, in_0, in_3);
	and (gm_n540, gm_n121, in_5, gm_n123, gm_n539, gm_n109);
	nand (gm_n541, gm_n118, in_15, in_11, gm_n540, gm_n297);
	nor (gm_n542, gm_n395, in_23, in_19, gm_n541, gm_n510);
	nand (gm_n543, gm_n306, gm_n50, gm_n133, gm_n542, gm_n455);
	nand (gm_n544, in_2, gm_n59, in_0, gm_n123, gm_n60);
	nor (gm_n545, gm_n544, gm_n246, in_8);
	nand (gm_n546, gm_n180, gm_n68, in_12, gm_n545, gm_n198);
	nor (gm_n547, gm_n84, gm_n52, gm_n72, gm_n546, gm_n103);
	nand (gm_n548, gm_n217, gm_n134, gm_n78, gm_n547);
	or (gm_n549, gm_n385, gm_n91, in_8);
	nor (gm_n550, gm_n504, in_16, gm_n157, gm_n549, gm_n253);
	nand (gm_n551, gm_n252, in_24, gm_n72, gm_n550, gm_n517);
	nor (gm_n552, gm_n80, gm_n229, gm_n78, gm_n551);
	nand (gm_n553, gm_n110, gm_n61, gm_n64);
	nor (gm_n554, gm_n106, gm_n68, in_12, gm_n553, gm_n245);
	nand (gm_n555, gm_n252, gm_n52, gm_n72, gm_n554, gm_n269);
	nor (gm_n556, gm_n216, gm_n176, in_28, gm_n555);
	nor (gm_n557, gm_n223, gm_n91, in_8);
	nand (gm_n558, gm_n189, in_16, in_12, gm_n557, gm_n346);
	nor (gm_n559, gm_n84, in_24, gm_n72, gm_n558, gm_n187);
	nand (gm_n560, gm_n492, gm_n134, gm_n78, gm_n559);
	not (gm_n561, gm_n209);
	nand (gm_n562, gm_n109, in_6, gm_n62);
	nor (gm_n563, gm_n160, gm_n562, in_8);
	nand (gm_n564, gm_n147, in_16, gm_n157, gm_n563, gm_n198);
	nor (gm_n565, gm_n187, gm_n52, in_20, gm_n564, gm_n561);
	nand (gm_n566, gm_n492, gm_n79, in_28, gm_n565);
	nor (gm_n567, in_2, in_1, gm_n90, in_4, gm_n60);
	nand (gm_n568, gm_n567, gm_n511, in_8);
	nor (gm_n569, gm_n504, gm_n68, in_12, gm_n568, gm_n245);
	nand (gm_n570, gm_n137, in_24, in_20, gm_n569, gm_n252);
	nor (gm_n571, gm_n475, gm_n260, gm_n78, gm_n570);
	and (gm_n572, gm_n188, in_16, in_12, gm_n348, gm_n146);
	nand (gm_n573, gm_n137, gm_n52, in_20, gm_n572, gm_n252);
	nor (gm_n574, gm_n371, gm_n229, gm_n78, gm_n573);
	not (gm_n575, gm_n392);
	not (gm_n576, gm_n311);
	nand (gm_n577, gm_n308, gm_n124, in_8);
	nor (gm_n578, gm_n576, gm_n222, gm_n105, gm_n577, gm_n453);
	nand (gm_n579, gm_n129, in_23, gm_n102, gm_n578, gm_n313);
	nor (gm_n580, gm_n575, gm_n50, in_27, gm_n579);
	not (gm_n581, gm_n393);
	nor (gm_n582, gm_n136, in_17, in_16);
	nand (gm_n583, in_6, in_5, gm_n123, gm_n539, in_7);
	nor (gm_n584, gm_n396, in_15, in_11, gm_n583, gm_n399);
	nand (gm_n585, gm_n582, gm_n195, in_19, gm_n584, gm_n126);
	nor (gm_n586, gm_n360, gm_n50, gm_n133, gm_n585, gm_n581);
	nor (gm_n587, gm_n199, in_1, gm_n90, in_4, gm_n60);
	nand (gm_n588, gm_n587, gm_n308, gm_n64);
	nor (gm_n589, gm_n139, gm_n68, gm_n157, gm_n588, gm_n245);
	nand (gm_n590, gm_n85, gm_n52, in_20, gm_n589, gm_n100);
	nor (gm_n591, gm_n176, gm_n80, gm_n78, gm_n590);
	nor (gm_n592, gm_n580, gm_n574, gm_n571, gm_n591, gm_n586);
	nand (gm_n593, in_2, in_1, gm_n90, gm_n123, in_3);
	nor (gm_n594, gm_n593, gm_n562, gm_n64);
	and (gm_n595, gm_n147, gm_n68, gm_n157, gm_n594, gm_n198);
	nand (gm_n596, gm_n137, gm_n52, gm_n72, gm_n595, gm_n196);
	nor (gm_n597, gm_n218, gm_n208, gm_n78, gm_n596);
	or (gm_n598, gm_n271, gm_n223);
	nor (gm_n599, gm_n159, in_12, gm_n64, gm_n598, gm_n168);
	nand (gm_n600, gm_n219, gm_n72, gm_n68, gm_n599, gm_n183);
	nor (gm_n601, gm_n216, in_28, gm_n52, gm_n600, gm_n206);
	not (gm_n602, gm_n472);
	nand (gm_n603, gm_n210, gm_n157, in_8, gm_n309, gm_n180);
	nor (gm_n604, gm_n504, in_20, gm_n68, gm_n603, gm_n602);
	nand (gm_n605, gm_n252, in_28, in_24, gm_n604, gm_n259);
	nor (gm_n606, gm_n605, gm_n176);
	nor (gm_n607, gm_n606, gm_n601, gm_n597);
	nor (gm_n608, gm_n88, gm_n68, in_12, gm_n264, gm_n504);
	nand (gm_n609, gm_n219, gm_n52, in_20, gm_n608, gm_n261);
	nor (gm_n610, gm_n260, gm_n218, in_28, gm_n609);
	not (gm_n611, gm_n339);
	nor (gm_n612, in_18, gm_n116, gm_n68);
	nor (gm_n613, gm_n347, gm_n224, in_8);
	and (gm_n614, gm_n188, gm_n333, gm_n105, gm_n613, gm_n612);
	nand (gm_n615, gm_n293, in_23, in_19, gm_n614, gm_n307);
	nor (gm_n616, gm_n611, in_31, in_27, gm_n615);
	not (gm_n617, gm_n307);
	not (gm_n618, gm_n425);
	nor (gm_n619, in_2, in_1, gm_n90, gm_n123, gm_n60);
	nand (gm_n620, gm_n619, gm_n210);
	nor (gm_n621, in_14, in_13, in_12);
	not (gm_n622, gm_n621);
	nor (gm_n623, gm_n618, in_15, in_11, gm_n622, gm_n620);
	nand (gm_n624, gm_n69, gm_n195, gm_n102, gm_n623, gm_n165);
	nor (gm_n625, gm_n303, in_31, gm_n133, gm_n624, gm_n617);
	nor (gm_n626, gm_n625, gm_n616, gm_n610);
	nand (gm_n627, gm_n592, gm_n566, gm_n560, gm_n626, gm_n607);
	not (gm_n628, gm_n261);
	nor (gm_n629, in_15, gm_n104, gm_n56);
	nor (gm_n630, gm_n347, gm_n91, in_8);
	nand (gm_n631, gm_n629, in_16, gm_n157, gm_n630, gm_n354);
	nor (gm_n632, gm_n628, in_24, gm_n72, gm_n631, gm_n413);
	nand (gm_n633, gm_n474, gm_n370, in_28, gm_n632);
	nor (gm_n634, gm_n65, gm_n64, in_7, gm_n530, in_10);
	nor (gm_n635, gm_n56, in_12, in_11);
	nand (gm_n636, gm_n482, gm_n136, gm_n104, gm_n635, gm_n634);
	nor (gm_n637, in_21, gm_n72, gm_n102);
	not (gm_n638, gm_n637);
	nor (gm_n639, gm_n53, in_24, gm_n195);
	not (gm_n640, gm_n639);
	nor (gm_n641, gm_n636, in_26, gm_n82, gm_n640, gm_n638);
	and (gm_n642, in_29, in_28);
	and (gm_n643, gm_n642, gm_n133);
	nand (gm_n644, gm_n641, gm_n50, in_30, gm_n643);
	and (gm_n645, gm_n403, gm_n210, gm_n64);
	nand (gm_n646, gm_n86, gm_n68, gm_n157, gm_n645, gm_n188);
	nor (gm_n647, gm_n187, gm_n52, in_20, gm_n646, gm_n101);
	nand (gm_n648, gm_n207, gm_n77, in_28, gm_n647);
	nand (gm_n649, gm_n648, gm_n644, gm_n633);
	nor (gm_n650, gm_n562, gm_n157, in_8, gm_n222, gm_n169);
	and (gm_n651, gm_n526, in_17, in_13, gm_n650, gm_n528);
	nor (gm_n652, in_24, gm_n195, gm_n82);
	and (gm_n653, gm_n409, in_25, gm_n81, gm_n652, gm_n651);
	nand (gm_n654, gm_n50, in_30, gm_n76, gm_n653);
	nand (gm_n655, gm_n200, gm_n110, gm_n64);
	or (gm_n656, gm_n245, gm_n139, in_12, gm_n655);
	nor (gm_n657, gm_n117, in_23, gm_n102, gm_n656, gm_n337);
	nor (gm_n658, in_26, gm_n53, in_24);
	nand (gm_n659, gm_n508, in_31, in_27, gm_n658, gm_n657);
	nand (gm_n660, gm_n146, in_16, gm_n157, gm_n594, gm_n232);
	nor (gm_n661, gm_n628, in_24, in_20, gm_n660, gm_n413);
	nand (gm_n662, gm_n177, gm_n194, gm_n78, gm_n661);
	nand (gm_n663, gm_n662, gm_n659, gm_n654);
	nor (gm_n664, gm_n627, gm_n556, gm_n552, gm_n663, gm_n649);
	and (gm_n665, in_10, in_9, in_8);
	not (gm_n666, gm_n665);
	nand (gm_n667, gm_n567, gm_n210);
	nor (gm_n668, gm_n366, gm_n105, in_11, gm_n667, gm_n666);
	nand (gm_n669, gm_n509, gm_n195, in_19, gm_n668, gm_n612);
	nor (gm_n670, gm_n51, gm_n50, in_27, gm_n669, gm_n581);
	not (gm_n671, gm_n455);
	nand (gm_n672, in_14, gm_n56, gm_n157);
	nand (gm_n673, in_10, gm_n65, gm_n64);
	nand (gm_n674, in_6, in_5, gm_n123, gm_n539, gm_n109);
	nor (gm_n675, gm_n672, in_15, in_11, gm_n674, gm_n673);
	nand (gm_n676, gm_n73, in_23, gm_n102, gm_n675, gm_n394);
	nor (gm_n677, in_30, in_29, gm_n78);
	not (gm_n678, gm_n677);
	nor (gm_n679, gm_n671, in_31, in_27, gm_n678, gm_n676);
	nor (gm_n680, gm_n319, in_15, gm_n58, gm_n433, gm_n366);
	nand (gm_n681, gm_n293, gm_n195, gm_n102, gm_n680, gm_n452);
	nor (gm_n682, gm_n51, gm_n50, in_27, gm_n681, gm_n617);
	nor (gm_n683, gm_n682, gm_n679, gm_n670);
	nor (gm_n684, gm_n88, in_16, gm_n157, gm_n287, gm_n221);
	nand (gm_n685, gm_n183, in_24, gm_n72, gm_n684, gm_n269);
	nor (gm_n686, gm_n208, gm_n268, in_28, gm_n685);
	not (gm_n687, gm_n492);
	nand (gm_n688, gm_n317, in_8, in_4, gm_n511);
	nor (gm_n689, gm_n167, gm_n68, in_12, gm_n688, gm_n179);
	nand (gm_n690, gm_n83, gm_n52, in_20, gm_n689, gm_n269);
	nor (gm_n691, gm_n687, gm_n371, gm_n78, gm_n690);
	nand (gm_n692, gm_n450, gm_n308, gm_n64);
	nor (gm_n693, gm_n106, in_16, gm_n157, gm_n692, gm_n167);
	nand (gm_n694, gm_n196, in_24, in_20, gm_n693, gm_n517);
	nor (gm_n695, gm_n132, gm_n216, in_28, gm_n694);
	nor (gm_n696, gm_n695, gm_n691, gm_n686);
	nand (gm_n697, gm_n664, gm_n548, gm_n543, gm_n696, gm_n683);
	or (gm_n698, gm_n168, in_16, in_12, gm_n688, gm_n222);
	nor (gm_n699, gm_n156, in_24, gm_n72, gm_n698, gm_n412);
	nand (gm_n700, gm_n259, gm_n217, in_28, gm_n699);
	or (gm_n701, gm_n254, gm_n562);
	or (gm_n702, gm_n673, gm_n105, gm_n58, gm_n701, gm_n366);
	nor (gm_n703, gm_n314, in_23, in_19, gm_n702, gm_n453);
	nand (gm_n704, gm_n173, gm_n50, gm_n133, gm_n703, gm_n339);
	nor (gm_n705, in_2, gm_n59, in_0, gm_n123, gm_n60);
	and (gm_n706, gm_n705, gm_n140, in_8);
	nand (gm_n707, gm_n86, gm_n68, in_12, gm_n706, gm_n346);
	nor (gm_n708, gm_n197, gm_n52, in_20, gm_n707, gm_n459);
	nand (gm_n709, gm_n492, gm_n259, in_28, gm_n708);
	nand (gm_n710, gm_n709, gm_n704, gm_n700);
	nor (gm_n711, in_7, in_6, gm_n62, gm_n224, in_8);
	nand (gm_n712, gm_n138, in_16, in_12, gm_n711, gm_n341);
	nor (gm_n713, gm_n561, gm_n52, in_20, gm_n712, gm_n459);
	nand (gm_n714, gm_n134, gm_n77, in_28, gm_n713);
	nor (gm_n715, in_7, in_6, gm_n62, gm_n544, in_8);
	nand (gm_n716, gm_n189, in_16, gm_n157, gm_n715, gm_n346);
	nor (gm_n717, gm_n156, gm_n52, gm_n72, gm_n716, gm_n412);
	nand (gm_n718, gm_n492, gm_n370, gm_n78, gm_n717);
	or (gm_n719, gm_n139, gm_n68, in_12, gm_n692, gm_n245);
	nor (gm_n720, gm_n156, in_24, gm_n72, gm_n719, gm_n197);
	nand (gm_n721, gm_n492, gm_n134, in_28, gm_n720);
	nand (gm_n722, gm_n721, gm_n718, gm_n714);
	nor (gm_n723, gm_n697, gm_n538, gm_n525, gm_n722, gm_n710);
	nor (gm_n724, gm_n106, in_16, gm_n157, gm_n287, gm_n107);
	nand (gm_n725, gm_n183, gm_n52, in_20, gm_n724, gm_n269);
	nor (gm_n726, gm_n475, gm_n216, gm_n78, gm_n725);
	nand (gm_n727, gm_n87, in_9, in_8);
	nand (gm_n728, gm_n200, gm_n122);
	nor (gm_n729, gm_n727, in_15, in_11, gm_n728, gm_n672);
	nand (gm_n730, gm_n582, gm_n195, in_19, gm_n729, gm_n509);
	nor (gm_n731, gm_n174, gm_n50, gm_n133, gm_n730, gm_n611);
	not (gm_n732, gm_n406);
	nand (gm_n733, in_2, gm_n59, gm_n90, gm_n123, gm_n60);
	or (gm_n734, gm_n223, in_13, gm_n58, gm_n733, gm_n666);
	nor (gm_n735, gm_n68, gm_n105, in_14);
	not (gm_n736, gm_n735);
	nor (gm_n737, gm_n732, gm_n116, gm_n157, gm_n736, gm_n734);
	nor (gm_n738, gm_n78, in_27, in_26);
	nand (gm_n739, gm_n408, in_25, in_21, gm_n738, gm_n737);
	nor (gm_n740, in_31, gm_n96, in_29, gm_n739);
	nor (gm_n741, gm_n740, gm_n731, gm_n726);
	not (gm_n742, gm_n517);
	nand (gm_n743, gm_n124, in_12, in_8, gm_n232, gm_n140);
	nor (gm_n744, gm_n158, gm_n72, gm_n68, gm_n743, gm_n742);
	nand (gm_n745, gm_n183, gm_n78, gm_n52, gm_n744, gm_n370);
	nor (gm_n746, gm_n745, gm_n132);
	nor (gm_n747, gm_n199, in_1, in_0, in_4, in_3);
	nand (gm_n748, gm_n747, gm_n262, gm_n64);
	nor (gm_n749, gm_n107, gm_n68, in_12, gm_n748, gm_n139);
	nand (gm_n750, gm_n137, gm_n52, gm_n72, gm_n749, gm_n261);
	nor (gm_n751, gm_n260, gm_n218, gm_n78, gm_n750);
	nand (gm_n752, gm_n87, in_9, gm_n64, gm_n308, gm_n211);
	nor (gm_n753, gm_n117, gm_n105, gm_n58, gm_n752, gm_n672);
	nand (gm_n754, gm_n55, in_23, gm_n102, gm_n753, gm_n126);
	nor (gm_n755, gm_n611, gm_n50, gm_n133, gm_n754);
	nor (gm_n756, gm_n755, gm_n751, gm_n746);
	nand (gm_n757, gm_n723, gm_n521, gm_n515, gm_n756, gm_n741);
	and (gm_n758, gm_n450, gm_n110, gm_n64);
	nand (gm_n759, gm_n146, gm_n68, gm_n157, gm_n758, gm_n147);
	nor (gm_n760, gm_n459, in_24, gm_n72, gm_n759, gm_n412);
	nand (gm_n761, gm_n205, gm_n134, gm_n78, gm_n760);
	nand (gm_n762, gm_n121, gm_n62, in_4, gm_n317, gm_n109);
	or (gm_n763, gm_n57, in_15, gm_n58, gm_n762, gm_n727);
	nor (gm_n764, gm_n423, in_23, in_19, gm_n763, gm_n300);
	nand (gm_n765, gm_n129, in_31, in_27, gm_n764, gm_n392);
	nor (gm_n766, gm_n105, in_14, gm_n56);
	nand (gm_n767, gm_n766, in_16, gm_n157, gm_n346, gm_n233);
	nor (gm_n768, gm_n101, gm_n52, gm_n72, gm_n767, gm_n103);
	nand (gm_n769, gm_n462, gm_n186, gm_n78, gm_n768);
	nand (gm_n770, gm_n769, gm_n765, gm_n761);
	or (gm_n771, in_7, in_6, gm_n62, gm_n91, gm_n64);
	nand (gm_n772, in_16, gm_n105, gm_n104);
	or (gm_n773, gm_n222, gm_n56, gm_n157, gm_n772, gm_n771);
	nor (gm_n774, gm_n151, gm_n81, gm_n116, gm_n773);
	nor (gm_n775, in_24, in_23, gm_n82);
	and (gm_n776, in_28, in_27, in_26);
	nand (gm_n777, gm_n774, in_29, in_25, gm_n776, gm_n775);
	nor (gm_n778, gm_n777, gm_n50, gm_n96);
	nor (out_1, gm_n770, gm_n757, gm_n507, gm_n778);
	not (gm_n780, gm_n462);
	or (gm_n781, gm_n544, gm_n246, gm_n64);
	nor (gm_n782, gm_n88, in_16, gm_n157, gm_n781, gm_n179);
	nand (gm_n783, gm_n85, gm_n52, in_20, gm_n782, gm_n183);
	nor (gm_n784, gm_n780, gm_n268, gm_n78, gm_n783);
	nor (gm_n785, in_7, in_6, gm_n62, gm_n160, gm_n64);
	nand (gm_n786, gm_n180, in_16, in_12, gm_n785, gm_n231);
	nor (gm_n787, gm_n156, in_24, in_20, gm_n786, gm_n516);
	nand (gm_n788, gm_n205, gm_n177, gm_n78, gm_n787);
	nor (gm_n789, gm_n271, gm_n562, gm_n64);
	nand (gm_n790, gm_n86, in_16, gm_n157, gm_n789, gm_n346);
	nor (gm_n791, gm_n84, gm_n52, gm_n72, gm_n790, gm_n742);
	nand (gm_n792, gm_n205, gm_n177, gm_n78, gm_n791);
	nand (gm_n793, gm_n140, in_12, gm_n64, gm_n705, gm_n147);
	nor (gm_n794, gm_n156, in_20, in_16, gm_n793, gm_n179);
	nand (gm_n795, gm_n252, in_28, gm_n52, gm_n794, gm_n259);
	nor (gm_n796, gm_n795, gm_n206);
	and (gm_n797, in_6, gm_n62, gm_n123, gm_n539, in_7);
	and (gm_n798, gm_n427, gm_n105, gm_n58, gm_n797, gm_n665);
	nand (gm_n799, gm_n313, in_23, in_19, gm_n798, gm_n362);
	nor (gm_n800, gm_n174, in_31, in_27, gm_n799, gm_n611);
	nand (gm_n801, gm_n333, in_15, in_11, gm_n334, gm_n66);
	nor (gm_n802, gm_n70, gm_n195, in_19, gm_n801, gm_n337);
	nand (gm_n803, gm_n339, in_31, gm_n133, gm_n802, gm_n658);
	not (gm_n804, gm_n183);
	nand (gm_n805, gm_n766, gm_n68, gm_n157, gm_n342, gm_n346);
	nor (gm_n806, gm_n156, gm_n52, in_20, gm_n805, gm_n804);
	nand (gm_n807, gm_n370, gm_n186, gm_n78, gm_n806);
	nand (gm_n808, gm_n498, gm_n210, gm_n64);
	nor (gm_n809, gm_n139, in_16, in_12, gm_n808, gm_n167);
	nand (gm_n810, gm_n83, gm_n52, in_20, gm_n809, gm_n237);
	nor (gm_n811, gm_n268, gm_n243, in_28, gm_n810);
	nor (gm_n812, gm_n111, gm_n157, gm_n64, gm_n222, gm_n221);
	nand (gm_n813, gm_n230, gm_n72, gm_n68, gm_n812, gm_n252);
	nor (gm_n814, gm_n216, in_28, in_24, gm_n813, gm_n268);
	nand (gm_n815, gm_n629, gm_n72, gm_n68, gm_n269, gm_n201);
	nor (gm_n816, gm_n135, gm_n78, gm_n52, gm_n815, gm_n628);
	nand (gm_n817, gm_n816, gm_n205);
	not (gm_n818, gm_n366);
	nand (gm_n819, gm_n120, in_15, in_11, gm_n818, gm_n334);
	nor (gm_n820, gm_n70, in_23, in_19, gm_n819, gm_n314);
	nand (gm_n821, gm_n173, in_31, in_27, gm_n820, gm_n339);
	or (gm_n822, gm_n88, in_12, in_8, gm_n254, gm_n246);
	nor (gm_n823, gm_n158, gm_n72, gm_n68, gm_n822, gm_n413);
	nand (gm_n824, gm_n83, in_28, gm_n52, gm_n823, gm_n259);
	nor (gm_n825, gm_n824, gm_n229);
	nand (gm_n826, gm_n262, gm_n124, gm_n64);
	nor (gm_n827, gm_n167, gm_n68, in_12, gm_n826, gm_n221);
	nand (gm_n828, gm_n183, in_24, gm_n72, gm_n827, gm_n230);
	nor (gm_n829, gm_n218, gm_n243, in_28, gm_n828);
	nor (gm_n830, gm_n727, gm_n105, gm_n58, gm_n762, gm_n576);
	nand (gm_n831, gm_n452, gm_n195, in_19, gm_n830, gm_n509);
	nor (gm_n832, gm_n54, in_31, gm_n133, gm_n831, gm_n436);
	nand (gm_n833, in_7, gm_n121, in_5, gm_n364, in_8);
	nor (gm_n834, gm_n106, in_16, in_12, gm_n833, gm_n159);
	nand (gm_n835, gm_n83, gm_n52, gm_n72, gm_n834, gm_n230);
	nor (gm_n836, gm_n80, gm_n229, in_28, gm_n835);
	or (gm_n837, gm_n562, in_12, in_8, gm_n271, gm_n253);
	nor (gm_n838, gm_n106, gm_n72, gm_n68, gm_n837, gm_n413);
	nand (gm_n839, gm_n100, gm_n78, gm_n52, gm_n838, gm_n134);
	nor (gm_n840, gm_n839, gm_n206);
	nor (gm_n841, gm_n832, gm_n829, gm_n825, gm_n840, gm_n836);
	not (gm_n842, gm_n508);
	nor (gm_n843, gm_n57, gm_n105, in_11, gm_n583, gm_n673);
	nand (gm_n844, gm_n313, in_23, in_19, gm_n843, gm_n394);
	nor (gm_n845, gm_n54, in_31, gm_n133, gm_n844, gm_n842);
	nand (gm_n846, gm_n511, gm_n61, in_8);
	nor (gm_n847, gm_n504, in_16, in_12, gm_n846, gm_n253);
	nand (gm_n848, gm_n209, gm_n52, gm_n72, gm_n847, gm_n230);
	nor (gm_n849, gm_n135, gm_n176, in_28, gm_n848);
	nor (gm_n850, in_9, gm_n64, gm_n109, gm_n479, gm_n87);
	nand (gm_n851, gm_n56, gm_n157, in_11, gm_n850, gm_n104);
	nor (gm_n852, in_17, in_16, gm_n105);
	not (gm_n853, gm_n852);
	nor (gm_n854, gm_n485, gm_n82, in_18, gm_n853, gm_n851);
	nand (gm_n855, gm_n639, gm_n96, in_26, gm_n854, gm_n643);
	nor (gm_n856, gm_n855, in_31);
	nor (gm_n857, gm_n856, gm_n849, gm_n845);
	or (gm_n858, gm_n562, gm_n157, gm_n64, gm_n286, gm_n160);
	nor (gm_n859, gm_n179, gm_n72, in_16, gm_n858, gm_n413);
	nand (gm_n860, gm_n99, in_28, in_24, gm_n859, gm_n183);
	nor (gm_n861, gm_n860, gm_n229);
	nand (gm_n862, gm_n122, gm_n120, gm_n58, gm_n427, gm_n309);
	nor (gm_n863, gm_n70, in_19, gm_n105, gm_n862, gm_n294);
	nand (gm_n864, gm_n115, gm_n133, gm_n195, gm_n863, gm_n173);
	nor (gm_n865, gm_n864, in_31);
	or (gm_n866, in_7, in_6, gm_n62, gm_n224, gm_n64);
	nor (gm_n867, gm_n88, gm_n68, in_12, gm_n866, gm_n504);
	nand (gm_n868, gm_n85, in_24, in_20, gm_n867, gm_n100);
	nor (gm_n869, gm_n135, gm_n176, in_28, gm_n868);
	nor (gm_n870, gm_n869, gm_n865, gm_n861);
	nand (gm_n871, gm_n841, gm_n821, gm_n817, gm_n870, gm_n857);
	and (gm_n872, gm_n238, gm_n122, gm_n64);
	nand (gm_n873, gm_n231, in_16, in_12, gm_n872, gm_n232);
	nor (gm_n874, gm_n84, gm_n52, in_20, gm_n873, gm_n156);
	nand (gm_n875, gm_n99, gm_n77, in_28, gm_n874);
	nor (gm_n876, gm_n271, gm_n246, gm_n64);
	nand (gm_n877, gm_n86, gm_n68, in_12, gm_n876, gm_n270);
	nor (gm_n878, gm_n156, gm_n52, in_20, gm_n877, gm_n561);
	nand (gm_n879, gm_n217, gm_n79, in_28, gm_n878);
	or (gm_n880, gm_n254, gm_n89);
	or (gm_n881, gm_n576, in_15, gm_n58, gm_n880, gm_n666);
	nor (gm_n882, gm_n117, gm_n195, in_19, gm_n881, gm_n294);
	nand (gm_n883, gm_n173, in_31, gm_n133, gm_n882, gm_n508);
	nand (gm_n884, gm_n883, gm_n879, gm_n875);
	nor (gm_n885, gm_n544, gm_n223, gm_n64);
	nand (gm_n886, gm_n138, in_16, in_12, gm_n885, gm_n147);
	nor (gm_n887, gm_n459, in_24, gm_n72, gm_n886, gm_n628);
	nand (gm_n888, gm_n462, gm_n186, in_28, gm_n887);
	and (gm_n889, gm_n64, gm_n123, gm_n60, gm_n511, gm_n141);
	nand (gm_n890, gm_n270, in_16, gm_n157, gm_n889, gm_n629);
	nor (gm_n891, gm_n804, gm_n52, in_20, gm_n890, gm_n742);
	nand (gm_n892, gm_n186, gm_n79, gm_n78, gm_n891);
	nor (gm_n893, gm_n544, gm_n562, gm_n64);
	nand (gm_n894, gm_n231, in_16, gm_n157, gm_n893, gm_n341);
	nor (gm_n895, gm_n197, in_24, gm_n72, gm_n894, gm_n602);
	nand (gm_n896, gm_n474, gm_n79, in_28, gm_n895);
	nand (gm_n897, gm_n896, gm_n892, gm_n888);
	nor (gm_n898, gm_n871, gm_n814, gm_n811, gm_n897, gm_n884);
	and (gm_n899, gm_n629, in_16, gm_n157, gm_n414, gm_n232);
	nand (gm_n900, gm_n83, in_24, gm_n72, gm_n899, gm_n219);
	nor (gm_n901, gm_n206, gm_n135, in_28, gm_n900);
	nand (gm_n902, gm_n309, gm_n210, gm_n64);
	nor (gm_n903, gm_n504, gm_n68, in_12, gm_n902, gm_n253);
	nand (gm_n904, gm_n220, in_24, in_20, gm_n903, gm_n517);
	nor (gm_n905, gm_n780, gm_n176, gm_n78, gm_n904);
	nand (gm_n906, gm_n567, gm_n110, in_8);
	nor (gm_n907, gm_n88, gm_n68, gm_n157, gm_n906, gm_n504);
	nand (gm_n908, gm_n219, gm_n52, gm_n72, gm_n907, gm_n209);
	nor (gm_n909, gm_n687, gm_n371, in_28, gm_n908);
	nor (gm_n910, gm_n909, gm_n905, gm_n901);
	not (gm_n911, gm_n612);
	nand (gm_n912, gm_n238, gm_n210, in_8);
	nor (gm_n913, gm_n399, gm_n222, gm_n105, gm_n912, gm_n911);
	nand (gm_n914, gm_n307, in_23, gm_n102, gm_n913, gm_n509);
	nor (gm_n915, gm_n360, in_31, in_27, gm_n914);
	nand (gm_n916, gm_n619, gm_n63, gm_n64);
	nor (gm_n917, gm_n88, in_16, in_12, gm_n916, gm_n139);
	nand (gm_n918, gm_n196, in_24, in_20, gm_n917, gm_n517);
	nor (gm_n919, gm_n475, gm_n208, in_28, gm_n918);
	nor (gm_n920, gm_n347, gm_n271, gm_n64);
	and (gm_n921, gm_n629, in_16, gm_n157, gm_n920, gm_n232);
	nand (gm_n922, gm_n209, gm_n52, gm_n72, gm_n921, gm_n269);
	nor (gm_n923, gm_n260, gm_n268, gm_n78, gm_n922);
	nor (gm_n924, gm_n923, gm_n919, gm_n915);
	nand (gm_n925, gm_n898, gm_n807, gm_n803, gm_n924, gm_n910);
	nand (gm_n926, gm_n138, in_16, in_12, gm_n354, gm_n212);
	nor (gm_n927, gm_n561, in_24, in_20, gm_n926, gm_n742);
	nand (gm_n928, gm_n217, gm_n99, in_28, gm_n927);
	nor (gm_n929, gm_n179, in_16, gm_n157, gm_n470, gm_n286);
	and (gm_n930, gm_n100, in_24, in_20, gm_n929, gm_n517);
	nand (gm_n931, gm_n205, gm_n79, gm_n78, gm_n930);
	nand (gm_n932, gm_n449, gm_n110, gm_n58, gm_n450);
	or (gm_n933, gm_n57, in_19, gm_n105, gm_n932, gm_n395);
	nor (gm_n934, gm_n54, gm_n133, in_23, gm_n933, gm_n127);
	nand (gm_n935, gm_n934, gm_n508, gm_n50);
	nand (gm_n936, gm_n935, gm_n931, gm_n928);
	not (gm_n937, gm_n432);
	nor (gm_n938, in_14, in_13, gm_n157);
	nand (gm_n939, gm_n937, gm_n105, in_11, gm_n540, gm_n938);
	nor (gm_n940, gm_n294, in_23, in_19, gm_n939, gm_n453);
	nand (gm_n941, gm_n455, in_31, gm_n133, gm_n940, gm_n677);
	nand (gm_n942, in_7, gm_n121, gm_n62);
	nor (gm_n943, gm_n107, gm_n157, gm_n64, gm_n942, gm_n254);
	nand (gm_n944, gm_n138, gm_n72, in_16, gm_n943, gm_n230);
	nor (gm_n945, gm_n216, gm_n78, gm_n52, gm_n944, gm_n197);
	nand (gm_n946, gm_n945, gm_n194);
	or (gm_n947, gm_n222, gm_n70, gm_n105, gm_n912, gm_n622);
	nor (gm_n948, gm_n174, gm_n195, gm_n102, gm_n947, gm_n510);
	nand (gm_n949, gm_n306, gm_n50, gm_n133, gm_n948);
	nand (gm_n950, gm_n949, gm_n946, gm_n941);
	nor (gm_n951, gm_n925, gm_n800, gm_n796, gm_n950, gm_n936);
	or (gm_n952, gm_n91, in_12, gm_n64, gm_n159, gm_n223);
	nor (gm_n953, gm_n158, in_20, in_16, gm_n952, gm_n459);
	nand (gm_n954, gm_n220, gm_n78, gm_n52, gm_n953, gm_n462);
	nor (gm_n955, gm_n954, gm_n475);
	and (gm_n956, gm_n122, gm_n123, gm_n60, gm_n297, gm_n141);
	and (gm_n957, gm_n582, in_15, in_11, gm_n956, gm_n118);
	nand (gm_n958, gm_n313, in_23, in_19, gm_n957, gm_n658);
	nor (gm_n959, gm_n51, gm_n50, in_27, gm_n958);
	nand (gm_n960, gm_n403, gm_n110, in_8);
	nor (gm_n961, gm_n139, gm_n68, gm_n157, gm_n960, gm_n286);
	nand (gm_n962, gm_n85, gm_n52, gm_n72, gm_n961, gm_n183);
	nor (gm_n963, gm_n475, gm_n135, in_28, gm_n962);
	nor (gm_n964, gm_n963, gm_n959, gm_n955);
	and (gm_n965, gm_n188, in_12, in_8, gm_n567, gm_n122);
	and (gm_n966, gm_n137, gm_n72, gm_n68, gm_n965, gm_n766);
	nand (gm_n967, gm_n79, gm_n78, in_24, gm_n966, gm_n83);
	nor (gm_n968, gm_n967, gm_n687);
	nor (gm_n969, gm_n347, gm_n169, gm_n64);
	and (gm_n970, gm_n629, gm_n68, gm_n157, gm_n969, gm_n354);
	nand (gm_n971, gm_n196, in_24, gm_n72, gm_n970, gm_n269);
	nor (gm_n972, gm_n132, gm_n80, gm_n78, gm_n971);
	nand (gm_n973, gm_n210, gm_n123, gm_n60, gm_n141);
	nor (gm_n974, gm_n107, gm_n157, gm_n64, gm_n973, gm_n221);
	nand (gm_n975, gm_n137, in_20, in_16, gm_n974, gm_n196);
	nor (gm_n976, gm_n371, in_28, in_24, gm_n975, gm_n687);
	nor (gm_n977, gm_n976, gm_n972, gm_n968);
	nand (gm_n978, gm_n951, gm_n792, gm_n788, gm_n977, gm_n964);
	nand (gm_n979, gm_n281, gm_n262, gm_n64);
	or (gm_n980, gm_n139, in_16, gm_n157, gm_n979, gm_n253);
	nor (gm_n981, gm_n561, in_24, gm_n72, gm_n980, gm_n459);
	nand (gm_n982, gm_n492, gm_n79, in_28, gm_n981);
	not (gm_n983, gm_n658);
	or (gm_n984, gm_n672, gm_n105, in_11, gm_n395, gm_n365);
	nor (gm_n985, gm_n337, in_23, gm_n102, gm_n984, gm_n983);
	nand (gm_n986, gm_n392, gm_n50, in_27, gm_n985);
	and (gm_n987, gm_n64, in_4, gm_n60, gm_n141, gm_n140);
	nand (gm_n988, gm_n188, in_16, in_12, gm_n987, gm_n146);
	nor (gm_n989, gm_n804, gm_n52, in_20, gm_n988, gm_n742);
	nand (gm_n990, gm_n207, gm_n186, gm_n78, gm_n989);
	nand (gm_n991, gm_n990, gm_n986, gm_n982);
	nand (gm_n992, gm_n121, in_5, gm_n123, gm_n539, in_7);
	nor (gm_n993, gm_n366, in_15, gm_n58, gm_n992, gm_n618);
	nand (gm_n994, gm_n361, in_23, in_19, gm_n993, gm_n452);
	nor (gm_n995, gm_n303, in_31, in_27, gm_n994, gm_n581);
	nor (out_2, gm_n991, gm_n978, gm_n784, gm_n995);
	nand (gm_n997, gm_n104, in_13, gm_n157);
	nor (gm_n998, gm_n119, in_15, in_11, gm_n997, gm_n880);
	nand (gm_n999, gm_n582, in_23, gm_n102, gm_n998, gm_n293);
	nor (gm_n1000, gm_n51, gm_n50, gm_n133, gm_n999, gm_n983);
	nand (gm_n1001, gm_n141, in_4, gm_n60, gm_n262);
	or (gm_n1002, gm_n319, in_15, gm_n58, gm_n1001, gm_n366);
	nor (gm_n1003, gm_n431, in_23, gm_n102, gm_n1002, gm_n911);
	nand (gm_n1004, gm_n455, gm_n50, in_27, gm_n1003, gm_n508);
	nand (gm_n1005, gm_n199, in_1, gm_n90, in_4, gm_n60);
	nor (gm_n1006, gm_n1005, gm_n223, gm_n64);
	nand (gm_n1007, gm_n766, in_16, in_12, gm_n1006, gm_n354);
	nor (gm_n1008, gm_n156, gm_n52, gm_n72, gm_n1007, gm_n412);
	nand (gm_n1009, gm_n474, gm_n370, in_28, gm_n1008);
	nand (gm_n1010, gm_n270, in_12, in_8, gm_n262, gm_n238);
	nor (gm_n1011, gm_n103, in_20, in_16, gm_n1010, gm_n168);
	nand (gm_n1012, gm_n79, in_28, in_24, gm_n1011, gm_n252);
	nor (gm_n1013, gm_n1012, gm_n132);
	nor (gm_n1014, gm_n167, in_16, gm_n157, gm_n522, gm_n168);
	nand (gm_n1015, gm_n209, gm_n52, in_20, gm_n1014, gm_n230);
	nor (gm_n1016, gm_n206, gm_n243, gm_n78, gm_n1015);
	nor (gm_n1017, gm_n347, gm_n160, in_8);
	nand (gm_n1018, gm_n188, in_16, gm_n157, gm_n1017, gm_n146);
	nor (gm_n1019, gm_n103, in_24, gm_n72, gm_n1018, gm_n412);
	nand (gm_n1020, gm_n462, gm_n186, in_28, gm_n1019);
	nor (gm_n1021, gm_n271, gm_n942, gm_n64);
	nand (gm_n1022, gm_n147, in_16, in_12, gm_n1021, gm_n766);
	nor (gm_n1023, gm_n178, gm_n52, in_20, gm_n1022, gm_n561);
	nand (gm_n1024, gm_n217, gm_n79, gm_n78, gm_n1023);
	nand (gm_n1025, gm_n308, gm_n211, in_8);
	nor (gm_n1026, gm_n168, in_16, gm_n157, gm_n1025, gm_n245);
	nand (gm_n1027, gm_n209, gm_n52, gm_n72, gm_n1026, gm_n230);
	nor (gm_n1028, gm_n475, gm_n371, in_28, gm_n1027);
	or (gm_n1029, gm_n109, gm_n121, in_5, gm_n465, gm_n64);
	nor (gm_n1030, gm_n504, gm_n68, gm_n157, gm_n1029, gm_n159);
	nand (gm_n1031, gm_n261, in_24, gm_n72, gm_n1030, gm_n472);
	nor (gm_n1032, gm_n176, gm_n80, gm_n78, gm_n1031);
	or (gm_n1033, gm_n179, gm_n157, in_11, gm_n762, gm_n673);
	nor (gm_n1034, gm_n459, in_20, in_16, gm_n1033, gm_n412);
	nand (gm_n1035, gm_n79, in_28, in_24, gm_n1034, gm_n492);
	or (gm_n1036, gm_n318, gm_n105, gm_n58, gm_n426, gm_n319);
	nor (gm_n1037, gm_n117, gm_n195, gm_n102, gm_n1036, gm_n314);
	nand (gm_n1038, gm_n302, gm_n50, in_27, gm_n1037, gm_n437);
	or (gm_n1039, gm_n169, gm_n223);
	nor (gm_n1040, gm_n88, in_12, gm_n64, gm_n1039, gm_n168);
	nand (gm_n1041, gm_n183, gm_n72, in_16, gm_n1040, gm_n269);
	nor (gm_n1042, gm_n208, gm_n78, in_24, gm_n1041, gm_n475);
	or (gm_n1043, gm_n385, gm_n169);
	nor (gm_n1044, gm_n319, in_15, gm_n58, gm_n1043, gm_n622);
	nand (gm_n1045, gm_n165, in_23, in_19, gm_n1044, gm_n362);
	nor (gm_n1046, gm_n303, gm_n50, in_27, gm_n1045, gm_n983);
	nor (gm_n1047, gm_n673, gm_n105, in_11, gm_n598, gm_n366);
	nand (gm_n1048, gm_n509, in_23, in_19, gm_n1047, gm_n612);
	nor (gm_n1049, gm_n617, gm_n50, in_27, gm_n1048, gm_n611);
	nand (gm_n1050, gm_n263, gm_n210, in_8);
	nor (gm_n1051, gm_n426, gm_n245, gm_n105, gm_n1050, gm_n453);
	nand (gm_n1052, gm_n455, gm_n195, gm_n102, gm_n1051, gm_n509);
	nor (gm_n1053, gm_n575, in_31, in_27, gm_n1052);
	nand (gm_n1054, in_28, in_27, gm_n98);
	not (gm_n1055, gm_n1054);
	nor (gm_n1056, gm_n320, gm_n81, gm_n116, gm_n736, gm_n527);
	nand (gm_n1057, gm_n325, in_29, in_25, gm_n1056, gm_n1055);
	nor (gm_n1058, gm_n1057, gm_n50, in_30);
	nor (gm_n1059, gm_n1049, gm_n1046, gm_n1042, gm_n1058, gm_n1053);
	nor (gm_n1060, gm_n942, gm_n91, gm_n64);
	and (gm_n1061, gm_n629, gm_n68, in_12, gm_n1060, gm_n341);
	nand (gm_n1062, gm_n85, gm_n52, gm_n72, gm_n1061, gm_n261);
	nor (gm_n1063, gm_n687, gm_n780, gm_n78, gm_n1062);
	or (gm_n1064, in_7, in_6, gm_n62, gm_n465, in_8);
	nor (gm_n1065, gm_n244, gm_n68, gm_n157, gm_n1064, gm_n159);
	nand (gm_n1066, gm_n83, in_24, in_20, gm_n1065, gm_n517);
	nor (gm_n1067, gm_n268, gm_n216, in_28, gm_n1066);
	or (gm_n1068, gm_n91, gm_n89, gm_n64);
	nor (gm_n1069, gm_n158, gm_n68, in_12, gm_n1068, gm_n253);
	nand (gm_n1070, gm_n85, in_24, in_20, gm_n1069, gm_n252);
	nor (gm_n1071, gm_n206, gm_n80, gm_n78, gm_n1070);
	nor (gm_n1072, gm_n1071, gm_n1067, gm_n1063);
	nand (gm_n1073, gm_n364, gm_n308, in_8);
	nor (gm_n1074, gm_n159, gm_n68, in_12, gm_n1073, gm_n221);
	nand (gm_n1075, gm_n261, gm_n52, in_20, gm_n1074, gm_n269);
	nor (gm_n1076, gm_n371, gm_n229, in_28, gm_n1075);
	nand (gm_n1077, gm_n270, in_12, gm_n64, gm_n498, gm_n511);
	nor (gm_n1078, gm_n103, gm_n72, gm_n68, gm_n1077, gm_n106);
	nand (gm_n1079, gm_n100, in_28, in_24, gm_n1078, gm_n462);
	nor (gm_n1080, gm_n1079, gm_n132);
	nor (gm_n1081, gm_n57, gm_n105, in_11, gm_n620, gm_n727);
	nand (gm_n1082, gm_n293, gm_n195, in_19, gm_n1081, gm_n362);
	nor (gm_n1083, gm_n360, in_31, gm_n133, gm_n1082, gm_n983);
	nor (gm_n1084, gm_n1083, gm_n1080, gm_n1076);
	nand (gm_n1085, gm_n1059, gm_n1038, gm_n1035, gm_n1084, gm_n1072);
	nand (gm_n1086, gm_n121, in_5, in_4, gm_n317, in_7);
	or (gm_n1087, gm_n57, in_15, gm_n58, gm_n1086, gm_n432);
	nor (gm_n1088, gm_n332, in_23, in_19, gm_n1087, gm_n294);
	nand (gm_n1089, gm_n392, in_31, in_27, gm_n1088, gm_n455);
	nor (gm_n1090, gm_n89, in_12, gm_n64, gm_n224, gm_n222);
	nand (gm_n1091, gm_n237, gm_n72, in_16, gm_n1090, gm_n189);
	nor (gm_n1092, gm_n101, in_28, in_24, gm_n1091, gm_n135);
	nand (gm_n1093, gm_n1092, gm_n474);
	and (gm_n1094, gm_n122, in_12, gm_n64, gm_n200, gm_n270);
	nand (gm_n1095, gm_n86, gm_n72, in_16, gm_n1094, gm_n219);
	nor (gm_n1096, gm_n101, gm_n78, gm_n52, gm_n1095, gm_n780);
	nand (gm_n1097, gm_n1096, gm_n97);
	nand (gm_n1098, gm_n1097, gm_n1093, gm_n1089);
	nand (gm_n1099, gm_n147, gm_n68, gm_n157, gm_n277, gm_n766);
	nor (gm_n1100, gm_n561, gm_n52, gm_n72, gm_n1099, gm_n742);
	nand (gm_n1101, gm_n492, gm_n207, in_28, gm_n1100);
	and (gm_n1102, gm_n450, gm_n122);
	nand (gm_n1103, gm_n297, gm_n105, gm_n58, gm_n1102, gm_n938);
	nor (gm_n1104, gm_n294, in_23, in_19, gm_n1103, gm_n363);
	nand (gm_n1105, gm_n115, gm_n50, gm_n133, gm_n1104, gm_n455);
	and (gm_n1106, in_8, gm_n123, gm_n60, gm_n511, gm_n141);
	nand (gm_n1107, gm_n138, gm_n68, in_12, gm_n1106, gm_n232);
	nor (gm_n1108, gm_n84, gm_n52, in_20, gm_n1107, gm_n742);
	nand (gm_n1109, gm_n474, gm_n79, gm_n78, gm_n1108);
	nand (gm_n1110, gm_n1109, gm_n1105, gm_n1101);
	nor (gm_n1111, gm_n1085, gm_n1032, gm_n1028, gm_n1110, gm_n1098);
	and (gm_n1112, gm_n346, gm_n629, gm_n157, gm_n419);
	nand (gm_n1113, gm_n73, in_23, gm_n102, gm_n1112, gm_n452);
	nor (gm_n1114, gm_n611, gm_n50, gm_n133, gm_n1113, gm_n983);
	nor (gm_n1115, gm_n727, in_15, in_11, gm_n499, gm_n672);
	nand (gm_n1116, gm_n69, in_23, in_19, gm_n1115, gm_n165);
	nor (gm_n1117, gm_n51, gm_n50, in_27, gm_n1116, gm_n671);
	not (gm_n1118, gm_n129);
	and (gm_n1119, gm_n310, in_15, in_11, gm_n665, gm_n818);
	nand (gm_n1120, gm_n166, in_23, in_19, gm_n1119, gm_n361);
	nor (gm_n1121, gm_n1118, gm_n50, gm_n133, gm_n1120, gm_n842);
	nor (gm_n1122, gm_n1121, gm_n1117, gm_n1114);
	nand (gm_n1123, gm_n511, gm_n309, gm_n64);
	nor (gm_n1124, gm_n179, in_16, gm_n157, gm_n1123, gm_n253);
	nand (gm_n1125, gm_n209, gm_n52, in_20, gm_n1124, gm_n517);
	nor (gm_n1126, gm_n206, gm_n135, gm_n78, gm_n1125);
	nand (gm_n1127, gm_n498, gm_n308);
	nor (gm_n1128, gm_n119, gm_n105, gm_n58, gm_n1127, gm_n426);
	nand (gm_n1129, gm_n126, gm_n195, in_19, gm_n1128, gm_n362);
	nor (gm_n1130, gm_n575, in_31, in_27, gm_n1129, gm_n581);
	nor (gm_n1131, in_20, gm_n102, gm_n136);
	nand (gm_n1132, gm_n122, gm_n65, gm_n64, gm_n403);
	nand (gm_n1133, in_12, gm_n58, gm_n87);
	nor (gm_n1134, gm_n529, gm_n116, gm_n56, gm_n1133, gm_n1132);
	nand (gm_n1135, gm_n534, gm_n53, gm_n81, gm_n1134, gm_n1131);
	nor (gm_n1136, in_31, gm_n96, in_29, gm_n1135, gm_n1054);
	nor (gm_n1137, gm_n1136, gm_n1130, gm_n1126);
	nand (gm_n1138, gm_n1111, gm_n1024, gm_n1020, gm_n1137, gm_n1122);
	nor (gm_n1139, gm_n733, gm_n246);
	nand (gm_n1140, gm_n120, in_15, in_11, gm_n1139, gm_n938);
	nor (gm_n1141, gm_n431, in_23, in_19, gm_n1140, gm_n395);
	nand (gm_n1142, gm_n306, gm_n50, in_27, gm_n1141, gm_n658);
	nand (gm_n1143, gm_n110, in_12, gm_n64, gm_n567, gm_n341);
	nor (gm_n1144, gm_n1143, gm_n158);
	and (gm_n1145, gm_n293, gm_n195, gm_n102, gm_n1144, gm_n299);
	nand (gm_n1146, gm_n55, in_31, gm_n133, gm_n1145, gm_n437);
	and (gm_n1147, gm_n511, gm_n211, in_8);
	nand (gm_n1148, gm_n86, gm_n68, gm_n157, gm_n1147, gm_n180);
	nor (gm_n1149, gm_n561, gm_n52, gm_n72, gm_n1148, gm_n459);
	nand (gm_n1150, gm_n134, gm_n77, in_28, gm_n1149);
	nand (gm_n1151, gm_n1150, gm_n1146, gm_n1142);
	nand (gm_n1152, gm_n198, in_16, gm_n157, gm_n920, gm_n354);
	nor (gm_n1153, gm_n187, in_24, in_20, gm_n1152, gm_n101);
	nand (gm_n1154, gm_n259, gm_n97, gm_n78, gm_n1153);
	nor (gm_n1155, gm_n271, gm_n942, in_8);
	nand (gm_n1156, gm_n629, gm_n68, gm_n157, gm_n1155, gm_n232);
	nor (gm_n1157, gm_n178, gm_n52, in_20, gm_n1156, gm_n197);
	nand (gm_n1158, gm_n207, gm_n194, in_28, gm_n1157);
	and (gm_n1159, gm_n122, in_12, gm_n64, gm_n567, gm_n232);
	nand (gm_n1160, gm_n237, in_20, in_16, gm_n1159, gm_n766);
	nor (gm_n1161, gm_n628, gm_n78, in_24, gm_n1160, gm_n371);
	nand (gm_n1162, gm_n1161, gm_n97);
	nand (gm_n1163, gm_n1162, gm_n1158, gm_n1154);
	nor (gm_n1164, gm_n1138, gm_n1016, gm_n1013, gm_n1163, gm_n1151);
	nand (gm_n1165, gm_n354, gm_n157, gm_n64, gm_n403, gm_n308);
	nor (gm_n1166, gm_n244, gm_n72, in_16, gm_n1165, gm_n602);
	nand (gm_n1167, gm_n207, in_28, gm_n52, gm_n1166, gm_n220);
	nor (gm_n1168, gm_n1167, gm_n475);
	nand (gm_n1169, gm_n210, gm_n157, gm_n64, gm_n450, gm_n354);
	nor (gm_n1170, gm_n504, in_20, in_16, gm_n1169, gm_n459);
	nand (gm_n1171, gm_n252, in_28, gm_n52, gm_n1170, gm_n259);
	nor (gm_n1172, gm_n1171, gm_n268);
	nor (gm_n1173, gm_n109, in_6, in_5, gm_n465, in_8);
	and (gm_n1174, gm_n198, gm_n68, gm_n157, gm_n1173, gm_n346);
	nand (gm_n1175, gm_n196, in_24, in_20, gm_n1174, gm_n517);
	nor (gm_n1176, gm_n243, gm_n229, in_28, gm_n1175);
	nor (gm_n1177, gm_n1176, gm_n1172, gm_n1168);
	nor (gm_n1178, gm_n385, gm_n224, gm_n64);
	and (gm_n1179, gm_n189, gm_n68, in_12, gm_n1178, gm_n147);
	nand (gm_n1180, gm_n85, gm_n52, gm_n72, gm_n1179, gm_n196);
	nor (gm_n1181, gm_n268, gm_n216, gm_n78, gm_n1180);
	nor (gm_n1182, gm_n222, gm_n56, gm_n157, gm_n771);
	nor (gm_n1183, gm_n68, in_15, gm_n104);
	and (gm_n1184, gm_n1182, gm_n81, gm_n116, gm_n1183, gm_n1131);
	nor (gm_n1185, in_24, gm_n195, in_22);
	nand (gm_n1186, gm_n738, in_29, gm_n53, gm_n1185, gm_n1184);
	nor (gm_n1187, gm_n1186, gm_n50, gm_n96);
	nor (gm_n1188, gm_n179, in_16, gm_n157, gm_n846, gm_n286);
	nand (gm_n1189, gm_n137, in_24, in_20, gm_n1188, gm_n252);
	nor (gm_n1190, gm_n780, gm_n206, in_28, gm_n1189);
	nor (gm_n1191, gm_n1190, gm_n1187, gm_n1181);
	nand (gm_n1192, gm_n1164, gm_n1009, gm_n1004, gm_n1191, gm_n1177);
	or (gm_n1193, gm_n159, in_16, gm_n157, gm_n264, gm_n168);
	nor (gm_n1194, gm_n178, gm_n52, in_20, gm_n1193, gm_n197);
	nand (gm_n1195, gm_n462, gm_n186, in_28, gm_n1194);
	and (gm_n1196, gm_n188, in_12, gm_n64, gm_n567, gm_n511);
	nand (gm_n1197, gm_n137, gm_n72, in_16, gm_n1196, gm_n146);
	nor (gm_n1198, gm_n80, in_28, in_24, gm_n1197, gm_n197);
	nand (gm_n1199, gm_n1198, gm_n194);
	nand (gm_n1200, gm_n199, gm_n59, in_0, in_4, in_3);
	nor (gm_n1201, gm_n1200, gm_n223);
	nand (gm_n1202, gm_n297, gm_n105, in_11, gm_n1201, gm_n427);
	nor (gm_n1203, gm_n70, gm_n195, in_19, gm_n1202, gm_n510);
	nand (gm_n1204, gm_n55, gm_n50, in_27, gm_n1203, gm_n508);
	nand (gm_n1205, gm_n1204, gm_n1199, gm_n1195);
	or (gm_n1206, gm_n366, gm_n942, in_11, gm_n1200, gm_n618);
	nor (gm_n1207, gm_n332, in_19, gm_n105, gm_n1206, gm_n314);
	nand (gm_n1208, gm_n302, gm_n133, gm_n195, gm_n1207, gm_n339);
	nor (gm_n1209, gm_n1208, in_31);
	nor (out_3, gm_n1205, gm_n1192, gm_n1000, gm_n1209);
	and (gm_n1211, gm_n198, in_20, gm_n68, gm_n1159, gm_n472);
	nand (gm_n1212, gm_n100, gm_n78, gm_n52, gm_n1211, gm_n462);
	nor (gm_n1213, gm_n1212, gm_n176);
	nand (gm_n1214, gm_n403, gm_n262);
	or (gm_n1215, gm_n244, in_12, gm_n64, gm_n1214, gm_n245);
	nor (gm_n1216, gm_n804, in_20, in_16, gm_n1215, gm_n742);
	nand (gm_n1217, gm_n177, in_28, in_24, gm_n1216, gm_n217);
	and (gm_n1218, gm_n270, in_12, in_8, gm_n511, gm_n238);
	nand (gm_n1219, gm_n138, gm_n72, in_16, gm_n1218, gm_n269);
	nor (gm_n1220, gm_n80, gm_n78, gm_n52, gm_n1219, gm_n84);
	nand (gm_n1221, gm_n1220, gm_n186);
	nand (gm_n1222, gm_n109, in_6, in_5, gm_n364, in_8);
	nor (gm_n1223, gm_n244, in_16, gm_n157, gm_n1222, gm_n245);
	nand (gm_n1224, gm_n85, gm_n52, gm_n72, gm_n1223, gm_n209);
	nor (gm_n1225, gm_n371, gm_n206, in_28, gm_n1224);
	nor (gm_n1226, gm_n199, gm_n59, in_0, in_4, gm_n60);
	nand (gm_n1227, gm_n1226, gm_n511);
	nor (gm_n1228, gm_n319, gm_n105, in_11, gm_n1227, gm_n426);
	nand (gm_n1229, gm_n166, in_23, in_19, gm_n1228, gm_n293);
	nor (gm_n1230, gm_n360, gm_n50, in_27, gm_n1229, gm_n581);
	not (gm_n1231, gm_n302);
	nor (gm_n1232, in_14, gm_n56, in_12);
	and (gm_n1233, gm_n63, gm_n61, in_11, gm_n1232, gm_n66);
	nand (gm_n1234, gm_n73, in_19, in_15, gm_n1233, gm_n394);
	nor (gm_n1235, gm_n1231, gm_n133, in_23, gm_n1234, gm_n611);
	nand (gm_n1236, gm_n1235, gm_n50);
	and (gm_n1237, gm_n238, gm_n110, in_8);
	nand (gm_n1238, gm_n86, gm_n68, gm_n157, gm_n1237, gm_n147);
	nor (gm_n1239, gm_n84, gm_n52, gm_n72, gm_n1238, gm_n178);
	nand (gm_n1240, gm_n207, gm_n77, gm_n78, gm_n1239);
	nand (gm_n1241, gm_n511, gm_n108, gm_n64);
	nor (gm_n1242, gm_n244, gm_n68, gm_n157, gm_n1241, gm_n107);
	nand (gm_n1243, gm_n196, in_24, in_20, gm_n1242, gm_n230);
	nor (gm_n1244, gm_n687, gm_n371, gm_n78, gm_n1243);
	nor (gm_n1245, gm_n88, gm_n157, gm_n64, gm_n973, gm_n504);
	nand (gm_n1246, gm_n219, in_20, in_16, gm_n1245, gm_n220);
	nor (gm_n1247, gm_n132, in_28, in_24, gm_n1246, gm_n260);
	nand (gm_n1248, gm_n180, in_16, in_12, gm_n1017, gm_n198);
	nor (gm_n1249, gm_n561, gm_n52, in_20, gm_n1248, gm_n742);
	nand (gm_n1250, gm_n217, gm_n134, gm_n78, gm_n1249);
	nand (gm_n1251, in_5, in_4, gm_n60, gm_n141, gm_n121);
	nor (gm_n1252, gm_n1251, in_8, in_7);
	nand (gm_n1253, gm_n231, in_16, in_12, gm_n1252, gm_n270);
	nor (gm_n1254, gm_n187, in_24, gm_n72, gm_n1253, gm_n197);
	nand (gm_n1255, gm_n462, gm_n186, gm_n78, gm_n1254);
	nor (gm_n1256, gm_n366, gm_n105, in_11, gm_n728, gm_n666);
	nand (gm_n1257, gm_n361, in_23, gm_n102, gm_n1256, gm_n362);
	nor (gm_n1258, gm_n617, in_31, gm_n133, gm_n1257, gm_n611);
	nand (gm_n1259, gm_n450, gm_n262);
	nor (gm_n1260, gm_n57, gm_n105, gm_n58, gm_n1259, gm_n666);
	nand (gm_n1261, gm_n126, in_23, in_19, gm_n1260, gm_n452);
	nor (gm_n1262, gm_n575, in_31, gm_n133, gm_n1261, gm_n983);
	nor (gm_n1263, gm_n504, gm_n68, in_12, gm_n549, gm_n222);
	nand (gm_n1264, gm_n183, gm_n52, gm_n72, gm_n1263, gm_n230);
	nor (gm_n1265, gm_n371, gm_n132, in_28, gm_n1264);
	or (gm_n1266, gm_n160, gm_n223);
	nor (gm_n1267, gm_n666, gm_n105, gm_n58, gm_n1266, gm_n997);
	nand (gm_n1268, gm_n165, gm_n195, in_19, gm_n1267, gm_n452);
	nor (gm_n1269, gm_n360, in_31, in_27, gm_n1268, gm_n581);
	nand (gm_n1270, gm_n262, gm_n108, in_8);
	nor (gm_n1271, gm_n221, in_16, in_12, gm_n1270, gm_n222);
	nand (gm_n1272, gm_n100, in_24, in_20, gm_n1271, gm_n237);
	nor (gm_n1273, gm_n260, gm_n206, in_28, gm_n1272);
	nor (gm_n1274, gm_n1265, gm_n1262, gm_n1258, gm_n1273, gm_n1269);
	nand (gm_n1275, gm_n238, gm_n63);
	nor (gm_n1276, gm_n672, in_15, in_11, gm_n1275, gm_n673);
	nand (gm_n1277, gm_n166, in_23, in_19, gm_n1276, gm_n313);
	nor (gm_n1278, gm_n581, gm_n50, gm_n133, gm_n1277, gm_n842);
	nand (gm_n1279, gm_n121, gm_n62, gm_n123, gm_n539, gm_n109);
	nor (gm_n1280, gm_n119, in_15, gm_n58, gm_n1279, gm_n576);
	nand (gm_n1281, gm_n73, gm_n195, in_19, gm_n1280, gm_n362);
	nor (gm_n1282, gm_n303, gm_n50, in_27, gm_n1281, gm_n983);
	nand (gm_n1283, gm_n124, in_12, in_8, gm_n511, gm_n232);
	nor (gm_n1284, gm_n1283, gm_n168);
	nand (gm_n1285, gm_n166, in_23, in_19, gm_n1284, gm_n361);
	nor (gm_n1286, gm_n1118, gm_n50, gm_n133, gm_n1285, gm_n611);
	nor (gm_n1287, gm_n1286, gm_n1282, gm_n1278);
	and (gm_n1288, gm_n189, in_16, gm_n157, gm_n893, gm_n346);
	nand (gm_n1289, gm_n237, in_24, in_20, gm_n1288, gm_n196);
	nor (gm_n1290, gm_n132, gm_n216, gm_n78, gm_n1289);
	nor (gm_n1291, gm_n139, gm_n68, in_12, gm_n912, gm_n245);
	nand (gm_n1292, gm_n85, in_24, gm_n72, gm_n1291, gm_n183);
	nor (gm_n1293, gm_n475, gm_n243, in_28, gm_n1292);
	nand (gm_n1294, in_7, gm_n121, gm_n62, gm_n364, gm_n64);
	nor (gm_n1295, gm_n158, gm_n68, gm_n157, gm_n1294, gm_n159);
	nand (gm_n1296, gm_n196, in_24, in_20, gm_n1295, gm_n472);
	nor (gm_n1297, gm_n216, gm_n229, in_28, gm_n1296);
	nor (gm_n1298, gm_n1297, gm_n1293, gm_n1290);
	nand (gm_n1299, gm_n1274, gm_n1255, gm_n1250, gm_n1298, gm_n1287);
	nand (gm_n1300, gm_n188, in_16, gm_n157, gm_n272, gm_n146);
	nor (gm_n1301, gm_n101, in_24, in_20, gm_n1300, gm_n178);
	nand (gm_n1302, gm_n462, gm_n217, in_28, gm_n1301);
	or (gm_n1303, gm_n544, gm_n942, gm_n64);
	or (gm_n1304, gm_n139, in_16, gm_n157, gm_n1303, gm_n253);
	nor (gm_n1305, gm_n84, gm_n52, in_20, gm_n1304, gm_n413);
	nand (gm_n1306, gm_n370, gm_n186, gm_n78, gm_n1305);
	nor (gm_n1307, gm_n246, gm_n157, in_8, gm_n286, gm_n355);
	nand (gm_n1308, gm_n137, gm_n72, gm_n68, gm_n1307, gm_n146);
	nor (gm_n1309, gm_n260, in_28, in_24, gm_n1308, gm_n628);
	nand (gm_n1310, gm_n1309, gm_n474);
	nand (gm_n1311, gm_n1310, gm_n1306, gm_n1302);
	nand (gm_n1312, gm_n86, in_16, gm_n157, gm_n512, gm_n188);
	nor (gm_n1313, gm_n101, in_24, gm_n72, gm_n1312, gm_n103);
	nand (gm_n1314, gm_n194, gm_n79, in_28, gm_n1313);
	and (gm_n1315, gm_n110, gm_n157, in_8, gm_n587, gm_n270);
	nand (gm_n1316, gm_n198, gm_n72, gm_n68, gm_n1315, gm_n230);
	nor (gm_n1317, gm_n516, gm_n78, gm_n52, gm_n1316, gm_n371);
	nand (gm_n1318, gm_n1317, gm_n217);
	and (gm_n1319, gm_n450, gm_n140);
	nand (gm_n1320, gm_n427, gm_n105, gm_n58, gm_n1319, gm_n665);
	nor (gm_n1321, gm_n117, in_23, gm_n102, gm_n1320, gm_n127);
	nand (gm_n1322, gm_n307, in_31, gm_n133, gm_n1321, gm_n508);
	nand (gm_n1323, gm_n1322, gm_n1318, gm_n1314);
	nor (gm_n1324, gm_n1299, gm_n1247, gm_n1244, gm_n1323, gm_n1311);
	nand (gm_n1325, gm_n210, gm_n61, in_8);
	nor (gm_n1326, gm_n88, in_16, in_12, gm_n1325, gm_n139);
	nand (gm_n1327, gm_n261, in_24, gm_n72, gm_n1326, gm_n517);
	nor (gm_n1328, gm_n243, gm_n229, in_28, gm_n1327);
	nand (gm_n1329, gm_n1226, gm_n110);
	nor (gm_n1330, gm_n576, gm_n105, in_11, gm_n1329, gm_n618);
	nand (gm_n1331, gm_n69, in_23, in_19, gm_n1330, gm_n73);
	nor (gm_n1332, gm_n51, gm_n50, gm_n133, gm_n1331, gm_n671);
	nor (gm_n1333, gm_n158, in_16, gm_n157, gm_n771, gm_n286);
	nand (gm_n1334, gm_n85, gm_n52, in_20, gm_n1333, gm_n252);
	nor (gm_n1335, gm_n208, gm_n229, gm_n78, gm_n1334);
	nor (gm_n1336, gm_n1335, gm_n1332, gm_n1328);
	nor (gm_n1337, in_7, gm_n121, in_5, gm_n465, in_8);
	and (gm_n1338, gm_n147, in_16, in_12, gm_n1337, gm_n198);
	nand (gm_n1339, gm_n252, gm_n52, in_20, gm_n1338, gm_n269);
	nor (gm_n1340, gm_n132, gm_n80, in_28, gm_n1339);
	nor (gm_n1341, gm_n221, gm_n68, gm_n157, gm_n568, gm_n253);
	nand (gm_n1342, gm_n183, in_24, gm_n72, gm_n1341, gm_n472);
	nor (gm_n1343, gm_n687, gm_n216, in_28, gm_n1342);
	nor (gm_n1344, gm_n318, in_15, gm_n58, gm_n426, gm_n432);
	nand (gm_n1345, gm_n582, gm_n195, gm_n102, gm_n1344, gm_n361);
	nor (gm_n1346, gm_n360, in_31, gm_n133, gm_n1345, gm_n983);
	nor (gm_n1347, gm_n1346, gm_n1343, gm_n1340);
	nand (gm_n1348, gm_n1324, gm_n1240, gm_n1236, gm_n1347, gm_n1336);
	or (gm_n1349, gm_n106, in_16, gm_n157, gm_n912, gm_n107);
	nor (gm_n1350, gm_n187, gm_n52, gm_n72, gm_n1349, gm_n804);
	nand (gm_n1351, gm_n207, gm_n97, gm_n78, gm_n1350);
	nor (gm_n1352, gm_n562, gm_n157, gm_n64, gm_n224, gm_n159);
	nand (gm_n1353, gm_n85, in_20, in_16, gm_n1352, gm_n86);
	nor (gm_n1354, gm_n216, in_28, in_24, gm_n1353, gm_n804);
	nand (gm_n1355, gm_n1354, gm_n97);
	nand (gm_n1356, gm_n498, gm_n262);
	or (gm_n1357, gm_n167, gm_n157, in_8, gm_n1356, gm_n221);
	nor (gm_n1358, gm_n516, gm_n72, in_16, gm_n1357, gm_n602);
	nand (gm_n1359, gm_n370, gm_n78, gm_n52, gm_n1358, gm_n474);
	nand (gm_n1360, gm_n1359, gm_n1355, gm_n1351);
	and (gm_n1361, gm_n262, gm_n238, gm_n64);
	nand (gm_n1362, gm_n766, in_16, gm_n157, gm_n1361, gm_n346);
	nor (gm_n1363, gm_n178, in_24, gm_n72, gm_n1362, gm_n516);
	nand (gm_n1364, gm_n99, gm_n77, gm_n78, gm_n1363);
	nand (gm_n1365, gm_n705, gm_n262, gm_n64);
	or (gm_n1366, gm_n107, in_16, gm_n157, gm_n1365, gm_n158);
	nor (gm_n1367, gm_n197, gm_n52, gm_n72, gm_n1366, gm_n459);
	nand (gm_n1368, gm_n134, gm_n77, gm_n78, gm_n1367);
	nor (gm_n1369, gm_n109, in_6, gm_n62, gm_n465, gm_n64);
	nand (gm_n1370, gm_n146, gm_n68, in_12, gm_n1369, gm_n341);
	nor (gm_n1371, gm_n101, gm_n52, gm_n72, gm_n1370, gm_n742);
	nand (gm_n1372, gm_n259, gm_n97, in_28, gm_n1371);
	nand (gm_n1373, gm_n1372, gm_n1368, gm_n1364);
	nor (gm_n1374, gm_n1348, gm_n1230, gm_n1225, gm_n1373, gm_n1360);
	nor (gm_n1375, gm_n179, in_12, gm_n64, gm_n286, gm_n282);
	nand (gm_n1376, gm_n137, gm_n72, in_16, gm_n1375, gm_n196);
	nor (gm_n1377, gm_n243, in_28, gm_n52, gm_n1376, gm_n218);
	nor (gm_n1378, gm_n168, in_16, gm_n157, gm_n655, gm_n253);
	nand (gm_n1379, gm_n183, in_24, in_20, gm_n1378, gm_n472);
	nor (gm_n1380, gm_n475, gm_n371, gm_n78, gm_n1379);
	and (gm_n1381, gm_n146, in_16, in_12, gm_n1106, gm_n346);
	nand (gm_n1382, gm_n85, in_24, gm_n72, gm_n1381, gm_n209);
	nor (gm_n1383, gm_n243, gm_n229, gm_n78, gm_n1382);
	nor (gm_n1384, gm_n1383, gm_n1380, gm_n1377);
	nand (gm_n1385, gm_n262, gm_n61, in_8);
	nor (gm_n1386, gm_n88, gm_n68, gm_n157, gm_n1385, gm_n168);
	nand (gm_n1387, gm_n261, in_24, in_20, gm_n1386, gm_n269);
	nor (gm_n1388, gm_n243, gm_n229, gm_n78, gm_n1387);
	or (gm_n1389, gm_n465, gm_n385, in_8);
	nor (gm_n1390, gm_n168, in_16, gm_n157, gm_n1389, gm_n253);
	nand (gm_n1391, gm_n261, gm_n52, in_20, gm_n1390, gm_n472);
	nor (gm_n1392, gm_n206, gm_n243, gm_n78, gm_n1391);
	nor (gm_n1393, gm_n355, gm_n562, in_8);
	and (gm_n1394, gm_n86, in_16, gm_n157, gm_n1393, gm_n270);
	nand (gm_n1395, gm_n219, in_24, gm_n72, gm_n1394, gm_n220);
	nor (gm_n1396, gm_n687, gm_n371, gm_n78, gm_n1395);
	nor (gm_n1397, gm_n1396, gm_n1392, gm_n1388);
	nand (gm_n1398, gm_n1374, gm_n1221, gm_n1217, gm_n1397, gm_n1384);
	and (gm_n1399, gm_n118, gm_n63, in_11, gm_n498, gm_n449);
	nand (gm_n1400, gm_n299, gm_n102, gm_n105, gm_n1399, gm_n336);
	nor (gm_n1401, gm_n575, in_27, in_23, gm_n1400, gm_n983);
	nand (gm_n1402, gm_n1401, in_31);
	nand (gm_n1403, gm_n937, gm_n105, in_11, gm_n797, gm_n427);
	nor (gm_n1404, gm_n70, in_23, gm_n102, gm_n1403, gm_n431);
	nand (gm_n1405, gm_n307, in_31, gm_n133, gm_n1404, gm_n339);
	nand (gm_n1406, gm_n309, gm_n140);
	or (gm_n1407, gm_n366, gm_n105, gm_n58, gm_n1406, gm_n618);
	nor (gm_n1408, gm_n117, gm_n195, in_19, gm_n1407, gm_n423);
	nand (gm_n1409, gm_n306, in_31, in_27, gm_n1408, gm_n658);
	nand (gm_n1410, gm_n1409, gm_n1405, gm_n1402);
	nor (gm_n1411, gm_n1005, gm_n89, in_8);
	and (gm_n1412, gm_n138, in_16, gm_n157, gm_n1411, gm_n147);
	nand (gm_n1413, gm_n219, in_24, gm_n72, gm_n1412, gm_n220);
	nor (gm_n1414, gm_n371, gm_n176, in_28, gm_n1413);
	nor (out_4, gm_n1410, gm_n1398, gm_n1213, gm_n1414);
	nand (gm_n1416, gm_n270, gm_n157, gm_n64, gm_n403, gm_n511);
	nor (gm_n1417, gm_n103, in_20, in_16, gm_n1416, gm_n168);
	nand (gm_n1418, gm_n261, gm_n78, gm_n52, gm_n1417, gm_n370);
	nor (gm_n1419, gm_n1418, gm_n132);
	nand (gm_n1420, gm_n237, in_20, gm_n68, gm_n965, gm_n138);
	nor (gm_n1421, gm_n80, gm_n78, gm_n52, gm_n1420, gm_n197);
	nand (gm_n1422, gm_n1421, gm_n474);
	nand (gm_n1423, gm_n148, gm_n68, gm_n157, gm_n766, gm_n270);
	nor (gm_n1424, gm_n178, in_24, gm_n72, gm_n1423, gm_n197);
	nand (gm_n1425, gm_n492, gm_n99, in_28, gm_n1424);
	nand (gm_n1426, gm_n180, in_12, gm_n64, gm_n238, gm_n110);
	nor (gm_n1427, gm_n158, gm_n72, in_16, gm_n1426, gm_n742);
	nand (gm_n1428, gm_n99, in_28, in_24, gm_n1427, gm_n220);
	nor (gm_n1429, gm_n1428, gm_n132);
	nand (gm_n1430, gm_n210, in_12, in_8, gm_n705, gm_n270);
	nor (gm_n1431, gm_n244, in_20, gm_n68, gm_n1430, gm_n602);
	nand (gm_n1432, gm_n100, gm_n78, in_24, gm_n1431, gm_n207);
	nor (gm_n1433, gm_n1432, gm_n268);
	or (gm_n1434, gm_n168, in_16, in_12, gm_n1068, gm_n245);
	nor (gm_n1435, gm_n101, gm_n52, gm_n72, gm_n1434, gm_n413);
	nand (gm_n1436, gm_n177, gm_n194, gm_n78, gm_n1435);
	and (gm_n1437, gm_n587, gm_n140, in_8);
	nand (gm_n1438, gm_n138, in_16, in_12, gm_n1437, gm_n232);
	nor (gm_n1439, gm_n103, in_24, gm_n72, gm_n1438, gm_n628);
	nand (gm_n1440, gm_n492, gm_n207, gm_n78, gm_n1439);
	nor (gm_n1441, gm_n504, gm_n68, gm_n157, gm_n1389, gm_n286);
	nand (gm_n1442, gm_n209, gm_n52, gm_n72, gm_n1441, gm_n269);
	nor (gm_n1443, gm_n268, gm_n243, in_28, gm_n1442);
	nand (gm_n1444, gm_n61, in_12, gm_n64, gm_n511, gm_n188);
	nor (gm_n1445, gm_n244, in_20, gm_n68, gm_n1444, gm_n103);
	nand (gm_n1446, gm_n79, gm_n78, in_24, gm_n1445, gm_n209);
	nor (gm_n1447, gm_n1446, gm_n268);
	nand (gm_n1448, gm_n612, in_15, gm_n58, gm_n1232, gm_n956);
	nor (gm_n1449, gm_n1118, in_23, gm_n102, gm_n1448, gm_n431);
	nand (gm_n1450, gm_n304, gm_n50, gm_n133, gm_n1449);
	nand (gm_n1451, gm_n629, in_16, in_12, gm_n348, gm_n354);
	nor (gm_n1452, gm_n84, gm_n52, gm_n72, gm_n1451, gm_n103);
	nand (gm_n1453, gm_n462, gm_n186, in_28, gm_n1452);
	nor (gm_n1454, gm_n139, in_16, gm_n157, gm_n1068, gm_n286);
	nand (gm_n1455, gm_n252, gm_n52, gm_n72, gm_n1454, gm_n517);
	nor (gm_n1456, gm_n208, gm_n206, gm_n78, gm_n1455);
	or (gm_n1457, gm_n167, gm_n139, gm_n157, gm_n588);
	or (gm_n1458, gm_n294, in_23, gm_n102, gm_n1457, gm_n911);
	nor (gm_n1459, gm_n436, in_31, in_27, gm_n1458, gm_n983);
	nor (gm_n1460, gm_n282, in_15, in_11, gm_n618, gm_n576);
	nand (gm_n1461, gm_n165, gm_n195, in_19, gm_n1460, gm_n394);
	nor (gm_n1462, gm_n303, in_31, gm_n133, gm_n1461, gm_n581);
	and (gm_n1463, gm_n180, in_16, gm_n157, gm_n889, gm_n198);
	nand (gm_n1464, gm_n83, gm_n52, in_20, gm_n1463, gm_n219);
	nor (gm_n1465, gm_n206, gm_n135, gm_n78, gm_n1464);
	nor (gm_n1466, gm_n244, gm_n68, gm_n157, gm_n1073, gm_n222);
	nand (gm_n1467, gm_n183, gm_n52, gm_n72, gm_n1466, gm_n517);
	nor (gm_n1468, gm_n260, gm_n132, in_28, gm_n1467);
	nor (gm_n1469, gm_n1462, gm_n1459, gm_n1456, gm_n1468, gm_n1465);
	nand (gm_n1470, gm_n308, gm_n341, gm_n64, gm_n747);
	nor (gm_n1471, gm_n426, in_19, gm_n105, gm_n1470, gm_n911);
	nand (gm_n1472, gm_n55, gm_n133, in_23, gm_n1471, gm_n293);
	nor (gm_n1473, gm_n1472, gm_n678, in_31);
	nor (gm_n1474, gm_n117, gm_n105, gm_n58, gm_n365, gm_n672);
	nand (gm_n1475, gm_n73, in_23, in_19, gm_n1474, gm_n393);
	nor (gm_n1476, gm_n51, gm_n50, in_27, gm_n1475);
	nor (gm_n1477, gm_n106, in_16, gm_n157, gm_n1241, gm_n167);
	nand (gm_n1478, gm_n220, gm_n52, in_20, gm_n1477, gm_n472);
	nor (gm_n1479, gm_n475, gm_n208, in_28, gm_n1478);
	nor (gm_n1480, gm_n1479, gm_n1476, gm_n1473);
	nand (gm_n1481, gm_n188, in_12, gm_n64, gm_n511, gm_n124);
	nor (gm_n1482, gm_n168, in_20, in_16, gm_n1481, gm_n413);
	nand (gm_n1483, gm_n134, gm_n78, gm_n52, gm_n1482, gm_n196);
	nor (gm_n1484, gm_n1483, gm_n475);
	nand (gm_n1485, gm_n211, gm_n122);
	nor (gm_n1486, gm_n319, gm_n105, in_11, gm_n1485, gm_n366);
	nand (gm_n1487, gm_n165, gm_n195, in_19, gm_n1486, gm_n612);
	nor (gm_n1488, gm_n174, in_31, in_27, gm_n1487, gm_n436);
	nor (gm_n1489, gm_n139, in_12, gm_n64, gm_n1214, gm_n167);
	nand (gm_n1490, gm_n209, in_20, gm_n68, gm_n1489, gm_n269);
	nor (gm_n1491, gm_n216, gm_n78, in_24, gm_n1490, gm_n475);
	nor (gm_n1492, gm_n1491, gm_n1488, gm_n1484);
	nand (gm_n1493, gm_n1469, gm_n1453, gm_n1450, gm_n1492, gm_n1480);
	nand (gm_n1494, gm_n311, gm_n147, in_15, gm_n1147, gm_n452);
	nor (gm_n1495, gm_n617, gm_n195, gm_n102, gm_n1494, gm_n314);
	nand (gm_n1496, gm_n392, gm_n50, in_27, gm_n1495);
	and (gm_n1497, gm_n262, gm_n61, gm_n64);
	nand (gm_n1498, gm_n188, in_16, in_12, gm_n1497, gm_n138);
	nor (gm_n1499, gm_n187, gm_n52, gm_n72, gm_n1498, gm_n412);
	nand (gm_n1500, gm_n462, gm_n217, gm_n78, gm_n1499);
	nand (gm_n1501, gm_n766, in_16, in_12, gm_n466, gm_n232);
	nor (gm_n1502, gm_n103, gm_n52, gm_n72, gm_n1501, gm_n628);
	nand (gm_n1503, gm_n99, gm_n77, in_28, gm_n1502);
	nand (gm_n1504, gm_n1503, gm_n1500, gm_n1496);
	nand (gm_n1505, gm_n450, gm_n140, gm_n64);
	or (gm_n1506, gm_n107, gm_n68, gm_n157, gm_n1505, gm_n504);
	nor (gm_n1507, gm_n516, in_24, in_20, gm_n1506, gm_n413);
	nand (gm_n1508, gm_n259, gm_n205, gm_n78, gm_n1507);
	or (gm_n1509, gm_n142, in_12, in_8, gm_n245, gm_n504);
	nor (gm_n1510, gm_n516, in_20, gm_n68, gm_n1509, gm_n602);
	nand (gm_n1511, gm_n194, in_28, gm_n52, gm_n1510, gm_n370);
	and (gm_n1512, gm_n270, in_12, in_8, gm_n308, gm_n238);
	nand (gm_n1513, gm_n198, gm_n72, gm_n68, gm_n1512, gm_n517);
	nor (gm_n1514, gm_n101, gm_n78, in_24, gm_n1513, gm_n780);
	nand (gm_n1515, gm_n1514, gm_n97);
	nand (gm_n1516, gm_n1515, gm_n1511, gm_n1508);
	nor (gm_n1517, gm_n1493, gm_n1447, gm_n1443, gm_n1516, gm_n1504);
	nand (gm_n1518, gm_n747, gm_n511);
	nor (gm_n1519, gm_n618, gm_n105, in_11, gm_n1518, gm_n622);
	nand (gm_n1520, gm_n73, gm_n195, gm_n102, gm_n1519, gm_n452);
	nor (gm_n1521, gm_n360, in_31, gm_n133, gm_n1520, gm_n617);
	nor (gm_n1522, gm_n103, in_20, gm_n68, gm_n822, gm_n504);
	nand (gm_n1523, gm_n79, in_28, in_24, gm_n1522, gm_n209);
	nor (gm_n1524, gm_n1523, gm_n268);
	or (gm_n1525, gm_n544, gm_n89, gm_n64);
	nor (gm_n1526, gm_n167, gm_n68, gm_n157, gm_n1525, gm_n168);
	nand (gm_n1527, gm_n83, gm_n52, gm_n72, gm_n1526, gm_n237);
	nor (gm_n1528, gm_n206, gm_n135, in_28, gm_n1527);
	nor (gm_n1529, gm_n1528, gm_n1524, gm_n1521);
	nor (gm_n1530, gm_n319, gm_n105, gm_n58, gm_n1001, gm_n997);
	nand (gm_n1531, gm_n361, in_23, gm_n102, gm_n1530, gm_n394);
	nor (gm_n1532, gm_n303, gm_n50, in_27, gm_n1531, gm_n983);
	nand (gm_n1533, gm_n308, gm_n397);
	nor (gm_n1534, gm_n672, gm_n105, gm_n64, gm_n1533, gm_n286);
	nand (gm_n1535, gm_n165, gm_n195, in_19, gm_n1534, gm_n452);
	nor (gm_n1536, gm_n671, gm_n50, in_27, gm_n1535, gm_n678);
	nand (gm_n1537, gm_n587, gm_n425, gm_n110);
	nor (gm_n1538, gm_n70, in_15, gm_n58, gm_n1537, gm_n672);
	nand (gm_n1539, gm_n126, in_23, gm_n102, gm_n1538, gm_n307);
	nor (gm_n1540, gm_n436, in_31, gm_n133, gm_n1539);
	nor (gm_n1541, gm_n1540, gm_n1536, gm_n1532);
	nand (gm_n1542, gm_n1517, gm_n1440, gm_n1436, gm_n1541, gm_n1529);
	nor (gm_n1543, gm_n109, in_6, in_5, gm_n465);
	nand (gm_n1544, gm_n333, in_15, gm_n58, gm_n1543, gm_n66);
	nor (gm_n1545, gm_n431, gm_n195, in_19, gm_n1544, gm_n363);
	nand (gm_n1546, gm_n658, in_31, in_27, gm_n1545, gm_n677);
	and (gm_n1547, gm_n64, gm_n123, gm_n60, gm_n141, gm_n210);
	nand (gm_n1548, gm_n138, gm_n68, gm_n157, gm_n1547, gm_n354);
	nor (gm_n1549, gm_n187, in_24, gm_n72, gm_n1548, gm_n628);
	nand (gm_n1550, gm_n474, gm_n134, gm_n78, gm_n1549);
	and (gm_n1551, gm_n665, gm_n308, gm_n200);
	nand (gm_n1552, gm_n582, gm_n105, gm_n58, gm_n1551, gm_n118);
	nor (gm_n1553, gm_n174, gm_n195, in_19, gm_n1552, gm_n510);
	nand (gm_n1554, gm_n306, gm_n50, gm_n133, gm_n1553);
	nand (gm_n1555, gm_n1554, gm_n1550, gm_n1546);
	or (gm_n1556, gm_n672, in_15, in_11, gm_n583, gm_n673);
	nor (gm_n1557, gm_n332, gm_n195, gm_n102, gm_n1556, gm_n337);
	nand (gm_n1558, gm_n304, gm_n50, gm_n133, gm_n1557, gm_n455);
	nor (gm_n1559, gm_n562, in_12, gm_n64, gm_n1200, gm_n222);
	nand (gm_n1560, gm_n86, in_20, gm_n68, gm_n1559, gm_n472);
	nor (gm_n1561, gm_n80, in_28, gm_n52, gm_n1560, gm_n561);
	nand (gm_n1562, gm_n1561, gm_n217);
	and (gm_n1563, gm_n63, in_9, in_8, gm_n450);
	nand (gm_n1564, gm_n157, gm_n58, gm_n87, gm_n1563, gm_n56);
	nor (gm_n1565, in_20, in_19, in_18);
	not (gm_n1566, gm_n1565);
	or (gm_n1567, gm_n772, gm_n81, gm_n116, gm_n1566, gm_n1564);
	nor (gm_n1568, gm_n326, in_29, in_25, gm_n1567, gm_n535);
	nand (gm_n1569, gm_n1568, gm_n50, in_30);
	nand (gm_n1570, gm_n1569, gm_n1562, gm_n1558);
	nor (gm_n1571, gm_n1542, gm_n1433, gm_n1429, gm_n1570, gm_n1555);
	nor (gm_n1572, gm_n363, gm_n245, in_15, gm_n1050, gm_n366);
	nand (gm_n1573, gm_n126, gm_n195, gm_n102, gm_n1572, gm_n173);
	nor (gm_n1574, gm_n436, in_31, in_27, gm_n1573);
	nand (gm_n1575, gm_n140, gm_n157, gm_n64, gm_n238, gm_n147);
	nor (gm_n1576, gm_n1575, gm_n179, in_16);
	nand (gm_n1577, gm_n220, gm_n52, gm_n72, gm_n1576, gm_n472);
	nor (gm_n1578, gm_n135, gm_n132, in_28, gm_n1577);
	or (gm_n1579, gm_n271, gm_n89, gm_n64);
	nor (gm_n1580, gm_n158, gm_n68, in_12, gm_n1579, gm_n159);
	nand (gm_n1581, gm_n252, in_24, gm_n72, gm_n1580, gm_n269);
	nor (gm_n1582, gm_n218, gm_n135, gm_n78, gm_n1581);
	nor (gm_n1583, gm_n1582, gm_n1578, gm_n1574);
	nor (gm_n1584, gm_n396, in_15, in_11, gm_n1518, gm_n426);
	nand (gm_n1585, gm_n73, gm_n195, gm_n102, gm_n1584, gm_n299);
	nor (gm_n1586, gm_n51, gm_n50, in_27, gm_n1585, gm_n174);
	nor (gm_n1587, gm_n167, in_16, in_12, gm_n1029, gm_n168);
	nand (gm_n1588, gm_n183, in_24, in_20, gm_n1587, gm_n517);
	nor (gm_n1589, gm_n475, gm_n243, gm_n78, gm_n1588);
	and (gm_n1590, gm_n766, in_16, in_12, gm_n630, gm_n341);
	nand (gm_n1591, gm_n85, gm_n52, gm_n72, gm_n1590, gm_n252);
	nor (gm_n1592, gm_n780, gm_n268, gm_n78, gm_n1591);
	nor (gm_n1593, gm_n1592, gm_n1589, gm_n1586);
	nand (gm_n1594, gm_n1571, gm_n1425, gm_n1422, gm_n1593, gm_n1583);
	nor (gm_n1595, in_7, in_6, gm_n62, gm_n169, gm_n64);
	nand (gm_n1596, gm_n180, in_16, in_12, gm_n1595, gm_n629);
	nor (gm_n1597, gm_n628, in_24, in_20, gm_n1596, gm_n742);
	nand (gm_n1598, gm_n134, gm_n194, gm_n78, gm_n1597);
	nand (gm_n1599, gm_n147, gm_n118, gm_n105, gm_n1147, gm_n166);
	nor (gm_n1600, gm_n337, gm_n195, gm_n102, gm_n1599, gm_n581);
	nand (gm_n1601, gm_n392, in_31, gm_n133, gm_n1600);
	and (gm_n1602, gm_n171, gm_n195, gm_n102, gm_n452, gm_n336);
	nand (gm_n1603, gm_n173, in_31, gm_n133, gm_n1602, gm_n508);
	nand (gm_n1604, gm_n1603, gm_n1601, gm_n1598);
	nor (gm_n1605, gm_n139, gm_n68, gm_n157, gm_n1325, gm_n159);
	nand (gm_n1606, gm_n196, in_24, in_20, gm_n1605, gm_n269);
	nor (gm_n1607, gm_n371, gm_n218, in_28, gm_n1606);
	nor (out_5, gm_n1604, gm_n1594, gm_n1419, gm_n1607);
	nor (gm_n1609, gm_n65, gm_n64, in_7);
	and (gm_n1610, in_5, in_4, gm_n60, gm_n141, gm_n121);
	nand (gm_n1611, gm_n635, gm_n1609, gm_n87, gm_n1610);
	nor (gm_n1612, gm_n529, gm_n81, in_17, gm_n1611, gm_n1566);
	nand (gm_n1613, gm_n325, gm_n76, gm_n53, gm_n1612, gm_n738);
	nor (gm_n1614, gm_n1613, gm_n50, gm_n96);
	nand (gm_n1615, gm_n189, in_16, in_12, gm_n1252, gm_n147);
	nor (gm_n1616, gm_n187, in_24, in_20, gm_n1615, gm_n804);
	nand (gm_n1617, gm_n177, gm_n77, in_28, gm_n1616);
	nand (gm_n1618, in_9, gm_n64, in_7);
	nor (gm_n1619, gm_n157, gm_n58, gm_n87, gm_n1618, gm_n1251);
	nand (gm_n1620, gm_n1619, gm_n146);
	nor (gm_n1621, gm_n332, gm_n195, gm_n102, gm_n1620, gm_n337);
	nand (gm_n1622, gm_n307, in_31, gm_n133, gm_n1621, gm_n339);
	or (gm_n1623, gm_n544, gm_n562, gm_n119);
	nor (gm_n1624, gm_n332, gm_n105, in_11, gm_n1623, gm_n622);
	nand (gm_n1625, gm_n165, in_23, in_19, gm_n1624, gm_n455);
	nor (gm_n1626, gm_n575, gm_n50, in_27, gm_n1625);
	nand (gm_n1627, gm_n108, gm_n210);
	nor (gm_n1628, gm_n319, in_15, in_11, gm_n1627, gm_n622);
	nand (gm_n1629, gm_n582, gm_n195, gm_n102, gm_n1628, gm_n336);
	nor (gm_n1630, gm_n611, gm_n50, gm_n133, gm_n1629, gm_n671);
	or (gm_n1631, gm_n432, gm_n223, gm_n58, gm_n593);
	or (gm_n1632, gm_n576, in_19, gm_n105, gm_n1631, gm_n363);
	nor (gm_n1633, gm_n174, in_27, gm_n195, gm_n1632, gm_n314);
	nand (gm_n1634, gm_n1633, gm_n304, in_31);
	nor (gm_n1635, gm_n246, gm_n91, in_8, gm_n159);
	nand (gm_n1636, gm_n299, gm_n102, gm_n105, gm_n1635, gm_n427);
	nor (gm_n1637, gm_n1118, in_27, gm_n195, gm_n1636, gm_n510);
	nand (gm_n1638, gm_n1637, gm_n677, in_31);
	nand (gm_n1639, gm_n397, gm_n262, gm_n64);
	nor (gm_n1640, gm_n158, gm_n68, in_12, gm_n1639, gm_n222);
	nand (gm_n1641, gm_n100, in_24, in_20, gm_n1640, gm_n472);
	nor (gm_n1642, gm_n135, gm_n176, in_28, gm_n1641);
	nand (gm_n1643, gm_n124, gm_n63, in_8);
	nor (gm_n1644, gm_n107, in_16, gm_n157, gm_n1643, gm_n158);
	nand (gm_n1645, gm_n209, in_24, in_20, gm_n1644, gm_n517);
	nor (gm_n1646, gm_n371, gm_n218, in_28, gm_n1645);
	nor (gm_n1647, gm_n593, gm_n942, in_8);
	nand (gm_n1648, gm_n147, gm_n68, in_12, gm_n1647, gm_n629);
	nor (gm_n1649, gm_n178, gm_n52, in_20, gm_n1648, gm_n804);
	nand (gm_n1650, gm_n207, gm_n97, gm_n78, gm_n1649);
	or (gm_n1651, gm_n88, gm_n157, in_8, gm_n1043, gm_n106);
	nor (gm_n1652, gm_n804, gm_n72, gm_n68, gm_n1651, gm_n413);
	nand (gm_n1653, gm_n370, gm_n78, in_24, gm_n1652, gm_n492);
	nor (gm_n1654, gm_n318, in_15, in_11, gm_n997, gm_n618);
	nand (gm_n1655, gm_n336, in_23, in_19, gm_n1654, gm_n362);
	nor (gm_n1656, gm_n51, in_31, gm_n133, gm_n1655, gm_n983);
	nand (gm_n1657, gm_n665, gm_n498, gm_n210);
	nor (gm_n1658, gm_n117, gm_n105, gm_n58, gm_n1657, gm_n997);
	nand (gm_n1659, gm_n55, gm_n195, gm_n102, gm_n1658, gm_n509);
	nor (gm_n1660, gm_n575, in_31, in_27, gm_n1659);
	nor (gm_n1661, gm_n244, in_12, gm_n64, gm_n1039, gm_n107);
	nand (gm_n1662, gm_n237, gm_n72, gm_n68, gm_n1661, gm_n196);
	nor (gm_n1663, gm_n243, gm_n78, gm_n52, gm_n1662, gm_n268);
	nand (gm_n1664, gm_n124, gm_n210);
	nor (gm_n1665, gm_n673, in_15, gm_n58, gm_n1664, gm_n366);
	nand (gm_n1666, gm_n69, in_23, gm_n102, gm_n1665, gm_n313);
	nor (gm_n1667, gm_n54, gm_n50, gm_n133, gm_n1666, gm_n611);
	nor (gm_n1668, gm_n672, gm_n105, in_11, gm_n396, gm_n142);
	nand (gm_n1669, gm_n69, in_23, gm_n102, gm_n1668, gm_n126);
	nor (gm_n1670, gm_n54, in_31, in_27, gm_n1669, gm_n575);
	nor (gm_n1671, gm_n1663, gm_n1660, gm_n1656, gm_n1670, gm_n1667);
	nor (gm_n1672, gm_n221, in_12, in_8, gm_n1043, gm_n245);
	nand (gm_n1673, gm_n237, gm_n72, gm_n68, gm_n1672, gm_n196);
	nor (gm_n1674, gm_n80, in_28, in_24, gm_n1673, gm_n475);
	nand (gm_n1675, gm_n262, gm_n124);
	nor (gm_n1676, gm_n426, gm_n105, in_11, gm_n1675, gm_n666);
	nand (gm_n1677, gm_n582, in_23, in_19, gm_n1676, gm_n293);
	nor (gm_n1678, gm_n174, in_31, gm_n133, gm_n1677, gm_n678);
	nor (gm_n1679, gm_n504, gm_n68, in_12, gm_n1303, gm_n245);
	nand (gm_n1680, gm_n219, gm_n52, gm_n72, gm_n1679, gm_n209);
	nor (gm_n1681, gm_n243, gm_n132, gm_n78, gm_n1680);
	nor (gm_n1682, gm_n1681, gm_n1678, gm_n1674);
	and (gm_n1683, in_6, gm_n62, gm_n123, gm_n539, gm_n109);
	nand (gm_n1684, gm_n56, in_12, gm_n58, gm_n1683, gm_n297);
	nor (gm_n1685, gm_n151, in_21, gm_n116, gm_n1684, gm_n772);
	nor (gm_n1686, in_28, gm_n133, gm_n98);
	nand (gm_n1687, gm_n534, gm_n76, gm_n53, gm_n1686, gm_n1685);
	nor (gm_n1688, gm_n1687, gm_n50, in_30);
	nand (gm_n1689, gm_n122, in_12, gm_n64, gm_n498, gm_n346);
	nor (gm_n1690, gm_n158, in_20, in_16, gm_n1689, gm_n602);
	nand (gm_n1691, gm_n99, gm_n78, gm_n52, gm_n1690, gm_n220);
	nor (gm_n1692, gm_n1691, gm_n687);
	nand (gm_n1693, gm_n403, gm_n140, in_8);
	nor (gm_n1694, gm_n244, in_16, in_12, gm_n1693, gm_n253);
	nand (gm_n1695, gm_n237, gm_n52, in_20, gm_n1694, gm_n252);
	nor (gm_n1696, gm_n260, gm_n176, gm_n78, gm_n1695);
	nor (gm_n1697, gm_n1696, gm_n1692, gm_n1688);
	nand (gm_n1698, gm_n1671, gm_n1653, gm_n1650, gm_n1697, gm_n1682);
	not (gm_n1699, gm_n1185);
	nand (gm_n1700, gm_n650, in_17, in_13, gm_n1131, gm_n735);
	nor (gm_n1701, gm_n535, gm_n53, gm_n81, gm_n1700, gm_n1699);
	nand (gm_n1702, gm_n50, gm_n96, gm_n76, gm_n1701);
	not (gm_n1703, gm_n73);
	nand (gm_n1704, gm_n66, in_15, in_11, gm_n621, gm_n540);
	nor (gm_n1705, gm_n1703, in_23, in_19, gm_n1704, gm_n911);
	nand (gm_n1706, gm_n173, gm_n50, gm_n133, gm_n1705, gm_n677);
	nor (gm_n1707, gm_n89, in_12, gm_n64, gm_n160, gm_n167);
	nand (gm_n1708, gm_n137, gm_n72, in_16, gm_n1707, gm_n198);
	nor (gm_n1709, gm_n101, in_28, gm_n52, gm_n1708, gm_n135);
	nand (gm_n1710, gm_n1709, gm_n186);
	nand (gm_n1711, gm_n1710, gm_n1706, gm_n1702);
	nand (gm_n1712, gm_n188, gm_n68, in_12, gm_n1173, gm_n146);
	nor (gm_n1713, gm_n516, in_24, in_20, gm_n1712, gm_n413);
	nand (gm_n1714, gm_n186, gm_n134, in_28, gm_n1713);
	nor (gm_n1715, in_7, in_6, gm_n62, gm_n254, in_8);
	nand (gm_n1716, gm_n188, gm_n69, in_15, gm_n1715, gm_n621);
	nor (gm_n1717, gm_n174, in_23, in_19, gm_n1716, gm_n510);
	nand (gm_n1718, gm_n304, in_31, gm_n133, gm_n1717);
	and (gm_n1719, gm_n121, gm_n62, gm_n123, gm_n539, in_7);
	nand (gm_n1720, gm_n120, gm_n105, in_11, gm_n1719, gm_n621);
	nor (gm_n1721, gm_n300, in_23, gm_n102, gm_n1720, gm_n314);
	nand (gm_n1722, gm_n129, in_31, gm_n133, gm_n1721, gm_n677);
	nand (gm_n1723, gm_n1722, gm_n1718, gm_n1714);
	nor (gm_n1724, gm_n1698, gm_n1646, gm_n1642, gm_n1723, gm_n1711);
	nor (gm_n1725, gm_n221, gm_n157, gm_n64, gm_n598, gm_n253);
	nand (gm_n1726, gm_n183, gm_n72, gm_n68, gm_n1725, gm_n472);
	nor (gm_n1727, gm_n80, in_28, gm_n52, gm_n1726, gm_n475);
	nand (gm_n1728, gm_n587, gm_n210, gm_n64);
	nor (gm_n1729, gm_n88, in_16, gm_n157, gm_n1728, gm_n168);
	nand (gm_n1730, gm_n219, in_24, in_20, gm_n1729, gm_n196);
	nor (gm_n1731, gm_n260, gm_n218, gm_n78, gm_n1730);
	nand (gm_n1732, gm_n705, gm_n63);
	nor (gm_n1733, gm_n366, gm_n105, gm_n58, gm_n1732, gm_n666);
	nand (gm_n1734, gm_n394, in_23, in_19, gm_n1733, gm_n509);
	nor (gm_n1735, gm_n174, gm_n50, gm_n133, gm_n1734, gm_n842);
	nor (gm_n1736, gm_n1735, gm_n1731, gm_n1727);
	nand (gm_n1737, gm_n140, gm_n124, gm_n64);
	nor (gm_n1738, gm_n88, gm_n68, gm_n157, gm_n1737, gm_n139);
	nand (gm_n1739, gm_n209, in_24, gm_n72, gm_n1738, gm_n230);
	nor (gm_n1740, gm_n687, gm_n216, gm_n78, gm_n1739);
	nand (gm_n1741, in_8, in_4, gm_n60, gm_n141, gm_n140);
	nor (gm_n1742, gm_n107, in_16, gm_n157, gm_n1741, gm_n139);
	nand (gm_n1743, gm_n219, in_24, in_20, gm_n1742, gm_n209);
	nor (gm_n1744, gm_n206, gm_n135, in_28, gm_n1743);
	nor (gm_n1745, gm_n88, in_16, in_12, gm_n1025, gm_n158);
	nand (gm_n1746, gm_n85, in_24, in_20, gm_n1745, gm_n261);
	nor (gm_n1747, gm_n132, gm_n216, in_28, gm_n1746);
	nor (gm_n1748, gm_n1747, gm_n1744, gm_n1740);
	nand (gm_n1749, gm_n1724, gm_n1638, gm_n1634, gm_n1748, gm_n1736);
	nor (gm_n1750, gm_n733, gm_n562, gm_n64);
	nand (gm_n1751, gm_n188, in_16, gm_n157, gm_n1750, gm_n198);
	nor (gm_n1752, gm_n156, in_24, in_20, gm_n1751, gm_n804);
	nand (gm_n1753, gm_n205, gm_n79, gm_n78, gm_n1752);
	and (gm_n1754, gm_n211, gm_n147, in_8, gm_n262);
	nand (gm_n1755, gm_n299, in_19, gm_n105, gm_n1754, gm_n1232);
	nor (gm_n1756, gm_n294, gm_n133, gm_n195, gm_n1755, gm_n1231);
	nand (gm_n1757, gm_n1756, gm_n304, in_31);
	and (gm_n1758, gm_n238, gm_n210);
	nand (gm_n1759, gm_n297, in_15, gm_n58, gm_n1758, gm_n427);
	nor (gm_n1760, gm_n117, gm_n195, gm_n102, gm_n1759, gm_n510);
	nand (gm_n1761, gm_n339, in_31, gm_n133, gm_n1760, gm_n455);
	nand (gm_n1762, gm_n1761, gm_n1757, gm_n1753);
	nand (gm_n1763, gm_n180, gm_n68, in_12, gm_n1337, gm_n198);
	nor (gm_n1764, gm_n156, in_24, gm_n72, gm_n1763, gm_n561);
	nand (gm_n1765, gm_n207, gm_n194, in_28, gm_n1764);
	and (gm_n1766, gm_n180, gm_n157, in_8, gm_n705, gm_n110);
	nand (gm_n1767, gm_n198, gm_n72, in_16, gm_n1766, gm_n269);
	nor (gm_n1768, gm_n216, in_28, gm_n52, gm_n1767, gm_n197);
	nand (gm_n1769, gm_n1768, gm_n186);
	and (gm_n1770, gm_n141, in_4, gm_n60, gm_n511);
	nand (gm_n1771, gm_n449, gm_n105, in_11, gm_n1770, gm_n938);
	nor (gm_n1772, gm_n70, in_23, gm_n102, gm_n1771, gm_n423);
	nand (gm_n1773, gm_n129, gm_n50, in_27, gm_n1772, gm_n508);
	nand (gm_n1774, gm_n1773, gm_n1769, gm_n1765);
	nor (gm_n1775, gm_n1749, gm_n1630, gm_n1626, gm_n1774, gm_n1762);
	and (gm_n1776, gm_n146, in_16, in_12, gm_n1361, gm_n147);
	nand (gm_n1777, gm_n261, in_24, gm_n72, gm_n1776, gm_n269);
	nor (gm_n1778, gm_n218, gm_n80, in_28, gm_n1777);
	nor (gm_n1779, gm_n106, gm_n68, in_12, gm_n1303, gm_n245);
	nand (gm_n1780, gm_n137, in_24, gm_n72, gm_n1779, gm_n209);
	nor (gm_n1781, gm_n218, gm_n208, in_28, gm_n1780);
	nand (gm_n1782, gm_n403, gm_n511, in_8);
	nor (gm_n1783, gm_n139, gm_n68, gm_n157, gm_n1782, gm_n159);
	nand (gm_n1784, gm_n220, in_24, in_20, gm_n1783, gm_n517);
	nor (gm_n1785, gm_n371, gm_n218, gm_n78, gm_n1784);
	nor (gm_n1786, gm_n1785, gm_n1781, gm_n1778);
	nand (gm_n1787, gm_n85, in_24, gm_n72, gm_n929, gm_n261);
	nor (gm_n1788, gm_n371, gm_n206, in_28, gm_n1787);
	nand (gm_n1789, gm_n262, gm_n157, gm_n64, gm_n309, gm_n341);
	nor (gm_n1790, gm_n244, gm_n72, in_16, gm_n1789, gm_n602);
	nand (gm_n1791, gm_n134, gm_n78, in_24, gm_n1790, gm_n196);
	nor (gm_n1792, gm_n1791, gm_n229);
	nor (gm_n1793, gm_n673, gm_n105, gm_n58, gm_n1214, gm_n426);
	nand (gm_n1794, gm_n165, in_23, in_19, gm_n1793, gm_n166);
	nor (gm_n1795, gm_n575, in_31, gm_n133, gm_n1794, gm_n671);
	nor (gm_n1796, gm_n1795, gm_n1792, gm_n1788);
	nand (gm_n1797, gm_n1775, gm_n1622, gm_n1617, gm_n1796, gm_n1786);
	nand (gm_n1798, gm_n189, gm_n68, in_12, gm_n512, gm_n232);
	nor (gm_n1799, gm_n178, gm_n52, gm_n72, gm_n1798, gm_n516);
	nand (gm_n1800, gm_n492, gm_n177, gm_n78, gm_n1799);
	nand (gm_n1801, gm_n199, gm_n59, gm_n90, gm_n123, in_3);
	nor (gm_n1802, gm_n385, gm_n1801);
	nand (gm_n1803, gm_n665, in_15, gm_n58, gm_n1802, gm_n1232);
	nor (gm_n1804, gm_n423, in_23, gm_n102, gm_n1803, gm_n453);
	nand (gm_n1805, gm_n129, in_31, in_27, gm_n1804, gm_n437);
	nand (gm_n1806, gm_n281, gm_n63);
	or (gm_n1807, gm_n158, gm_n157, in_8, gm_n1806, gm_n159);
	nor (gm_n1808, gm_n84, in_20, gm_n68, gm_n1807, gm_n187);
	nand (gm_n1809, gm_n134, in_28, in_24, gm_n1808, gm_n492);
	nand (gm_n1810, gm_n1809, gm_n1805, gm_n1800);
	nand (gm_n1811, gm_n200, gm_n140, gm_n64);
	nor (gm_n1812, gm_n179, in_16, gm_n157, gm_n1811, gm_n245);
	nand (gm_n1813, gm_n100, in_24, in_20, gm_n1812, gm_n137);
	nor (gm_n1814, gm_n475, gm_n243, in_28, gm_n1813);
	nor (out_6, gm_n1810, gm_n1797, gm_n1614, gm_n1814);
	nor (gm_n1816, gm_n593, gm_n89, in_8);
	and (gm_n1817, gm_n138, in_16, in_12, gm_n1816, gm_n341);
	nand (gm_n1818, gm_n83, in_24, in_20, gm_n1817, gm_n269);
	nor (gm_n1819, gm_n268, gm_n135, gm_n78, gm_n1818);
	or (gm_n1820, gm_n244, gm_n68, gm_n157, gm_n225, gm_n88);
	nor (gm_n1821, gm_n187, gm_n52, in_20, gm_n1820, gm_n101);
	nand (gm_n1822, gm_n205, gm_n134, in_28, gm_n1821);
	nand (gm_n1823, gm_n629, in_16, in_12, gm_n1369, gm_n354);
	nor (gm_n1824, gm_n187, gm_n52, gm_n72, gm_n1823, gm_n804);
	nand (gm_n1825, gm_n186, gm_n177, in_28, gm_n1824);
	nor (gm_n1826, gm_n57, gm_n105, gm_n58, gm_n1279, gm_n396);
	nand (gm_n1827, gm_n509, in_23, gm_n102, gm_n1826, gm_n612);
	nor (gm_n1828, gm_n1231, gm_n50, gm_n133, gm_n1827, gm_n303);
	nor (gm_n1829, gm_n576, in_15, gm_n58, gm_n1001, gm_n396);
	nand (gm_n1830, gm_n361, in_23, in_19, gm_n1829, gm_n612);
	nor (gm_n1831, gm_n617, gm_n50, in_27, gm_n1830, gm_n436);
	nand (gm_n1832, gm_n333, gm_n102, gm_n105, gm_n1754, gm_n166);
	nor (gm_n1833, gm_n423, in_27, in_23, gm_n1832, gm_n174);
	nand (gm_n1834, gm_n1833, gm_n115, gm_n50);
	nor (gm_n1835, gm_n169, in_12, in_8, gm_n347, gm_n245);
	nand (gm_n1836, gm_n85, gm_n72, in_16, gm_n1835, gm_n189);
	nor (gm_n1837, gm_n197, gm_n78, in_24, gm_n1836, gm_n371);
	nand (gm_n1838, gm_n1837, gm_n77);
	nand (gm_n1839, gm_n705, gm_n308, gm_n64);
	nor (gm_n1840, gm_n167, gm_n68, gm_n157, gm_n1839, gm_n168);
	nand (gm_n1841, gm_n183, in_24, in_20, gm_n1840, gm_n472);
	nor (gm_n1842, gm_n218, gm_n243, gm_n78, gm_n1841);
	nor (gm_n1843, gm_n504, gm_n157, in_8, gm_n499, gm_n286);
	nand (gm_n1844, gm_n83, gm_n72, in_16, gm_n1843, gm_n85);
	nor (gm_n1845, gm_n216, gm_n78, in_24, gm_n1844, gm_n475);
	nor (gm_n1846, gm_n224, gm_n223, in_8);
	nand (gm_n1847, gm_n766, in_16, gm_n157, gm_n1846, gm_n346);
	nor (gm_n1848, gm_n187, in_24, in_20, gm_n1847, gm_n628);
	nand (gm_n1849, gm_n217, gm_n79, gm_n78, gm_n1848);
	nor (gm_n1850, gm_n347, gm_n65, gm_n64, gm_n544);
	nor (gm_n1851, gm_n157, gm_n58, in_10);
	and (gm_n1852, gm_n321, in_17, in_13, gm_n1851, gm_n1850);
	and (gm_n1853, gm_n408, in_25, gm_n81, gm_n1852, gm_n526);
	nand (gm_n1854, gm_n50, gm_n96, in_29, gm_n1853, gm_n738);
	nor (gm_n1855, gm_n106, in_16, gm_n157, gm_n826, gm_n222);
	nand (gm_n1856, gm_n209, gm_n52, in_20, gm_n1855, gm_n230);
	nor (gm_n1857, gm_n135, gm_n132, in_28, gm_n1856);
	nor (gm_n1858, gm_n159, in_12, gm_n64, gm_n386, gm_n168);
	nand (gm_n1859, gm_n219, in_20, in_16, gm_n1858, gm_n252);
	nor (gm_n1860, gm_n132, gm_n78, in_24, gm_n1859, gm_n780);
	nor (gm_n1861, gm_n167, gm_n157, gm_n64, gm_n1533, gm_n179);
	nand (gm_n1862, gm_n219, gm_n72, in_16, gm_n1861, gm_n183);
	nor (gm_n1863, gm_n132, gm_n78, in_24, gm_n1862, gm_n135);
	nand (gm_n1864, gm_n61, gm_n157, in_8, gm_n270, gm_n140);
	nor (gm_n1865, gm_n244, gm_n72, gm_n68, gm_n1864, gm_n742);
	nand (gm_n1866, gm_n79, in_28, in_24, gm_n1865, gm_n252);
	nor (gm_n1867, gm_n1866, gm_n475);
	nor (gm_n1868, gm_n244, gm_n68, gm_n157, gm_n170, gm_n107);
	nand (gm_n1869, gm_n137, gm_n52, gm_n72, gm_n1868, gm_n196);
	nor (gm_n1870, gm_n260, gm_n218, gm_n78, gm_n1869);
	nor (gm_n1871, gm_n1863, gm_n1860, gm_n1857, gm_n1870, gm_n1867);
	nor (gm_n1872, gm_n142, gm_n105, in_11, gm_n399, gm_n319);
	nand (gm_n1873, gm_n313, in_23, in_19, gm_n1872, gm_n394);
	nor (gm_n1874, gm_n1118, gm_n50, in_27, gm_n1873, gm_n575);
	nor (gm_n1875, gm_n673, in_15, in_11, gm_n398, gm_n366);
	nand (gm_n1876, gm_n582, gm_n195, gm_n102, gm_n1875, gm_n165);
	nor (gm_n1877, gm_n671, in_31, gm_n133, gm_n1876, gm_n678);
	or (gm_n1878, gm_n223, in_12, in_8, gm_n544, gm_n245);
	nor (gm_n1879, gm_n106, in_20, in_16, gm_n1878, gm_n742);
	nand (gm_n1880, gm_n177, in_28, gm_n52, gm_n1879, gm_n261);
	nor (gm_n1881, gm_n1880, gm_n218);
	nor (gm_n1882, gm_n1881, gm_n1877, gm_n1874);
	nor (gm_n1883, gm_n672, gm_n105, gm_n58, gm_n598, gm_n673);
	nand (gm_n1884, gm_n69, gm_n195, in_19, gm_n1883, gm_n336);
	nor (gm_n1885, gm_n617, gm_n50, in_27, gm_n1884, gm_n575);
	nor (gm_n1886, gm_n106, gm_n68, gm_n157, gm_n287, gm_n167);
	nand (gm_n1887, gm_n219, in_24, gm_n72, gm_n1886, gm_n220);
	nor (gm_n1888, gm_n260, gm_n229, in_28, gm_n1887);
	or (gm_n1889, gm_n385, gm_n224, in_8);
	nor (gm_n1890, gm_n168, in_16, in_12, gm_n1889, gm_n253);
	nand (gm_n1891, gm_n230, in_24, in_20, gm_n1890, gm_n252);
	nor (gm_n1892, gm_n260, gm_n218, in_28, gm_n1891);
	nor (gm_n1893, gm_n1892, gm_n1888, gm_n1885);
	nand (gm_n1894, gm_n1871, gm_n1854, gm_n1849, gm_n1893, gm_n1882);
	and (gm_n1895, gm_n511, gm_n238, gm_n64);
	nand (gm_n1896, gm_n147, in_16, in_12, gm_n1895, gm_n766);
	nor (gm_n1897, gm_n187, in_24, in_20, gm_n1896, gm_n516);
	nand (gm_n1898, gm_n217, gm_n134, in_28, gm_n1897);
	or (gm_n1899, in_21, in_20);
	nor (gm_n1900, gm_n253, gm_n157, in_8, gm_n385, gm_n355);
	nand (gm_n1901, gm_n136, in_14, in_13, gm_n1900, gm_n482);
	nor (gm_n1902, in_25, in_24, gm_n195);
	not (gm_n1903, gm_n1902);
	nor (gm_n1904, gm_n1899, in_22, gm_n102, gm_n1903, gm_n1901);
	nor (gm_n1905, in_29, gm_n78, in_27);
	nand (gm_n1906, gm_n50, gm_n96, gm_n98, gm_n1905, gm_n1904);
	and (gm_n1907, gm_n109, in_6, gm_n62, gm_n364);
	nand (gm_n1908, gm_n138, in_12, gm_n64, gm_n1907, gm_n232);
	nor (gm_n1909, gm_n84, gm_n72, in_16, gm_n1908, gm_n103);
	nand (gm_n1910, gm_n177, in_28, gm_n52, gm_n1909, gm_n186);
	nand (gm_n1911, gm_n1910, gm_n1906, gm_n1898);
	nor (gm_n1912, gm_n245, in_8, in_7, gm_n530);
	nand (gm_n1913, gm_n362, in_19, gm_n105, gm_n1912, gm_n938);
	nor (gm_n1914, gm_n1703, in_27, in_23, gm_n1913, gm_n617);
	nand (gm_n1915, gm_n1914, gm_n306, in_31);
	nand (gm_n1916, gm_n180, in_16, gm_n157, gm_n557, gm_n766);
	nor (gm_n1917, gm_n103, in_24, gm_n72, gm_n1916, gm_n412);
	nand (gm_n1918, gm_n99, gm_n77, in_28, gm_n1917);
	nand (gm_n1919, gm_n270, in_16, gm_n157, gm_n1547, gm_n629);
	nor (gm_n1920, gm_n84, in_24, gm_n72, gm_n1919, gm_n413);
	nand (gm_n1921, gm_n207, gm_n186, in_28, gm_n1920);
	nand (gm_n1922, gm_n1921, gm_n1918, gm_n1915);
	nor (gm_n1923, gm_n1894, gm_n1845, gm_n1842, gm_n1922, gm_n1911);
	and (gm_n1924, gm_n189, gm_n68, in_12, gm_n356, gm_n147);
	nand (gm_n1925, gm_n237, in_24, gm_n72, gm_n1924, gm_n220);
	nor (gm_n1926, gm_n780, gm_n206, in_28, gm_n1925);
	nand (gm_n1927, gm_n270, in_12, gm_n64, gm_n587, gm_n511);
	nor (gm_n1928, gm_n103, in_20, in_16, gm_n1927, gm_n179);
	nand (gm_n1929, gm_n220, gm_n78, gm_n52, gm_n1928, gm_n462);
	nor (gm_n1930, gm_n1929, gm_n206);
	nor (gm_n1931, gm_n168, gm_n157, in_8, gm_n1806, gm_n253);
	nand (gm_n1932, gm_n219, gm_n72, gm_n68, gm_n1931, gm_n183);
	nor (gm_n1933, gm_n371, gm_n78, in_24, gm_n1932, gm_n475);
	nor (gm_n1934, gm_n1933, gm_n1930, gm_n1926);
	nor (gm_n1935, gm_n221, in_16, gm_n157, gm_n1123, gm_n253);
	nand (gm_n1936, gm_n237, gm_n52, gm_n72, gm_n1935, gm_n183);
	nor (gm_n1937, gm_n218, gm_n243, in_28, gm_n1936);
	and (gm_n1938, gm_n147, gm_n68, in_12, gm_n987, gm_n629);
	nand (gm_n1939, gm_n100, in_24, in_20, gm_n1938, gm_n219);
	nor (gm_n1940, gm_n260, gm_n218, gm_n78, gm_n1939);
	and (gm_n1941, gm_n66, in_15, gm_n58, gm_n540, gm_n938);
	nand (gm_n1942, gm_n126, gm_n195, in_19, gm_n1941, gm_n299);
	nor (gm_n1943, gm_n54, in_31, in_27, gm_n1942, gm_n611);
	nor (gm_n1944, gm_n1943, gm_n1940, gm_n1937);
	nand (gm_n1945, gm_n1923, gm_n1838, gm_n1834, gm_n1944, gm_n1934);
	nand (gm_n1946, gm_n619, gm_n511);
	or (gm_n1947, gm_n119, in_15, gm_n58, gm_n1946, gm_n997);
	nor (gm_n1948, gm_n294, in_23, in_19, gm_n1947, gm_n395);
	nand (gm_n1949, gm_n55, gm_n50, in_27, gm_n1948, gm_n677);
	or (gm_n1950, gm_n396, in_15, gm_n58, gm_n1806, gm_n399);
	nor (gm_n1951, gm_n294, in_23, in_19, gm_n1950, gm_n300);
	nand (gm_n1952, gm_n455, gm_n50, gm_n133, gm_n1951, gm_n677);
	nor (gm_n1953, gm_n295, gm_n223);
	nand (gm_n1954, gm_n189, in_12, gm_n64, gm_n1953, gm_n354);
	nor (gm_n1955, gm_n412, gm_n72, gm_n68, gm_n1954, gm_n413);
	nand (gm_n1956, gm_n259, in_28, gm_n52, gm_n1955, gm_n474);
	nand (gm_n1957, gm_n1956, gm_n1952, gm_n1949);
	nand (gm_n1958, gm_n766, gm_n68, gm_n157, gm_n377, gm_n341);
	nor (gm_n1959, gm_n156, gm_n52, in_20, gm_n1958, gm_n561);
	nand (gm_n1960, gm_n492, gm_n462, gm_n78, gm_n1959);
	nand (gm_n1961, gm_n333, gm_n105, gm_n58, gm_n1201, gm_n665);
	nor (gm_n1962, gm_n117, in_23, gm_n102, gm_n1961, gm_n314);
	nand (gm_n1963, gm_n173, gm_n50, gm_n133, gm_n1962, gm_n677);
	nand (gm_n1964, gm_n146, in_16, in_12, gm_n758, gm_n354);
	nor (gm_n1965, gm_n459, in_24, gm_n72, gm_n1964, gm_n628);
	nand (gm_n1966, gm_n205, gm_n177, in_28, gm_n1965);
	nand (gm_n1967, gm_n1966, gm_n1963, gm_n1960);
	nor (gm_n1968, gm_n1945, gm_n1831, gm_n1828, gm_n1967, gm_n1957);
	nor (gm_n1969, gm_n673, in_15, in_11, gm_n583, gm_n426);
	nand (gm_n1970, gm_n293, gm_n195, in_19, gm_n1969, gm_n299);
	nor (gm_n1971, gm_n54, in_31, gm_n133, gm_n1970, gm_n303);
	nand (gm_n1972, gm_n110, in_12, gm_n64, gm_n498, gm_n232);
	nor (gm_n1973, gm_n244, in_20, in_16, gm_n1972, gm_n602);
	nand (gm_n1974, gm_n79, in_28, gm_n52, gm_n1973, gm_n220);
	nor (gm_n1975, gm_n1974, gm_n475);
	nor (gm_n1976, gm_n432, in_15, gm_n58, gm_n1259, gm_n366);
	nand (gm_n1977, gm_n165, in_23, gm_n102, gm_n1976, gm_n452);
	nor (gm_n1978, gm_n51, gm_n50, gm_n133, gm_n1977, gm_n174);
	nor (gm_n1979, gm_n1978, gm_n1975, gm_n1971);
	nor (gm_n1980, gm_n244, gm_n68, gm_n157, gm_n1294, gm_n253);
	nand (gm_n1981, gm_n261, in_24, in_20, gm_n1980, gm_n269);
	nor (gm_n1982, gm_n475, gm_n216, gm_n78, gm_n1981);
	nor (gm_n1983, gm_n395, gm_n102, gm_n105, gm_n932, gm_n399);
	nand (gm_n1984, gm_n126, gm_n133, gm_n195, gm_n1983, gm_n393);
	nor (gm_n1985, gm_n1984, gm_n360, gm_n50);
	nand (gm_n1986, gm_n109, in_6, in_5, gm_n364, gm_n64);
	nor (gm_n1987, gm_n179, gm_n68, gm_n157, gm_n1986, gm_n245);
	nand (gm_n1988, gm_n237, gm_n52, gm_n72, gm_n1987, gm_n209);
	nor (gm_n1989, gm_n218, gm_n208, gm_n78, gm_n1988);
	nor (gm_n1990, gm_n1989, gm_n1985, gm_n1982);
	nand (gm_n1991, gm_n1968, gm_n1825, gm_n1822, gm_n1990, gm_n1979);
	nand (gm_n1992, gm_n86, in_16, in_12, gm_n789, gm_n354);
	nor (gm_n1993, gm_n178, in_24, gm_n72, gm_n1992, gm_n804);
	nand (gm_n1994, gm_n99, gm_n97, in_28, gm_n1993);
	or (gm_n1995, in_9, in_8, in_7);
	nor (gm_n1996, gm_n87, gm_n121, gm_n62, gm_n1995, gm_n355);
	nand (gm_n1997, gm_n582, in_15, in_11, gm_n1996, gm_n118);
	nor (gm_n1998, gm_n617, gm_n195, gm_n102, gm_n1997, gm_n510);
	nand (gm_n1999, gm_n508, gm_n50, in_27, gm_n1998);
	and (gm_n2000, gm_n587, gm_n262, in_8);
	nand (gm_n2001, gm_n189, in_16, gm_n157, gm_n2000, gm_n341);
	nor (gm_n2002, gm_n197, gm_n52, in_20, gm_n2001, gm_n742);
	nand (gm_n2003, gm_n207, gm_n205, gm_n78, gm_n2002);
	nand (gm_n2004, gm_n2003, gm_n1999, gm_n1994);
	and (gm_n2005, gm_n511, gm_n232, gm_n64, gm_n705);
	and (gm_n2006, gm_n333, gm_n102, gm_n105, gm_n2005, gm_n394);
	nand (gm_n2007, gm_n126, in_27, in_23, gm_n2006, gm_n173);
	nor (gm_n2008, gm_n2007, gm_n360, gm_n50);
	nor (out_7, gm_n2004, gm_n1991, gm_n1819, gm_n2008);
	nor (gm_n2010, gm_n244, gm_n68, in_12, gm_n902, gm_n107);
	nand (gm_n2011, gm_n209, in_24, in_20, gm_n2010, gm_n230);
	nor (gm_n2012, gm_n260, gm_n218, gm_n78, gm_n2011);
	nor (gm_n2013, in_12, in_11, gm_n87);
	nand (gm_n2014, gm_n528, gm_n116, gm_n56, gm_n2013, gm_n1850);
	nand (gm_n2015, in_24, gm_n195, gm_n82);
	nor (gm_n2016, gm_n151, in_25, in_21, gm_n2015, gm_n2014);
	nand (gm_n2017, gm_n50, in_30, gm_n76, gm_n2016, gm_n1686);
	and (gm_n2018, gm_n587, gm_n122, gm_n64);
	nand (gm_n2019, gm_n189, in_16, in_12, gm_n2018, gm_n147);
	nor (gm_n2020, gm_n804, gm_n52, gm_n72, gm_n2019, gm_n413);
	nand (gm_n2021, gm_n259, gm_n194, gm_n78, gm_n2020);
	nand (gm_n2022, gm_n110, gm_n157, gm_n64, gm_n498, gm_n232);
	nor (gm_n2023, gm_n168, gm_n72, gm_n68, gm_n2022, gm_n602);
	nand (gm_n2024, gm_n261, in_28, in_24, gm_n2023, gm_n370);
	nor (gm_n2025, gm_n2024, gm_n176);
	and (gm_n2026, gm_n937, in_15, in_11, gm_n1139, gm_n427);
	nand (gm_n2027, gm_n166, gm_n195, gm_n102, gm_n2026, gm_n361);
	nor (gm_n2028, gm_n54, in_31, gm_n133, gm_n2027, gm_n303);
	and (gm_n2029, gm_n122, gm_n61);
	nand (gm_n2030, gm_n66, in_15, in_11, gm_n427, gm_n2029);
	nor (gm_n2031, gm_n70, gm_n195, gm_n102, gm_n2030, gm_n127);
	nand (gm_n2032, gm_n455, gm_n50, gm_n133, gm_n2031, gm_n508);
	nand (gm_n2033, gm_n231, gm_n68, gm_n157, gm_n630, gm_n354);
	nor (gm_n2034, gm_n459, gm_n52, gm_n72, gm_n2033, gm_n628);
	nand (gm_n2035, gm_n217, gm_n79, gm_n78, gm_n2034);
	and (gm_n2036, gm_n146, gm_n68, in_12, gm_n1547, gm_n147);
	nand (gm_n2037, gm_n219, gm_n52, gm_n72, gm_n2036, gm_n220);
	nor (gm_n2038, gm_n475, gm_n216, in_28, gm_n2037);
	or (gm_n2039, in_7, in_6, gm_n62, gm_n544, gm_n64);
	nor (gm_n2040, gm_n107, in_16, in_12, gm_n2039, gm_n139);
	nand (gm_n2041, gm_n85, in_24, gm_n72, gm_n2040, gm_n252);
	nor (gm_n2042, gm_n260, gm_n268, in_28, gm_n2041);
	nand (gm_n2043, gm_n629, gm_n68, gm_n157, gm_n1155, gm_n354);
	nor (gm_n2044, gm_n561, in_24, in_20, gm_n2043, gm_n742);
	nand (gm_n2045, gm_n217, gm_n79, gm_n78, gm_n2044);
	nor (gm_n2046, gm_n465, gm_n385, gm_n64);
	nand (gm_n2047, gm_n188, in_16, in_12, gm_n2046, gm_n766);
	nor (gm_n2048, gm_n412, gm_n52, gm_n72, gm_n2047, gm_n413);
	nand (gm_n2049, gm_n370, gm_n194, gm_n78, gm_n2048);
	nor (gm_n2050, gm_n106, gm_n68, in_12, gm_n1050, gm_n253);
	nand (gm_n2051, gm_n83, in_24, in_20, gm_n2050, gm_n472);
	nor (gm_n2052, gm_n268, gm_n216, gm_n78, gm_n2051);
	nand (gm_n2053, gm_n450, gm_n511, in_8);
	nor (gm_n2054, gm_n504, gm_n68, gm_n157, gm_n2053, gm_n245);
	nand (gm_n2055, gm_n83, gm_n52, gm_n72, gm_n2054, gm_n85);
	nor (gm_n2056, gm_n206, gm_n216, in_28, gm_n2055);
	nor (gm_n2057, gm_n395, gm_n102, gm_n105, gm_n932, gm_n622);
	nand (gm_n2058, gm_n165, gm_n133, gm_n195, gm_n2057, gm_n658);
	nor (gm_n2059, gm_n2058, gm_n303, gm_n50);
	nand (gm_n2060, gm_n309, gm_n140, in_8);
	nor (gm_n2061, gm_n107, gm_n68, in_12, gm_n2060, gm_n158);
	nand (gm_n2062, gm_n237, gm_n52, in_20, gm_n2061, gm_n252);
	nor (gm_n2063, gm_n268, gm_n243, gm_n78, gm_n2062);
	and (gm_n2064, gm_n362, gm_n354, in_15, gm_n645, gm_n621);
	nand (gm_n2065, gm_n126, gm_n195, gm_n102, gm_n2064, gm_n455);
	nor (gm_n2066, gm_n575, gm_n50, gm_n133, gm_n2065);
	nor (gm_n2067, gm_n2059, gm_n2056, gm_n2052, gm_n2066, gm_n2063);
	nor (gm_n2068, gm_n139, gm_n157, in_11, gm_n762, gm_n673);
	nand (gm_n2069, gm_n137, in_20, gm_n68, gm_n2068, gm_n209);
	nor (gm_n2070, gm_n216, in_28, in_24, gm_n2069, gm_n687);
	nor (gm_n2071, gm_n167, in_16, gm_n157, gm_n1365, gm_n158);
	nand (gm_n2072, gm_n83, gm_n52, gm_n72, gm_n2071, gm_n472);
	nor (gm_n2073, gm_n687, gm_n243, gm_n78, gm_n2072);
	nand (gm_n2074, gm_n293, in_23, in_19, gm_n1144, gm_n612);
	nor (gm_n2075, gm_n575, gm_n50, in_27, gm_n2074, gm_n671);
	nor (gm_n2076, gm_n2075, gm_n2073, gm_n2070);
	nand (gm_n2077, gm_n308, gm_n61, in_8);
	nor (gm_n2078, gm_n167, gm_n672, in_15, gm_n2077, gm_n911);
	nand (gm_n2079, gm_n302, gm_n195, in_19, gm_n2078, gm_n509);
	nor (gm_n2080, gm_n575, gm_n50, gm_n133, gm_n2079);
	nand (gm_n2081, gm_n403, gm_n63);
	nor (gm_n2082, gm_n396, in_15, in_11, gm_n2081, gm_n399);
	nand (gm_n2083, gm_n73, in_23, gm_n102, gm_n2082, gm_n362);
	nor (gm_n2084, gm_n842, in_31, gm_n133, gm_n2083, gm_n983);
	nand (gm_n2085, gm_n1226, gm_n210);
	nor (gm_n2086, gm_n666, gm_n105, in_11, gm_n2085, gm_n997);
	nand (gm_n2087, gm_n293, gm_n195, in_19, gm_n2086, gm_n299);
	nor (gm_n2088, gm_n1231, gm_n50, in_27, gm_n2087, gm_n436);
	nor (gm_n2089, gm_n2088, gm_n2084, gm_n2080);
	nand (gm_n2090, gm_n2067, gm_n2049, gm_n2045, gm_n2089, gm_n2076);
	nand (gm_n2091, gm_n86, gm_n72, gm_n68, gm_n472, gm_n239);
	nor (gm_n2092, gm_n197, in_28, gm_n52, gm_n2091, gm_n780);
	nand (gm_n2093, gm_n2092, gm_n492);
	nand (gm_n2094, gm_n146, in_16, in_12, gm_n1895, gm_n232);
	nor (gm_n2095, gm_n156, gm_n52, gm_n72, gm_n2094, gm_n628);
	nand (gm_n2096, gm_n99, gm_n97, gm_n78, gm_n2095);
	nand (gm_n2097, gm_n938, gm_n105, in_11, gm_n1683, gm_n425);
	nor (gm_n2098, gm_n70, gm_n195, gm_n102, gm_n2097, gm_n314);
	nand (gm_n2099, gm_n339, gm_n50, gm_n133, gm_n2098, gm_n455);
	nand (gm_n2100, gm_n2099, gm_n2096, gm_n2093);
	nand (gm_n2101, gm_n66, in_15, gm_n58, gm_n1319, gm_n427);
	nor (gm_n2102, gm_n70, gm_n195, in_19, gm_n2101, gm_n314);
	nand (gm_n2103, gm_n393, in_31, in_27, gm_n2102, gm_n677);
	and (gm_n2104, gm_n587, gm_n63, in_8);
	nand (gm_n2105, gm_n146, in_16, in_12, gm_n2104, gm_n346);
	nor (gm_n2106, gm_n101, in_24, gm_n72, gm_n2105, gm_n156);
	nand (gm_n2107, gm_n177, gm_n194, gm_n78, gm_n2106);
	or (gm_n2108, gm_n57, in_15, gm_n58, gm_n762, gm_n119);
	nor (gm_n2109, gm_n1703, gm_n195, in_19, gm_n2108, gm_n117);
	nand (gm_n2110, gm_n115, gm_n50, in_27, gm_n2109, gm_n173);
	nand (gm_n2111, gm_n2110, gm_n2107, gm_n2103);
	nor (gm_n2112, gm_n2090, gm_n2042, gm_n2038, gm_n2111, gm_n2100);
	nor (gm_n2113, gm_n672, gm_n105, gm_n58, gm_n673, gm_n282);
	nand (gm_n2114, gm_n582, gm_n195, gm_n102, gm_n2113, gm_n165);
	nor (gm_n2115, gm_n1118, gm_n50, in_27, gm_n2114, gm_n436);
	and (gm_n2116, gm_n188, gm_n333, gm_n105, gm_n889, gm_n166);
	nand (gm_n2117, gm_n455, in_23, gm_n102, gm_n2116, gm_n509);
	nor (gm_n2118, gm_n678, in_31, in_27, gm_n2117);
	nand (gm_n2119, gm_n180, gm_n157, gm_n64, gm_n403, gm_n140);
	nor (gm_n2120, gm_n179, gm_n72, gm_n68, gm_n2119, gm_n742);
	nand (gm_n2121, gm_n259, in_28, gm_n52, gm_n2120, gm_n261);
	nor (gm_n2122, gm_n2121, gm_n268);
	nor (gm_n2123, gm_n2122, gm_n2118, gm_n2115);
	nand (gm_n2124, gm_n140, gm_n61, gm_n64);
	nor (gm_n2125, gm_n159, gm_n68, in_12, gm_n2124, gm_n179);
	nand (gm_n2126, gm_n209, gm_n52, gm_n72, gm_n2125, gm_n472);
	nor (gm_n2127, gm_n780, gm_n268, in_28, gm_n2126);
	or (gm_n2128, gm_n169, gm_n246, in_8);
	nor (gm_n2129, gm_n244, in_16, gm_n157, gm_n2128, gm_n253);
	nand (gm_n2130, gm_n237, gm_n52, gm_n72, gm_n2129, gm_n261);
	nor (gm_n2131, gm_n218, gm_n80, gm_n78, gm_n2130);
	nor (gm_n2132, gm_n622, in_15, in_11, gm_n762, gm_n666);
	nand (gm_n2133, gm_n313, gm_n195, gm_n102, gm_n2132, gm_n452);
	nor (gm_n2134, gm_n1118, in_31, gm_n133, gm_n2133, gm_n575);
	nor (gm_n2135, gm_n2134, gm_n2131, gm_n2127);
	nand (gm_n2136, gm_n2112, gm_n2035, gm_n2032, gm_n2135, gm_n2123);
	nand (gm_n2137, gm_n118, in_15, gm_n58, gm_n1102, gm_n665);
	nor (gm_n2138, gm_n1703, gm_n195, gm_n102, gm_n2137, gm_n363);
	nand (gm_n2139, gm_n129, gm_n50, in_27, gm_n2138, gm_n306);
	and (gm_n2140, gm_n122, gm_n157, in_8, gm_n567, gm_n270);
	nand (gm_n2141, gm_n146, in_20, in_16, gm_n2140, gm_n517);
	nor (gm_n2142, gm_n216, in_28, gm_n52, gm_n2141, gm_n197);
	nand (gm_n2143, gm_n2142, gm_n77);
	nor (gm_n2144, gm_n465, gm_n223, gm_n64);
	and (gm_n2145, gm_n138, in_16, gm_n157, gm_n2144, gm_n232);
	and (gm_n2146, gm_n83, in_24, gm_n72, gm_n2145, gm_n230);
	nand (gm_n2147, gm_n217, gm_n79, gm_n78, gm_n2146);
	nand (gm_n2148, gm_n2147, gm_n2143, gm_n2139);
	nor (gm_n2149, gm_n347, gm_n1005);
	nand (gm_n2150, gm_n449, in_15, in_11, gm_n2149, gm_n1232);
	nor (gm_n2151, gm_n127, gm_n195, gm_n102, gm_n2150, gm_n395);
	nand (gm_n2152, gm_n173, in_31, in_27, gm_n2151, gm_n677);
	or (gm_n2153, gm_n504, in_16, in_12, gm_n1639, gm_n253);
	nor (gm_n2154, gm_n197, in_24, in_20, gm_n2153, gm_n602);
	nand (gm_n2155, gm_n370, gm_n77, in_28, gm_n2154);
	and (gm_n2156, gm_n120, gm_n63, in_11, gm_n498);
	nand (gm_n2157, gm_n299, in_19, in_15, gm_n2156, gm_n938);
	nor (gm_n2158, gm_n581, in_27, gm_n195, gm_n2157, gm_n510);
	nand (gm_n2159, gm_n2158, gm_n306, in_31);
	nand (gm_n2160, gm_n2159, gm_n2155, gm_n2152);
	nor (gm_n2161, gm_n2136, gm_n2028, gm_n2025, gm_n2160, gm_n2148);
	nand (gm_n2162, gm_n308, gm_n238, gm_n64);
	nor (gm_n2163, gm_n221, in_16, gm_n157, gm_n2162, gm_n245);
	nand (gm_n2164, gm_n100, in_24, gm_n72, gm_n2163, gm_n517);
	nor (gm_n2165, gm_n218, gm_n135, gm_n78, gm_n2164);
	nand (gm_n2166, gm_n308, gm_n263, in_8);
	nor (gm_n2167, gm_n158, in_16, in_12, gm_n2166, gm_n159);
	nand (gm_n2168, gm_n237, gm_n52, in_20, gm_n2167, gm_n183);
	nor (gm_n2169, gm_n260, gm_n229, in_28, gm_n2168);
	nand (gm_n2170, gm_n147, gm_n63, in_8, gm_n1226);
	nor (gm_n2171, gm_n117, gm_n102, in_15, gm_n2170, gm_n576);
	nand (gm_n2172, gm_n165, gm_n133, gm_n195, gm_n2171, gm_n307);
	nor (gm_n2173, gm_n2172, gm_n436, in_31);
	nor (gm_n2174, gm_n2173, gm_n2169, gm_n2165);
	nor (gm_n2175, gm_n106, in_16, in_12, gm_n781, gm_n167);
	nand (gm_n2176, gm_n83, gm_n52, gm_n72, gm_n2175, gm_n219);
	nor (gm_n2177, gm_n475, gm_n260, gm_n78, gm_n2176);
	nand (gm_n2178, gm_n705, gm_n210, gm_n64);
	nor (gm_n2179, gm_n221, gm_n68, in_12, gm_n2178, gm_n222);
	nand (gm_n2180, gm_n261, gm_n52, in_20, gm_n2179, gm_n517);
	nor (gm_n2181, gm_n243, gm_n229, gm_n78, gm_n2180);
	and (gm_n2182, gm_n146, in_16, gm_n157, gm_n377, gm_n270);
	nand (gm_n2183, gm_n196, in_24, gm_n72, gm_n2182, gm_n472);
	nor (gm_n2184, gm_n687, gm_n780, gm_n78, gm_n2183);
	nor (gm_n2185, gm_n2184, gm_n2181, gm_n2177);
	nand (gm_n2186, gm_n2161, gm_n2021, gm_n2017, gm_n2185, gm_n2174);
	or (gm_n2187, gm_n244, in_16, in_12, gm_n264, gm_n253);
	nor (gm_n2188, gm_n101, gm_n52, in_20, gm_n2187, gm_n103);
	nand (gm_n2189, gm_n177, gm_n194, gm_n78, gm_n2188);
	nor (gm_n2190, in_9, gm_n64, gm_n109, gm_n530);
	nor (gm_n2191, in_12, gm_n58, in_10);
	nand (gm_n2192, gm_n405, gm_n116, in_13, gm_n2191, gm_n2190);
	nor (gm_n2193, gm_n1699, gm_n53, in_21, gm_n2192, gm_n1566);
	nand (gm_n2194, gm_n50, gm_n96, in_29, gm_n2193, gm_n409);
	nand (gm_n2195, gm_n200, gm_n122, gm_n64);
	or (gm_n2196, gm_n139, gm_n68, in_12, gm_n2195, gm_n286);
	nor (gm_n2197, gm_n516, in_24, in_20, gm_n2196, gm_n413);
	nand (gm_n2198, gm_n79, gm_n77, in_28, gm_n2197);
	nand (gm_n2199, gm_n2198, gm_n2194, gm_n2189);
	nand (gm_n2200, gm_n140, gm_n157, in_8, gm_n211, gm_n270);
	nor (gm_n2201, gm_n103, in_20, gm_n68, gm_n2200, gm_n106);
	nand (gm_n2202, gm_n134, gm_n78, in_24, gm_n2201, gm_n261);
	nor (gm_n2203, gm_n2202, gm_n176);
	nor (out_8, gm_n2199, gm_n2186, gm_n2012, gm_n2203);
	and (gm_n2205, gm_n188, in_12, in_8, gm_n587, gm_n262);
	and (gm_n2206, gm_n405, in_17, gm_n56, gm_n2205, gm_n1565);
	nand (gm_n2207, gm_n327, in_25, in_21, gm_n2206, gm_n534);
	nor (gm_n2208, gm_n50, gm_n96, gm_n76, gm_n2207);
	nand (gm_n2209, gm_n231, in_16, gm_n157, gm_n2144, gm_n346);
	nor (gm_n2210, gm_n103, gm_n52, gm_n72, gm_n2209, gm_n516);
	nand (gm_n2211, gm_n492, gm_n79, gm_n78, gm_n2210);
	and (gm_n2212, gm_n587, gm_n262, gm_n64);
	nand (gm_n2213, gm_n189, gm_n68, in_12, gm_n2212, gm_n341);
	nor (gm_n2214, gm_n103, in_24, in_20, gm_n2213, gm_n804);
	nand (gm_n2215, gm_n177, gm_n97, in_28, gm_n2214);
	not (gm_n2216, gm_n738);
	nor (gm_n2217, gm_n531, gm_n116, in_13, gm_n1132, gm_n772);
	nand (gm_n2218, gm_n652, gm_n53, in_21, gm_n2217, gm_n1565);
	nor (gm_n2219, gm_n50, gm_n96, gm_n76, gm_n2218, gm_n2216);
	and (gm_n2220, gm_n188, gm_n68, in_12, gm_n1895, gm_n629);
	nand (gm_n2221, gm_n137, gm_n52, in_20, gm_n2220, gm_n261);
	nor (gm_n2222, gm_n780, gm_n132, in_28, gm_n2221);
	and (gm_n2223, gm_n63, in_12, in_8, gm_n263, gm_n188);
	nand (gm_n2224, gm_n137, in_20, gm_n68, gm_n2223, gm_n629);
	nor (gm_n2225, gm_n135, gm_n78, in_24, gm_n2224, gm_n804);
	nand (gm_n2226, gm_n2225, gm_n492);
	nand (gm_n2227, in_14, in_13, in_12, gm_n1393, gm_n147);
	nor (gm_n2228, in_17, gm_n68, in_15, gm_n2227, in_18);
	nor (gm_n2229, gm_n81, in_20, in_19);
	and (gm_n2230, gm_n639, gm_n98, gm_n82, gm_n2229, gm_n2228);
	nor (gm_n2231, in_29, gm_n78, gm_n133);
	nand (gm_n2232, gm_n2230, in_31, gm_n96, gm_n2231);
	nand (gm_n2233, gm_n567, gm_n63);
	nor (gm_n2234, gm_n672, in_15, in_11, gm_n2233, gm_n432);
	nand (gm_n2235, gm_n582, in_23, gm_n102, gm_n2234, gm_n293);
	nor (gm_n2236, gm_n1118, gm_n50, gm_n133, gm_n2235, gm_n575);
	nor (gm_n2237, gm_n1200, gm_n319, gm_n942);
	and (gm_n2238, gm_n938, gm_n105, gm_n58, gm_n2237, gm_n612);
	nand (gm_n2239, gm_n302, gm_n195, in_19, gm_n2238, gm_n336);
	nor (gm_n2240, gm_n842, in_31, in_27, gm_n2239);
	or (gm_n2241, gm_n168, gm_n68, in_12, gm_n1123, gm_n253);
	nor (gm_n2242, gm_n84, gm_n52, gm_n72, gm_n2241, gm_n459);
	nand (gm_n2243, gm_n134, gm_n77, in_28, gm_n2242);
	nor (gm_n2244, gm_n355, gm_n942, gm_n64);
	nand (gm_n2245, gm_n147, gm_n68, gm_n157, gm_n2244, gm_n766);
	nor (gm_n2246, gm_n156, gm_n52, in_20, gm_n2245, gm_n804);
	nand (gm_n2247, gm_n205, gm_n99, in_28, gm_n2246);
	nor (gm_n2248, gm_n88, gm_n68, gm_n157, gm_n1505, gm_n158);
	nand (gm_n2249, gm_n85, in_24, gm_n72, gm_n2248, gm_n183);
	nor (gm_n2250, gm_n780, gm_n229, gm_n78, gm_n2249);
	and (gm_n2251, gm_n231, in_16, gm_n157, gm_n557, gm_n354);
	nand (gm_n2252, gm_n196, gm_n52, in_20, gm_n2251, gm_n269);
	nor (gm_n2253, gm_n243, gm_n229, in_28, gm_n2252);
	or (gm_n2254, gm_n254, gm_n223, gm_n64);
	nor (gm_n2255, gm_n107, gm_n244, gm_n157, gm_n2254);
	nand (gm_n2256, gm_n293, in_23, gm_n102, gm_n2255, gm_n612);
	nor (gm_n2257, gm_n617, in_31, gm_n133, gm_n2256, gm_n575);
	nor (gm_n2258, gm_n363, gm_n105, gm_n58, gm_n1623, gm_n426);
	nand (gm_n2259, gm_n55, gm_n195, in_19, gm_n2258, gm_n293);
	nor (gm_n2260, gm_n51, in_31, gm_n133, gm_n2259);
	nor (gm_n2261, gm_n107, gm_n157, gm_n64, gm_n1533, gm_n221);
	nand (gm_n2262, gm_n85, gm_n72, gm_n68, gm_n2261, gm_n252);
	nor (gm_n2263, gm_n216, gm_n78, gm_n52, gm_n2262, gm_n687);
	nor (gm_n2264, gm_n2257, gm_n2253, gm_n2250, gm_n2263, gm_n2260);
	nand (gm_n2265, gm_n122, gm_n66, in_11, gm_n124);
	nor (gm_n2266, gm_n453, in_19, gm_n105, gm_n2265, gm_n622);
	nand (gm_n2267, gm_n361, in_27, gm_n195, gm_n2266, gm_n658);
	nor (gm_n2268, gm_n2267, gm_n360, gm_n50);
	nor (gm_n2269, gm_n319, gm_n105, gm_n58, gm_n1001, gm_n426);
	nand (gm_n2270, gm_n361, in_23, in_19, gm_n2269, gm_n362);
	nor (gm_n2271, gm_n617, gm_n50, gm_n133, gm_n2270, gm_n611);
	nand (gm_n2272, gm_n238, gm_n140, in_8, gm_n346);
	nor (gm_n2273, gm_n70, in_19, gm_n105, gm_n2272, gm_n426);
	nand (gm_n2274, gm_n129, in_27, gm_n195, gm_n2273, gm_n509);
	nor (gm_n2275, gm_n2274, gm_n303, gm_n50);
	nor (gm_n2276, gm_n2275, gm_n2271, gm_n2268);
	nor (gm_n2277, gm_n70, in_15, in_11, gm_n1657, gm_n399);
	nand (gm_n2278, gm_n302, in_23, gm_n102, gm_n2277, gm_n313);
	nor (gm_n2279, gm_n360, gm_n50, gm_n133, gm_n2278);
	nor (gm_n2280, gm_n363, gm_n105, in_11, gm_n752, gm_n426);
	nand (gm_n2281, gm_n73, gm_n195, in_19, gm_n2280, gm_n129);
	nor (gm_n2282, gm_n303, in_31, in_27, gm_n2281);
	or (gm_n2283, gm_n544, gm_n385);
	nor (gm_n2284, gm_n426, in_15, gm_n58, gm_n2283, gm_n666);
	nand (gm_n2285, gm_n166, in_23, gm_n102, gm_n2284, gm_n336);
	nor (gm_n2286, gm_n51, in_31, gm_n133, gm_n2285, gm_n1231);
	nor (gm_n2287, gm_n2286, gm_n2282, gm_n2279);
	nand (gm_n2288, gm_n2264, gm_n2247, gm_n2243, gm_n2287, gm_n2276);
	nand (gm_n2289, gm_n198, gm_n68, in_12, gm_n987, gm_n232);
	nor (gm_n2290, gm_n187, in_24, gm_n72, gm_n2289, gm_n804);
	nand (gm_n2291, gm_n217, gm_n177, gm_n78, gm_n2290);
	nand (gm_n2292, gm_n166, in_19, gm_n105, gm_n2005, gm_n1232);
	nor (gm_n2293, gm_n127, in_27, gm_n195, gm_n2292, gm_n983);
	nand (gm_n2294, gm_n2293, gm_n437, gm_n50);
	nand (gm_n2295, gm_n180, in_16, in_12, gm_n876, gm_n629);
	nor (gm_n2296, gm_n516, gm_n52, in_20, gm_n2295, gm_n459);
	nand (gm_n2297, gm_n134, gm_n77, in_28, gm_n2296);
	nand (gm_n2298, gm_n2297, gm_n2294, gm_n2291);
	or (gm_n2299, gm_n139, gm_n68, in_12, gm_n781, gm_n159);
	nor (gm_n2300, gm_n187, gm_n52, gm_n72, gm_n2299, gm_n628);
	nand (gm_n2301, gm_n259, gm_n77, in_28, gm_n2300);
	nand (gm_n2302, gm_n270, in_16, gm_n157, gm_n512, gm_n629);
	nor (gm_n2303, gm_n101, in_24, in_20, gm_n2302, gm_n459);
	nand (gm_n2304, gm_n492, gm_n99, in_28, gm_n2303);
	nand (gm_n2305, gm_n138, in_16, in_12, gm_n920, gm_n341);
	nor (gm_n2306, gm_n84, gm_n52, in_20, gm_n2305, gm_n187);
	nand (gm_n2307, gm_n205, gm_n134, in_28, gm_n2306);
	nand (gm_n2308, gm_n2307, gm_n2304, gm_n2301);
	nor (gm_n2309, gm_n2288, gm_n2240, gm_n2236, gm_n2308, gm_n2298);
	and (gm_n2310, gm_n118, gm_n102, gm_n105, gm_n2156, gm_n394);
	nand (gm_n2311, gm_n293, gm_n133, gm_n195, gm_n2310, gm_n393);
	nor (gm_n2312, gm_n2311, gm_n360, in_31);
	nor (gm_n2313, gm_n583, gm_n105, gm_n58, gm_n666, gm_n622);
	nand (gm_n2314, gm_n582, gm_n195, in_19, gm_n2313, gm_n336);
	nor (gm_n2315, gm_n54, gm_n50, in_27, gm_n2314, gm_n360);
	nand (gm_n2316, gm_n180, in_12, in_8, gm_n511, gm_n200);
	nor (gm_n2317, gm_n139, gm_n72, gm_n68, gm_n2316, gm_n602);
	nand (gm_n2318, gm_n83, in_28, in_24, gm_n2317, gm_n462);
	nor (gm_n2319, gm_n2318, gm_n206);
	nor (gm_n2320, gm_n2319, gm_n2315, gm_n2312);
	and (gm_n2321, gm_n189, in_16, gm_n157, gm_n1237, gm_n232);
	nand (gm_n2322, gm_n83, in_24, gm_n72, gm_n2321, gm_n269);
	nor (gm_n2323, gm_n475, gm_n780, in_28, gm_n2322);
	nor (gm_n2324, gm_n179, in_16, in_12, gm_n1025, gm_n222);
	nand (gm_n2325, gm_n237, in_24, gm_n72, gm_n2324, gm_n220);
	nor (gm_n2326, gm_n687, gm_n208, in_28, gm_n2325);
	and (gm_n2327, gm_n231, gm_n68, in_12, gm_n1647, gm_n341);
	nand (gm_n2328, gm_n183, in_24, gm_n72, gm_n2327, gm_n517);
	nor (gm_n2329, gm_n687, gm_n216, gm_n78, gm_n2328);
	nor (gm_n2330, gm_n2329, gm_n2326, gm_n2323);
	nand (gm_n2331, gm_n2309, gm_n2232, gm_n2226, gm_n2330, gm_n2320);
	nor (gm_n2332, gm_n593, gm_n385);
	nand (gm_n2333, gm_n621, in_15, in_11, gm_n2332, gm_n665);
	nor (gm_n2334, gm_n363, gm_n195, in_19, gm_n2333, gm_n510);
	nand (gm_n2335, gm_n55, gm_n50, gm_n133, gm_n2334, gm_n339);
	and (gm_n2336, gm_n567, gm_n262, gm_n64);
	nand (gm_n2337, gm_n189, in_16, in_12, gm_n2336, gm_n147);
	nor (gm_n2338, gm_n178, in_24, gm_n72, gm_n2337, gm_n804);
	nand (gm_n2339, gm_n462, gm_n186, gm_n78, gm_n2338);
	nand (gm_n2340, gm_n189, gm_n68, gm_n157, gm_n789, gm_n341);
	nor (gm_n2341, gm_n101, in_24, gm_n72, gm_n2340, gm_n156);
	nand (gm_n2342, gm_n370, gm_n97, gm_n78, gm_n2341);
	nand (gm_n2343, gm_n2342, gm_n2339, gm_n2335);
	nor (gm_n2344, gm_n150, gm_n53, in_21, gm_n2015, gm_n527);
	nand (gm_n2345, gm_n50, gm_n96, gm_n76, gm_n2344, gm_n776);
	nand (gm_n2346, gm_n146, in_16, gm_n157, gm_n1178, gm_n232);
	nor (gm_n2347, gm_n103, in_24, gm_n72, gm_n2346, gm_n412);
	nand (gm_n2348, gm_n492, gm_n99, in_28, gm_n2347);
	nand (gm_n2349, gm_n198, in_16, gm_n157, gm_n711, gm_n346);
	nor (gm_n2350, gm_n178, in_24, in_20, gm_n2349, gm_n804);
	nand (gm_n2351, gm_n134, gm_n77, gm_n78, gm_n2350);
	nand (gm_n2352, gm_n2351, gm_n2348, gm_n2345);
	nor (gm_n2353, gm_n2331, gm_n2222, gm_n2219, gm_n2352, gm_n2343);
	nand (gm_n2354, gm_n210, in_12, in_8, gm_n587, gm_n232);
	nor (gm_n2355, gm_n244, in_20, in_16, gm_n2354, gm_n103);
	nand (gm_n2356, gm_n207, in_28, in_24, gm_n2355, gm_n220);
	nor (gm_n2357, gm_n2356, gm_n206);
	nand (gm_n2358, gm_n137, gm_n52, gm_n72, gm_n2145, gm_n252);
	nor (gm_n2359, gm_n206, gm_n80, gm_n78, gm_n2358);
	and (gm_n2360, gm_n118, gm_n105, in_11, gm_n1543, gm_n665);
	nand (gm_n2361, gm_n299, in_23, gm_n102, gm_n2360, gm_n361);
	nor (gm_n2362, gm_n1118, gm_n50, in_27, gm_n2361, gm_n611);
	nor (gm_n2363, gm_n2362, gm_n2359, gm_n2357);
	and (gm_n2364, gm_n237, in_20, gm_n68, gm_n1315, gm_n189);
	nand (gm_n2365, gm_n83, gm_n78, gm_n52, gm_n2364, gm_n462);
	nor (gm_n2366, gm_n2365, gm_n206);
	nor (gm_n2367, gm_n106, in_16, gm_n157, gm_n2039, gm_n159);
	nand (gm_n2368, gm_n83, gm_n52, in_20, gm_n2367, gm_n219);
	nor (gm_n2369, gm_n687, gm_n243, in_28, gm_n2368);
	nand (gm_n2370, in_6, in_5, in_4, gm_n317, in_7);
	nor (gm_n2371, gm_n622, gm_n105, gm_n58, gm_n2370, gm_n666);
	nand (gm_n2372, gm_n73, in_23, gm_n102, gm_n2371, gm_n299);
	nor (gm_n2373, gm_n51, in_31, in_27, gm_n2372, gm_n617);
	nor (gm_n2374, gm_n2373, gm_n2369, gm_n2366);
	nand (gm_n2375, gm_n2353, gm_n2215, gm_n2211, gm_n2374, gm_n2363);
	nor (gm_n2376, gm_n222, gm_n157, gm_n64, gm_n593, gm_n942);
	nand (gm_n2377, gm_n237, in_20, in_16, gm_n2376, gm_n146);
	nor (gm_n2378, gm_n208, in_28, gm_n52, gm_n2377, gm_n628);
	nand (gm_n2379, gm_n2378, gm_n474);
	or (gm_n2380, gm_n57, in_15, in_11, gm_n1275, gm_n319);
	nor (gm_n2381, gm_n70, gm_n195, gm_n102, gm_n2380, gm_n337);
	nand (gm_n2382, gm_n173, in_31, in_27, gm_n2381, gm_n508);
	nand (gm_n2383, gm_n2029, in_15, in_11, gm_n665, gm_n621);
	nor (gm_n2384, gm_n423, gm_n195, in_19, gm_n2383, gm_n300);
	nand (gm_n2385, gm_n173, gm_n50, gm_n133, gm_n2384, gm_n339);
	nand (gm_n2386, gm_n2385, gm_n2382, gm_n2379);
	nand (gm_n2387, gm_n137, in_24, gm_n72, gm_n1576, gm_n220);
	nor (gm_n2388, gm_n371, gm_n176, in_28, gm_n2387);
	nor (out_9, gm_n2386, gm_n2375, gm_n2208, gm_n2388);
	nand (gm_n2390, gm_n449, gm_n309, gm_n122);
	nor (gm_n2391, gm_n300, gm_n105, in_11, gm_n2390, gm_n576);
	nand (gm_n2392, gm_n126, in_23, in_19, gm_n2391, gm_n658);
	nor (gm_n2393, gm_n678, gm_n50, gm_n133, gm_n2392);
	or (gm_n2394, gm_n139, gm_n157, in_8, gm_n386, gm_n286);
	nor (gm_n2395, gm_n412, gm_n72, gm_n68, gm_n2394, gm_n602);
	nand (gm_n2396, gm_n77, in_28, gm_n52, gm_n2395, gm_n207);
	nand (gm_n2397, gm_n308, gm_n354, gm_n64, gm_n619);
	or (gm_n2398, gm_n117, in_19, in_15, gm_n2397, gm_n366);
	nor (gm_n2399, gm_n431, gm_n133, in_23, gm_n2398, gm_n983);
	nand (gm_n2400, gm_n2399, gm_n304, in_31);
	and (gm_n2401, gm_n138, gm_n72, in_16, gm_n1094, gm_n219);
	nand (gm_n2402, gm_n183, in_28, in_24, gm_n2401, gm_n462);
	nor (gm_n2403, gm_n2402, gm_n268);
	and (gm_n2404, gm_n180, gm_n68, gm_n157, gm_n885, gm_n198);
	nand (gm_n2405, gm_n137, gm_n52, gm_n72, gm_n2404, gm_n183);
	nor (gm_n2406, gm_n260, gm_n218, in_28, gm_n2405);
	or (gm_n2407, gm_n168, in_16, gm_n157, gm_n445, gm_n286);
	nor (gm_n2408, gm_n178, in_24, in_20, gm_n2407, gm_n412);
	nand (gm_n2409, gm_n194, gm_n79, in_28, gm_n2408);
	nor (gm_n2410, in_7, gm_n121, gm_n62, gm_n465, gm_n64);
	nand (gm_n2411, gm_n188, in_16, in_12, gm_n2410, gm_n189);
	nor (gm_n2412, gm_n516, gm_n52, gm_n72, gm_n2411, gm_n413);
	nand (gm_n2413, gm_n492, gm_n462, in_28, gm_n2412);
	nor (gm_n2414, gm_n159, gm_n68, in_12, gm_n916, gm_n179);
	nand (gm_n2415, gm_n237, in_24, gm_n72, gm_n2414, gm_n261);
	nor (gm_n2416, gm_n687, gm_n243, in_28, gm_n2415);
	or (gm_n2417, gm_n70, in_23, gm_n102, gm_n656, gm_n423);
	nor (gm_n2418, gm_n174, gm_n50, gm_n133, gm_n2417, gm_n842);
	or (gm_n2419, gm_n672, gm_n105, in_11, gm_n1485, gm_n396);
	nor (gm_n2420, gm_n510, gm_n195, gm_n102, gm_n2419, gm_n911);
	nand (gm_n2421, gm_n173, in_31, in_27, gm_n2420, gm_n508);
	nand (gm_n2422, gm_n629, in_16, in_12, gm_n1895, gm_n232);
	nor (gm_n2423, gm_n197, in_24, gm_n72, gm_n2422, gm_n459);
	nand (gm_n2424, gm_n259, gm_n194, in_28, gm_n2423);
	and (gm_n2425, gm_n341, gm_n69, gm_n105, gm_n512, gm_n818);
	nand (gm_n2426, gm_n509, gm_n195, gm_n102, gm_n2425, gm_n658);
	nor (gm_n2427, gm_n436, in_31, in_27, gm_n2426);
	nor (gm_n2428, gm_n319, in_15, in_11, gm_n1329, gm_n366);
	nand (gm_n2429, gm_n69, in_23, in_19, gm_n2428, gm_n361);
	nor (gm_n2430, gm_n436, in_31, in_27, gm_n2429, gm_n671);
	nand (gm_n2431, gm_n747, gm_n110, in_8);
	nor (gm_n2432, gm_n139, in_16, gm_n157, gm_n2431, gm_n167);
	nand (gm_n2433, gm_n100, gm_n52, in_20, gm_n2432, gm_n219);
	nor (gm_n2434, gm_n218, gm_n208, gm_n78, gm_n2433);
	nor (gm_n2435, gm_n106, gm_n68, gm_n157, gm_n2178, gm_n286);
	nand (gm_n2436, gm_n183, gm_n52, gm_n72, gm_n2435, gm_n230);
	nor (gm_n2437, gm_n475, gm_n216, in_28, gm_n2436);
	nor (gm_n2438, gm_n576, in_15, in_11, gm_n701, gm_n618);
	nand (gm_n2439, gm_n73, in_23, gm_n102, gm_n2438, gm_n394);
	nor (gm_n2440, gm_n54, gm_n50, in_27, gm_n2439, gm_n360);
	nor (gm_n2441, gm_n2434, gm_n2430, gm_n2427, gm_n2440, gm_n2437);
	or (gm_n2442, gm_n223, gm_n727, in_11, gm_n593, gm_n366);
	nor (gm_n2443, gm_n127, in_19, in_15, gm_n2442, gm_n395);
	nand (gm_n2444, gm_n339, gm_n133, gm_n195, gm_n2443, gm_n658);
	nor (gm_n2445, gm_n2444, in_31);
	nor (gm_n2446, gm_n673, gm_n105, gm_n58, gm_n2081, gm_n622);
	nand (gm_n2447, gm_n313, gm_n195, gm_n102, gm_n2446, gm_n612);
	nor (gm_n2448, gm_n983, gm_n50, gm_n133, gm_n2447, gm_n678);
	and (gm_n2449, gm_n146, in_16, gm_n157, gm_n2018, gm_n270);
	nand (gm_n2450, gm_n219, in_24, in_20, gm_n2449, gm_n252);
	nor (gm_n2451, gm_n135, gm_n132, in_28, gm_n2450);
	nor (gm_n2452, gm_n2451, gm_n2448, gm_n2445);
	nor (gm_n2453, gm_n116, gm_n68, gm_n105, gm_n2227, gm_n136);
	nor (gm_n2454, gm_n81, gm_n72, in_19);
	nor (gm_n2455, in_25, gm_n52, gm_n195);
	nand (gm_n2456, gm_n2453, in_26, gm_n82, gm_n2455, gm_n2454);
	nor (gm_n2457, in_29, in_28, in_27);
	not (gm_n2458, gm_n2457);
	nor (gm_n2459, gm_n2456, gm_n50, in_30, gm_n2458);
	nor (gm_n2460, gm_n159, gm_n68, gm_n157, gm_n1050, gm_n168);
	nand (gm_n2461, gm_n220, in_24, gm_n72, gm_n2460, gm_n230);
	nor (gm_n2462, gm_n243, gm_n132, gm_n78, gm_n2461);
	nand (gm_n2463, gm_n124, gm_n110);
	nor (gm_n2464, gm_n432, in_15, gm_n58, gm_n2463, gm_n366);
	nand (gm_n2465, gm_n582, in_23, in_19, gm_n2464, gm_n313);
	nor (gm_n2466, gm_n575, in_31, in_27, gm_n2465, gm_n581);
	nor (gm_n2467, gm_n2466, gm_n2462, gm_n2459);
	nand (gm_n2468, gm_n2441, gm_n2424, gm_n2421, gm_n2467, gm_n2452);
	nor (gm_n2469, gm_n107, gm_n157, gm_n64, gm_n385, gm_n254);
	nand (gm_n2470, gm_n86, gm_n72, in_16, gm_n2469, gm_n230);
	nor (gm_n2471, gm_n101, gm_n78, gm_n52, gm_n2470, gm_n780);
	nand (gm_n2472, gm_n2471, gm_n194);
	nand (gm_n2473, gm_n629, gm_n68, gm_n157, gm_n1411, gm_n341);
	nor (gm_n2474, gm_n561, gm_n52, in_20, gm_n2473, gm_n742);
	nand (gm_n2475, gm_n134, gm_n97, in_28, gm_n2474);
	nor (gm_n2476, gm_n56, gm_n157, in_11);
	nor (gm_n2477, gm_n116, in_16, gm_n105);
	nand (gm_n2478, gm_n480, in_18, in_14, gm_n2477, gm_n2476);
	nor (gm_n2479, gm_n486, in_26, gm_n82, gm_n2478, gm_n638);
	nand (gm_n2480, gm_n1905, in_31, gm_n96, gm_n2479);
	nand (gm_n2481, gm_n2480, gm_n2475, gm_n2472);
	nand (gm_n2482, gm_n198, gm_n68, in_12, gm_n872, gm_n341);
	nor (gm_n2483, gm_n516, gm_n52, gm_n72, gm_n2482, gm_n413);
	nand (gm_n2484, gm_n207, gm_n77, in_28, gm_n2483);
	nand (gm_n2485, gm_n219, gm_n72, gm_n68, gm_n2376, gm_n629);
	nor (gm_n2486, gm_n216, in_28, gm_n52, gm_n2485, gm_n561);
	nand (gm_n2487, gm_n2486, gm_n77);
	nand (gm_n2488, gm_n86, gm_n68, gm_n157, gm_n872, gm_n354);
	nor (gm_n2489, gm_n561, gm_n52, gm_n72, gm_n2488, gm_n459);
	nand (gm_n2490, gm_n134, gm_n97, gm_n78, gm_n2489);
	nand (gm_n2491, gm_n2490, gm_n2487, gm_n2484);
	nor (gm_n2492, gm_n2468, gm_n2418, gm_n2416, gm_n2491, gm_n2481);
	nor (gm_n2493, gm_n88, in_16, gm_n157, gm_n2166, gm_n221);
	nand (gm_n2494, gm_n230, gm_n52, gm_n72, gm_n2493, gm_n261);
	nor (gm_n2495, gm_n475, gm_n216, gm_n78, gm_n2494);
	and (gm_n2496, gm_n198, in_16, gm_n157, gm_n1411, gm_n346);
	nand (gm_n2497, gm_n85, gm_n52, in_20, gm_n2496, gm_n261);
	nor (gm_n2498, gm_n371, gm_n206, gm_n78, gm_n2497);
	nand (gm_n2499, gm_n747, gm_n308, in_8);
	nor (gm_n2500, gm_n159, in_16, in_12, gm_n2499, gm_n168);
	nand (gm_n2501, gm_n137, gm_n52, in_20, gm_n2500, gm_n196);
	nor (gm_n2502, gm_n687, gm_n135, gm_n78, gm_n2501);
	nor (gm_n2503, gm_n2502, gm_n2498, gm_n2495);
	nand (gm_n2504, gm_n141, in_4, gm_n60, gm_n308);
	nor (gm_n2505, gm_n672, in_15, gm_n58, gm_n2504, gm_n319);
	nand (gm_n2506, gm_n69, gm_n195, gm_n102, gm_n2505, gm_n126);
	nor (gm_n2507, gm_n303, gm_n50, gm_n133, gm_n2506, gm_n617);
	nor (gm_n2508, gm_n159, gm_n68, in_12, gm_n2195, gm_n168);
	nand (gm_n2509, gm_n137, gm_n52, gm_n72, gm_n2508, gm_n196);
	nor (gm_n2510, gm_n268, gm_n80, in_28, gm_n2509);
	nor (gm_n2511, gm_n161, gm_n68, in_12, gm_n253, gm_n221);
	nand (gm_n2512, gm_n137, in_24, gm_n72, gm_n2511, gm_n196);
	nor (gm_n2513, gm_n687, gm_n243, in_28, gm_n2512);
	nor (gm_n2514, gm_n2513, gm_n2510, gm_n2507);
	nand (gm_n2515, gm_n2492, gm_n2413, gm_n2409, gm_n2514, gm_n2503);
	nand (gm_n2516, gm_n629, in_16, gm_n157, gm_n348, gm_n346);
	nor (gm_n2517, gm_n178, in_24, in_20, gm_n2516, gm_n197);
	nand (gm_n2518, gm_n205, gm_n177, in_28, gm_n2517);
	or (gm_n2519, gm_n88, in_15, in_8, gm_n1039, gm_n576);
	nor (gm_n2520, gm_n332, gm_n195, gm_n102, gm_n2519, gm_n337);
	nand (gm_n2521, gm_n55, gm_n50, gm_n133, gm_n2520, gm_n437);
	nor (gm_n2522, gm_n562, in_12, in_8, gm_n733, gm_n222);
	nand (gm_n2523, gm_n86, in_20, in_16, gm_n2522, gm_n517);
	nor (gm_n2524, gm_n561, in_28, gm_n52, gm_n2523, gm_n260);
	nand (gm_n2525, gm_n2524, gm_n492);
	nand (gm_n2526, gm_n2525, gm_n2521, gm_n2518);
	and (gm_n2527, in_7, gm_n121, in_5, gm_n364, gm_n64);
	nand (gm_n2528, gm_n86, gm_n68, gm_n157, gm_n2527, gm_n354);
	nor (gm_n2529, gm_n101, gm_n52, gm_n72, gm_n2528, gm_n459);
	nand (gm_n2530, gm_n462, gm_n205, gm_n78, gm_n2529);
	nand (gm_n2531, gm_n189, gm_n72, gm_n68, gm_n1307, gm_n269);
	nor (gm_n2532, gm_n84, gm_n78, in_24, gm_n2531, gm_n135);
	nand (gm_n2533, gm_n2532, gm_n217);
	nand (gm_n2534, gm_n64, in_4, gm_n60, gm_n141, gm_n122);
	or (gm_n2535, gm_n106, gm_n68, in_12, gm_n2534, gm_n159);
	nor (gm_n2536, gm_n156, gm_n52, in_20, gm_n2535, gm_n804);
	nand (gm_n2537, gm_n99, gm_n97, gm_n78, gm_n2536);
	nand (gm_n2538, gm_n2537, gm_n2533, gm_n2530);
	nor (gm_n2539, gm_n2515, gm_n2406, gm_n2403, gm_n2538, gm_n2526);
	and (gm_n2540, gm_n237, gm_n72, gm_n68, gm_n2140, gm_n766);
	nand (gm_n2541, gm_n209, in_28, in_24, gm_n2540, gm_n462);
	nor (gm_n2542, gm_n2541, gm_n176);
	nor (gm_n2543, gm_n727, gm_n105, gm_n58, gm_n997, gm_n762);
	nand (gm_n2544, gm_n336, gm_n195, gm_n102, gm_n2543, gm_n362);
	nor (gm_n2545, gm_n51, in_31, gm_n133, gm_n2544, gm_n54);
	nor (gm_n2546, gm_n244, in_12, in_8, gm_n1356, gm_n107);
	nand (gm_n2547, gm_n252, gm_n72, in_16, gm_n2546, gm_n472);
	nor (gm_n2548, gm_n135, gm_n78, gm_n52, gm_n2547, gm_n268);
	nor (gm_n2549, gm_n2548, gm_n2545, gm_n2542);
	nor (gm_n2550, gm_n672, gm_n105, in_11, gm_n1086, gm_n396);
	nand (gm_n2551, gm_n165, gm_n195, gm_n102, gm_n2550, gm_n452);
	nor (gm_n2552, gm_n51, gm_n50, gm_n133, gm_n2551, gm_n174);
	and (gm_n2553, gm_n118, gm_n105, in_11, gm_n1770, gm_n937);
	nand (gm_n2554, gm_n336, gm_n195, in_19, gm_n2553, gm_n612);
	nor (gm_n2555, gm_n51, gm_n50, in_27, gm_n2554, gm_n54);
	nand (gm_n2556, gm_n567, gm_n308, gm_n64);
	nor (gm_n2557, gm_n106, in_16, in_12, gm_n2556, gm_n253);
	nand (gm_n2558, gm_n85, in_24, in_20, gm_n2557, gm_n261);
	nor (gm_n2559, gm_n243, gm_n132, gm_n78, gm_n2558);
	nor (gm_n2560, gm_n2559, gm_n2555, gm_n2552);
	nand (gm_n2561, gm_n2539, gm_n2400, gm_n2396, gm_n2560, gm_n2549);
	nand (gm_n2562, gm_n118, gm_n188, gm_n105, gm_n613, gm_n394);
	nor (gm_n2563, gm_n671, in_23, in_19, gm_n2562, gm_n510);
	nand (gm_n2564, gm_n437, in_31, in_27, gm_n2563);
	or (gm_n2565, gm_n286, in_15, gm_n64, gm_n1533, gm_n366);
	nor (gm_n2566, gm_n423, in_23, in_19, gm_n2565, gm_n300);
	nand (gm_n2567, gm_n173, in_31, gm_n133, gm_n2566, gm_n306);
	or (gm_n2568, gm_n942, gm_n169, gm_n64);
	or (gm_n2569, gm_n158, in_16, in_12, gm_n2568, gm_n286);
	nor (gm_n2570, gm_n628, in_24, gm_n72, gm_n2569, gm_n742);
	nand (gm_n2571, gm_n217, gm_n99, gm_n78, gm_n2570);
	nand (gm_n2572, gm_n2571, gm_n2567, gm_n2564);
	and (gm_n2573, gm_n118, gm_n105, in_11, gm_n1551, gm_n612);
	nand (gm_n2574, gm_n165, gm_n195, gm_n102, gm_n2573, gm_n455);
	nor (gm_n2575, gm_n360, in_31, in_27, gm_n2574);
	nor (out_10, gm_n2572, gm_n2561, gm_n2393, gm_n2575);
	and (gm_n2577, gm_n147, in_16, gm_n157, gm_n1816, gm_n629);
	nand (gm_n2578, gm_n137, in_24, gm_n72, gm_n2577, gm_n261);
	nor (gm_n2579, gm_n371, gm_n206, gm_n78, gm_n2578);
	nor (gm_n2580, gm_n385, gm_n355, gm_n64);
	nand (gm_n2581, gm_n188, gm_n68, gm_n157, gm_n2580, gm_n629);
	nor (gm_n2582, gm_n178, gm_n52, in_20, gm_n2581, gm_n516);
	nand (gm_n2583, gm_n259, gm_n194, gm_n78, gm_n2582);
	nand (gm_n2584, gm_n311, gm_n354, gm_n105, gm_n645, gm_n362);
	nor (gm_n2585, gm_n127, gm_n195, in_19, gm_n2584, gm_n581);
	nand (gm_n2586, gm_n508, gm_n50, in_27, gm_n2585);
	nor (gm_n2587, gm_n139, gm_n68, in_12, gm_n1693, gm_n286);
	nand (gm_n2588, gm_n83, gm_n52, gm_n72, gm_n2587, gm_n85);
	nor (gm_n2589, gm_n218, gm_n135, in_28, gm_n2588);
	nand (gm_n2590, gm_n297, gm_n263, gm_n122);
	nor (gm_n2591, gm_n366, in_15, in_11, gm_n2590, gm_n453);
	nand (gm_n2592, gm_n293, gm_n195, in_19, gm_n2591, gm_n658);
	nor (gm_n2593, gm_n303, in_31, in_27, gm_n2592);
	nor (gm_n2594, gm_n223, gm_n1801);
	nand (gm_n2595, gm_n818, gm_n105, gm_n58, gm_n2594, gm_n425);
	nor (gm_n2596, gm_n294, in_23, in_19, gm_n2595, gm_n453);
	nand (gm_n2597, gm_n455, in_31, in_27, gm_n2596, gm_n508);
	nor (gm_n2598, gm_n222, gm_n157, gm_n64, gm_n385, gm_n224);
	and (gm_n2599, gm_n1183, gm_n116, gm_n56, gm_n2598, gm_n1565);
	and (gm_n2600, gm_n327, gm_n53, gm_n81, gm_n2599, gm_n775);
	nand (gm_n2601, in_31, gm_n96, in_29, gm_n2600);
	or (gm_n2602, gm_n479, gm_n109);
	nor (gm_n2603, gm_n119, gm_n105, gm_n58, gm_n2602, gm_n399);
	nand (gm_n2604, gm_n336, in_23, in_19, gm_n2603, gm_n394);
	nor (gm_n2605, gm_n360, in_31, gm_n133, gm_n2604, gm_n617);
	and (gm_n2606, gm_n270, in_16, in_12, gm_n2336, gm_n766);
	nand (gm_n2607, gm_n100, in_24, gm_n72, gm_n2606, gm_n237);
	nor (gm_n2608, gm_n208, gm_n206, gm_n78, gm_n2607);
	or (gm_n2609, gm_n221, gm_n68, gm_n157, gm_n688, gm_n286);
	nor (gm_n2610, gm_n84, in_24, in_20, gm_n2609, gm_n156);
	nand (gm_n2611, gm_n462, gm_n205, gm_n78, gm_n2610);
	nor (gm_n2612, gm_n295, gm_n562, in_8);
	nand (gm_n2613, gm_n188, in_16, gm_n157, gm_n2612, gm_n138);
	nor (gm_n2614, gm_n101, in_24, in_20, gm_n2613, gm_n178);
	nand (gm_n2615, gm_n134, gm_n77, in_28, gm_n2614);
	nor (gm_n2616, gm_n57, gm_n105, in_11, gm_n674, gm_n727);
	nand (gm_n2617, gm_n165, gm_n195, gm_n102, gm_n2616, gm_n394);
	nor (gm_n2618, gm_n174, gm_n50, gm_n133, gm_n2617, gm_n436);
	nand (gm_n2619, gm_n361, in_23, gm_n102, gm_n1284, gm_n362);
	nor (gm_n2620, gm_n617, gm_n50, gm_n133, gm_n2619, gm_n436);
	nor (gm_n2621, gm_n244, gm_n68, in_12, gm_n2195, gm_n167);
	nand (gm_n2622, gm_n183, gm_n52, gm_n72, gm_n2621, gm_n472);
	nor (gm_n2623, gm_n475, gm_n80, gm_n78, gm_n2622);
	nor (gm_n2624, gm_n366, gm_n105, in_11, gm_n1279, gm_n666);
	nand (gm_n2625, gm_n126, gm_n195, gm_n102, gm_n2624, gm_n362);
	nor (gm_n2626, gm_n174, in_31, gm_n133, gm_n2625, gm_n611);
	nand (gm_n2627, gm_n346, in_12, in_8, gm_n1226, gm_n262);
	nor (gm_n2628, gm_n504, in_20, gm_n68, gm_n2627, gm_n459);
	nand (gm_n2629, gm_n134, gm_n78, gm_n52, gm_n2628, gm_n183);
	nor (gm_n2630, gm_n2629, gm_n206);
	nor (gm_n2631, gm_n2623, gm_n2620, gm_n2618, gm_n2630, gm_n2626);
	nor (gm_n2632, gm_n168, gm_n68, in_12, gm_n1270, gm_n286);
	nand (gm_n2633, gm_n230, gm_n52, gm_n72, gm_n2632, gm_n261);
	nor (gm_n2634, gm_n268, gm_n135, in_28, gm_n2633);
	nor (gm_n2635, gm_n88, in_12, in_8, gm_n1806, gm_n139);
	nand (gm_n2636, gm_n252, in_20, in_16, gm_n2635, gm_n269);
	nor (gm_n2637, gm_n206, gm_n78, in_24, gm_n2636, gm_n780);
	nand (gm_n2638, gm_n210, in_12, in_8, gm_n587, gm_n346);
	nor (gm_n2639, gm_n221, gm_n72, gm_n68, gm_n2638, gm_n602);
	nand (gm_n2640, gm_n83, gm_n78, in_24, gm_n2639, gm_n99);
	nor (gm_n2641, gm_n2640, gm_n176);
	nor (gm_n2642, gm_n2641, gm_n2637, gm_n2634);
	nand (gm_n2643, gm_n511, gm_n200, gm_n64);
	nor (gm_n2644, gm_n244, in_16, in_12, gm_n2643, gm_n88);
	nand (gm_n2645, gm_n100, in_24, in_20, gm_n2644, gm_n230);
	nor (gm_n2646, gm_n208, gm_n229, gm_n78, gm_n2645);
	nor (gm_n2647, gm_n159, gm_n68, gm_n157, gm_n1303, gm_n168);
	nand (gm_n2648, gm_n183, gm_n52, in_20, gm_n2647, gm_n230);
	nor (gm_n2649, gm_n268, gm_n135, gm_n78, gm_n2648);
	nand (gm_n2650, gm_n180, gm_n157, in_8, gm_n122, gm_n108);
	nor (gm_n2651, gm_n178, in_20, in_16, gm_n2650, gm_n221);
	nand (gm_n2652, gm_n99, in_28, in_24, gm_n2651, gm_n100);
	nor (gm_n2653, gm_n2652, gm_n268);
	nor (gm_n2654, gm_n2653, gm_n2649, gm_n2646);
	nand (gm_n2655, gm_n2631, gm_n2615, gm_n2611, gm_n2654, gm_n2642);
	nand (gm_n2656, gm_n86, in_16, in_12, gm_n356, gm_n341);
	nor (gm_n2657, gm_n178, in_24, gm_n72, gm_n2656, gm_n804);
	nand (gm_n2658, gm_n217, gm_n207, gm_n78, gm_n2657);
	nor (gm_n2659, gm_n107, gm_n157, in_8, gm_n942, gm_n160);
	nand (gm_n2660, gm_n189, gm_n72, gm_n68, gm_n2659, gm_n517);
	nor (gm_n2661, gm_n243, in_28, gm_n52, gm_n2660, gm_n412);
	nand (gm_n2662, gm_n2661, gm_n97);
	nand (gm_n2663, gm_n86, in_16, gm_n157, gm_n2000, gm_n354);
	nor (gm_n2664, gm_n187, in_24, in_20, gm_n2663, gm_n804);
	nand (gm_n2665, gm_n370, gm_n97, gm_n78, gm_n2664);
	nand (gm_n2666, gm_n2665, gm_n2662, gm_n2658);
	nor (gm_n2667, gm_n355, gm_n89);
	nand (gm_n2668, gm_n66, in_15, in_11, gm_n2667, gm_n938);
	nor (gm_n2669, gm_n431, in_23, gm_n102, gm_n2668, gm_n453);
	nand (gm_n2670, gm_n304, in_31, gm_n133, gm_n2669, gm_n455);
	or (gm_n2671, gm_n319, gm_n105, gm_n58, gm_n2233, gm_n366);
	nor (gm_n2672, gm_n127, gm_n195, in_19, gm_n2671, gm_n300);
	nand (gm_n2673, gm_n302, in_31, gm_n133, gm_n2672, gm_n339);
	nand (gm_n2674, gm_n188, gm_n68, gm_n157, gm_n1060, gm_n231);
	nor (gm_n2675, gm_n412, in_24, in_20, gm_n2674, gm_n742);
	nand (gm_n2676, gm_n259, gm_n194, in_28, gm_n2675);
	nand (gm_n2677, gm_n2676, gm_n2673, gm_n2670);
	nor (gm_n2678, gm_n2655, gm_n2608, gm_n2605, gm_n2677, gm_n2666);
	nor (gm_n2679, gm_n168, gm_n68, gm_n157, gm_n1025, gm_n253);
	nand (gm_n2680, gm_n196, in_24, in_20, gm_n2679, gm_n269);
	nor (gm_n2681, gm_n206, gm_n243, in_28, gm_n2680);
	nand (gm_n2682, gm_n109, gm_n121, in_5, gm_n364, gm_n64);
	nor (gm_n2683, gm_n88, in_16, in_12, gm_n2682, gm_n139);
	nand (gm_n2684, gm_n83, in_24, gm_n72, gm_n2683, gm_n237);
	nor (gm_n2685, gm_n780, gm_n176, gm_n78, gm_n2684);
	nor (gm_n2686, gm_n88, in_16, gm_n157, gm_n960, gm_n504);
	nand (gm_n2687, gm_n100, gm_n52, in_20, gm_n2686, gm_n472);
	nor (gm_n2688, gm_n475, gm_n135, gm_n78, gm_n2687);
	nor (gm_n2689, gm_n2688, gm_n2685, gm_n2681);
	nor (gm_n2690, gm_n282, in_15, in_11, gm_n426, gm_n673);
	nand (gm_n2691, gm_n69, in_23, gm_n102, gm_n2690, gm_n165);
	nor (gm_n2692, gm_n360, gm_n50, in_27, gm_n2691, gm_n617);
	or (gm_n2693, gm_n544, gm_n89);
	nor (gm_n2694, gm_n432, gm_n105, gm_n58, gm_n2693, gm_n426);
	nand (gm_n2695, gm_n126, in_23, in_19, gm_n2694, gm_n452);
	nor (gm_n2696, gm_n174, in_31, in_27, gm_n2695, gm_n303);
	or (gm_n2697, gm_n942, gm_n224);
	nor (gm_n2698, gm_n319, in_15, in_11, gm_n2697, gm_n366);
	nand (gm_n2699, gm_n126, gm_n195, in_19, gm_n2698, gm_n452);
	nor (gm_n2700, gm_n1231, gm_n50, in_27, gm_n2699, gm_n436);
	nor (gm_n2701, gm_n2700, gm_n2696, gm_n2692);
	nand (gm_n2702, gm_n2678, gm_n2601, gm_n2597, gm_n2701, gm_n2689);
	nor (gm_n2703, gm_n385, gm_n91);
	nand (gm_n2704, gm_n311, in_15, in_11, gm_n2703, gm_n449);
	nor (gm_n2705, gm_n395, gm_n195, in_19, gm_n2704, gm_n510);
	nand (gm_n2706, gm_n115, in_31, in_27, gm_n2705, gm_n302);
	nor (gm_n2707, gm_n91, gm_n157, in_8, gm_n942, gm_n253);
	nand (gm_n2708, gm_n189, gm_n72, in_16, gm_n2707, gm_n230);
	nor (gm_n2709, gm_n243, in_28, in_24, gm_n2708, gm_n628);
	nand (gm_n2710, gm_n2709, gm_n474);
	or (gm_n2711, gm_n672, gm_n102, gm_n105, gm_n1631, gm_n332);
	nor (gm_n2712, gm_n127, in_27, gm_n195, gm_n2711, gm_n174);
	nand (gm_n2713, gm_n2712, gm_n677, gm_n50);
	nand (gm_n2714, gm_n2713, gm_n2710, gm_n2706);
	nor (gm_n2715, gm_n942, in_12, in_8, gm_n544, gm_n286);
	nand (gm_n2716, gm_n137, gm_n72, gm_n68, gm_n2715, gm_n231);
	nor (gm_n2717, gm_n197, gm_n78, in_24, gm_n2716, gm_n780);
	nand (gm_n2718, gm_n2717, gm_n97);
	nand (gm_n2719, gm_n394, gm_n188, in_15, gm_n889, gm_n621);
	nor (gm_n2720, gm_n1118, in_23, in_19, gm_n2719, gm_n337);
	nand (gm_n2721, gm_n115, in_31, gm_n133, gm_n2720);
	nand (gm_n2722, gm_n231, gm_n68, in_12, gm_n613, gm_n232);
	nor (gm_n2723, gm_n103, gm_n52, in_20, gm_n2722, gm_n412);
	nand (gm_n2724, gm_n474, gm_n370, gm_n78, gm_n2723);
	nand (gm_n2725, gm_n2724, gm_n2721, gm_n2718);
	nor (gm_n2726, gm_n2702, gm_n2593, gm_n2589, gm_n2725, gm_n2714);
	or (gm_n2727, gm_n245, in_12, in_8, gm_n544, gm_n942);
	nor (gm_n2728, gm_n504, gm_n72, gm_n68, gm_n2727, gm_n156);
	nand (gm_n2729, gm_n177, in_28, gm_n52, gm_n2728, gm_n183);
	nor (gm_n2730, gm_n2729, gm_n176);
	and (gm_n2731, gm_n189, gm_n68, in_12, gm_n1106, gm_n270);
	nand (gm_n2732, gm_n100, gm_n52, in_20, gm_n2731, gm_n230);
	nor (gm_n2733, gm_n216, gm_n229, in_28, gm_n2732);
	and (gm_n2734, gm_n86, in_16, in_12, gm_n758, gm_n232);
	nand (gm_n2735, gm_n220, gm_n52, gm_n72, gm_n2734, gm_n472);
	nor (gm_n2736, gm_n218, gm_n208, in_28, gm_n2735);
	nor (gm_n2737, gm_n2736, gm_n2733, gm_n2730);
	nor (gm_n2738, in_16, in_15, gm_n104);
	and (gm_n2739, gm_n406, in_17, gm_n56, gm_n2738, gm_n2205);
	nand (gm_n2740, gm_n775, gm_n53, in_21, gm_n2739, gm_n1055);
	nor (gm_n2741, in_31, in_30, gm_n76, gm_n2740);
	nand (gm_n2742, gm_n321, gm_n116, in_13, gm_n2013, gm_n1563);
	or (gm_n2743, gm_n152, gm_n53, in_21, gm_n2742, gm_n323);
	nor (gm_n2744, in_31, gm_n96, gm_n76, gm_n2743, gm_n328);
	nor (gm_n2745, gm_n119, in_15, gm_n58, gm_n1259, gm_n426);
	nand (gm_n2746, gm_n126, gm_n195, in_19, gm_n2745, gm_n452);
	nor (gm_n2747, gm_n54, in_31, gm_n133, gm_n2746, gm_n303);
	nor (gm_n2748, gm_n2747, gm_n2744, gm_n2741);
	nand (gm_n2749, gm_n2726, gm_n2586, gm_n2583, gm_n2748, gm_n2737);
	nand (gm_n2750, gm_n120, in_15, in_11, gm_n1770, gm_n818);
	nor (gm_n2751, gm_n423, gm_n195, gm_n102, gm_n2750, gm_n453);
	nand (gm_n2752, gm_n129, gm_n50, in_27, gm_n2751, gm_n392);
	or (gm_n2753, gm_n139, in_16, gm_n157, gm_n1241, gm_n222);
	nor (gm_n2754, gm_n84, in_24, in_20, gm_n2753, gm_n187);
	nand (gm_n2755, gm_n259, gm_n97, in_28, gm_n2754);
	or (gm_n2756, gm_n504, gm_n68, in_12, gm_n1639, gm_n286);
	nor (gm_n2757, gm_n178, in_24, gm_n72, gm_n2756, gm_n412);
	nand (gm_n2758, gm_n207, gm_n186, gm_n78, gm_n2757);
	nand (gm_n2759, gm_n2758, gm_n2755, gm_n2752);
	nor (gm_n2760, gm_n88, in_16, gm_n157, gm_n2178, gm_n504);
	nand (gm_n2761, gm_n83, in_24, in_20, gm_n2760, gm_n472);
	nor (gm_n2762, gm_n260, gm_n268, in_28, gm_n2761);
	nor (out_11, gm_n2759, gm_n2749, gm_n2579, gm_n2762);
	nor (gm_n2764, gm_n167, gm_n68, gm_n157, gm_n1064, gm_n158);
	and (gm_n2765, gm_n100, in_24, gm_n72, gm_n2764, gm_n219);
	and (gm_n2766, gm_n370, gm_n77, in_28, gm_n2765);
	nand (gm_n2767, gm_n629, in_16, gm_n157, gm_n1252, gm_n341);
	or (gm_n2768, gm_n628, in_24, gm_n72, gm_n2767, gm_n413);
	nor (gm_n2769, gm_n208, gm_n229, in_28, gm_n2768);
	and (gm_n2770, gm_n180, in_16, in_12, gm_n1021, gm_n146);
	and (gm_n2771, gm_n183, gm_n52, in_20, gm_n2770, gm_n472);
	and (gm_n2772, gm_n259, gm_n97, gm_n78, gm_n2771);
	nor (gm_n2773, gm_n244, gm_n72, gm_n68, gm_n2727, gm_n742);
	nand (gm_n2774, gm_n79, gm_n78, gm_n52, gm_n2773, gm_n83);
	nor (gm_n2775, gm_n2774, gm_n687);
	not (gm_n2776, gm_n319);
	and (gm_n2777, gm_n311, gm_n105, gm_n58, gm_n2703, gm_n2776);
	nand (gm_n2778, gm_n293, gm_n195, in_19, gm_n2777, gm_n612);
	nor (gm_n2779, gm_n54, gm_n50, gm_n133, gm_n2778, gm_n436);
	or (gm_n2780, gm_n366, in_15, in_11, gm_n2463, gm_n396);
	nor (gm_n2781, gm_n300, gm_n195, gm_n102, gm_n2780, gm_n337);
	nand (gm_n2782, gm_n173, gm_n50, gm_n133, gm_n2781, gm_n508);
	and (gm_n2783, gm_n120, in_15, in_11, gm_n2667, gm_n311);
	nand (gm_n2784, gm_n165, in_23, in_19, gm_n2783, gm_n452);
	or (gm_n2785, gm_n1118, in_31, in_27, gm_n2784, gm_n575);
	nor (gm_n2786, gm_n88, gm_n68, gm_n157, gm_n1639, gm_n504);
	nand (gm_n2787, gm_n100, in_24, gm_n72, gm_n2786, gm_n219);
	nor (gm_n2788, gm_n687, gm_n371, in_28, gm_n2787);
	nor (gm_n2789, gm_n727, in_15, in_11, gm_n1279, gm_n997);
	nand (gm_n2790, gm_n165, gm_n195, gm_n102, gm_n2789, gm_n362);
	nor (gm_n2791, gm_n611, in_31, in_27, gm_n2790, gm_n671);
	nor (gm_n2792, gm_n253, gm_n105, gm_n64, gm_n997, gm_n386);
	and (gm_n2793, gm_n73, in_23, in_19, gm_n2792, gm_n452);
	nand (gm_n2794, gm_n307, gm_n50, in_27, gm_n2793, gm_n677);
	nor (gm_n2795, gm_n167, gm_n68, in_12, gm_n1782, gm_n179);
	nand (gm_n2796, gm_n237, gm_n52, gm_n72, gm_n2795, gm_n196);
	or (gm_n2797, gm_n687, gm_n243, gm_n78, gm_n2796);
	and (gm_n2798, gm_n138, gm_n68, gm_n157, gm_n1147, gm_n354);
	nand (gm_n2799, gm_n137, in_24, gm_n72, gm_n2798, gm_n261);
	nor (gm_n2800, gm_n687, gm_n208, in_28, gm_n2799);
	nor (gm_n2801, gm_n151, gm_n81, in_17, gm_n1611, gm_n736);
	nand (gm_n2802, gm_n1055, gm_n76, in_25, gm_n2801, gm_n1185);
	nor (gm_n2803, gm_n2802, gm_n50, in_30);
	or (gm_n2804, gm_n254, gm_n246, gm_n64);
	nor (gm_n2805, gm_n107, in_16, gm_n157, gm_n2804, gm_n221);
	nand (gm_n2806, gm_n261, in_24, gm_n72, gm_n2805, gm_n472);
	nor (gm_n2807, gm_n260, gm_n229, in_28, gm_n2806);
	nor (gm_n2808, gm_n622, in_15, in_11, gm_n1664, gm_n666);
	nand (gm_n2809, gm_n165, gm_n195, gm_n102, gm_n2808, gm_n612);
	nor (gm_n2810, gm_n575, in_31, gm_n133, gm_n2809, gm_n581);
	nor (gm_n2811, gm_n673, in_15, gm_n58, gm_n1732, gm_n399);
	nand (gm_n2812, gm_n509, in_23, gm_n102, gm_n2811, gm_n612);
	nor (gm_n2813, gm_n303, gm_n50, gm_n133, gm_n2812, gm_n581);
	nor (gm_n2814, gm_n2807, gm_n2803, gm_n2800, gm_n2813, gm_n2810);
	nand (gm_n2815, gm_n63, gm_n157, gm_n64, gm_n747, gm_n232);
	nor (gm_n2816, gm_n179, gm_n72, in_16, gm_n2815, gm_n742);
	nand (gm_n2817, gm_n100, gm_n78, gm_n52, gm_n2816, gm_n207);
	nor (gm_n2818, gm_n2817, gm_n268);
	nor (gm_n2819, gm_n504, in_16, gm_n157, gm_n1123, gm_n159);
	nand (gm_n2820, gm_n85, gm_n52, in_20, gm_n2819, gm_n261);
	nor (gm_n2821, gm_n206, gm_n80, gm_n78, gm_n2820);
	nor (gm_n2822, gm_n727, in_15, gm_n58, gm_n499, gm_n672);
	nand (gm_n2823, gm_n299, in_23, gm_n102, gm_n2822, gm_n361);
	nor (gm_n2824, gm_n617, gm_n50, gm_n133, gm_n2823, gm_n611);
	nor (gm_n2825, gm_n2824, gm_n2821, gm_n2818);
	nor (gm_n2826, gm_n727, in_15, gm_n58, gm_n1675, gm_n366);
	nand (gm_n2827, gm_n293, in_23, gm_n102, gm_n2826, gm_n362);
	nor (gm_n2828, gm_n611, in_31, in_27, gm_n2827, gm_n671);
	nor (gm_n2829, gm_n672, in_15, gm_n58, gm_n1485, gm_n673);
	nand (gm_n2830, gm_n166, gm_n195, in_19, gm_n2829, gm_n336);
	nor (gm_n2831, gm_n575, gm_n50, gm_n133, gm_n2830, gm_n581);
	nand (gm_n2832, gm_n425, gm_n309, gm_n110);
	nor (gm_n2833, gm_n117, gm_n105, in_11, gm_n2832, gm_n426);
	nand (gm_n2834, gm_n73, in_23, gm_n102, gm_n2833, gm_n455);
	nor (gm_n2835, gm_n436, gm_n50, gm_n133, gm_n2834);
	nor (gm_n2836, gm_n2835, gm_n2831, gm_n2828);
	nand (gm_n2837, gm_n2814, gm_n2797, gm_n2794, gm_n2836, gm_n2825);
	or (gm_n2838, gm_n453, in_15, gm_n58, gm_n2590, gm_n997);
	nor (gm_n2839, gm_n510, gm_n195, in_19, gm_n2838, gm_n983);
	nand (gm_n2840, gm_n306, in_31, gm_n133, gm_n2839);
	or (gm_n2841, gm_n89, in_12, gm_n64, gm_n286, gm_n160);
	or (gm_n2842, gm_n106, gm_n72, gm_n68, gm_n2841, gm_n178);
	nor (gm_n2843, gm_n216, gm_n78, in_24, gm_n2842, gm_n412);
	nand (gm_n2844, gm_n2843, gm_n97);
	and (gm_n2845, gm_n118, gm_n105, in_8, gm_n1907, gm_n346);
	nand (gm_n2846, gm_n166, gm_n195, in_19, gm_n2845, gm_n313);
	or (gm_n2847, gm_n51, gm_n50, in_27, gm_n2846, gm_n983);
	nand (gm_n2848, gm_n2847, gm_n2844, gm_n2840);
	nand (gm_n2849, gm_n425, in_15, gm_n58, gm_n797, gm_n427);
	nor (gm_n2850, gm_n127, gm_n195, in_19, gm_n2849, gm_n395);
	nand (gm_n2851, gm_n115, in_31, gm_n133, gm_n2850, gm_n173);
	nand (gm_n2852, gm_n189, in_16, in_12, gm_n893, gm_n180);
	nor (gm_n2853, gm_n187, gm_n52, gm_n72, gm_n2852, gm_n804);
	nand (gm_n2854, gm_n462, gm_n217, in_28, gm_n2853);
	or (gm_n2855, gm_n109, gm_n121, in_5, gm_n465);
	or (gm_n2856, gm_n672, in_15, in_11, gm_n2855, gm_n618);
	nor (gm_n2857, gm_n117, gm_n195, gm_n102, gm_n2856, gm_n127);
	nand (gm_n2858, gm_n173, gm_n50, gm_n133, gm_n2857, gm_n392);
	nand (gm_n2859, gm_n2858, gm_n2854, gm_n2851);
	nor (gm_n2860, gm_n2837, gm_n2791, gm_n2788, gm_n2859, gm_n2848);
	nor (gm_n2861, gm_n319, gm_n105, gm_n58, gm_n992, gm_n399);
	nand (gm_n2862, gm_n509, gm_n195, in_19, gm_n2861, gm_n612);
	nor (gm_n2863, gm_n174, gm_n50, in_27, gm_n2862, gm_n303);
	nor (gm_n2864, gm_n106, gm_n68, gm_n157, gm_n1029, gm_n159);
	nand (gm_n2865, gm_n252, gm_n52, gm_n72, gm_n2864, gm_n472);
	nor (gm_n2866, gm_n216, gm_n176, gm_n78, gm_n2865);
	nor (gm_n2867, gm_n253, in_15, gm_n64, gm_n997, gm_n386);
	nand (gm_n2868, gm_n73, gm_n195, gm_n102, gm_n2867, gm_n582);
	nor (gm_n2869, gm_n575, gm_n50, in_27, gm_n2868, gm_n671);
	nor (gm_n2870, gm_n2869, gm_n2866, gm_n2863);
	nor (gm_n2871, gm_n107, in_16, gm_n157, gm_n2804, gm_n179);
	nand (gm_n2872, gm_n85, in_24, in_20, gm_n2871, gm_n183);
	nor (gm_n2873, gm_n268, gm_n80, in_28, gm_n2872);
	nor (gm_n2874, gm_n399, gm_n105, in_11, gm_n2697, gm_n618);
	nand (gm_n2875, gm_n582, gm_n195, gm_n102, gm_n2874, gm_n509);
	nor (gm_n2876, gm_n51, gm_n50, in_27, gm_n2875, gm_n54);
	nor (gm_n2877, gm_n88, gm_n68, in_12, gm_n2039, gm_n221);
	nand (gm_n2878, gm_n100, in_24, in_20, gm_n2877, gm_n472);
	nor (gm_n2879, gm_n780, gm_n176, gm_n78, gm_n2878);
	nor (gm_n2880, gm_n2879, gm_n2876, gm_n2873);
	nand (gm_n2881, gm_n2860, gm_n2785, gm_n2782, gm_n2880, gm_n2870);
	or (gm_n2882, in_7, in_6, gm_n62, gm_n160, in_8);
	nor (gm_n2883, gm_n221, in_16, in_12, gm_n2882, gm_n253);
	nand (gm_n2884, gm_n219, in_24, gm_n72, gm_n2883, gm_n220);
	nor (gm_n2885, gm_n132, gm_n216, gm_n78, gm_n2884);
	and (gm_n2886, gm_n766, gm_n68, gm_n157, gm_n2104, gm_n341);
	nand (gm_n2887, gm_n252, in_24, gm_n72, gm_n2886, gm_n269);
	nor (gm_n2888, gm_n780, gm_n229, gm_n78, gm_n2887);
	nor (gm_n2889, gm_n106, in_16, in_12, gm_n1525, gm_n286);
	nand (gm_n2890, gm_n85, gm_n52, gm_n72, gm_n2889, gm_n252);
	nor (gm_n2891, gm_n218, gm_n216, in_28, gm_n2890);
	or (gm_n2892, gm_n2885, gm_n2881, gm_n2779, gm_n2891, gm_n2888);
	not (gm_n2893, gm_n488);
	and (gm_n2894, gm_n87, gm_n65, in_8, gm_n200, gm_n210);
	nor (gm_n2895, in_13, gm_n157, in_11);
	and (gm_n2896, gm_n482, in_18, in_14, gm_n2895, gm_n2894);
	nand (gm_n2897, gm_n637, gm_n98, in_22, gm_n2896, gm_n1902);
	nor (gm_n2898, gm_n2893, in_31, in_30, gm_n2897);
	nor (gm_n2899, gm_n179, in_16, in_12, gm_n1728, gm_n245);
	nand (gm_n2900, gm_n237, in_24, gm_n72, gm_n2899, gm_n183);
	nor (gm_n2901, gm_n218, gm_n243, in_28, gm_n2900);
	and (gm_n2902, gm_n120, gm_n105, in_11, gm_n1683, gm_n311);
	and (gm_n2903, gm_n299, gm_n195, gm_n102, gm_n2902, gm_n361);
	and (gm_n2904, gm_n55, gm_n50, in_27, gm_n2903, gm_n508);
	nor (gm_n2905, gm_n2904, gm_n2901, gm_n2898);
	not (gm_n2906, gm_n2905);
	and (gm_n2907, gm_n270, in_16, gm_n157, gm_n1497, gm_n766);
	nand (gm_n2908, gm_n85, gm_n52, in_20, gm_n2907, gm_n220);
	nor (gm_n2909, gm_n208, gm_n206, in_28, gm_n2908);
	and (gm_n2910, gm_n66, gm_n105, gm_n58, gm_n1232, gm_n540);
	and (gm_n2911, gm_n166, gm_n195, gm_n102, gm_n2910, gm_n336);
	and (gm_n2912, gm_n307, gm_n50, in_27, gm_n2911, gm_n677);
	and (gm_n2913, gm_n138, gm_n157, in_8, gm_n1953, gm_n341);
	nand (gm_n2914, gm_n85, gm_n72, gm_n68, gm_n2913, gm_n100);
	nor (gm_n2915, gm_n243, gm_n78, gm_n52, gm_n2914, gm_n268);
	nor (gm_n2916, gm_n2915, gm_n2912, gm_n2909);
	not (gm_n2917, gm_n2916);
	or (gm_n2918, gm_n2892, gm_n2775, gm_n2772, gm_n2917, gm_n2906);
	nor (gm_n2919, gm_n57, gm_n102, in_15, gm_n2265, gm_n332);
	nand (gm_n2920, gm_n173, gm_n133, in_23, gm_n2919, gm_n361);
	nor (gm_n2921, gm_n2920, gm_n360, gm_n50);
	nor (gm_n2922, gm_n167, in_16, in_12, gm_n1050, gm_n221);
	and (gm_n2923, gm_n183, in_24, gm_n72, gm_n2922, gm_n472);
	and (gm_n2924, gm_n99, gm_n77, in_28, gm_n2923);
	and (gm_n2925, gm_n818, in_15, gm_n58, gm_n540, gm_n449);
	nand (gm_n2926, gm_n336, gm_n195, gm_n102, gm_n2925, gm_n452);
	nor (gm_n2927, gm_n360, gm_n50, in_27, gm_n2926, gm_n983);
	nor (gm_n2928, gm_n2927, gm_n2924, gm_n2921);
	not (gm_n2929, gm_n2928);
	nor (gm_n2930, gm_n673, gm_n105, gm_n58, gm_n762, gm_n622);
	nand (gm_n2931, gm_n509, gm_n195, in_19, gm_n2930, gm_n612);
	nor (gm_n2932, gm_n575, gm_n50, in_27, gm_n2931, gm_n581);
	or (gm_n2933, gm_n167, in_12, gm_n64, gm_n347, gm_n160);
	or (gm_n2934, gm_n139, gm_n72, in_16, gm_n2933, gm_n459);
	or (gm_n2935, gm_n208, gm_n78, gm_n52, gm_n2934, gm_n561);
	nor (gm_n2936, gm_n2935, gm_n268);
	nor (gm_n2937, gm_n727, gm_n105, in_11, gm_n701, gm_n622);
	and (gm_n2938, gm_n582, gm_n195, in_19, gm_n2937, gm_n336);
	and (gm_n2939, gm_n115, gm_n50, gm_n133, gm_n2938, gm_n455);
	nor (gm_n2940, gm_n2939, gm_n2936, gm_n2932);
	not (gm_n2941, gm_n2940);
	or (gm_n2942, gm_n2918, gm_n2769, gm_n2766, gm_n2941, gm_n2929);
	nor (gm_n2943, gm_n107, in_12, in_8, gm_n1043, gm_n158);
	nand (gm_n2944, gm_n230, in_20, in_16, gm_n2943, gm_n261);
	nor (gm_n2945, gm_n176, in_28, in_24, gm_n2944, gm_n260);
	and (gm_n2946, gm_n297, gm_n105, gm_n58, gm_n2332, gm_n1232);
	nand (gm_n2947, gm_n361, in_23, in_19, gm_n2946, gm_n362);
	nor (gm_n2948, gm_n436, gm_n50, in_27, gm_n2947, gm_n983);
	nor (gm_n2949, gm_n221, in_16, gm_n157, gm_n549, gm_n245);
	and (gm_n2950, gm_n196, in_24, in_20, gm_n2949, gm_n472);
	and (gm_n2951, gm_n492, gm_n370, gm_n78, gm_n2950);
	and (gm_n2952, gm_n180, gm_n68, in_12, gm_n645, gm_n138);
	and (gm_n2953, gm_n219, in_24, in_20, gm_n2952, gm_n209);
	and (gm_n2954, gm_n194, gm_n79, gm_n78, gm_n2953);
	nor (gm_n2955, gm_n672, in_15, gm_n58, gm_n1127, gm_n396);
	nand (gm_n2956, gm_n126, in_23, gm_n102, gm_n2955, gm_n612);
	nor (gm_n2957, gm_n54, in_31, gm_n133, gm_n2956, gm_n436);
	nor (gm_n2958, gm_n244, in_12, gm_n64, gm_n1039, gm_n245);
	nand (gm_n2959, gm_n219, in_20, in_16, gm_n2958, gm_n196);
	nor (gm_n2960, gm_n216, gm_n78, gm_n52, gm_n2959, gm_n475);
	and (gm_n2961, gm_n138, in_12, in_8, gm_n1953, gm_n346);
	nand (gm_n2962, gm_n196, gm_n72, gm_n68, gm_n2961, gm_n472);
	or (gm_n2963, gm_n371, gm_n78, in_24, gm_n2962, gm_n475);
	nor (gm_n2964, gm_n139, in_16, in_12, gm_n833, gm_n253);
	nand (gm_n2965, gm_n219, gm_n52, in_20, gm_n2964, gm_n196);
	or (gm_n2966, gm_n268, gm_n216, gm_n78, gm_n2965);
	nand (gm_n2967, gm_n146, gm_n68, in_12, gm_n876, gm_n147);
	or (gm_n2968, gm_n156, in_24, gm_n72, gm_n2967, gm_n561);
	nor (gm_n2969, gm_n780, gm_n229, in_28, gm_n2968);
	and (gm_n2970, gm_n309, gm_n110, in_8);
	nand (gm_n2971, gm_n189, in_16, gm_n157, gm_n2970, gm_n180);
	or (gm_n2972, gm_n84, gm_n52, in_20, gm_n2971, gm_n742);
	nor (gm_n2973, gm_n218, gm_n208, gm_n78, gm_n2972);
	nor (gm_n2974, gm_n319, in_15, gm_n58, gm_n2081, gm_n622);
	nand (gm_n2975, gm_n313, gm_n195, in_19, gm_n2974, gm_n612);
	nor (gm_n2976, gm_n303, in_31, in_27, gm_n2975, gm_n983);
	and (gm_n2977, gm_n425, gm_n105, gm_n58, gm_n1232, gm_n540);
	nand (gm_n2978, gm_n362, gm_n195, in_19, gm_n2977, gm_n509);
	nor (gm_n2979, gm_n360, in_31, gm_n133, gm_n2978, gm_n983);
	nor (gm_n2980, gm_n396, gm_n105, gm_n58, gm_n1001, gm_n426);
	nand (gm_n2981, gm_n69, in_23, gm_n102, gm_n2980, gm_n165);
	nor (gm_n2982, gm_n360, gm_n50, in_27, gm_n2981, gm_n617);
	and (gm_n2983, gm_n449, in_15, gm_n58, gm_n1719, gm_n1232);
	nand (gm_n2984, gm_n336, in_23, in_19, gm_n2983, gm_n452);
	nor (gm_n2985, gm_n575, gm_n50, gm_n133, gm_n2984, gm_n983);
	and (gm_n2986, gm_n180, in_16, in_12, gm_n1750, gm_n231);
	nand (gm_n2987, gm_n230, in_24, gm_n72, gm_n2986, gm_n252);
	nor (gm_n2988, gm_n218, gm_n208, gm_n78, gm_n2987);
	nor (gm_n2989, gm_n399, in_15, in_11, gm_n1664, gm_n618);
	nand (gm_n2990, gm_n313, in_23, gm_n102, gm_n2989, gm_n362);
	nor (gm_n2991, gm_n51, in_31, in_27, gm_n2990, gm_n174);
	nor (gm_n2992, gm_n179, gm_n68, in_12, gm_n255, gm_n245);
	nand (gm_n2993, gm_n100, gm_n52, in_20, gm_n2992, gm_n137);
	nor (gm_n2994, gm_n243, gm_n176, gm_n78, gm_n2993);
	or (gm_n2995, gm_n2988, gm_n2985, gm_n2982, gm_n2994, gm_n2991);
	and (gm_n2996, gm_n346, gm_n157, in_8, gm_n450, gm_n308);
	and (gm_n2997, gm_n219, gm_n72, gm_n68, gm_n2996, gm_n766);
	nand (gm_n2998, gm_n177, gm_n78, gm_n52, gm_n2997, gm_n209);
	nor (gm_n2999, gm_n2998, gm_n687);
	nor (gm_n3000, gm_n106, in_16, in_12, gm_n1029, gm_n253);
	nand (gm_n3001, gm_n261, gm_n52, gm_n72, gm_n3000, gm_n472);
	nor (gm_n3002, gm_n218, gm_n243, gm_n78, gm_n3001);
	or (gm_n3003, gm_n179, gm_n68, in_12, gm_n2162, gm_n253);
	or (gm_n3004, gm_n516, in_24, gm_n72, gm_n3003, gm_n742);
	nor (gm_n3005, gm_n80, gm_n229, in_28, gm_n3004);
	or (gm_n3006, gm_n3005, gm_n3002, gm_n2999);
	nor (gm_n3007, gm_n622, gm_n105, gm_n58, gm_n762, gm_n666);
	nand (gm_n3008, gm_n313, in_23, gm_n102, gm_n3007, gm_n452);
	nor (gm_n3009, gm_n1118, in_31, in_27, gm_n3008, gm_n360);
	nand (gm_n3010, gm_n118, in_15, in_11, gm_n1319, gm_n665);
	or (gm_n3011, gm_n1703, gm_n195, in_19, gm_n3010, gm_n911);
	nor (gm_n3012, gm_n575, gm_n50, gm_n133, gm_n3011, gm_n983);
	nand (gm_n3013, gm_n231, in_16, gm_n157, gm_n1006, gm_n270);
	or (gm_n3014, gm_n101, in_24, in_20, gm_n3013, gm_n178);
	nor (gm_n3015, gm_n780, gm_n229, gm_n78, gm_n3014);
	or (gm_n3016, gm_n3015, gm_n3012, gm_n3009);
	or (gm_n3017, gm_n2995, gm_n2979, gm_n2976, gm_n3016, gm_n3006);
	nand (gm_n3018, gm_n188, gm_n68, in_12, gm_n1237, gm_n231);
	or (gm_n3019, gm_n101, gm_n52, gm_n72, gm_n3018, gm_n103);
	nor (gm_n3020, gm_n268, gm_n80, in_28, gm_n3019);
	and (gm_n3021, gm_n341, gm_n157, in_8, gm_n511, gm_n309);
	and (gm_n3022, gm_n86, gm_n72, gm_n68, gm_n3021, gm_n237);
	and (gm_n3023, gm_n196, in_28, gm_n52, gm_n3022, gm_n462);
	and (gm_n3024, gm_n3023, gm_n474);
	nor (gm_n3025, gm_n106, in_16, gm_n157, gm_n688, gm_n253);
	and (gm_n3026, gm_n85, in_24, gm_n72, gm_n3025, gm_n196);
	and (gm_n3027, gm_n492, gm_n177, in_28, gm_n3026);
	or (gm_n3028, gm_n3027, gm_n3024, gm_n3020);
	nor (gm_n3029, gm_n244, in_16, in_12, gm_n2534, gm_n253);
	and (gm_n3030, gm_n252, in_24, in_20, gm_n3029, gm_n517);
	and (gm_n3031, gm_n207, gm_n186, gm_n78, gm_n3030);
	nor (gm_n3032, gm_n179, gm_n68, in_12, gm_n577, gm_n286);
	nand (gm_n3033, gm_n83, gm_n52, gm_n72, gm_n3032, gm_n230);
	nor (gm_n3034, gm_n475, gm_n216, in_28, gm_n3033);
	or (gm_n3035, gm_n57, gm_n105, gm_n58, gm_n1329, gm_n673);
	or (gm_n3036, gm_n70, gm_n195, in_19, gm_n3035, gm_n510);
	nor (gm_n3037, gm_n1118, gm_n50, gm_n133, gm_n3036, gm_n303);
	or (gm_n3038, gm_n3037, gm_n3034, gm_n3031);
	nor (gm_n3039, gm_n3017, gm_n2973, gm_n2969, gm_n3038, gm_n3028);
	and (gm_n3040, gm_n612, gm_n102, in_15, gm_n1912, gm_n1232);
	and (gm_n3041, gm_n165, gm_n133, in_23, gm_n3040, gm_n307);
	and (gm_n3042, gm_n3041, gm_n677, gm_n50);
	and (gm_n3043, gm_n198, in_16, gm_n157, gm_n1547, gm_n346);
	nand (gm_n3044, gm_n137, gm_n52, in_20, gm_n3043, gm_n220);
	nor (gm_n3045, gm_n260, gm_n206, in_28, gm_n3044);
	and (gm_n3046, gm_n124, gm_n157, gm_n64, gm_n308, gm_n147);
	and (gm_n3047, gm_n231, gm_n72, gm_n68, gm_n3046, gm_n269);
	and (gm_n3048, gm_n252, gm_n78, in_24, gm_n3047, gm_n259);
	and (gm_n3049, gm_n3048, gm_n217);
	nor (gm_n3050, gm_n3049, gm_n3045, gm_n3042);
	nand (gm_n3051, gm_n146, gm_n68, in_12, gm_n1178, gm_n341);
	or (gm_n3052, gm_n84, gm_n52, in_20, gm_n3051, gm_n602);
	nor (gm_n3053, gm_n216, gm_n229, in_28, gm_n3052);
	and (gm_n3054, gm_n147, in_16, gm_n157, gm_n1437, gm_n629);
	nand (gm_n3055, gm_n83, in_24, in_20, gm_n3054, gm_n237);
	nor (gm_n3056, gm_n218, gm_n216, gm_n78, gm_n3055);
	nor (gm_n3057, gm_n179, in_16, gm_n157, gm_n2431, gm_n253);
	nand (gm_n3058, gm_n237, in_24, in_20, gm_n3057, gm_n261);
	nor (gm_n3059, gm_n268, gm_n243, gm_n78, gm_n3058);
	nor (gm_n3060, gm_n3059, gm_n3056, gm_n3053);
	nand (gm_n3061, gm_n3039, gm_n2966, gm_n2963, gm_n3060, gm_n3050);
	and (gm_n3062, gm_n140, gm_n157, in_8, gm_n341, gm_n238);
	nand (gm_n3063, gm_n138, gm_n72, gm_n68, gm_n3062, gm_n472);
	nor (gm_n3064, gm_n804, in_28, in_24, gm_n3063, gm_n260);
	nand (gm_n3065, gm_n3064, gm_n205);
	nor (gm_n3066, gm_n432, in_15, gm_n58, gm_n992, gm_n622);
	nand (gm_n3067, gm_n73, gm_n195, in_19, gm_n3066, gm_n582);
	or (gm_n3068, gm_n51, gm_n50, in_27, gm_n3067, gm_n581);
	nand (gm_n3069, gm_n86, gm_n68, gm_n157, gm_n1173, gm_n232);
	nor (gm_n3070, gm_n628, in_24, in_20, gm_n3069, gm_n742);
	nand (gm_n3071, gm_n97, gm_n79, gm_n78, gm_n3070);
	nand (gm_n3072, gm_n3071, gm_n3068, gm_n3065);
	nand (gm_n3073, gm_n180, in_16, gm_n157, gm_n2244, gm_n231);
	nor (gm_n3074, gm_n84, gm_n52, in_20, gm_n3073, gm_n602);
	nand (gm_n3075, gm_n79, gm_n77, gm_n78, gm_n3074);
	or (gm_n3076, gm_n57, in_15, in_11, gm_n1732, gm_n727);
	nor (gm_n3077, gm_n127, in_23, in_19, gm_n3076, gm_n363);
	nand (gm_n3078, gm_n55, gm_n50, gm_n133, gm_n3077, gm_n392);
	nor (gm_n3079, gm_n106, in_16, gm_n157, gm_n245, gm_n170);
	nand (gm_n3080, gm_n196, gm_n52, in_20, gm_n3079, gm_n472);
	or (gm_n3081, gm_n780, gm_n132, in_28, gm_n3080);
	nand (gm_n3082, gm_n3081, gm_n3078, gm_n3075);
	or (gm_n3083, gm_n3061, gm_n2960, gm_n2957, gm_n3082, gm_n3072);
	nor (gm_n3084, gm_n57, in_15, gm_n58, gm_n618, gm_n282);
	nand (gm_n3085, gm_n361, in_23, in_19, gm_n3084, gm_n612);
	nor (gm_n3086, gm_n617, gm_n50, gm_n133, gm_n3085, gm_n611);
	nor (gm_n3087, gm_n107, in_16, gm_n157, gm_n2643, gm_n158);
	and (gm_n3088, gm_n83, gm_n52, gm_n72, gm_n3087, gm_n237);
	and (gm_n3089, gm_n492, gm_n79, in_28, gm_n3088);
	nor (gm_n3090, gm_n504, gm_n68, gm_n157, gm_n1525, gm_n222);
	nand (gm_n3091, gm_n83, in_24, gm_n72, gm_n3090, gm_n230);
	nor (gm_n3092, gm_n371, gm_n218, in_28, gm_n3091);
	or (gm_n3093, gm_n3086, gm_n3083, gm_n2954, gm_n3092, gm_n3089);
	and (gm_n3094, gm_n333, in_15, in_11, gm_n2237, gm_n166);
	and (gm_n3095, gm_n313, in_23, gm_n102, gm_n3094, gm_n455);
	and (gm_n3096, gm_n677, in_31, gm_n133, gm_n3095);
	and (gm_n3097, gm_n198, in_16, in_12, gm_n987, gm_n341);
	and (gm_n3098, gm_n183, gm_n52, in_20, gm_n3097, gm_n269);
	and (gm_n3099, gm_n492, gm_n462, in_28, gm_n3098);
	nand (gm_n3100, gm_n188, in_12, gm_n64, gm_n705, gm_n511);
	or (gm_n3101, gm_n221, gm_n72, in_16, gm_n3100, gm_n459);
	or (gm_n3102, gm_n628, in_28, in_24, gm_n3101, gm_n780);
	nor (gm_n3103, gm_n3102, gm_n206);
	nor (gm_n3104, gm_n3103, gm_n3099, gm_n3096);
	not (gm_n3105, gm_n3104);
	nand (gm_n3106, gm_n66, in_15, gm_n58, gm_n1102, gm_n938);
	nor (gm_n3107, gm_n294, gm_n195, in_19, gm_n3106, gm_n300);
	and (gm_n3108, gm_n455, in_31, in_27, gm_n3107, gm_n508);
	nor (gm_n3109, gm_n504, in_16, in_12, gm_n1811, gm_n286);
	nand (gm_n3110, gm_n220, gm_n52, gm_n72, gm_n3109, gm_n230);
	nor (gm_n3111, gm_n268, gm_n135, in_28, gm_n3110);
	and (gm_n3112, gm_n188, in_16, in_12, gm_n1106, gm_n231);
	and (gm_n3113, gm_n230, in_24, gm_n72, gm_n3112, gm_n261);
	and (gm_n3114, gm_n134, gm_n194, gm_n78, gm_n3113);
	nor (gm_n3115, gm_n3114, gm_n3111, gm_n3108);
	not (gm_n3116, gm_n3115);
	or (gm_n3117, gm_n3093, gm_n2951, gm_n2948, gm_n3116, gm_n3105);
	or (gm_n3118, gm_n347, gm_n254, in_8);
	nor (gm_n3119, gm_n244, in_16, gm_n157, gm_n3118, gm_n222);
	and (gm_n3120, gm_n220, gm_n52, gm_n72, gm_n3119, gm_n517);
	and (gm_n3121, gm_n259, gm_n77, gm_n78, gm_n3120);
	nor (new_out2, gm_n3117, gm_n2945, gm_n2942, gm_n3121);
	nor (gm_n3123, gm_n221, gm_n68, in_12, gm_n1986, gm_n253);
	nand (gm_n3124, gm_n83, gm_n52, gm_n72, gm_n3123, gm_n472);
	nor (gm_n3125, gm_n260, gm_n206, gm_n78, gm_n3124);
	and (gm_n3126, gm_n66, in_15, in_11, gm_n334, gm_n118);
	nand (gm_n3127, gm_n452, in_23, in_19, gm_n3126, gm_n509);
	nor (gm_n3128, gm_n51, in_31, in_27, gm_n3127, gm_n983);
	and (gm_n3129, gm_n180, in_16, gm_n157, gm_n233, gm_n629);
	and (gm_n3130, gm_n261, in_24, gm_n72, gm_n3129, gm_n472);
	and (gm_n3131, gm_n370, gm_n217, gm_n78, gm_n3130);
	and (gm_n3132, gm_n2776, in_15, in_11, gm_n2594, gm_n1232);
	nand (gm_n3133, gm_n126, in_23, in_19, gm_n3132, gm_n166);
	or (gm_n3134, gm_n617, gm_n50, in_27, gm_n3133, gm_n436);
	nor (gm_n3135, gm_n167, gm_n68, in_12, gm_n179, gm_n170);
	nand (gm_n3136, gm_n220, in_24, gm_n72, gm_n3135, gm_n517);
	or (gm_n3137, gm_n206, gm_n216, gm_n78, gm_n3136);
	nor (gm_n3138, gm_n221, gm_n68, gm_n157, gm_n2077, gm_n245);
	nand (gm_n3139, gm_n196, in_24, in_20, gm_n3138, gm_n472);
	nor (gm_n3140, gm_n208, gm_n268, gm_n78, gm_n3139);
	nand (gm_n3141, gm_n747, gm_n210, in_8);
	nor (gm_n3142, gm_n167, gm_n68, gm_n157, gm_n3141, gm_n221);
	nand (gm_n3143, gm_n83, gm_n52, gm_n72, gm_n3142, gm_n85);
	nor (gm_n3144, gm_n371, gm_n229, in_28, gm_n3143);
	nor (gm_n3145, gm_n179, in_16, in_12, gm_n577, gm_n245);
	nand (gm_n3146, gm_n230, gm_n52, gm_n72, gm_n3145, gm_n261);
	or (gm_n3147, gm_n260, gm_n176, in_28, gm_n3146);
	nor (gm_n3148, gm_n159, gm_n68, in_12, gm_n2431, gm_n168);
	nand (gm_n3149, gm_n100, in_24, gm_n72, gm_n3148, gm_n237);
	or (gm_n3150, gm_n206, gm_n243, gm_n78, gm_n3149);
	nand (gm_n3151, gm_n63, in_12, in_8, gm_n1226, gm_n270);
	nor (gm_n3152, gm_n187, in_20, in_16, gm_n3151, gm_n106);
	nand (gm_n3153, gm_n99, gm_n78, gm_n52, gm_n3152, gm_n209);
	nor (gm_n3154, gm_n3153, gm_n229);
	nor (gm_n3155, gm_n167, in_16, in_12, gm_n1505, gm_n158);
	nand (gm_n3156, gm_n183, gm_n52, gm_n72, gm_n3155, gm_n472);
	nor (gm_n3157, gm_n208, gm_n229, in_28, gm_n3156);
	or (gm_n3158, gm_n432, in_15, in_11, gm_n997, gm_n880);
	nor (gm_n3159, gm_n337, in_23, in_19, gm_n3158, gm_n453);
	and (gm_n3160, gm_n302, gm_n50, gm_n133, gm_n3159, gm_n508);
	nor (gm_n3161, gm_n253, in_15, gm_n64, gm_n386, gm_n366);
	nand (gm_n3162, gm_n73, in_23, gm_n102, gm_n3161, gm_n362);
	nor (gm_n3163, gm_n581, gm_n50, in_27, gm_n3162, gm_n842);
	nor (gm_n3164, gm_n244, gm_n68, gm_n157, gm_n2077, gm_n88);
	nand (gm_n3165, gm_n237, gm_n52, gm_n72, gm_n3164, gm_n183);
	nor (gm_n3166, gm_n687, gm_n135, in_28, gm_n3165);
	and (gm_n3167, gm_n189, in_12, gm_n64, gm_n1907, gm_n232);
	nand (gm_n3168, gm_n137, in_20, in_16, gm_n3167, gm_n183);
	nor (gm_n3169, gm_n206, in_28, gm_n52, gm_n3168, gm_n780);
	and (gm_n3170, gm_n189, in_16, gm_n157, gm_n190, gm_n147);
	nand (gm_n3171, gm_n137, gm_n52, gm_n72, gm_n3170, gm_n209);
	nor (gm_n3172, gm_n176, gm_n80, gm_n78, gm_n3171);
	or (gm_n3173, gm_n3166, gm_n3163, gm_n3160, gm_n3172, gm_n3169);
	or (gm_n3174, gm_n107, in_16, gm_n157, gm_n568, gm_n139);
	nor (gm_n3175, gm_n84, gm_n52, in_20, gm_n3174, gm_n413);
	nand (gm_n3176, gm_n205, gm_n177, in_28, gm_n3175);
	and (gm_n3177, gm_n198, in_16, in_12, gm_n1715, gm_n354);
	and (gm_n3178, gm_n209, in_24, in_20, gm_n3177, gm_n472);
	nand (gm_n3179, gm_n492, gm_n370, in_28, gm_n3178);
	or (gm_n3180, gm_n672, gm_n105, gm_n58, gm_n1214, gm_n618);
	nor (gm_n3181, gm_n332, gm_n195, in_19, gm_n3180, gm_n337);
	nand (gm_n3182, gm_n302, gm_n50, gm_n133, gm_n3181, gm_n677);
	nand (gm_n3183, gm_n3182, gm_n3179, gm_n3176);
	or (gm_n3184, gm_n167, gm_n68, in_12, gm_n781, gm_n179);
	nor (gm_n3185, gm_n103, in_24, gm_n72, gm_n3184, gm_n804);
	nand (gm_n3186, gm_n492, gm_n99, in_28, gm_n3185);
	nor (gm_n3187, gm_n119, gm_n105, gm_n58, gm_n2504, gm_n622);
	nand (gm_n3188, gm_n166, in_23, gm_n102, gm_n3187, gm_n313);
	or (gm_n3189, gm_n303, in_31, gm_n133, gm_n3188, gm_n983);
	nor (gm_n3190, gm_n117, gm_n195, in_19, gm_n1620, gm_n337);
	nand (gm_n3191, gm_n393, in_31, gm_n133, gm_n3190, gm_n508);
	nand (gm_n3192, gm_n3191, gm_n3189, gm_n3186);
	nor (gm_n3193, gm_n3173, gm_n3157, gm_n3154, gm_n3192, gm_n3183);
	nor (gm_n3194, gm_n672, in_15, in_11, gm_n1279, gm_n319);
	nand (gm_n3195, gm_n69, gm_n195, in_19, gm_n3194, gm_n313);
	nor (gm_n3196, gm_n54, gm_n50, gm_n133, gm_n3195, gm_n303);
	nor (gm_n3197, gm_n139, in_16, in_12, gm_n2568, gm_n222);
	nand (gm_n3198, gm_n137, in_24, in_20, gm_n3197, gm_n252);
	nor (gm_n3199, gm_n687, gm_n780, in_28, gm_n3198);
	nand (gm_n3200, gm_n333, gm_n105, in_11, gm_n1996, gm_n166);
	or (gm_n3201, gm_n337, gm_n195, in_19, gm_n3200, gm_n983);
	nor (gm_n3202, gm_n303, gm_n50, gm_n133, gm_n3201);
	nor (gm_n3203, gm_n3202, gm_n3199, gm_n3196);
	nor (gm_n3204, gm_n57, in_15, in_11, gm_n2602, gm_n432);
	nand (gm_n3205, gm_n165, in_23, in_19, gm_n3204, gm_n452);
	nor (gm_n3206, gm_n54, gm_n50, gm_n133, gm_n3205, gm_n436);
	nor (gm_n3207, gm_n167, gm_n68, gm_n157, gm_n2254, gm_n221);
	nand (gm_n3208, gm_n237, gm_n52, gm_n72, gm_n3207, gm_n220);
	nor (gm_n3209, gm_n206, gm_n216, gm_n78, gm_n3208);
	and (gm_n3210, gm_n449, gm_n105, in_11, gm_n2703, gm_n427);
	nand (gm_n3211, gm_n299, gm_n195, gm_n102, gm_n3210, gm_n336);
	nor (gm_n3212, gm_n303, in_31, gm_n133, gm_n3211, gm_n671);
	nor (gm_n3213, gm_n3212, gm_n3209, gm_n3206);
	nand (gm_n3214, gm_n3193, gm_n3150, gm_n3147, gm_n3213, gm_n3203);
	nor (gm_n3215, gm_n562, in_12, in_8, gm_n169, gm_n167);
	nand (gm_n3216, gm_n231, gm_n72, gm_n68, gm_n3215, gm_n472);
	nor (gm_n3217, gm_n243, gm_n78, in_24, gm_n3216, gm_n412);
	nand (gm_n3218, gm_n3217, gm_n492);
	nor (gm_n3219, in_7, in_6, gm_n62, gm_n271, gm_n64);
	nand (gm_n3220, gm_n138, gm_n68, in_12, gm_n3219, gm_n341);
	nor (gm_n3221, gm_n156, gm_n52, gm_n72, gm_n3220, gm_n197);
	nand (gm_n3222, gm_n474, gm_n134, gm_n78, gm_n3221);
	nor (gm_n3223, gm_n244, in_16, gm_n157, gm_n2882, gm_n245);
	and (gm_n3224, gm_n237, gm_n52, in_20, gm_n3223, gm_n261);
	nand (gm_n3225, gm_n205, gm_n79, gm_n78, gm_n3224);
	nand (gm_n3226, gm_n3225, gm_n3222, gm_n3218);
	nand (gm_n3227, gm_n188, gm_n68, gm_n157, gm_n1595, gm_n198);
	nor (gm_n3228, gm_n804, gm_n52, in_20, gm_n3227, gm_n602);
	nand (gm_n3229, gm_n186, gm_n99, gm_n78, gm_n3228);
	nand (gm_n3230, gm_n2776, gm_n105, gm_n58, gm_n2149, gm_n818);
	nor (gm_n3231, gm_n337, in_23, in_19, gm_n3230, gm_n363);
	nand (gm_n3232, gm_n115, in_31, gm_n133, gm_n3231, gm_n55);
	and (gm_n3233, gm_n146, in_16, gm_n157, gm_n1750, gm_n346);
	and (gm_n3234, gm_n137, in_24, gm_n72, gm_n3233, gm_n220);
	nand (gm_n3235, gm_n217, gm_n99, in_28, gm_n3234);
	nand (gm_n3236, gm_n3235, gm_n3232, gm_n3229);
	nor (gm_n3237, gm_n3214, gm_n3144, gm_n3140, gm_n3236, gm_n3226);
	nand (gm_n3238, gm_n63, gm_n157, in_8, gm_n200, gm_n270);
	nor (gm_n3239, gm_n504, in_20, in_16, gm_n3238, gm_n602);
	nand (gm_n3240, gm_n99, in_28, in_24, gm_n3239, gm_n261);
	nor (gm_n3241, gm_n3240, gm_n176);
	nor (gm_n3242, gm_n244, in_16, gm_n157, gm_n553, gm_n167);
	nand (gm_n3243, gm_n83, in_24, in_20, gm_n3242, gm_n230);
	nor (gm_n3244, gm_n475, gm_n780, in_28, gm_n3243);
	nor (gm_n3245, gm_n666, gm_n105, in_11, gm_n997, gm_n880);
	and (gm_n3246, gm_n293, gm_n195, gm_n102, gm_n3245, gm_n452);
	and (gm_n3247, gm_n302, in_31, in_27, gm_n3246, gm_n508);
	nor (gm_n3248, gm_n3247, gm_n3244, gm_n3241);
	nor (gm_n3249, gm_n179, in_16, in_12, gm_n2804, gm_n253);
	nand (gm_n3250, gm_n209, gm_n52, in_20, gm_n3249, gm_n269);
	nor (gm_n3251, gm_n687, gm_n260, in_28, gm_n3250);
	and (gm_n3252, gm_n136, in_14, in_13, gm_n2477, gm_n1900);
	nor (gm_n3253, in_21, gm_n72, in_19);
	nand (gm_n3254, gm_n639, in_26, in_22, gm_n3253, gm_n3252);
	nor (gm_n3255, gm_n2458, gm_n50, in_30, gm_n3254);
	nor (gm_n3256, gm_n727, in_15, gm_n58, gm_n2085, gm_n672);
	nand (gm_n3257, gm_n582, in_23, gm_n102, gm_n3256, gm_n361);
	nor (gm_n3258, gm_n1231, in_31, in_27, gm_n3257, gm_n611);
	nor (gm_n3259, gm_n3258, gm_n3255, gm_n3251);
	nand (gm_n3260, gm_n3237, gm_n3137, gm_n3134, gm_n3259, gm_n3248);
	and (gm_n3261, gm_n198, gm_n68, in_12, gm_n545, gm_n346);
	nand (gm_n3262, gm_n83, in_24, in_20, gm_n3261, gm_n472);
	nor (gm_n3263, gm_n218, gm_n135, in_28, gm_n3262);
	and (gm_n3264, gm_n629, gm_n68, in_12, gm_n1750, gm_n232);
	nand (gm_n3265, gm_n261, in_24, in_20, gm_n3264, gm_n269);
	nor (gm_n3266, gm_n687, gm_n216, gm_n78, gm_n3265);
	nor (gm_n3267, gm_n159, in_16, gm_n157, gm_n225, gm_n221);
	nand (gm_n3268, gm_n196, gm_n52, gm_n72, gm_n3267, gm_n517);
	nor (gm_n3269, gm_n132, gm_n216, in_28, gm_n3268);
	nor (gm_n3270, gm_n3269, gm_n3266, gm_n3263);
	not (gm_n3271, gm_n3270);
	nor (gm_n3272, gm_n167, gm_n68, gm_n157, gm_n1579, gm_n221);
	nand (gm_n3273, gm_n230, gm_n52, in_20, gm_n3272, gm_n261);
	nor (gm_n3274, gm_n780, gm_n268, in_28, gm_n3273);
	nor (gm_n3275, gm_n88, gm_n68, gm_n157, gm_n2053, gm_n139);
	nand (gm_n3276, gm_n219, gm_n52, gm_n72, gm_n3275, gm_n183);
	nor (gm_n3277, gm_n208, gm_n206, gm_n78, gm_n3276);
	nand (gm_n3278, gm_n1635, gm_n333, gm_n105);
	or (gm_n3279, gm_n332, gm_n195, in_19, gm_n3278, gm_n314);
	nor (gm_n3280, gm_n54, in_31, in_27, gm_n3279, gm_n678);
	nor (gm_n3281, gm_n3280, gm_n3277, gm_n3274);
	not (gm_n3282, gm_n3281);
	or (gm_n3283, gm_n3260, gm_n3131, gm_n3128, gm_n3282, gm_n3271);
	and (gm_n3284, gm_n188, gm_n333, in_15, gm_n1715, gm_n452);
	nand (gm_n3285, gm_n55, in_23, gm_n102, gm_n3284, gm_n165);
	nor (gm_n3286, gm_n575, in_31, in_27, gm_n3285);
	nand (gm_n3287, gm_n210, in_12, in_8, gm_n450, gm_n346);
	or (gm_n3288, gm_n244, in_20, gm_n68, gm_n3287, gm_n459);
	or (gm_n3289, gm_n80, gm_n78, gm_n52, gm_n3288, gm_n628);
	nor (gm_n3290, gm_n3289, gm_n229);
	nor (gm_n3291, gm_n139, gm_n68, gm_n157, gm_n568, gm_n222);
	and (gm_n3292, gm_n220, in_24, in_20, gm_n3291, gm_n230);
	and (gm_n3293, gm_n370, gm_n97, gm_n78, gm_n3292);
	or (gm_n3294, gm_n3286, gm_n3283, gm_n3125, gm_n3293, gm_n3290);
	nor (gm_n3295, gm_n107, in_12, in_8, gm_n733, gm_n223);
	and (gm_n3296, gm_n766, in_20, in_16, gm_n3295, gm_n230);
	nand (gm_n3297, gm_n79, gm_n78, in_24, gm_n3296, gm_n183);
	nor (gm_n3298, gm_n3297, gm_n268);
	nor (gm_n3299, gm_n88, in_16, in_12, gm_n1811, gm_n168);
	nand (gm_n3300, gm_n261, gm_n52, gm_n72, gm_n3299, gm_n517);
	nor (gm_n3301, gm_n780, gm_n206, gm_n78, gm_n3300);
	and (gm_n3302, gm_n449, gm_n105, in_11, gm_n621, gm_n424);
	nand (gm_n3303, gm_n126, in_23, gm_n102, gm_n3302, gm_n612);
	nor (gm_n3304, gm_n54, in_31, in_27, gm_n3303, gm_n611);
	and (gm_n3305, gm_n86, gm_n68, in_12, gm_n414, gm_n346);
	and (gm_n3306, gm_n183, gm_n52, gm_n72, gm_n3305, gm_n517);
	and (gm_n3307, gm_n134, gm_n77, in_28, gm_n3306);
	nand (gm_n3308, gm_n147, gm_n157, gm_n64, gm_n403, gm_n511);
	nor (gm_n3309, in_16, in_15, in_14);
	not (gm_n3310, gm_n3309);
	or (gm_n3311, gm_n732, gm_n116, gm_n56, gm_n3310, gm_n3308);
	nor (gm_n3312, gm_n326, gm_n53, gm_n81, gm_n3311, gm_n535);
	nand (gm_n3313, in_31, in_30, gm_n76, gm_n3312);
	nand (gm_n3314, gm_n180, in_16, in_12, gm_n706, gm_n231);
	nor (gm_n3315, gm_n178, in_24, gm_n72, gm_n3314, gm_n516);
	nand (gm_n3316, gm_n370, gm_n97, gm_n78, gm_n3315);
	nor (gm_n3317, gm_n727, in_15, in_11, gm_n1664, gm_n366);
	nand (gm_n3318, gm_n293, in_23, in_19, gm_n3317, gm_n612);
	nor (gm_n3319, gm_n1231, gm_n50, gm_n133, gm_n3318, gm_n303);
	nand (gm_n3320, gm_n63, gm_n61, in_11, gm_n427, gm_n120);
	nor (gm_n3321, gm_n337, gm_n102, gm_n105, gm_n3320, gm_n453);
	nand (gm_n3322, gm_n302, gm_n133, gm_n195, gm_n3321, gm_n392);
	nor (gm_n3323, gm_n3322, in_31);
	nand (gm_n3324, gm_n86, in_16, in_12, gm_n969, gm_n180);
	nor (gm_n3325, gm_n516, in_24, gm_n72, gm_n3324, gm_n742);
	nand (gm_n3326, gm_n207, gm_n97, gm_n78, gm_n3325);
	and (gm_n3327, gm_n180, gm_n68, in_12, gm_n613, gm_n766);
	and (gm_n3328, gm_n100, gm_n52, gm_n72, gm_n3327, gm_n517);
	nand (gm_n3329, gm_n462, gm_n205, gm_n78, gm_n3328);
	nor (gm_n3330, gm_n319, in_15, in_11, gm_n1043, gm_n399);
	nand (gm_n3331, gm_n299, gm_n195, in_19, gm_n3330, gm_n313);
	nor (gm_n3332, gm_n1118, in_31, gm_n133, gm_n3331, gm_n436);
	and (gm_n3333, gm_n118, in_15, in_8, gm_n1907, gm_n346);
	nand (gm_n3334, gm_n165, in_23, gm_n102, gm_n3333, gm_n299);
	nor (gm_n3335, gm_n1231, gm_n50, gm_n133, gm_n3334, gm_n611);
	or (gm_n3336, gm_n119, in_15, gm_n58, gm_n2463, gm_n622);
	nor (gm_n3337, gm_n337, in_23, gm_n102, gm_n3336, gm_n363);
	nand (gm_n3338, gm_n302, gm_n50, in_27, gm_n3337, gm_n306);
	nand (gm_n3339, gm_n629, gm_n68, gm_n157, gm_n1816, gm_n232);
	nor (gm_n3340, gm_n561, in_24, gm_n72, gm_n3339, gm_n602);
	nand (gm_n3341, gm_n492, gm_n99, gm_n78, gm_n3340);
	nor (gm_n3342, gm_n244, in_16, in_12, gm_n2053, gm_n286);
	nand (gm_n3343, gm_n237, gm_n52, gm_n72, gm_n3342, gm_n220);
	or (gm_n3344, gm_n371, gm_n218, in_28, gm_n3343);
	nand (gm_n3345, gm_n766, gm_n68, gm_n157, gm_n1361, gm_n341);
	nor (gm_n3346, gm_n84, in_24, in_20, gm_n3345, gm_n742);
	nand (gm_n3347, gm_n474, gm_n79, gm_n78, gm_n3346);
	nor (gm_n3348, gm_n88, gm_n157, in_8, gm_n733, gm_n385);
	nand (gm_n3349, gm_n189, gm_n72, in_16, gm_n3348, gm_n517);
	nor (gm_n3350, gm_n208, gm_n78, in_24, gm_n3349, gm_n561);
	nand (gm_n3351, gm_n3350, gm_n205);
	nand (gm_n3352, gm_n3344, gm_n3341, gm_n3338, gm_n3351, gm_n3347);
	nor (gm_n3353, gm_n127, in_23, in_19, gm_n1457, gm_n453);
	nand (gm_n3354, gm_n339, gm_n50, in_27, gm_n3353, gm_n393);
	and (gm_n3355, gm_n341, gm_n582, in_15, gm_n1715, gm_n938);
	nand (gm_n3356, gm_n302, gm_n195, in_19, gm_n3355, gm_n313);
	or (gm_n3357, gm_n51, in_31, in_27, gm_n3356);
	nand (gm_n3358, gm_n189, gm_n68, gm_n157, gm_n557, gm_n354);
	nor (gm_n3359, gm_n156, in_24, gm_n72, gm_n3358, gm_n804);
	nand (gm_n3360, gm_n492, gm_n462, in_28, gm_n3359);
	nand (gm_n3361, gm_n3360, gm_n3357, gm_n3354);
	nand (gm_n3362, gm_n85, gm_n72, gm_n68, gm_n3295, gm_n198);
	nor (gm_n3363, gm_n628, gm_n78, gm_n52, gm_n3362, gm_n780);
	nand (gm_n3364, gm_n3363, gm_n194);
	nor (gm_n3365, gm_n106, in_12, in_8, gm_n1533, gm_n107);
	nand (gm_n3366, gm_n196, in_20, gm_n68, gm_n3365, gm_n517);
	or (gm_n3367, gm_n243, in_28, gm_n52, gm_n3366, gm_n206);
	nor (gm_n3368, gm_n107, gm_n157, in_8, gm_n254, gm_n246);
	nand (gm_n3369, gm_n766, in_20, gm_n68, gm_n3368, gm_n472);
	nor (gm_n3370, gm_n804, gm_n78, gm_n52, gm_n3369, gm_n208);
	nand (gm_n3371, gm_n3370, gm_n186);
	nand (gm_n3372, gm_n3371, gm_n3367, gm_n3364);
	nor (gm_n3373, gm_n3352, gm_n3335, gm_n3332, gm_n3372, gm_n3361);
	nor (gm_n3374, gm_n119, gm_n105, in_11, gm_n1627, gm_n622);
	nand (gm_n3375, gm_n582, in_23, in_19, gm_n3374, gm_n293);
	nor (gm_n3376, gm_n174, gm_n50, gm_n133, gm_n3375, gm_n611);
	nand (gm_n3377, gm_n100, in_24, in_20, gm_n1855, gm_n517);
	nor (gm_n3378, gm_n206, gm_n243, in_28, gm_n3377);
	nand (gm_n3379, gm_n180, gm_n157, gm_n64, gm_n281, gm_n110);
	nor (gm_n3380, gm_n244, in_20, in_16, gm_n3379, gm_n178);
	nand (gm_n3381, gm_n177, gm_n78, in_24, gm_n3380, gm_n196);
	nor (gm_n3382, gm_n3381, gm_n176);
	nor (gm_n3383, gm_n3382, gm_n3378, gm_n3376);
	nor (gm_n3384, gm_n672, gm_n105, gm_n58, gm_n1356, gm_n319);
	nand (gm_n3385, gm_n165, gm_n195, in_19, gm_n3384, gm_n394);
	nor (gm_n3386, gm_n51, in_31, in_27, gm_n3385, gm_n983);
	nor (gm_n3387, gm_n107, in_16, in_12, gm_n979, gm_n158);
	nand (gm_n3388, gm_n209, gm_n52, in_20, gm_n3387, gm_n269);
	nor (gm_n3389, gm_n780, gm_n206, in_28, gm_n3388);
	nand (gm_n3390, gm_n567, gm_n140, in_8);
	nor (gm_n3391, gm_n244, gm_n68, gm_n157, gm_n3390, gm_n107);
	nand (gm_n3392, gm_n83, in_24, in_20, gm_n3391, gm_n269);
	nor (gm_n3393, gm_n206, gm_n216, in_28, gm_n3392);
	nor (gm_n3394, gm_n3393, gm_n3389, gm_n3386);
	nand (gm_n3395, gm_n3373, gm_n3329, gm_n3326, gm_n3394, gm_n3383);
	nor (gm_n3396, gm_n618, gm_n105, gm_n58, gm_n1266, gm_n426);
	nand (gm_n3397, gm_n361, in_23, in_19, gm_n3396, gm_n452);
	or (gm_n3398, gm_n54, in_31, gm_n133, gm_n3397, gm_n575);
	nor (gm_n3399, gm_n366, gm_n102, in_15, gm_n2272, gm_n911);
	and (gm_n3400, gm_n313, in_27, gm_n195, gm_n3399, gm_n455);
	nand (gm_n3401, gm_n3400, gm_n508, gm_n50);
	or (gm_n3402, gm_n88, gm_n68, in_12, gm_n1294, gm_n179);
	nor (gm_n3403, gm_n84, gm_n52, gm_n72, gm_n3402, gm_n459);
	nand (gm_n3404, gm_n462, gm_n217, gm_n78, gm_n3403);
	nand (gm_n3405, gm_n3404, gm_n3401, gm_n3398);
	and (gm_n3406, gm_n210, gm_n157, in_8, gm_n450, gm_n180);
	nand (gm_n3407, gm_n321, in_17, in_13, gm_n3406, gm_n526);
	nor (gm_n3408, gm_n535, in_25, gm_n81, gm_n3407, gm_n2015);
	nand (gm_n3409, in_31, in_30, in_29, gm_n3408);
	or (gm_n3410, gm_n107, in_16, in_12, gm_n1064, gm_n168);
	nor (gm_n3411, gm_n187, in_24, in_20, gm_n3410, gm_n628);
	nand (gm_n3412, gm_n177, gm_n194, in_28, gm_n3411);
	nand (gm_n3413, gm_n818, in_15, in_11, gm_n1758, gm_n425);
	nor (gm_n3414, gm_n300, in_23, in_19, gm_n3413, gm_n510);
	nand (gm_n3415, gm_n302, gm_n50, gm_n133, gm_n3414, gm_n339);
	nand (gm_n3416, gm_n3415, gm_n3412, gm_n3409);
	nor (gm_n3417, gm_n3395, gm_n3323, gm_n3319, gm_n3416, gm_n3405);
	nor (gm_n3418, gm_n426, in_15, in_11, gm_n880, gm_n666);
	nand (gm_n3419, gm_n299, gm_n195, gm_n102, gm_n3418, gm_n361);
	nor (gm_n3420, gm_n303, in_31, gm_n133, gm_n3419, gm_n617);
	nor (gm_n3421, gm_n107, gm_n68, in_12, gm_n2128, gm_n158);
	nand (gm_n3422, gm_n83, in_24, gm_n72, gm_n3421, gm_n269);
	nor (gm_n3423, gm_n687, gm_n208, in_28, gm_n3422);
	nand (gm_n3424, gm_n110, gm_n157, gm_n64, gm_n403, gm_n232);
	nor (gm_n3425, gm_n221, in_20, in_16, gm_n3424, gm_n459);
	nand (gm_n3426, gm_n83, in_28, gm_n52, gm_n3425, gm_n259);
	nor (gm_n3427, gm_n3426, gm_n218);
	nor (gm_n3428, gm_n3427, gm_n3423, gm_n3420);
	nand (gm_n3429, gm_n270, in_12, gm_n64, gm_n567, gm_n511);
	nor (gm_n3430, gm_n168, gm_n72, in_16, gm_n3429, gm_n459);
	nand (gm_n3431, gm_n252, in_28, gm_n52, gm_n3430, gm_n462);
	nor (gm_n3432, gm_n3431, gm_n475);
	nor (gm_n3433, gm_n88, in_16, gm_n157, gm_n2124, gm_n139);
	nand (gm_n3434, gm_n237, gm_n52, in_20, gm_n3433, gm_n252);
	nor (gm_n3435, gm_n371, gm_n229, gm_n78, gm_n3434);
	nor (gm_n3436, gm_n504, gm_n157, in_8, gm_n1533, gm_n222);
	nand (gm_n3437, gm_n237, gm_n72, in_16, gm_n3436, gm_n252);
	nor (gm_n3438, gm_n229, in_28, gm_n52, gm_n3437, gm_n371);
	nor (gm_n3439, gm_n3438, gm_n3435, gm_n3432);
	nand (gm_n3440, gm_n3417, gm_n3316, gm_n3313, gm_n3439, gm_n3428);
	and (gm_n3441, gm_n146, gm_n68, in_12, gm_n2970, gm_n341);
	nand (gm_n3442, gm_n220, in_24, in_20, gm_n3441, gm_n230);
	nor (gm_n3443, gm_n371, gm_n132, in_28, gm_n3442);
	nand (gm_n3444, gm_n263, gm_n110, in_8);
	nor (gm_n3445, gm_n106, in_16, in_12, gm_n3444, gm_n167);
	nand (gm_n3446, gm_n100, gm_n52, in_20, gm_n3445, gm_n219);
	nor (gm_n3447, gm_n371, gm_n268, gm_n78, gm_n3446);
	and (gm_n3448, gm_n333, in_15, gm_n58, gm_n797, gm_n120);
	and (gm_n3449, gm_n313, gm_n195, in_19, gm_n3448, gm_n362);
	and (gm_n3450, gm_n129, gm_n50, gm_n133, gm_n3449, gm_n339);
	nor (gm_n3451, gm_n3450, gm_n3447, gm_n3443);
	not (gm_n3452, gm_n3451);
	nor (gm_n3453, gm_n672, gm_n105, in_11, gm_n433, gm_n673);
	and (gm_n3454, gm_n582, gm_n195, gm_n102, gm_n3453, gm_n509);
	and (gm_n3455, gm_n55, in_31, gm_n133, gm_n3454, gm_n677);
	and (gm_n3456, gm_n118, in_15, gm_n58, gm_n2149, gm_n297);
	nand (gm_n3457, gm_n126, in_23, gm_n102, gm_n3456, gm_n394);
	nor (gm_n3458, gm_n174, gm_n50, in_27, gm_n3457, gm_n575);
	nor (gm_n3459, gm_n159, gm_n68, in_12, gm_n2804, gm_n168);
	nand (gm_n3460, gm_n209, in_24, gm_n72, gm_n3459, gm_n472);
	nor (gm_n3461, gm_n371, gm_n229, in_28, gm_n3460);
	nor (gm_n3462, gm_n3461, gm_n3458, gm_n3455);
	not (gm_n3463, gm_n3462);
	or (gm_n3464, gm_n3440, gm_n3307, gm_n3304, gm_n3463, gm_n3452);
	nand (gm_n3465, gm_n263, gm_n140, gm_n64);
	nor (gm_n3466, gm_n244, in_16, gm_n157, gm_n3465, gm_n167);
	and (gm_n3467, gm_n83, in_24, in_20, gm_n3466, gm_n269);
	and (gm_n3468, gm_n370, gm_n97, gm_n78, gm_n3467);
	nor (gm_n3469, gm_n168, gm_n68, in_12, gm_n3141, gm_n222);
	nand (gm_n3470, gm_n100, gm_n52, gm_n72, gm_n3469, gm_n230);
	nor (gm_n3471, gm_n243, gm_n229, gm_n78, gm_n3470);
	nor (gm_n3472, gm_n244, in_16, gm_n157, gm_n2060, gm_n286);
	and (gm_n3473, gm_n209, gm_n52, in_20, gm_n3472, gm_n517);
	and (gm_n3474, gm_n259, gm_n194, gm_n78, gm_n3473);
	or (gm_n3475, gm_n3468, gm_n3464, gm_n3301, gm_n3474, gm_n3471);
	nor (gm_n3476, gm_n618, gm_n105, in_11, gm_n997, gm_n667);
	and (gm_n3477, gm_n73, gm_n195, gm_n102, gm_n3476, gm_n166);
	and (gm_n3478, gm_n302, gm_n50, gm_n133, gm_n3477, gm_n306);
	nor (new_out3, gm_n3475, gm_n3298, gm_n3294, gm_n3478);
	or (gm_n3480, new_out3, new_out2);
	or (gm_n3481, gm_n300, gm_n222, in_15, gm_n622, gm_n577);
	nor (gm_n3482, gm_n617, in_23, in_19, gm_n3481, gm_n431);
	and (gm_n3483, gm_n508, in_31, gm_n133, gm_n3482);
	nand (gm_n3484, gm_n87, in_9, gm_n64, gm_n705, gm_n122);
	or (gm_n3485, gm_n117, gm_n105, gm_n58, gm_n3484, gm_n576);
	nor (gm_n3486, gm_n423, gm_n195, gm_n102, gm_n3485, gm_n671);
	nand (gm_n3487, gm_n392, gm_n50, in_27, gm_n3486);
	nand (gm_n3488, gm_n189, in_16, gm_n157, gm_n2336, gm_n232);
	nor (gm_n3489, gm_n178, in_24, gm_n72, gm_n3488, gm_n561);
	nand (gm_n3490, gm_n194, gm_n79, gm_n78, gm_n3489);
	nor (gm_n3491, gm_n426, gm_n105, gm_n58, gm_n701, gm_n666);
	nand (gm_n3492, gm_n166, in_23, gm_n102, gm_n3491, gm_n313);
	nor (gm_n3493, gm_n1231, in_31, gm_n133, gm_n3492, gm_n611);
	not (gm_n3494, gm_n152);
	nand (gm_n3495, gm_n72, in_19, gm_n136);
	nor (gm_n3496, gm_n529, gm_n81, in_17, gm_n3495, gm_n1684);
	nand (gm_n3497, gm_n3494, in_29, gm_n53, gm_n3496, gm_n1686);
	nor (gm_n3498, gm_n3497, gm_n50, gm_n96);
	nand (gm_n3499, gm_n188, gm_n68, gm_n157, gm_n212, gm_n198);
	nor (gm_n3500, gm_n804, gm_n52, in_20, gm_n3499, gm_n413);
	nand (gm_n3501, gm_n462, gm_n186, gm_n78, gm_n3500);
	nor (gm_n3502, gm_n139, in_16, in_12, gm_n906, gm_n167);
	and (gm_n3503, gm_n196, in_24, gm_n72, gm_n3502, gm_n472);
	nand (gm_n3504, gm_n370, gm_n217, in_28, gm_n3503);
	nor (gm_n3505, gm_n672, in_15, in_11, gm_n1406, gm_n673);
	nand (gm_n3506, gm_n313, gm_n195, gm_n102, gm_n3505, gm_n612);
	nor (gm_n3507, gm_n1118, gm_n50, in_27, gm_n3506, gm_n842);
	and (gm_n3508, gm_n766, gm_n68, gm_n157, gm_n2527, gm_n341);
	nand (gm_n3509, gm_n220, in_24, in_20, gm_n3508, gm_n269);
	nor (gm_n3510, gm_n268, gm_n243, gm_n78, gm_n3509);
	nand (gm_n3511, gm_n180, in_16, gm_n157, gm_n1106, gm_n766);
	nor (gm_n3512, gm_n197, gm_n52, in_20, gm_n3511, gm_n459);
	nand (gm_n3513, gm_n370, gm_n97, gm_n78, gm_n3512);
	nand (gm_n3514, gm_n189, gm_n68, in_12, gm_n2580, gm_n180);
	nor (gm_n3515, gm_n187, gm_n52, gm_n72, gm_n3514, gm_n101);
	nand (gm_n3516, gm_n492, gm_n462, in_28, gm_n3515);
	nor (gm_n3517, gm_n504, in_16, in_12, gm_n906, gm_n286);
	nand (gm_n3518, gm_n100, gm_n52, gm_n72, gm_n3517, gm_n517);
	nor (gm_n3519, gm_n687, gm_n135, in_28, gm_n3518);
	and (gm_n3520, gm_n452, gm_n341, gm_n105, gm_n1715, gm_n621);
	nand (gm_n3521, gm_n165, gm_n195, gm_n102, gm_n3520, gm_n173);
	nor (gm_n3522, gm_n303, gm_n50, in_27, gm_n3521);
	nor (gm_n3523, gm_n319, gm_n105, gm_n58, gm_n433, gm_n399);
	nand (gm_n3524, gm_n73, gm_n195, gm_n102, gm_n3523, gm_n452);
	nor (gm_n3525, gm_n1118, gm_n50, gm_n133, gm_n3524, gm_n678);
	nor (gm_n3526, gm_n106, gm_n68, gm_n157, gm_n960, gm_n253);
	nand (gm_n3527, gm_n220, gm_n52, gm_n72, gm_n3526, gm_n517);
	nor (gm_n3528, gm_n218, gm_n208, gm_n78, gm_n3527);
	nor (gm_n3529, gm_n179, gm_n68, gm_n157, gm_n286, gm_n247);
	nand (gm_n3530, gm_n209, gm_n52, in_20, gm_n3529, gm_n269);
	nor (gm_n3531, gm_n216, gm_n229, gm_n78, gm_n3530);
	nor (gm_n3532, gm_n3525, gm_n3522, gm_n3519, gm_n3531, gm_n3528);
	and (gm_n3533, gm_n297, in_15, gm_n58, gm_n1802, gm_n938);
	nand (gm_n3534, gm_n582, gm_n195, gm_n102, gm_n3533, gm_n126);
	nor (gm_n3535, gm_n51, in_31, in_27, gm_n3534, gm_n983);
	and (gm_n3536, gm_n118, gm_n105, in_11, gm_n1102, gm_n665);
	nand (gm_n3537, gm_n361, gm_n195, in_19, gm_n3536, gm_n362);
	nor (gm_n3538, gm_n611, gm_n50, gm_n133, gm_n3537, gm_n983);
	nand (gm_n3539, gm_n587, gm_n122);
	nor (gm_n3540, gm_n396, gm_n105, gm_n58, gm_n3539, gm_n622);
	nand (gm_n3541, gm_n126, in_23, in_19, gm_n3540, gm_n299);
	nor (gm_n3542, gm_n51, gm_n50, in_27, gm_n3541, gm_n617);
	nor (gm_n3543, gm_n3542, gm_n3538, gm_n3535);
	and (gm_n3544, gm_n705, gm_n122, in_8);
	and (gm_n3545, gm_n270, in_16, in_12, gm_n3544, gm_n629);
	nand (gm_n3546, gm_n183, gm_n52, gm_n72, gm_n3545, gm_n472);
	nor (gm_n3547, gm_n216, gm_n176, gm_n78, gm_n3546);
	and (gm_n3548, gm_n180, in_16, in_12, gm_n563, gm_n138);
	nand (gm_n3549, gm_n196, gm_n52, gm_n72, gm_n3548, gm_n472);
	nor (gm_n3550, gm_n208, gm_n229, gm_n78, gm_n3549);
	nor (gm_n3551, gm_n88, in_16, in_12, gm_n2499, gm_n158);
	nand (gm_n3552, gm_n209, in_24, gm_n72, gm_n3551, gm_n472);
	nor (gm_n3553, gm_n371, gm_n176, gm_n78, gm_n3552);
	nor (gm_n3554, gm_n3553, gm_n3550, gm_n3547);
	nand (gm_n3555, gm_n3532, gm_n3516, gm_n3513, gm_n3554, gm_n3543);
	nor (gm_n3556, gm_n57, gm_n105, in_11, gm_n1259, gm_n119);
	nand (gm_n3557, gm_n73, in_23, gm_n102, gm_n3556, gm_n612);
	or (gm_n3558, gm_n174, in_31, in_27, gm_n3557, gm_n303);
	nand (gm_n3559, gm_n189, gm_n68, gm_n157, gm_n630, gm_n270);
	nor (gm_n3560, gm_n156, gm_n52, gm_n72, gm_n3559, gm_n804);
	nand (gm_n3561, gm_n177, gm_n194, in_28, gm_n3560);
	nor (gm_n3562, gm_n158, gm_n68, gm_n157, gm_n1303, gm_n245);
	nand (gm_n3563, gm_n100, in_24, gm_n72, gm_n3562, gm_n269);
	or (gm_n3564, gm_n780, gm_n218, in_28, gm_n3563);
	nand (gm_n3565, gm_n3564, gm_n3561, gm_n3558);
	nand (gm_n3566, gm_n231, gm_n72, gm_n68, gm_n1094, gm_n517);
	nor (gm_n3567, gm_n197, in_28, gm_n52, gm_n3566, gm_n208);
	nand (gm_n3568, gm_n3567, gm_n186);
	nand (gm_n3569, gm_n180, in_16, gm_n157, gm_n1173, gm_n146);
	nor (gm_n3570, gm_n84, gm_n52, gm_n72, gm_n3569, gm_n103);
	nand (gm_n3571, gm_n492, gm_n79, in_28, gm_n3570);
	nor (gm_n3572, gm_n504, gm_n68, gm_n157, gm_n3118, gm_n159);
	and (gm_n3573, gm_n137, in_24, in_20, gm_n3572, gm_n261);
	nand (gm_n3574, gm_n370, gm_n97, gm_n78, gm_n3573);
	nand (gm_n3575, gm_n3574, gm_n3571, gm_n3568);
	nor (gm_n3576, gm_n3555, gm_n3510, gm_n3507, gm_n3575, gm_n3565);
	nor (gm_n3577, gm_n57, gm_n105, in_11, gm_n1946, gm_n727);
	nand (gm_n3578, gm_n293, in_23, in_19, gm_n3577, gm_n362);
	nor (gm_n3579, gm_n1231, gm_n50, in_27, gm_n3578, gm_n303);
	nor (gm_n3580, gm_n366, gm_n105, gm_n58, gm_n1356, gm_n396);
	nand (gm_n3581, gm_n299, in_23, in_19, gm_n3580, gm_n509);
	nor (gm_n3582, gm_n581, gm_n50, gm_n133, gm_n3581, gm_n436);
	or (gm_n3583, in_12, in_8, in_7, gm_n530, gm_n167);
	nor (gm_n3584, gm_n139, in_20, gm_n68, gm_n3583, gm_n459);
	nand (gm_n3585, gm_n99, gm_n78, gm_n52, gm_n3584, gm_n220);
	nor (gm_n3586, gm_n3585, gm_n687);
	nor (gm_n3587, gm_n3586, gm_n3582, gm_n3579);
	and (gm_n3588, gm_n146, in_16, in_12, gm_n872, gm_n270);
	nand (gm_n3589, gm_n252, in_24, gm_n72, gm_n3588, gm_n517);
	nor (gm_n3590, gm_n80, gm_n229, gm_n78, gm_n3589);
	or (gm_n3591, gm_n246, gm_n157, in_8, gm_n286, gm_n224);
	nor (gm_n3592, gm_n106, in_20, gm_n68, gm_n3591, gm_n459);
	nand (gm_n3593, gm_n100, in_28, gm_n52, gm_n3592, gm_n134);
	nor (gm_n3594, gm_n3593, gm_n176);
	nor (gm_n3595, gm_n221, in_20, in_16, gm_n2841, gm_n413);
	nand (gm_n3596, gm_n209, in_28, in_24, gm_n3595, gm_n370);
	nor (gm_n3597, gm_n3596, gm_n268);
	nor (gm_n3598, gm_n3597, gm_n3594, gm_n3590);
	nand (gm_n3599, gm_n3576, gm_n3504, gm_n3501, gm_n3598, gm_n3587);
	or (gm_n3600, gm_n244, gm_n68, gm_n157, gm_n2039, gm_n245);
	nor (gm_n3601, gm_n804, gm_n52, in_20, gm_n3600, gm_n413);
	nand (gm_n3602, gm_n79, gm_n77, gm_n78, gm_n3601);
	nor (gm_n3603, gm_n300, in_23, gm_n102, gm_n3278, gm_n337);
	nand (gm_n3604, gm_n307, gm_n50, gm_n133, gm_n3603, gm_n392);
	nand (gm_n3605, gm_n629, in_16, in_12, gm_n3544, gm_n354);
	nor (gm_n3606, gm_n101, gm_n52, in_20, gm_n3605, gm_n459);
	nand (gm_n3607, gm_n462, gm_n205, gm_n78, gm_n3606);
	nand (gm_n3608, gm_n3607, gm_n3604, gm_n3602);
	nand (gm_n3609, gm_n198, in_16, in_12, gm_n2970, gm_n354);
	nor (gm_n3610, gm_n84, in_24, gm_n72, gm_n3609, gm_n156);
	nand (gm_n3611, gm_n134, gm_n194, in_28, gm_n3610);
	nor (gm_n3612, gm_n139, in_16, gm_n157, gm_n1123, gm_n222);
	nand (gm_n3613, gm_n220, in_24, in_20, gm_n3612, gm_n517);
	or (gm_n3614, gm_n135, gm_n132, gm_n78, gm_n3613);
	nor (gm_n3615, gm_n142, gm_n105, gm_n58, gm_n997, gm_n396);
	and (gm_n3616, gm_n166, in_23, gm_n102, gm_n3615, gm_n361);
	nand (gm_n3617, gm_n455, in_31, gm_n133, gm_n3616, gm_n677);
	nand (gm_n3618, gm_n3617, gm_n3614, gm_n3611);
	nor (gm_n3619, gm_n3599, gm_n3498, gm_n3493, gm_n3618, gm_n3608);
	nand (gm_n3620, gm_n354, in_12, gm_n64, gm_n308, gm_n263);
	nor (gm_n3621, gm_n179, gm_n72, gm_n68, gm_n3620, gm_n742);
	nand (gm_n3622, gm_n79, in_28, in_24, gm_n3621, gm_n100);
	nor (gm_n3623, gm_n3622, gm_n176);
	nor (gm_n3624, gm_n576, gm_n167, gm_n105, gm_n2077, gm_n911);
	nand (gm_n3625, gm_n55, in_23, in_19, gm_n3624, gm_n126);
	nor (gm_n3626, gm_n575, gm_n50, in_27, gm_n3625);
	nand (gm_n3627, gm_n511, gm_n397, in_8);
	nor (gm_n3628, gm_n504, in_16, in_12, gm_n3627, gm_n167);
	nand (gm_n3629, gm_n83, in_24, gm_n72, gm_n3628, gm_n517);
	nor (gm_n3630, gm_n475, gm_n260, gm_n78, gm_n3629);
	nor (gm_n3631, gm_n3630, gm_n3626, gm_n3623);
	nor (gm_n3632, gm_n504, in_16, in_12, gm_n245, gm_n161);
	nand (gm_n3633, gm_n196, gm_n52, gm_n72, gm_n3632, gm_n230);
	nor (gm_n3634, gm_n475, gm_n260, in_28, gm_n3633);
	nor (gm_n3635, gm_n117, gm_n102, in_15, gm_n2170, gm_n672);
	nand (gm_n3636, gm_n293, gm_n133, in_23, gm_n3635, gm_n307);
	nor (gm_n3637, gm_n3636, gm_n360, gm_n50);
	nor (gm_n3638, gm_n139, gm_n68, gm_n157, gm_n588, gm_n222);
	nand (gm_n3639, gm_n220, gm_n52, gm_n72, gm_n3638, gm_n472);
	nor (gm_n3640, gm_n208, gm_n132, gm_n78, gm_n3639);
	nor (gm_n3641, gm_n3640, gm_n3637, gm_n3634);
	nand (gm_n3642, gm_n3619, gm_n3490, gm_n3487, gm_n3641, gm_n3631);
	nor (gm_n3643, gm_n319, in_15, in_11, gm_n1043, gm_n622);
	and (gm_n3644, gm_n73, gm_n195, in_19, gm_n3643, gm_n166);
	and (gm_n3645, gm_n302, in_31, in_27, gm_n3644, gm_n677);
	nand (gm_n3646, gm_n747, gm_n63, in_8);
	nor (gm_n3647, gm_n504, gm_n68, in_12, gm_n3646, gm_n159);
	nand (gm_n3648, gm_n83, in_24, in_20, gm_n3647, gm_n219);
	nor (gm_n3649, gm_n135, gm_n132, gm_n78, gm_n3648);
	and (gm_n3650, gm_n180, gm_n68, gm_n157, gm_n2144, gm_n138);
	nand (gm_n3651, gm_n230, in_24, gm_n72, gm_n3650, gm_n261);
	nor (gm_n3652, gm_n218, gm_n135, in_28, gm_n3651);
	or (gm_n3653, gm_n3645, gm_n3642, gm_n3483, gm_n3652, gm_n3649);
	nor (gm_n3654, gm_n396, gm_n105, gm_n58, gm_n2504, gm_n426);
	and (gm_n3655, gm_n73, in_23, gm_n102, gm_n3654, gm_n582);
	and (gm_n3656, gm_n129, gm_n50, gm_n133, gm_n3655, gm_n677);
	nor (gm_n3657, gm_n179, gm_n68, in_12, gm_n1737, gm_n245);
	nand (gm_n3658, gm_n209, gm_n52, in_20, gm_n3657, gm_n517);
	nor (gm_n3659, gm_n475, gm_n208, in_28, gm_n3658);
	nor (gm_n3660, gm_n168, gm_n68, gm_n157, gm_n253, gm_n247);
	and (gm_n3661, gm_n196, in_24, in_20, gm_n3660, gm_n517);
	and (gm_n3662, gm_n462, gm_n217, in_28, gm_n3661);
	and (gm_n3663, gm_n138, in_16, gm_n157, gm_n1437, gm_n346);
	and (gm_n3664, gm_n85, in_24, in_20, gm_n3663, gm_n100);
	and (gm_n3665, gm_n474, gm_n462, gm_n78, gm_n3664);
	nor (gm_n3666, gm_n504, in_16, in_12, gm_n1525, gm_n286);
	nand (gm_n3667, gm_n83, in_24, gm_n72, gm_n3666, gm_n137);
	nor (gm_n3668, gm_n475, gm_n260, in_28, gm_n3667);
	nor (gm_n3669, gm_n319, gm_n105, gm_n58, gm_n2081, gm_n366);
	nand (gm_n3670, gm_n582, gm_n195, in_19, gm_n3669, gm_n509);
	nor (gm_n3671, gm_n360, in_31, in_27, gm_n3670, gm_n617);
	nor (gm_n3672, gm_n363, gm_n102, gm_n105, gm_n1631, gm_n997);
	and (gm_n3673, gm_n55, in_27, gm_n195, gm_n3672, gm_n336);
	nand (gm_n3674, gm_n3673, gm_n437, gm_n50);
	or (gm_n3675, gm_n57, gm_n105, gm_n58, gm_n2693, gm_n119);
	nor (gm_n3676, gm_n423, in_23, gm_n102, gm_n3675, gm_n300);
	nand (gm_n3677, gm_n115, gm_n50, gm_n133, gm_n3676, gm_n658);
	or (gm_n3678, gm_n396, gm_n105, in_11, gm_n2697, gm_n997);
	or (gm_n3679, gm_n127, in_23, in_19, gm_n3678, gm_n332);
	nor (gm_n3680, gm_n1118, gm_n50, gm_n133, gm_n3679, gm_n842);
	and (gm_n3681, gm_n63, in_12, gm_n64, gm_n397, gm_n188);
	and (gm_n3682, gm_n137, gm_n72, gm_n68, gm_n3681, gm_n146);
	and (gm_n3683, gm_n99, in_28, in_24, gm_n3682, gm_n196);
	and (gm_n3684, gm_n3683, gm_n205);
	nand (gm_n3685, gm_n231, in_16, in_12, gm_n233, gm_n270);
	or (gm_n3686, gm_n84, in_24, in_20, gm_n3685, gm_n742);
	nor (gm_n3687, gm_n260, gm_n132, in_28, gm_n3686);
	or (gm_n3688, gm_n244, gm_n72, in_16, gm_n2638, gm_n459);
	or (gm_n3689, gm_n208, in_28, in_24, gm_n3688, gm_n412);
	nor (gm_n3690, gm_n3689, gm_n229);
	nor (gm_n3691, gm_n106, in_16, gm_n157, gm_n1325, gm_n222);
	nand (gm_n3692, gm_n196, gm_n52, in_20, gm_n3691, gm_n472);
	nor (gm_n3693, gm_n475, gm_n80, in_28, gm_n3692);
	or (gm_n3694, gm_n57, in_15, gm_n58, gm_n2693, gm_n432);
	or (gm_n3695, gm_n1703, in_23, gm_n102, gm_n3694, gm_n911);
	nor (gm_n3696, gm_n51, gm_n50, gm_n133, gm_n3695, gm_n1118);
	or (gm_n3697, gm_n168, in_16, in_12, gm_n3627, gm_n245);
	or (gm_n3698, gm_n412, gm_n52, gm_n72, gm_n3697, gm_n413);
	nor (gm_n3699, gm_n135, gm_n229, in_28, gm_n3698);
	nor (gm_n3700, gm_n107, gm_n68, in_12, gm_n1385, gm_n168);
	nand (gm_n3701, gm_n85, gm_n52, gm_n72, gm_n3700, gm_n196);
	nor (gm_n3702, gm_n208, gm_n176, in_28, gm_n3701);
	or (gm_n3703, gm_n159, gm_n68, gm_n157, gm_n808, gm_n179);
	or (gm_n3704, gm_n101, in_24, in_20, gm_n3703, gm_n459);
	nor (gm_n3705, gm_n371, gm_n268, in_28, gm_n3704);
	or (gm_n3706, gm_n3699, gm_n3696, gm_n3693, gm_n3705, gm_n3702);
	or (gm_n3707, gm_n221, gm_n68, in_12, gm_n3444, gm_n222);
	or (gm_n3708, gm_n187, in_24, in_20, gm_n3707, gm_n197);
	nor (gm_n3709, gm_n687, gm_n208, in_28, gm_n3708);
	nor (gm_n3710, gm_n562, gm_n157, gm_n64, gm_n1200, gm_n159);
	nand (gm_n3711, gm_n189, in_20, gm_n68, gm_n3710, gm_n137);
	or (gm_n3712, gm_n804, in_28, gm_n52, gm_n3711, gm_n371);
	nor (gm_n3713, gm_n3712, gm_n475);
	and (gm_n3714, gm_n66, in_15, gm_n58, gm_n1802, gm_n311);
	nand (gm_n3715, gm_n293, gm_n195, gm_n102, gm_n3714, gm_n452);
	nor (gm_n3716, gm_n51, in_31, in_27, gm_n3715, gm_n617);
	or (gm_n3717, gm_n3716, gm_n3713, gm_n3709);
	and (gm_n3718, gm_n118, gm_n105, in_11, gm_n1802, gm_n297);
	nand (gm_n3719, gm_n73, in_23, gm_n102, gm_n3718, gm_n362);
	nor (gm_n3720, gm_n617, in_31, gm_n133, gm_n3719, gm_n678);
	nor (gm_n3721, gm_n106, in_16, gm_n157, gm_n372, gm_n159);
	nand (gm_n3722, gm_n230, gm_n52, in_20, gm_n3721, gm_n252);
	nor (gm_n3723, gm_n260, gm_n176, in_28, gm_n3722);
	nor (gm_n3724, gm_n159, gm_n68, in_12, gm_n381, gm_n168);
	nand (gm_n3725, gm_n83, in_24, in_20, gm_n3724, gm_n137);
	nor (gm_n3726, gm_n687, gm_n243, in_28, gm_n3725);
	or (gm_n3727, gm_n3726, gm_n3723, gm_n3720);
	or (gm_n3728, gm_n3706, gm_n3690, gm_n3687, gm_n3727, gm_n3717);
	nor (gm_n3729, gm_n244, gm_n68, gm_n157, gm_n1839, gm_n286);
	nand (gm_n3730, gm_n100, in_24, in_20, gm_n3729, gm_n237);
	nor (gm_n3731, gm_n135, gm_n132, gm_n78, gm_n3730);
	or (gm_n3732, gm_n319, in_15, in_11, gm_n3539, gm_n622);
	or (gm_n3733, gm_n300, gm_n195, in_19, gm_n3732, gm_n431);
	nor (gm_n3734, gm_n51, in_31, gm_n133, gm_n3733, gm_n1231);
	nand (gm_n3735, gm_n189, in_16, gm_n157, gm_n1846, gm_n341);
	or (gm_n3736, gm_n101, gm_n52, in_20, gm_n3735, gm_n459);
	nor (gm_n3737, gm_n208, gm_n229, in_28, gm_n3736);
	or (gm_n3738, gm_n3737, gm_n3734, gm_n3731);
	or (gm_n3739, gm_n673, gm_n105, gm_n58, gm_n1086, gm_n399);
	or (gm_n3740, gm_n300, in_23, in_19, gm_n3739, gm_n431);
	nor (gm_n3741, gm_n174, in_31, gm_n133, gm_n3740, gm_n842);
	nand (gm_n3742, gm_n346, gm_n582, in_15, gm_n758, gm_n938);
	or (gm_n3743, gm_n127, gm_n195, gm_n102, gm_n3742, gm_n174);
	nor (gm_n3744, gm_n303, gm_n50, in_27, gm_n3743);
	or (gm_n3745, gm_n91, in_12, in_8, gm_n167, gm_n562);
	nor (gm_n3746, gm_n156, in_20, gm_n68, gm_n3745, gm_n168);
	nand (gm_n3747, gm_n252, gm_n78, in_24, gm_n3746, gm_n462);
	nor (gm_n3748, gm_n3747, gm_n229);
	or (gm_n3749, gm_n3748, gm_n3744, gm_n3741);
	nor (gm_n3750, gm_n3728, gm_n3684, gm_n3680, gm_n3749, gm_n3738);
	nand (gm_n3751, gm_n189, gm_n68, in_12, gm_n920, gm_n341);
	or (gm_n3752, gm_n156, gm_n52, in_20, gm_n3751, gm_n804);
	nor (gm_n3753, gm_n206, gm_n80, in_28, gm_n3752);
	and (gm_n3754, gm_n140, gm_n157, gm_n64, gm_n587, gm_n232);
	and (gm_n3755, gm_n189, gm_n72, in_16, gm_n3754, gm_n230);
	and (gm_n3756, gm_n220, in_28, gm_n52, gm_n3755, gm_n370);
	and (gm_n3757, gm_n3756, gm_n77);
	nand (gm_n3758, gm_n198, gm_n68, gm_n157, gm_n2336, gm_n354);
	or (gm_n3759, gm_n103, in_24, gm_n72, gm_n3758, gm_n412);
	nor (gm_n3760, gm_n268, gm_n243, gm_n78, gm_n3759);
	nor (gm_n3761, gm_n3760, gm_n3757, gm_n3753);
	or (gm_n3762, gm_n322, in_17, gm_n157, gm_n734, gm_n323);
	or (gm_n3763, gm_n152, in_25, gm_n81, gm_n3762, gm_n1054);
	nor (gm_n3764, gm_n50, in_30, gm_n76, gm_n3763);
	or (gm_n3765, gm_n396, gm_n105, gm_n58, gm_n2233, gm_n622);
	or (gm_n3766, gm_n337, gm_n195, in_19, gm_n3765, gm_n911);
	nor (gm_n3767, gm_n617, in_31, in_27, gm_n3766, gm_n842);
	nor (gm_n3768, gm_n89, gm_n157, in_8, gm_n224, gm_n159);
	and (gm_n3769, gm_n237, in_20, gm_n68, gm_n3768, gm_n138);
	and (gm_n3770, gm_n100, gm_n78, gm_n52, gm_n3769, gm_n134);
	and (gm_n3771, gm_n3770, gm_n492);
	nor (gm_n3772, gm_n3771, gm_n3767, gm_n3764);
	nand (gm_n3773, gm_n3750, gm_n3677, gm_n3674, gm_n3772, gm_n3761);
	nor (gm_n3774, in_17, gm_n68, gm_n105);
	and (gm_n3775, gm_n1996, gm_n136, gm_n104, gm_n3774, gm_n2476);
	nor (gm_n3776, gm_n81, in_20, gm_n102);
	nor (gm_n3777, gm_n53, gm_n52, in_23);
	nand (gm_n3778, gm_n3775, in_26, in_22, gm_n3777, gm_n3776);
	nand (gm_n3779, in_29, gm_n78, in_27);
	nor (gm_n3780, gm_n3778, gm_n50, gm_n96, gm_n3779);
	nor (gm_n3781, gm_n70, in_15, in_11, gm_n3484, gm_n576);
	nand (gm_n3782, gm_n361, in_23, gm_n102, gm_n3781, gm_n658);
	nor (gm_n3783, gm_n575, in_31, gm_n133, gm_n3782);
	nand (gm_n3784, gm_n309, gm_n63, gm_n64);
	nor (gm_n3785, gm_n106, gm_n68, gm_n157, gm_n3784, gm_n286);
	nand (gm_n3786, gm_n83, in_24, gm_n72, gm_n3785, gm_n137);
	nor (gm_n3787, gm_n208, gm_n176, gm_n78, gm_n3786);
	or (gm_n3788, gm_n3780, gm_n3773, gm_n3671, gm_n3787, gm_n3783);
	or (gm_n3789, in_10, gm_n121, gm_n62, gm_n1995, gm_n355);
	nor (gm_n3790, in_13, gm_n157, gm_n58);
	not (gm_n3791, gm_n3790);
	nor (gm_n3792, gm_n853, gm_n136, gm_n104, gm_n3791, gm_n3789);
	and (gm_n3793, in_25, in_24, in_23);
	nand (gm_n3794, gm_n2229, in_26, gm_n82, gm_n3793, gm_n3792);
	nor (gm_n3795, gm_n2458, in_31, gm_n96, gm_n3794);
	nor (gm_n3796, gm_n221, in_16, gm_n157, gm_n553, gm_n222);
	nand (gm_n3797, gm_n196, in_24, in_20, gm_n3796, gm_n472);
	nor (gm_n3798, gm_n475, gm_n260, in_28, gm_n3797);
	nor (gm_n3799, gm_n103, gm_n72, in_16, gm_n1972, gm_n158);
	nand (gm_n3800, gm_n99, in_28, gm_n52, gm_n3799, gm_n220);
	nor (gm_n3801, gm_n3800, gm_n687);
	nor (gm_n3802, gm_n3801, gm_n3798, gm_n3795);
	not (gm_n3803, gm_n3802);
	nor (gm_n3804, gm_n244, gm_n68, in_12, gm_n2039, gm_n253);
	nand (gm_n3805, gm_n220, in_24, gm_n72, gm_n3804, gm_n230);
	nor (gm_n3806, gm_n687, gm_n80, in_28, gm_n3805);
	nand (gm_n3807, gm_n140, in_12, in_8, gm_n200, gm_n270);
	nor (gm_n3808, gm_n178, in_20, gm_n68, gm_n3807, gm_n179);
	nand (gm_n3809, gm_n220, in_28, in_24, gm_n3808, gm_n259);
	nor (gm_n3810, gm_n3809, gm_n268);
	and (gm_n3811, gm_n66, in_15, gm_n58, gm_n1543, gm_n938);
	and (gm_n3812, gm_n165, in_23, gm_n102, gm_n3811, gm_n299);
	and (gm_n3813, gm_n304, gm_n50, in_27, gm_n3812, gm_n393);
	nor (gm_n3814, gm_n3813, gm_n3810, gm_n3806);
	not (gm_n3815, gm_n3814);
	or (gm_n3816, gm_n3788, gm_n3668, gm_n3665, gm_n3815, gm_n3803);
	nand (gm_n3817, gm_n180, gm_n157, in_8, gm_n567, gm_n262);
	or (gm_n3818, gm_n504, in_20, in_16, gm_n3817, gm_n742);
	or (gm_n3819, gm_n84, in_28, gm_n52, gm_n3818, gm_n260);
	nor (gm_n3820, gm_n3819, gm_n268);
	and (gm_n3821, gm_n146, in_16, in_12, gm_n1337, gm_n147);
	and (gm_n3822, gm_n252, in_24, gm_n72, gm_n3821, gm_n269);
	and (gm_n3823, gm_n194, gm_n79, gm_n78, gm_n3822);
	and (gm_n3824, gm_n270, in_16, in_12, gm_n2970, gm_n198);
	and (gm_n3825, gm_n196, gm_n52, in_20, gm_n3824, gm_n517);
	and (gm_n3826, gm_n194, gm_n79, gm_n78, gm_n3825);
	nor (gm_n3827, gm_n3826, gm_n3823, gm_n3820);
	not (gm_n3828, gm_n3827);
	or (gm_n3829, in_17, gm_n68, in_15, gm_n851, gm_n136);
	nor (gm_n3830, gm_n485, in_26, in_22, gm_n3829, gm_n1903);
	nand (gm_n3831, gm_n50, in_30, in_27, gm_n3830, gm_n642);
	nand (gm_n3832, gm_n210, in_12, in_8, gm_n211, gm_n180);
	or (gm_n3833, gm_n504, gm_n72, in_16, gm_n3832, gm_n156);
	or (gm_n3834, gm_n216, gm_n78, gm_n52, gm_n3833, gm_n516);
	nor (gm_n3835, gm_n3834, gm_n132);
	nor (gm_n3836, gm_n57, in_15, gm_n58, gm_n2832, gm_n332);
	and (gm_n3837, gm_n173, in_23, gm_n102, gm_n3836, gm_n509);
	and (gm_n3838, gm_n339, in_31, in_27, gm_n3837);
	nor (gm_n3839, gm_n3838, gm_n3835);
	nand (gm_n3840, gm_n3839, gm_n3831);
	or (gm_n3841, gm_n3816, gm_n3662, gm_n3659, gm_n3840, gm_n3828);
	nor (gm_n3842, gm_n167, gm_n68, gm_n157, gm_n2556, gm_n168);
	nand (gm_n3843, gm_n219, in_24, gm_n72, gm_n3842, gm_n209);
	nor (gm_n3844, gm_n260, gm_n206, gm_n78, gm_n3843);
	nor (new_out4, gm_n3841, gm_n3656, gm_n3653, gm_n3844);
	and (gm_n3846, gm_n427, in_19, gm_n105, gm_n2005, gm_n452);
	and (gm_n3847, gm_n73, in_27, in_23, gm_n3846, gm_n173);
	and (gm_n3848, gm_n3847, gm_n677, gm_n50);
	and (gm_n3849, gm_n86, gm_n68, gm_n157, gm_n969, gm_n270);
	and (gm_n3850, gm_n220, gm_n52, gm_n72, gm_n3849, gm_n517);
	and (gm_n3851, gm_n207, gm_n194, in_28, gm_n3850);
	or (gm_n3852, gm_n57, gm_n105, gm_n58, gm_n880, gm_n432);
	nor (gm_n3853, gm_n300, gm_n195, in_19, gm_n3852, gm_n431);
	and (gm_n3854, gm_n455, gm_n50, in_27, gm_n3853, gm_n508);
	nor (gm_n3855, gm_n672, in_15, in_11, gm_n666, gm_n318);
	and (gm_n3856, gm_n361, gm_n195, in_19, gm_n3855, gm_n394);
	and (gm_n3857, gm_n55, gm_n50, in_27, gm_n3856, gm_n306);
	nor (gm_n3858, gm_n139, gm_n157, in_8, gm_n1533, gm_n167);
	nand (gm_n3859, gm_n219, gm_n72, gm_n68, gm_n3858, gm_n261);
	nor (gm_n3860, gm_n216, in_28, gm_n52, gm_n3859, gm_n687);
	or (gm_n3861, gm_n673, gm_n105, in_11, gm_n1214, gm_n576);
	or (gm_n3862, gm_n300, in_23, in_19, gm_n3861, gm_n337);
	nor (gm_n3863, gm_n51, in_31, gm_n133, gm_n3862, gm_n671);
	or (gm_n3864, gm_n119, in_15, gm_n58, gm_n2233, gm_n576);
	nor (gm_n3865, gm_n70, gm_n195, gm_n102, gm_n3864, gm_n1703);
	nand (gm_n3866, gm_n302, in_31, gm_n133, gm_n3865, gm_n508);
	nor (gm_n3867, gm_n57, gm_n105, gm_n58, gm_n992, gm_n618);
	nand (gm_n3868, gm_n293, in_23, gm_n102, gm_n3867, gm_n362);
	nor (gm_n3869, gm_n51, in_31, in_27, gm_n3868, gm_n983);
	or (gm_n3870, gm_n57, gm_n105, gm_n58, gm_n1227, gm_n119);
	or (gm_n3871, gm_n294, in_23, in_19, gm_n3870, gm_n395);
	nor (gm_n3872, gm_n575, gm_n50, in_27, gm_n3871, gm_n983);
	nor (gm_n3873, gm_n57, gm_n105, gm_n58, gm_n1266, gm_n673);
	nand (gm_n3874, gm_n293, in_23, gm_n102, gm_n3873, gm_n612);
	nor (gm_n3875, gm_n51, in_31, in_27, gm_n3874, gm_n1118);
	nor (gm_n3876, gm_n672, in_15, gm_n58, gm_n2390, gm_n363);
	nand (gm_n3877, gm_n165, in_23, in_19, gm_n3876, gm_n658);
	nor (gm_n3878, gm_n575, in_31, gm_n133, gm_n3877);
	or (gm_n3879, gm_n119, gm_n105, gm_n58, gm_n2283, gm_n576);
	or (gm_n3880, gm_n453, gm_n195, in_19, gm_n3879, gm_n510);
	nor (gm_n3881, gm_n581, in_31, gm_n133, gm_n3880, gm_n842);
	nor (gm_n3882, gm_n167, gm_n157, gm_n64, gm_n386, gm_n179);
	nand (gm_n3883, gm_n252, gm_n72, in_16, gm_n3882, gm_n269);
	nor (gm_n3884, gm_n243, gm_n78, in_24, gm_n3883, gm_n268);
	or (gm_n3885, gm_n673, gm_n105, in_11, gm_n620, gm_n399);
	or (gm_n3886, gm_n1703, in_23, in_19, gm_n3885, gm_n911);
	nor (gm_n3887, gm_n1118, gm_n50, in_27, gm_n3886, gm_n575);
	nand (gm_n3888, gm_n86, in_16, in_12, gm_n2018, gm_n341);
	or (gm_n3889, gm_n459, gm_n52, in_20, gm_n3888, gm_n412);
	nor (gm_n3890, gm_n176, gm_n80, in_28, gm_n3889);
	nand (gm_n3891, gm_n69, in_23, in_19, gm_n1112, gm_n73);
	nor (gm_n3892, gm_n983, in_31, gm_n133, gm_n3891, gm_n678);
	or (gm_n3893, gm_n3887, gm_n3884, gm_n3881, gm_n3892, gm_n3890);
	and (gm_n3894, gm_n1565, in_17, gm_n56, gm_n3309, gm_n2598);
	nand (gm_n3895, gm_n325, gm_n53, gm_n81, gm_n3894, gm_n1686);
	nor (gm_n3896, gm_n50, in_30, gm_n76, gm_n3895);
	nor (gm_n3897, gm_n432, in_15, in_11, gm_n583, gm_n366);
	nand (gm_n3898, gm_n293, in_23, in_19, gm_n3897, gm_n612);
	nor (gm_n3899, gm_n360, in_31, in_27, gm_n3898, gm_n983);
	nor (gm_n3900, gm_n295, gm_n942, gm_n64);
	nand (gm_n3901, gm_n146, gm_n68, gm_n157, gm_n3900, gm_n270);
	or (gm_n3902, gm_n804, gm_n52, gm_n72, gm_n3901, gm_n413);
	nor (gm_n3903, gm_n208, gm_n176, in_28, gm_n3902);
	or (gm_n3904, gm_n3903, gm_n3899, gm_n3896);
	nor (gm_n3905, gm_n504, gm_n68, in_12, gm_n3465, gm_n159);
	nand (gm_n3906, gm_n137, gm_n52, in_20, gm_n3905, gm_n209);
	nor (gm_n3907, gm_n243, gm_n229, in_28, gm_n3906);
	and (gm_n3908, gm_n146, in_12, in_8, gm_n1953, gm_n346);
	nand (gm_n3909, gm_n237, gm_n72, in_16, gm_n3908, gm_n183);
	nor (gm_n3910, gm_n208, in_28, in_24, gm_n3909, gm_n218);
	and (gm_n3911, gm_n231, gm_n68, gm_n157, gm_n2527, gm_n354);
	nand (gm_n3912, gm_n252, in_24, in_20, gm_n3911, gm_n269);
	nor (gm_n3913, gm_n687, gm_n208, in_28, gm_n3912);
	or (gm_n3914, gm_n3913, gm_n3910, gm_n3907);
	or (gm_n3915, gm_n3893, gm_n3878, gm_n3875, gm_n3914, gm_n3904);
	nand (gm_n3916, gm_n296, gm_n105, in_11, gm_n449, gm_n818);
	or (gm_n3917, gm_n117, gm_n195, gm_n102, gm_n3916, gm_n314);
	nor (gm_n3918, gm_n575, gm_n50, gm_n133, gm_n3917, gm_n983);
	and (gm_n3919, gm_n190, in_16, gm_n157, gm_n341, gm_n198);
	nand (gm_n3920, gm_n220, in_24, in_20, gm_n3919, gm_n269);
	nor (gm_n3921, gm_n371, gm_n268, gm_n78, gm_n3920);
	nor (gm_n3922, gm_n89, gm_n157, gm_n64, gm_n286, gm_n160);
	and (gm_n3923, gm_n86, gm_n72, gm_n68, gm_n3922, gm_n230);
	and (gm_n3924, gm_n177, gm_n78, in_24, gm_n3923, gm_n261);
	and (gm_n3925, gm_n3924, gm_n186);
	or (gm_n3926, gm_n3925, gm_n3921, gm_n3918);
	nor (gm_n3927, gm_n221, in_16, gm_n157, gm_n1889, gm_n286);
	nand (gm_n3928, gm_n261, gm_n52, in_20, gm_n3927, gm_n472);
	nor (gm_n3929, gm_n216, gm_n176, gm_n78, gm_n3928);
	and (gm_n3930, in_7, gm_n121, gm_n62, gm_n364, in_8);
	and (gm_n3931, gm_n147, gm_n68, in_12, gm_n3930, gm_n629);
	and (gm_n3932, gm_n196, in_24, gm_n72, gm_n3931, gm_n472);
	and (gm_n3933, gm_n462, gm_n205, gm_n78, gm_n3932);
	nor (gm_n3934, gm_n88, in_16, gm_n157, gm_n3390, gm_n158);
	nand (gm_n3935, gm_n219, gm_n52, in_20, gm_n3934, gm_n252);
	nor (gm_n3936, gm_n475, gm_n243, in_28, gm_n3935);
	or (gm_n3937, gm_n3936, gm_n3933, gm_n3929);
	nor (gm_n3938, gm_n3915, gm_n3872, gm_n3869, gm_n3937, gm_n3926);
	nand (gm_n3939, gm_n198, in_20, gm_n68, gm_n3710, gm_n230);
	nor (gm_n3940, gm_n80, in_28, in_24, gm_n3939, gm_n561);
	nand (gm_n3941, gm_n3940, gm_n186);
	nor (gm_n3942, gm_n396, in_15, gm_n58, gm_n2463, gm_n399);
	and (gm_n3943, gm_n73, gm_n195, gm_n102, gm_n3942, gm_n394);
	nand (gm_n3944, gm_n302, in_31, gm_n133, gm_n3943, gm_n392);
	nor (gm_n3945, gm_n395, gm_n102, in_15, gm_n2397, gm_n997);
	and (gm_n3946, gm_n313, gm_n133, gm_n195, gm_n3945, gm_n455);
	nand (gm_n3947, gm_n3946, gm_n115, gm_n50);
	nand (gm_n3948, gm_n3941, gm_n3938, gm_n3866, gm_n3947, gm_n3944);
	nor (gm_n3949, gm_n139, in_16, in_12, gm_n2077, gm_n159);
	nand (gm_n3950, gm_n237, gm_n52, in_20, gm_n3949, gm_n261);
	or (gm_n3951, gm_n206, gm_n80, gm_n78, gm_n3950);
	and (gm_n3952, gm_n333, gm_n105, gm_n58, gm_n449, gm_n334);
	nand (gm_n3953, gm_n126, gm_n195, in_19, gm_n3952, gm_n612);
	or (gm_n3954, gm_n581, gm_n50, gm_n133, gm_n3953, gm_n678);
	and (gm_n3955, gm_n63, in_12, in_8, gm_n232, gm_n211);
	nand (gm_n3956, gm_n629, in_20, gm_n68, gm_n3955, gm_n230);
	nor (gm_n3957, gm_n135, in_28, gm_n52, gm_n3956, gm_n561);
	nand (gm_n3958, gm_n3957, gm_n474);
	nand (gm_n3959, gm_n3958, gm_n3954, gm_n3951);
	or (gm_n3960, gm_n70, gm_n105, in_11, gm_n1537, gm_n366);
	nor (gm_n3961, gm_n1703, gm_n195, in_19, gm_n3960, gm_n617);
	nand (gm_n3962, gm_n392, gm_n50, in_27, gm_n3961);
	nand (gm_n3963, gm_n766, gm_n68, in_12, gm_n706, gm_n341);
	nor (gm_n3964, gm_n561, in_24, in_20, gm_n3963, gm_n602);
	nand (gm_n3965, gm_n474, gm_n462, gm_n78, gm_n3964);
	nand (gm_n3966, gm_n766, in_20, in_16, gm_n1619, gm_n472);
	nor (gm_n3967, gm_n84, in_28, in_24, gm_n3966, gm_n243);
	nand (gm_n3968, gm_n3967, gm_n186);
	nand (gm_n3969, gm_n3968, gm_n3965, gm_n3962);
	or (gm_n3970, gm_n3948, gm_n3863, gm_n3860, gm_n3969, gm_n3959);
	nor (gm_n3971, gm_n88, in_15, in_8, gm_n1039, gm_n622);
	nand (gm_n3972, gm_n582, gm_n195, gm_n102, gm_n3971, gm_n165);
	nor (gm_n3973, gm_n1118, in_31, gm_n133, gm_n3972, gm_n611);
	and (gm_n3974, gm_n333, gm_n105, gm_n58, gm_n2594, gm_n2776);
	nand (gm_n3975, gm_n293, gm_n195, in_19, gm_n3974, gm_n362);
	nor (gm_n3976, gm_n1231, gm_n50, gm_n133, gm_n3975, gm_n303);
	nand (gm_n3977, gm_n118, gm_n66, in_11, gm_n263, gm_n122);
	nor (gm_n3978, gm_n70, in_19, in_15, gm_n3977, gm_n314);
	nand (gm_n3979, gm_n304, in_27, in_23, gm_n3978, gm_n658);
	nor (gm_n3980, gm_n3979, gm_n50);
	nor (gm_n3981, gm_n3980, gm_n3976, gm_n3973);
	not (gm_n3982, gm_n3981);
	and (gm_n3983, gm_n612, gm_n346, in_15, gm_n758, gm_n621);
	nand (gm_n3984, gm_n173, gm_n195, in_19, gm_n3983, gm_n336);
	nor (gm_n3985, gm_n436, in_31, in_27, gm_n3984);
	nor (gm_n3986, gm_n88, gm_n68, in_12, gm_n2556, gm_n168);
	nand (gm_n3987, gm_n230, in_24, in_20, gm_n3986, gm_n261);
	nor (gm_n3988, gm_n206, gm_n80, gm_n78, gm_n3987);
	and (gm_n3989, gm_n147, gm_n157, gm_n64, gm_n403, gm_n511);
	nand (gm_n3990, gm_n1131, gm_n116, in_13, gm_n3989, gm_n2738);
	or (gm_n3991, gm_n2216, in_25, in_21, gm_n3990, gm_n1699);
	nor (gm_n3992, in_31, in_30, in_29, gm_n3991);
	nor (gm_n3993, gm_n3992, gm_n3988, gm_n3985);
	not (gm_n3994, gm_n3993);
	or (gm_n3995, gm_n3970, gm_n3857, gm_n3854, gm_n3994, gm_n3982);
	nand (gm_n3996, gm_n140, gm_n157, gm_n64, gm_n747, gm_n270);
	or (gm_n3997, gm_n187, in_20, gm_n68, gm_n3996, gm_n168);
	or (gm_n3998, gm_n243, gm_n78, in_24, gm_n3997, gm_n628);
	nor (gm_n3999, gm_n3998, gm_n229);
	nand (gm_n4000, gm_n231, in_20, gm_n68, gm_n1196, gm_n230);
	or (gm_n4001, gm_n628, in_28, gm_n52, gm_n4000, gm_n371);
	nor (gm_n4002, gm_n4001, gm_n132);
	nor (gm_n4003, gm_n244, gm_n68, in_12, gm_n588, gm_n88);
	and (gm_n4004, gm_n219, in_24, in_20, gm_n4003, gm_n220);
	and (gm_n4005, gm_n462, gm_n186, gm_n78, gm_n4004);
	nor (gm_n4006, gm_n4005, gm_n4002, gm_n3999);
	not (gm_n4007, gm_n4006);
	nor (gm_n4008, gm_n666, in_15, gm_n58, gm_n1664, gm_n997);
	nand (gm_n4009, gm_n69, gm_n195, gm_n102, gm_n4008, gm_n336);
	nor (gm_n4010, gm_n1118, gm_n50, gm_n133, gm_n4009, gm_n436);
	and (gm_n4011, gm_n333, gm_n105, gm_n58, gm_n1719, gm_n2776);
	and (gm_n4012, gm_n582, in_23, in_19, gm_n4011, gm_n361);
	and (gm_n4013, gm_n339, gm_n50, in_27, gm_n4012, gm_n455);
	nor (gm_n4014, gm_n504, in_12, in_8, gm_n1039, gm_n286);
	nand (gm_n4015, gm_n230, in_20, gm_n68, gm_n4014, gm_n252);
	nor (gm_n4016, gm_n176, in_28, in_24, gm_n4015, gm_n260);
	nor (gm_n4017, gm_n4016, gm_n4013, gm_n4010);
	not (gm_n4018, gm_n4017);
	or (gm_n4019, gm_n3995, gm_n3851, gm_n3848, gm_n4018, gm_n4007);
	and (gm_n4020, gm_n629, in_16, in_12, gm_n2212, gm_n354);
	nand (gm_n4021, gm_n220, in_24, in_20, gm_n4020, gm_n230);
	nor (gm_n4022, gm_n371, gm_n206, in_28, gm_n4021);
	or (gm_n4023, gm_n727, gm_n105, gm_n58, gm_n992, gm_n366);
	nor (gm_n4024, gm_n453, in_23, in_19, gm_n4023, gm_n510);
	nand (gm_n4025, gm_n339, in_31, gm_n133, gm_n4024, gm_n455);
	nand (gm_n4026, gm_n354, gm_n157, in_8, gm_n263, gm_n262);
	nor (gm_n4027, gm_n178, gm_n72, in_16, gm_n4026, gm_n139);
	nand (gm_n4028, gm_n207, in_28, in_24, gm_n4027, gm_n209);
	nor (gm_n4029, gm_n4028, gm_n229);
	nor (gm_n4030, gm_n106, in_16, gm_n157, gm_n1385, gm_n253);
	nand (gm_n4031, gm_n237, in_24, in_20, gm_n4030, gm_n183);
	nor (gm_n4032, gm_n206, gm_n80, gm_n78, gm_n4031);
	or (gm_n4033, gm_n618, gm_n105, gm_n58, gm_n1485, gm_n622);
	nor (gm_n4034, gm_n332, in_23, in_19, gm_n4033, gm_n314);
	nand (gm_n4035, gm_n306, in_31, gm_n133, gm_n4034, gm_n658);
	and (gm_n4036, gm_n63, in_12, in_8, gm_n619, gm_n180);
	nand (gm_n4037, gm_n85, gm_n72, gm_n68, gm_n4036, gm_n146);
	nor (gm_n4038, gm_n516, gm_n78, in_24, gm_n4037, gm_n371);
	nand (gm_n4039, gm_n4038, gm_n474);
	nor (gm_n4040, gm_n576, gm_n105, in_11, gm_n1806, gm_n319);
	nand (gm_n4041, gm_n165, in_23, in_19, gm_n4040, gm_n362);
	nor (gm_n4042, gm_n575, gm_n50, in_27, gm_n4041, gm_n983);
	nor (gm_n4043, gm_n106, gm_n68, gm_n157, gm_n3784, gm_n167);
	nand (gm_n4044, gm_n137, in_24, in_20, gm_n4043, gm_n196);
	nor (gm_n4045, gm_n475, gm_n135, gm_n78, gm_n4044);
	nor (gm_n4046, gm_n106, gm_n157, gm_n64, gm_n286, gm_n111);
	and (gm_n4047, gm_n237, gm_n72, in_16, gm_n4046, gm_n220);
	nand (gm_n4048, gm_n79, gm_n78, gm_n52, gm_n4047, gm_n492);
	nor (gm_n4049, gm_n57, gm_n102, gm_n105, gm_n1470, gm_n453);
	and (gm_n4050, gm_n293, gm_n133, in_23, gm_n4049, gm_n302);
	nand (gm_n4051, gm_n4050, gm_n304, gm_n50);
	or (gm_n4052, gm_n88, gm_n105, in_8, gm_n1039, gm_n576);
	nor (gm_n4053, gm_n300, in_23, gm_n102, gm_n4052, gm_n314);
	nand (gm_n4054, gm_n302, in_31, gm_n133, gm_n4053, gm_n508);
	or (gm_n4055, gm_n179, gm_n68, in_12, gm_n2060, gm_n253);
	nor (gm_n4056, gm_n156, in_24, in_20, gm_n4055, gm_n516);
	nand (gm_n4057, gm_n97, gm_n79, gm_n78, gm_n4056);
	and (gm_n4058, gm_n86, in_20, gm_n68, gm_n518, gm_n230);
	nand (gm_n4059, gm_n196, in_28, gm_n52, gm_n4058, gm_n259);
	nor (gm_n4060, gm_n4059, gm_n687);
	nor (gm_n4061, gm_n396, gm_n105, in_11, gm_n2233, gm_n426);
	nand (gm_n4062, gm_n69, in_23, gm_n102, gm_n4061, gm_n126);
	nor (gm_n4063, gm_n1118, in_31, gm_n133, gm_n4062, gm_n678);
	nor (gm_n4064, gm_n504, in_16, gm_n157, gm_n247, gm_n167);
	nand (gm_n4065, gm_n137, in_24, in_20, gm_n4064, gm_n220);
	nor (gm_n4066, gm_n260, gm_n218, gm_n78, gm_n4065);
	and (gm_n4067, gm_n498, gm_n511, in_8);
	and (gm_n4068, gm_n231, gm_n68, in_12, gm_n4067, gm_n346);
	nand (gm_n4069, gm_n196, in_24, in_20, gm_n4068, gm_n517);
	nor (gm_n4070, gm_n176, gm_n80, in_28, gm_n4069);
	and (gm_n4071, gm_n333, in_15, in_11, gm_n1683, gm_n665);
	and (gm_n4072, gm_n165, in_23, gm_n102, gm_n4071, gm_n362);
	and (gm_n4073, gm_n455, gm_n50, gm_n133, gm_n4072, gm_n677);
	nor (gm_n4074, gm_n4066, gm_n4063, gm_n4060, gm_n4073, gm_n4070);
	and (gm_n4075, gm_n482, gm_n136, in_14, gm_n3790, gm_n2894);
	nand (gm_n4076, gm_n2455, in_26, in_22, gm_n4075, gm_n3253);
	nor (gm_n4077, gm_n3779, in_31, gm_n96, gm_n4076);
	nor (gm_n4078, gm_n673, gm_n105, in_11, gm_n2855, gm_n622);
	nand (gm_n4079, gm_n165, in_23, gm_n102, gm_n4078, gm_n452);
	nor (gm_n4080, gm_n1231, gm_n50, gm_n133, gm_n4079, gm_n575);
	nor (gm_n4081, gm_n88, in_16, gm_n157, gm_n3646, gm_n106);
	nand (gm_n4082, gm_n83, in_24, gm_n72, gm_n4081, gm_n269);
	nor (gm_n4083, gm_n176, gm_n80, gm_n78, gm_n4082);
	nor (gm_n4084, gm_n4083, gm_n4080, gm_n4077);
	nand (gm_n4085, gm_n63, gm_n157, gm_n64, gm_n108, gm_n180);
	nor (gm_n4086, gm_n244, in_20, in_16, gm_n4085, gm_n103);
	nand (gm_n4087, gm_n196, gm_n78, in_24, gm_n4086, gm_n462);
	nor (gm_n4088, gm_n4087, gm_n229);
	nor (gm_n4089, gm_n396, gm_n105, in_11, gm_n997, gm_n583);
	nand (gm_n4090, gm_n166, in_23, in_19, gm_n4089, gm_n509);
	nor (gm_n4091, gm_n54, gm_n50, gm_n133, gm_n4090, gm_n678);
	nor (gm_n4092, gm_n156, in_20, gm_n68, gm_n1481, gm_n158);
	nand (gm_n4093, gm_n79, in_28, gm_n52, gm_n4092, gm_n252);
	nor (gm_n4094, gm_n4093, gm_n132);
	nor (gm_n4095, gm_n4094, gm_n4091, gm_n4088);
	and (gm_n4096, gm_n4074, gm_n4057, gm_n4054, gm_n4095, gm_n4084);
	nor (gm_n4097, gm_n426, in_15, in_11, gm_n1266, gm_n666);
	nand (gm_n4098, gm_n73, gm_n195, gm_n102, gm_n4097, gm_n299);
	nor (gm_n4099, gm_n54, gm_n50, in_27, gm_n4098, gm_n360);
	nor (gm_n4100, gm_n167, gm_n68, in_12, gm_n445, gm_n179);
	nand (gm_n4101, gm_n83, in_24, in_20, gm_n4100, gm_n269);
	nor (gm_n4102, gm_n132, gm_n216, gm_n78, gm_n4101);
	nor (gm_n4103, gm_n179, gm_n68, in_12, gm_n3118, gm_n286);
	nand (gm_n4104, gm_n261, gm_n52, in_20, gm_n4103, gm_n269);
	nor (gm_n4105, gm_n260, gm_n218, gm_n78, gm_n4104);
	nor (gm_n4106, gm_n4105, gm_n4102, gm_n4099);
	and (gm_n4107, gm_n189, gm_n68, in_12, gm_n2000, gm_n147);
	nand (gm_n4108, gm_n209, gm_n52, gm_n72, gm_n4107, gm_n517);
	nor (gm_n4109, gm_n268, gm_n135, gm_n78, gm_n4108);
	nor (gm_n4110, gm_n167, gm_n68, in_12, gm_n168, gm_n161);
	nand (gm_n4111, gm_n83, in_24, in_20, gm_n4110, gm_n269);
	nor (gm_n4112, gm_n216, gm_n176, gm_n78, gm_n4111);
	or (gm_n4113, gm_n159, gm_n157, in_8, gm_n347, gm_n271);
	nor (gm_n4114, gm_n103, gm_n72, gm_n68, gm_n4113, gm_n158);
	nand (gm_n4115, gm_n261, in_28, in_24, gm_n4114, gm_n370);
	nor (gm_n4116, gm_n4115, gm_n176);
	nor (gm_n4117, gm_n4116, gm_n4112, gm_n4109);
	nand (gm_n4118, gm_n4096, gm_n4051, gm_n4048, gm_n4117, gm_n4106);
	or (gm_n4119, gm_n88, gm_n68, in_12, gm_n748, gm_n504);
	nor (gm_n4120, gm_n197, gm_n52, in_20, gm_n4119, gm_n459);
	nand (gm_n4121, gm_n79, gm_n77, in_28, gm_n4120);
	or (gm_n4122, gm_n432, gm_n105, gm_n58, gm_n1086, gm_n366);
	nor (gm_n4123, gm_n117, gm_n195, in_19, gm_n4122, gm_n337);
	nand (gm_n4124, gm_n306, in_31, gm_n133, gm_n4123, gm_n393);
	nand (gm_n4125, gm_n86, gm_n68, gm_n157, gm_n3900, gm_n346);
	nor (gm_n4126, gm_n178, gm_n52, gm_n72, gm_n4125, gm_n628);
	nand (gm_n4127, gm_n207, gm_n205, in_28, gm_n4126);
	nand (gm_n4128, gm_n4127, gm_n4124, gm_n4121);
	nand (gm_n4129, gm_n405, gm_n116, in_13, gm_n3406, gm_n406);
	nor (gm_n4130, gm_n152, gm_n53, gm_n81, gm_n4129, gm_n328);
	nand (gm_n4131, in_31, in_30, gm_n76, gm_n4130);
	nand (gm_n4132, gm_n147, in_16, gm_n157, gm_n630, gm_n198);
	nor (gm_n4133, gm_n187, gm_n52, gm_n72, gm_n4132, gm_n804);
	nand (gm_n4134, gm_n492, gm_n99, in_28, gm_n4133);
	nand (gm_n4135, gm_n188, gm_n68, in_12, gm_n758, gm_n766);
	nor (gm_n4136, gm_n187, in_24, gm_n72, gm_n4135, gm_n561);
	nand (gm_n4137, gm_n186, gm_n177, gm_n78, gm_n4136);
	nand (gm_n4138, gm_n4137, gm_n4134, gm_n4131);
	nor (gm_n4139, gm_n4118, gm_n4045, gm_n4042, gm_n4138, gm_n4128);
	nor (gm_n4140, gm_n159, in_16, gm_n157, gm_n902, gm_n221);
	nand (gm_n4141, gm_n230, in_24, in_20, gm_n4140, gm_n261);
	nor (gm_n4142, gm_n218, gm_n135, gm_n78, gm_n4141);
	nand (gm_n4143, gm_n188, gm_n157, in_8, gm_n747, gm_n262);
	nor (gm_n4144, gm_n179, gm_n72, in_16, gm_n4143, gm_n413);
	nand (gm_n4145, gm_n83, gm_n78, gm_n52, gm_n4144, gm_n134);
	nor (gm_n4146, gm_n4145, gm_n475);
	nor (gm_n4147, gm_n88, gm_n68, in_12, gm_n1643, gm_n221);
	nand (gm_n4148, gm_n85, in_24, in_20, gm_n4147, gm_n196);
	nor (gm_n4149, gm_n687, gm_n80, in_28, gm_n4148);
	nor (gm_n4150, gm_n4149, gm_n4146, gm_n4142);
	nand (gm_n4151, gm_n361, in_23, in_19, gm_n2255, gm_n362);
	nor (gm_n4152, gm_n1118, in_31, in_27, gm_n4151, gm_n575);
	and (gm_n4153, gm_n297, in_15, in_11, gm_n1758, gm_n621);
	nand (gm_n4154, gm_n166, in_23, gm_n102, gm_n4153, gm_n313);
	nor (gm_n4155, gm_n1231, in_31, gm_n133, gm_n4154, gm_n842);
	nor (gm_n4156, gm_n139, gm_n68, gm_n157, gm_n692, gm_n222);
	nand (gm_n4157, gm_n137, in_24, gm_n72, gm_n4156, gm_n252);
	nor (gm_n4158, gm_n206, gm_n216, gm_n78, gm_n4157);
	nor (gm_n4159, gm_n4158, gm_n4155, gm_n4152);
	nand (gm_n4160, gm_n4139, gm_n4039, gm_n4035, gm_n4159, gm_n4150);
	nand (gm_n4161, gm_n188, in_16, in_12, gm_n414, gm_n629);
	nor (gm_n4162, gm_n101, gm_n52, in_20, gm_n4161, gm_n178);
	nand (gm_n4163, gm_n194, gm_n99, gm_n78, gm_n4162);
	or (gm_n4164, gm_n672, gm_n105, in_11, gm_n318, gm_n119);
	nor (gm_n4165, gm_n423, gm_n195, gm_n102, gm_n4164, gm_n911);
	nand (gm_n4166, gm_n129, in_31, gm_n133, gm_n4165, gm_n392);
	nand (gm_n4167, gm_n86, in_16, gm_n157, gm_n2612, gm_n180);
	nor (gm_n4168, gm_n804, in_24, gm_n72, gm_n4167, gm_n742);
	nand (gm_n4169, gm_n134, gm_n194, gm_n78, gm_n4168);
	nand (gm_n4170, gm_n4169, gm_n4166, gm_n4163);
	nand (gm_n4171, gm_n231, in_16, gm_n157, gm_n4067, gm_n341);
	nor (gm_n4172, gm_n156, in_24, in_20, gm_n4171, gm_n516);
	nand (gm_n4173, gm_n207, gm_n97, gm_n78, gm_n4172);
	nor (gm_n4174, gm_n119, in_15, in_11, gm_n1001, gm_n426);
	nand (gm_n4175, gm_n293, gm_n195, gm_n102, gm_n4174, gm_n299);
	or (gm_n4176, gm_n617, gm_n50, gm_n133, gm_n4175, gm_n436);
	and (gm_n4177, gm_n147, gm_n68, in_12, gm_n785, gm_n629);
	nand (gm_n4178, gm_n237, gm_n52, in_20, gm_n4177, gm_n220);
	or (gm_n4179, gm_n260, gm_n268, gm_n78, gm_n4178);
	nand (gm_n4180, gm_n4179, gm_n4176, gm_n4173);
	nor (gm_n4181, gm_n4160, gm_n4032, gm_n4029, gm_n4180, gm_n4170);
	or (gm_n4182, gm_n67, in_19, in_15, gm_n399, gm_n332);
	nor (gm_n4183, gm_n617, gm_n133, in_23, gm_n4182, gm_n314);
	nand (gm_n4184, gm_n4183, gm_n508, gm_n50);
	nor (gm_n4185, gm_n179, in_16, gm_n157, gm_n287, gm_n222);
	nand (gm_n4186, gm_n137, gm_n52, in_20, gm_n4185, gm_n261);
	or (gm_n4187, gm_n208, gm_n176, in_28, gm_n4186);
	nand (gm_n4188, gm_n231, in_16, gm_n157, gm_n466, gm_n346);
	nor (gm_n4189, gm_n516, gm_n52, in_20, gm_n4188, gm_n602);
	nand (gm_n4190, gm_n370, gm_n97, in_28, gm_n4189);
	nand (gm_n4191, gm_n4184, gm_n4181, gm_n4025, gm_n4190, gm_n4187);
	and (gm_n4192, gm_n404, in_17, gm_n56, gm_n1183, gm_n406);
	and (gm_n4193, gm_n3494, gm_n53, gm_n81, gm_n4192, gm_n738);
	and (gm_n4194, in_31, in_30, in_29, gm_n4193);
	nor (new_out5, gm_n4191, gm_n4022, gm_n4019, gm_n4194);
	or (gm_n4196, new_out5, new_out4);
	nand (new_out1, gm_n4196, gm_n3480);
endmodule
